module basic_5000_50000_5000_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_1543,In_31);
nor U1 (N_1,In_2535,In_4440);
nand U2 (N_2,In_4422,In_3043);
or U3 (N_3,In_3329,In_3522);
and U4 (N_4,In_2008,In_731);
nor U5 (N_5,In_2023,In_3352);
or U6 (N_6,In_4643,In_2701);
nor U7 (N_7,In_4070,In_249);
and U8 (N_8,In_4009,In_1575);
or U9 (N_9,In_2926,In_2239);
and U10 (N_10,In_3242,In_4095);
xnor U11 (N_11,In_3478,In_3519);
and U12 (N_12,In_614,In_3729);
and U13 (N_13,In_3597,In_2253);
and U14 (N_14,In_587,In_3592);
nand U15 (N_15,In_1091,In_2897);
nand U16 (N_16,In_2922,In_180);
nor U17 (N_17,In_601,In_357);
nand U18 (N_18,In_1950,In_910);
xnor U19 (N_19,In_4029,In_2295);
and U20 (N_20,In_4937,In_2579);
nor U21 (N_21,In_2268,In_4894);
nand U22 (N_22,In_1327,In_1560);
nand U23 (N_23,In_1992,In_1365);
or U24 (N_24,In_4186,In_2000);
nor U25 (N_25,In_4544,In_3145);
nand U26 (N_26,In_4997,In_3573);
or U27 (N_27,In_2675,In_632);
nand U28 (N_28,In_3792,In_2123);
nor U29 (N_29,In_128,In_3552);
xor U30 (N_30,In_2471,In_45);
nand U31 (N_31,In_3765,In_4063);
or U32 (N_32,In_4588,In_2717);
nand U33 (N_33,In_3001,In_3927);
nand U34 (N_34,In_1624,In_2519);
xor U35 (N_35,In_2198,In_2248);
nor U36 (N_36,In_3018,In_2040);
nor U37 (N_37,In_1240,In_1746);
nand U38 (N_38,In_1810,In_4781);
and U39 (N_39,In_2937,In_1233);
nand U40 (N_40,In_4494,In_774);
nor U41 (N_41,In_4188,In_941);
nand U42 (N_42,In_1069,In_87);
nor U43 (N_43,In_4858,In_2709);
or U44 (N_44,In_2284,In_7);
or U45 (N_45,In_1200,In_4496);
nor U46 (N_46,In_257,In_695);
and U47 (N_47,In_4832,In_3159);
xnor U48 (N_48,In_3098,In_3425);
or U49 (N_49,In_426,In_531);
nand U50 (N_50,In_2467,In_3095);
nor U51 (N_51,In_3545,In_1550);
nand U52 (N_52,In_3643,In_3735);
nor U53 (N_53,In_1863,In_4108);
nor U54 (N_54,In_2898,In_942);
and U55 (N_55,In_1479,In_2447);
nor U56 (N_56,In_1786,In_562);
and U57 (N_57,In_3548,In_3977);
nand U58 (N_58,In_276,In_2732);
nand U59 (N_59,In_550,In_1457);
nor U60 (N_60,In_4033,In_1370);
or U61 (N_61,In_584,In_2708);
or U62 (N_62,In_3233,In_4181);
nor U63 (N_63,In_3166,In_3534);
nor U64 (N_64,In_2165,In_3035);
and U65 (N_65,In_4110,In_501);
nor U66 (N_66,In_3564,In_1164);
nor U67 (N_67,In_1683,In_103);
nand U68 (N_68,In_4721,In_1274);
and U69 (N_69,In_2992,In_1173);
nand U70 (N_70,In_3569,In_1596);
or U71 (N_71,In_4048,In_4268);
nor U72 (N_72,In_1836,In_3361);
nand U73 (N_73,In_4003,In_311);
and U74 (N_74,In_3997,In_2084);
or U75 (N_75,In_681,In_3720);
or U76 (N_76,In_2612,In_3669);
nor U77 (N_77,In_4325,In_1617);
nand U78 (N_78,In_2729,In_2779);
nor U79 (N_79,In_3746,In_3183);
nor U80 (N_80,In_2644,In_4207);
and U81 (N_81,In_3324,In_2416);
or U82 (N_82,In_838,In_1696);
nor U83 (N_83,In_341,In_3533);
nand U84 (N_84,In_2459,In_4375);
xor U85 (N_85,In_1237,In_860);
and U86 (N_86,In_736,In_3126);
nor U87 (N_87,In_2391,In_3524);
nand U88 (N_88,In_4730,In_1954);
and U89 (N_89,In_2403,In_4983);
xnor U90 (N_90,In_56,In_3815);
or U91 (N_91,In_4550,In_3882);
nor U92 (N_92,In_3933,In_4545);
and U93 (N_93,In_1217,In_3479);
nand U94 (N_94,In_592,In_3827);
nand U95 (N_95,In_1480,In_4501);
nor U96 (N_96,In_42,In_4819);
nor U97 (N_97,In_145,In_168);
and U98 (N_98,In_793,In_2134);
and U99 (N_99,In_3283,In_4514);
nand U100 (N_100,In_3468,In_1724);
or U101 (N_101,In_189,In_4265);
xnor U102 (N_102,In_1887,In_4384);
nor U103 (N_103,In_2113,In_1962);
nand U104 (N_104,In_1466,In_298);
xnor U105 (N_105,In_856,In_3794);
and U106 (N_106,In_2027,In_1459);
nor U107 (N_107,In_210,In_205);
nand U108 (N_108,In_2370,In_1875);
or U109 (N_109,In_4951,In_797);
nand U110 (N_110,In_2074,In_89);
nor U111 (N_111,In_1559,In_2563);
or U112 (N_112,In_1495,In_4124);
nand U113 (N_113,In_2028,In_1698);
and U114 (N_114,In_4910,In_1305);
nand U115 (N_115,In_2648,In_229);
nor U116 (N_116,In_214,In_3508);
nor U117 (N_117,In_2301,In_4293);
nand U118 (N_118,In_1901,In_1022);
nand U119 (N_119,In_3893,In_1941);
xnor U120 (N_120,In_783,In_1717);
and U121 (N_121,In_256,In_980);
or U122 (N_122,In_1801,In_381);
nor U123 (N_123,In_3038,In_3347);
xnor U124 (N_124,In_3976,In_4764);
or U125 (N_125,In_561,In_4513);
and U126 (N_126,In_2322,In_3574);
nor U127 (N_127,In_325,In_3915);
xor U128 (N_128,In_4974,In_4453);
nor U129 (N_129,In_3682,In_4470);
and U130 (N_130,In_4150,In_2182);
nand U131 (N_131,In_4465,In_1910);
and U132 (N_132,In_1018,In_4392);
and U133 (N_133,In_96,In_4237);
or U134 (N_134,In_3611,In_3202);
or U135 (N_135,In_2629,In_261);
and U136 (N_136,In_2397,In_4649);
xnor U137 (N_137,In_4799,In_2367);
or U138 (N_138,In_2196,In_2238);
xnor U139 (N_139,In_4370,In_1672);
nor U140 (N_140,In_4895,In_2410);
and U141 (N_141,In_2394,In_2858);
nand U142 (N_142,In_3481,In_3435);
and U143 (N_143,In_3723,In_369);
and U144 (N_144,In_4787,In_2161);
nand U145 (N_145,In_3620,In_484);
nor U146 (N_146,In_4510,In_2310);
and U147 (N_147,In_1636,In_1158);
nor U148 (N_148,In_901,In_4835);
or U149 (N_149,In_3251,In_643);
nor U150 (N_150,In_4023,In_1354);
and U151 (N_151,In_1519,In_3871);
nand U152 (N_152,In_1730,In_1140);
nand U153 (N_153,In_1947,In_4404);
or U154 (N_154,In_1278,In_861);
and U155 (N_155,In_4930,In_4248);
or U156 (N_156,In_3424,In_4612);
and U157 (N_157,In_4230,In_1774);
and U158 (N_158,In_894,In_3045);
and U159 (N_159,In_3239,In_2057);
and U160 (N_160,In_2460,In_480);
nor U161 (N_161,In_641,In_2334);
or U162 (N_162,In_1852,In_1264);
nand U163 (N_163,In_30,In_2090);
or U164 (N_164,In_3998,In_3231);
nor U165 (N_165,In_613,In_2339);
nor U166 (N_166,In_1858,In_599);
nand U167 (N_167,In_2044,In_4302);
nand U168 (N_168,In_905,In_4251);
or U169 (N_169,In_3816,In_20);
nand U170 (N_170,In_2250,In_4802);
or U171 (N_171,In_3865,In_2792);
and U172 (N_172,In_230,In_1433);
xor U173 (N_173,In_4255,In_1716);
nand U174 (N_174,In_2808,In_1361);
and U175 (N_175,In_3559,In_2225);
and U176 (N_176,In_2585,In_4814);
and U177 (N_177,In_4319,In_3858);
and U178 (N_178,In_3078,In_4776);
or U179 (N_179,In_3629,In_3623);
nor U180 (N_180,In_2895,In_4449);
nor U181 (N_181,In_78,In_1690);
nand U182 (N_182,In_1899,In_1455);
nor U183 (N_183,In_3172,In_945);
and U184 (N_184,In_4932,In_589);
nor U185 (N_185,In_1651,In_2480);
or U186 (N_186,In_4722,In_4693);
or U187 (N_187,In_1053,In_2744);
nand U188 (N_188,In_3909,In_1854);
nand U189 (N_189,In_2829,In_2303);
nand U190 (N_190,In_4523,In_2277);
or U191 (N_191,In_3773,In_4542);
nor U192 (N_192,In_1300,In_3897);
nand U193 (N_193,In_2029,In_1921);
nor U194 (N_194,In_760,In_3455);
nand U195 (N_195,In_3895,In_3475);
and U196 (N_196,In_2313,In_1086);
or U197 (N_197,In_3550,In_1824);
nand U198 (N_198,In_3614,In_383);
nor U199 (N_199,In_3843,In_4535);
and U200 (N_200,In_1039,In_799);
xor U201 (N_201,In_2135,In_3512);
nand U202 (N_202,In_3171,In_2032);
nand U203 (N_203,In_687,In_4130);
nand U204 (N_204,In_3131,In_2521);
or U205 (N_205,In_102,In_2879);
nor U206 (N_206,In_2620,In_4236);
or U207 (N_207,In_3841,In_2826);
nor U208 (N_208,In_1268,In_519);
xor U209 (N_209,In_1750,In_2232);
nand U210 (N_210,In_1833,In_4675);
or U211 (N_211,In_4143,In_2331);
and U212 (N_212,In_4843,In_2107);
xor U213 (N_213,In_3802,In_3096);
nor U214 (N_214,In_663,In_1190);
or U215 (N_215,In_4847,In_1007);
nor U216 (N_216,In_3007,In_2414);
nor U217 (N_217,In_1737,In_4196);
and U218 (N_218,In_404,In_367);
nor U219 (N_219,In_4264,In_1449);
or U220 (N_220,In_3063,In_4120);
and U221 (N_221,In_326,In_2933);
xnor U222 (N_222,In_3907,In_3293);
nand U223 (N_223,In_2121,In_4398);
nand U224 (N_224,In_4304,In_4443);
or U225 (N_225,In_3103,In_2260);
and U226 (N_226,In_127,In_594);
or U227 (N_227,In_4957,In_3327);
nor U228 (N_228,In_1520,In_1827);
nor U229 (N_229,In_242,In_224);
or U230 (N_230,In_2589,In_4041);
and U231 (N_231,In_4706,In_4679);
and U232 (N_232,In_2236,In_3889);
nand U233 (N_233,In_1556,In_4518);
or U234 (N_234,In_3292,In_4968);
nor U235 (N_235,In_883,In_3957);
nor U236 (N_236,In_3396,In_2346);
nand U237 (N_237,In_3679,In_4429);
or U238 (N_238,In_4272,In_4418);
nand U239 (N_239,In_1676,In_302);
nor U240 (N_240,In_1333,In_604);
or U241 (N_241,In_3453,In_694);
and U242 (N_242,In_4849,In_2466);
nor U243 (N_243,In_3608,In_50);
and U244 (N_244,In_4378,In_1679);
nor U245 (N_245,In_2559,In_285);
or U246 (N_246,In_2674,In_4395);
and U247 (N_247,In_3951,In_1630);
and U248 (N_248,In_3141,In_204);
xor U249 (N_249,In_2477,In_2944);
xnor U250 (N_250,In_2246,In_2583);
and U251 (N_251,In_3551,In_1882);
nor U252 (N_252,In_977,In_4360);
xor U253 (N_253,In_1198,In_824);
nor U254 (N_254,In_958,In_4623);
nor U255 (N_255,In_3437,In_1869);
and U256 (N_256,In_585,In_4493);
and U257 (N_257,In_473,In_407);
and U258 (N_258,In_1095,In_837);
xnor U259 (N_259,In_3111,In_4235);
or U260 (N_260,In_3199,In_263);
nand U261 (N_261,In_3780,In_672);
or U262 (N_262,In_4636,In_4328);
and U263 (N_263,In_2386,In_4482);
or U264 (N_264,In_4904,In_17);
nor U265 (N_265,In_4936,In_2622);
or U266 (N_266,In_1471,In_1841);
and U267 (N_267,In_76,In_4618);
and U268 (N_268,In_4458,In_1865);
nand U269 (N_269,In_999,In_1631);
nor U270 (N_270,In_1031,In_3644);
nand U271 (N_271,In_4401,In_2125);
nand U272 (N_272,In_4277,In_3579);
and U273 (N_273,In_4833,In_2691);
nand U274 (N_274,In_4317,In_1891);
xor U275 (N_275,In_260,In_4890);
nor U276 (N_276,In_468,In_4354);
and U277 (N_277,In_2288,In_676);
nor U278 (N_278,In_548,In_1171);
nand U279 (N_279,In_3712,In_1736);
and U280 (N_280,In_2593,In_90);
or U281 (N_281,In_4955,In_4755);
or U282 (N_282,In_4363,In_379);
or U283 (N_283,In_1979,In_2124);
nand U284 (N_284,In_1501,In_122);
xor U285 (N_285,In_1502,In_1983);
nor U286 (N_286,In_829,In_2813);
or U287 (N_287,In_1016,In_3822);
or U288 (N_288,In_2531,In_1915);
and U289 (N_289,In_3866,In_2856);
xnor U290 (N_290,In_2984,In_105);
nor U291 (N_291,In_3959,In_679);
and U292 (N_292,In_979,In_2538);
nor U293 (N_293,In_3394,In_2671);
and U294 (N_294,In_4024,In_1211);
and U295 (N_295,In_3810,In_3986);
or U296 (N_296,In_823,In_2417);
and U297 (N_297,In_2553,In_2876);
nand U298 (N_298,In_3404,In_4123);
nor U299 (N_299,In_1082,In_1371);
or U300 (N_300,In_343,In_795);
nor U301 (N_301,In_4768,In_1425);
and U302 (N_302,In_4362,In_3116);
and U303 (N_303,In_524,In_2696);
or U304 (N_304,In_1710,In_1830);
nor U305 (N_305,In_2363,In_4498);
nor U306 (N_306,In_2734,In_2643);
nor U307 (N_307,In_3743,In_3916);
or U308 (N_308,In_3681,In_2490);
nor U309 (N_309,In_2603,In_2037);
or U310 (N_310,In_857,In_2136);
nor U311 (N_311,In_3088,In_4943);
and U312 (N_312,In_1911,In_904);
nor U313 (N_313,In_2050,In_3408);
nor U314 (N_314,In_1285,In_2966);
and U315 (N_315,In_3304,In_3776);
and U316 (N_316,In_401,In_4775);
nor U317 (N_317,In_4221,In_3747);
nor U318 (N_318,In_4146,In_3006);
nor U319 (N_319,In_665,In_2081);
and U320 (N_320,In_4558,In_4083);
and U321 (N_321,In_4045,In_3835);
nand U322 (N_322,In_1959,In_259);
and U323 (N_323,In_2989,In_2968);
or U324 (N_324,In_3325,In_4305);
or U325 (N_325,In_3617,In_2349);
or U326 (N_326,In_953,In_4137);
nand U327 (N_327,In_3092,In_2633);
and U328 (N_328,In_1020,In_464);
and U329 (N_329,In_1689,In_395);
xnor U330 (N_330,In_2767,In_1430);
nand U331 (N_331,In_3788,In_3060);
nor U332 (N_332,In_3008,In_408);
xnor U333 (N_333,In_2783,In_218);
nand U334 (N_334,In_3728,In_3232);
nor U335 (N_335,In_2690,In_2951);
nor U336 (N_336,In_37,In_4871);
nor U337 (N_337,In_738,In_3590);
nor U338 (N_338,In_606,In_4416);
and U339 (N_339,In_2427,In_2833);
or U340 (N_340,In_3384,In_3253);
nand U341 (N_341,In_1837,In_3647);
and U342 (N_342,In_745,In_1493);
nor U343 (N_343,In_130,In_2372);
nor U344 (N_344,In_4313,In_4244);
nor U345 (N_345,In_1044,In_845);
or U346 (N_346,In_3848,In_1913);
or U347 (N_347,In_4187,In_2104);
nand U348 (N_348,In_339,In_833);
nor U349 (N_349,In_3108,In_4393);
nor U350 (N_350,In_4134,In_471);
nor U351 (N_351,In_2980,In_1212);
or U352 (N_352,In_2264,In_4719);
nand U353 (N_353,In_4477,In_1613);
and U354 (N_354,In_669,In_988);
nor U355 (N_355,In_4136,In_4076);
and U356 (N_356,In_110,In_792);
and U357 (N_357,In_1666,In_3488);
nor U358 (N_358,In_1360,In_2814);
xor U359 (N_359,In_3932,In_1350);
and U360 (N_360,In_616,In_216);
xnor U361 (N_361,In_2927,In_2375);
nand U362 (N_362,In_418,In_3892);
nor U363 (N_363,In_3264,In_2498);
nand U364 (N_364,In_3021,In_3138);
or U365 (N_365,In_3279,In_1450);
or U366 (N_366,In_2591,In_3791);
or U367 (N_367,In_577,In_27);
nor U368 (N_368,In_3881,In_2166);
and U369 (N_369,In_1778,In_2619);
or U370 (N_370,In_2496,In_3803);
nand U371 (N_371,In_3817,In_1184);
nand U372 (N_372,In_3041,In_2736);
nor U373 (N_373,In_3595,In_2442);
or U374 (N_374,In_4850,In_314);
and U375 (N_375,In_3527,In_3276);
and U376 (N_376,In_95,In_3255);
or U377 (N_377,In_545,In_2906);
and U378 (N_378,In_1551,In_3888);
nand U379 (N_379,In_1318,In_4778);
and U380 (N_380,In_3715,In_2598);
or U381 (N_381,In_3499,In_3302);
or U382 (N_382,In_2321,In_4281);
xor U383 (N_383,In_1826,In_4984);
nor U384 (N_384,In_2474,In_1168);
or U385 (N_385,In_826,In_382);
nand U386 (N_386,In_1831,In_771);
nor U387 (N_387,In_516,In_2841);
or U388 (N_388,In_2302,In_3646);
nand U389 (N_389,In_3901,In_1050);
nand U390 (N_390,In_44,In_1435);
nor U391 (N_391,In_4297,In_162);
and U392 (N_392,In_2625,In_4674);
or U393 (N_393,In_491,In_2673);
nor U394 (N_394,In_1374,In_3645);
nor U395 (N_395,In_4665,In_902);
or U396 (N_396,In_2497,In_1423);
nor U397 (N_397,In_459,In_2790);
or U398 (N_398,In_6,In_2365);
nand U399 (N_399,In_926,In_3105);
nand U400 (N_400,In_4352,In_855);
and U401 (N_401,In_3049,In_207);
nor U402 (N_402,In_1150,In_4026);
nor U403 (N_403,In_441,In_2602);
nand U404 (N_404,In_1533,In_4089);
and U405 (N_405,In_363,In_2835);
nor U406 (N_406,In_4232,In_807);
nand U407 (N_407,In_2065,In_965);
nand U408 (N_408,In_2749,In_3365);
nor U409 (N_409,In_898,In_847);
xnor U410 (N_410,In_2069,In_754);
and U411 (N_411,In_1186,In_3401);
or U412 (N_412,In_1578,In_1598);
nand U413 (N_413,In_1581,In_2942);
or U414 (N_414,In_115,In_4011);
nor U415 (N_415,In_3149,In_4896);
xnor U416 (N_416,In_3767,In_4807);
or U417 (N_417,In_1605,In_3785);
nor U418 (N_418,In_1013,In_1194);
and U419 (N_419,In_2621,In_3946);
xnor U420 (N_420,In_3017,In_1848);
and U421 (N_421,In_4901,In_3502);
or U422 (N_422,In_3867,In_1092);
or U423 (N_423,In_2382,In_2282);
or U424 (N_424,In_1110,In_2839);
or U425 (N_425,In_4096,In_4864);
xor U426 (N_426,In_36,In_1484);
nor U427 (N_427,In_3062,In_2796);
and U428 (N_428,In_2594,In_2635);
xnor U429 (N_429,In_3459,In_1195);
nor U430 (N_430,In_2969,In_2351);
nand U431 (N_431,In_332,In_3358);
or U432 (N_432,In_2094,In_2290);
nand U433 (N_433,In_4891,In_3616);
or U434 (N_434,In_1342,In_4050);
nand U435 (N_435,In_1603,In_2706);
xor U436 (N_436,In_3194,In_3245);
or U437 (N_437,In_729,In_2784);
nand U438 (N_438,In_213,In_1106);
xor U439 (N_439,In_1059,In_1974);
nand U440 (N_440,In_1375,In_1135);
or U441 (N_441,In_758,In_2011);
and U442 (N_442,In_2838,In_3683);
xor U443 (N_443,In_876,In_4999);
nand U444 (N_444,In_2507,In_3718);
or U445 (N_445,In_3982,In_1832);
or U446 (N_446,In_4691,In_1440);
or U447 (N_447,In_3263,In_3371);
nand U448 (N_448,In_3772,In_3412);
nor U449 (N_449,In_2994,In_3570);
nand U450 (N_450,In_4065,In_3553);
and U451 (N_451,In_291,In_1406);
xor U452 (N_452,In_3197,In_2005);
and U453 (N_453,In_2546,In_3709);
or U454 (N_454,In_3870,In_2751);
and U455 (N_455,In_3000,In_990);
or U456 (N_456,In_1482,In_234);
or U457 (N_457,In_3262,In_1469);
xor U458 (N_458,In_4341,In_503);
nand U459 (N_459,In_1614,In_4229);
nand U460 (N_460,In_3082,In_4824);
nor U461 (N_461,In_4872,In_3167);
or U462 (N_462,In_2097,In_921);
nor U463 (N_463,In_3985,In_1096);
nand U464 (N_464,In_664,In_4042);
xor U465 (N_465,In_4876,In_843);
nor U466 (N_466,In_618,In_2383);
nand U467 (N_467,In_1756,In_2388);
and U468 (N_468,In_4223,In_4817);
or U469 (N_469,In_4001,In_542);
or U470 (N_470,In_1409,In_1668);
and U471 (N_471,In_209,In_4756);
xor U472 (N_472,In_2482,In_2340);
nor U473 (N_473,In_4147,In_4348);
nor U474 (N_474,In_57,In_1635);
and U475 (N_475,In_2186,In_3537);
nor U476 (N_476,In_1369,In_3168);
and U477 (N_477,In_1294,In_1105);
and U478 (N_478,In_1973,In_3080);
or U479 (N_479,In_2806,In_4758);
nor U480 (N_480,In_2568,In_198);
or U481 (N_481,In_174,In_4502);
and U482 (N_482,In_3156,In_3447);
nor U483 (N_483,In_831,In_1052);
or U484 (N_484,In_4812,In_3055);
and U485 (N_485,In_3594,In_19);
or U486 (N_486,In_2974,In_4680);
nor U487 (N_487,In_4028,In_1846);
xnor U488 (N_488,In_2529,In_4972);
and U489 (N_489,In_2586,In_4073);
and U490 (N_490,In_2430,In_4668);
and U491 (N_491,In_569,In_3762);
nor U492 (N_492,In_4438,In_2857);
xor U493 (N_493,In_2923,In_4785);
and U494 (N_494,In_3529,In_3831);
nor U495 (N_495,In_971,In_324);
nor U496 (N_496,In_289,In_3600);
and U497 (N_497,In_2925,In_2893);
or U498 (N_498,In_368,In_2170);
nor U499 (N_499,In_1647,In_4642);
nand U500 (N_500,In_267,In_4918);
or U501 (N_501,In_109,In_3355);
and U502 (N_502,In_4818,In_3217);
and U503 (N_503,In_2797,In_3993);
nand U504 (N_504,In_3072,In_3676);
and U505 (N_505,In_4049,In_1664);
nor U506 (N_506,In_4877,In_2722);
nor U507 (N_507,In_22,In_2574);
nor U508 (N_508,In_2399,In_430);
and U509 (N_509,In_1427,In_3994);
nand U510 (N_510,In_2667,In_1707);
nor U511 (N_511,In_1989,In_711);
xnor U512 (N_512,In_3813,In_2009);
nor U513 (N_513,In_1993,In_485);
or U514 (N_514,In_4640,In_2762);
nand U515 (N_515,In_1553,In_1623);
nor U516 (N_516,In_2520,In_454);
nor U517 (N_517,In_4125,In_1045);
or U518 (N_518,In_854,In_3031);
nand U519 (N_519,In_3650,In_1969);
nand U520 (N_520,In_2173,In_3342);
or U521 (N_521,In_1844,In_99);
nor U522 (N_522,In_2501,In_1994);
nand U523 (N_523,In_3235,In_3722);
or U524 (N_524,In_2218,In_2472);
and U525 (N_525,In_1758,In_4356);
or U526 (N_526,In_2,In_526);
xnor U527 (N_527,In_3148,In_1917);
or U528 (N_528,In_2448,In_3809);
and U529 (N_529,In_4525,In_4579);
nand U530 (N_530,In_3787,In_4434);
and U531 (N_531,In_79,In_3825);
nor U532 (N_532,In_1267,In_3387);
nand U533 (N_533,In_3317,In_1662);
and U534 (N_534,In_2434,In_3980);
nand U535 (N_535,In_3910,In_2567);
nor U536 (N_536,In_1151,In_2319);
and U537 (N_537,In_4086,In_3996);
nor U538 (N_538,In_3350,In_3393);
xor U539 (N_539,In_4782,In_1693);
and U540 (N_540,In_185,In_816);
nor U541 (N_541,In_3706,In_3641);
xnor U542 (N_542,In_2745,In_2304);
or U543 (N_543,In_2827,In_4869);
nand U544 (N_544,In_2102,In_2483);
and U545 (N_545,In_1143,In_3414);
nand U546 (N_546,In_4650,In_1665);
nand U547 (N_547,In_2828,In_2830);
xnor U548 (N_548,In_1289,In_3161);
nor U549 (N_549,In_4667,In_2961);
or U550 (N_550,In_3410,In_3561);
or U551 (N_551,In_2788,In_4822);
nand U552 (N_552,In_1055,In_3497);
nand U553 (N_553,In_3484,In_2424);
or U554 (N_554,In_4982,In_477);
and U555 (N_555,In_504,In_1080);
and U556 (N_556,In_2465,In_2852);
nand U557 (N_557,In_3717,In_879);
or U558 (N_558,In_704,In_4531);
nand U559 (N_559,In_1531,In_3100);
nor U560 (N_560,In_3578,In_3212);
or U561 (N_561,In_2243,In_4165);
nor U562 (N_562,In_1000,In_4726);
nand U563 (N_563,In_1236,In_4015);
or U564 (N_564,In_4900,In_4059);
or U565 (N_565,In_3924,In_4540);
nand U566 (N_566,In_1588,In_2177);
xor U567 (N_567,In_3536,In_2765);
or U568 (N_568,In_4840,In_4991);
nor U569 (N_569,In_3582,In_3398);
or U570 (N_570,In_2769,In_4607);
nor U571 (N_571,In_940,In_3370);
and U572 (N_572,In_4645,In_3775);
or U573 (N_573,In_1656,In_3940);
nand U574 (N_574,In_1302,In_4777);
nand U575 (N_575,In_2451,In_3955);
nand U576 (N_576,In_630,In_3240);
nand U577 (N_577,In_3047,In_2584);
and U578 (N_578,In_1661,In_1741);
xnor U579 (N_579,In_4810,In_4546);
nor U580 (N_580,In_2659,In_4431);
nor U581 (N_581,In_3127,In_3806);
and U582 (N_582,In_455,In_2169);
nor U583 (N_583,In_1152,In_97);
nand U584 (N_584,In_2015,In_2114);
nand U585 (N_585,In_1250,In_4701);
and U586 (N_586,In_3849,In_2463);
nor U587 (N_587,In_4556,In_1372);
nand U588 (N_588,In_467,In_2016);
nor U589 (N_589,In_3670,In_554);
and U590 (N_590,In_3413,In_4017);
or U591 (N_591,In_1272,In_3200);
or U592 (N_592,In_2713,In_507);
nand U593 (N_593,In_463,In_3671);
xnor U594 (N_594,In_2429,In_3160);
nand U595 (N_595,In_2775,In_756);
or U596 (N_596,In_4704,In_512);
nor U597 (N_597,In_4105,In_3121);
or U598 (N_598,In_1775,In_1132);
nand U599 (N_599,In_4092,In_4102);
nand U600 (N_600,In_2938,In_4007);
nor U601 (N_601,In_1395,In_846);
and U602 (N_602,In_4303,In_1367);
and U603 (N_603,In_3227,In_2440);
or U604 (N_604,In_2931,In_380);
nand U605 (N_605,In_208,In_2229);
xnor U606 (N_606,In_3299,In_840);
or U607 (N_607,In_3270,In_1968);
or U608 (N_608,In_147,In_3236);
nor U609 (N_609,In_18,In_3944);
nor U610 (N_610,In_1782,In_782);
nor U611 (N_611,In_619,In_4025);
nand U612 (N_612,In_3050,In_2866);
nor U613 (N_613,In_3019,In_1606);
or U614 (N_614,In_386,In_2278);
or U615 (N_615,In_2241,In_3196);
nand U616 (N_616,In_3298,In_2997);
and U617 (N_617,In_3296,In_2245);
or U618 (N_618,In_949,In_445);
nand U619 (N_619,In_1379,In_1547);
and U620 (N_620,In_71,In_1043);
xor U621 (N_621,In_4881,In_639);
nand U622 (N_622,In_3637,In_918);
nand U623 (N_623,In_1384,In_1130);
nand U624 (N_624,In_1443,In_2700);
and U625 (N_625,In_4560,In_4669);
and U626 (N_626,In_3978,In_4171);
or U627 (N_627,In_4892,In_348);
and U628 (N_628,In_3555,In_2254);
nor U629 (N_629,In_2422,In_539);
or U630 (N_630,In_1859,In_1538);
nand U631 (N_631,In_2130,In_1447);
or U632 (N_632,In_4821,In_532);
and U633 (N_633,In_265,In_1126);
xor U634 (N_634,In_319,In_338);
and U635 (N_635,In_3385,In_3833);
nand U636 (N_636,In_3386,In_2511);
and U637 (N_637,In_262,In_374);
xnor U638 (N_638,In_3686,In_874);
nor U639 (N_639,In_2617,In_3213);
and U640 (N_640,In_2766,In_2075);
and U641 (N_641,In_850,In_766);
and U642 (N_642,In_4177,In_1075);
nand U643 (N_643,In_3962,In_4113);
nand U644 (N_644,In_1735,In_2139);
and U645 (N_645,In_3503,In_1040);
or U646 (N_646,In_3381,In_2660);
nand U647 (N_647,In_3113,In_4018);
or U648 (N_648,In_4606,In_2212);
xnor U649 (N_649,In_839,In_3960);
xnor U650 (N_650,In_195,In_4122);
and U651 (N_651,In_2601,In_2971);
nand U652 (N_652,In_2127,In_739);
nor U653 (N_653,In_1642,In_1652);
nor U654 (N_654,In_728,In_4786);
xor U655 (N_655,In_4156,In_3069);
nand U656 (N_656,In_4906,In_1407);
or U657 (N_657,In_967,In_3464);
nor U658 (N_658,In_3795,In_3917);
nand U659 (N_659,In_4068,In_1712);
xnor U660 (N_660,In_1314,In_4069);
and U661 (N_661,In_3542,In_3124);
or U662 (N_662,In_2600,In_4442);
xnor U663 (N_663,In_844,In_2689);
and U664 (N_664,In_1937,In_3950);
nor U665 (N_665,In_2366,In_3139);
or U666 (N_666,In_2269,In_2428);
and U667 (N_667,In_1748,In_2395);
and U668 (N_668,In_3842,In_2335);
nor U669 (N_669,In_2996,In_269);
nor U670 (N_670,In_1702,In_1402);
nor U671 (N_671,In_4423,In_1527);
nor U672 (N_672,In_1377,In_3373);
nor U673 (N_673,In_3029,In_2995);
or U674 (N_674,In_1753,In_4426);
nand U675 (N_675,In_529,In_4376);
nand U676 (N_676,In_2794,In_3364);
xor U677 (N_677,In_4087,In_929);
nor U678 (N_678,In_841,In_1768);
xor U679 (N_679,In_1952,In_4329);
nand U680 (N_680,In_2330,In_333);
nor U681 (N_681,In_2332,In_3838);
and U682 (N_682,In_135,In_3144);
or U683 (N_683,In_3333,In_4956);
or U684 (N_684,In_3030,In_1991);
nand U685 (N_685,In_4499,In_3760);
nor U686 (N_686,In_2802,In_2325);
or U687 (N_687,In_3309,In_1199);
or U688 (N_688,In_703,In_2006);
nor U689 (N_689,In_2446,In_4225);
and U690 (N_690,In_2555,In_1114);
or U691 (N_691,In_1926,In_3777);
xor U692 (N_692,In_2523,In_2624);
or U693 (N_693,In_3819,In_132);
nor U694 (N_694,In_3135,In_3409);
or U695 (N_695,In_457,In_49);
and U696 (N_696,In_1535,In_4155);
nor U697 (N_697,In_1902,In_3678);
or U698 (N_698,In_4884,In_2572);
and U699 (N_699,In_3494,In_4262);
and U700 (N_700,In_2720,In_3828);
or U701 (N_701,In_296,In_1655);
and U702 (N_702,In_3726,In_1692);
nand U703 (N_703,In_547,In_3267);
or U704 (N_704,In_4382,In_1638);
xnor U705 (N_705,In_1916,In_3230);
nor U706 (N_706,In_1871,In_2972);
or U707 (N_707,In_3457,In_2018);
nand U708 (N_708,In_1112,In_2204);
nor U709 (N_709,In_1474,In_1982);
nand U710 (N_710,In_1589,In_1823);
and U711 (N_711,In_4859,In_2499);
nor U712 (N_712,In_1048,In_2715);
and U713 (N_713,In_157,In_3067);
xor U714 (N_714,In_4486,In_300);
and U715 (N_715,In_2657,In_726);
and U716 (N_716,In_911,In_983);
or U717 (N_717,In_1776,In_1860);
nor U718 (N_718,In_3739,In_3090);
and U719 (N_719,In_4613,In_722);
or U720 (N_720,In_46,In_1475);
nor U721 (N_721,In_2051,In_1536);
or U722 (N_722,In_3793,In_645);
nor U723 (N_723,In_3811,In_3089);
or U724 (N_724,In_1188,In_2126);
and U725 (N_725,In_1512,In_500);
nand U726 (N_726,In_867,In_3274);
and U727 (N_727,In_3257,In_4452);
nand U728 (N_728,In_389,In_3705);
or U729 (N_729,In_3860,In_1101);
nand U730 (N_730,In_1783,In_4973);
or U731 (N_731,In_4206,In_3618);
and U732 (N_732,In_1847,In_1009);
nor U733 (N_733,In_2692,In_3184);
nor U734 (N_734,In_2609,In_438);
or U735 (N_735,In_4708,In_4190);
and U736 (N_736,In_674,In_1260);
nor U737 (N_737,In_481,In_4414);
nand U738 (N_738,In_1317,In_2411);
or U739 (N_739,In_3829,In_1658);
and U740 (N_740,In_1078,In_3884);
and U741 (N_741,In_4377,In_3493);
or U742 (N_742,In_4260,In_437);
nor U743 (N_743,In_1172,In_3758);
nor U744 (N_744,In_2661,In_3869);
and U745 (N_745,In_4336,In_2001);
nand U746 (N_746,In_2163,In_1678);
and U747 (N_747,In_3411,In_4217);
nor U748 (N_748,In_200,In_1805);
or U749 (N_749,In_118,In_1003);
or U750 (N_750,In_1814,In_2853);
xor U751 (N_751,In_2171,In_3824);
and U752 (N_752,In_4176,In_2145);
and U753 (N_753,In_2412,In_3700);
and U754 (N_754,In_2867,In_194);
nor U755 (N_755,In_3624,In_4723);
nor U756 (N_756,In_1633,In_2289);
nor U757 (N_757,In_4813,In_1908);
xnor U758 (N_758,In_3942,In_1397);
and U759 (N_759,In_423,In_4439);
nand U760 (N_760,In_1442,In_3308);
nor U761 (N_761,In_4767,In_281);
and U762 (N_762,In_140,In_3970);
and U763 (N_763,In_2393,In_3259);
or U764 (N_764,In_356,In_2012);
or U765 (N_765,In_2408,In_2882);
xor U766 (N_766,In_241,In_3420);
nor U767 (N_767,In_2547,In_1806);
and U768 (N_768,In_3649,In_4436);
xor U769 (N_769,In_3741,In_2899);
nor U770 (N_770,In_274,In_246);
or U771 (N_771,In_3778,In_143);
and U772 (N_772,In_525,In_2781);
and U773 (N_773,In_3465,In_402);
or U774 (N_774,In_4457,In_653);
nand U775 (N_775,In_3157,In_944);
or U776 (N_776,In_4437,In_4227);
xnor U777 (N_777,In_1102,In_450);
or U778 (N_778,In_116,In_3530);
and U779 (N_779,In_4624,In_518);
nor U780 (N_780,In_2283,In_2921);
and U781 (N_781,In_2918,In_1682);
or U782 (N_782,In_4861,In_1304);
nand U783 (N_783,In_1585,In_1248);
nand U784 (N_784,In_3591,In_186);
xor U785 (N_785,In_2216,In_163);
or U786 (N_786,In_69,In_1249);
nand U787 (N_787,In_1597,In_2076);
nor U788 (N_788,In_1686,In_1454);
or U789 (N_789,In_212,In_3395);
and U790 (N_790,In_54,In_2569);
or U791 (N_791,In_4605,In_1970);
or U792 (N_792,In_957,In_3024);
or U793 (N_793,In_1749,In_4210);
nand U794 (N_794,In_998,In_3753);
nor U795 (N_795,In_1711,In_3422);
xnor U796 (N_796,In_391,In_303);
nand U797 (N_797,In_4780,In_284);
nand U798 (N_798,In_2374,In_670);
and U799 (N_799,In_907,In_4682);
and U800 (N_800,In_434,In_3286);
and U801 (N_801,In_917,In_1943);
nand U802 (N_802,In_537,In_2222);
or U803 (N_803,In_780,In_4094);
nor U804 (N_804,In_565,In_1070);
nor U805 (N_805,In_4552,In_2710);
and U806 (N_806,In_4067,In_4744);
or U807 (N_807,In_2280,In_173);
nor U808 (N_808,In_3781,In_211);
and U809 (N_809,In_3483,In_413);
or U810 (N_810,In_3695,In_1169);
nor U811 (N_811,In_2651,In_4351);
and U812 (N_812,In_2401,In_4985);
nor U813 (N_813,In_2369,In_3046);
or U814 (N_814,In_2495,In_1584);
and U815 (N_815,In_1494,In_3539);
or U816 (N_816,In_3054,In_3313);
or U817 (N_817,In_4646,In_32);
nor U818 (N_818,In_3416,In_1273);
or U819 (N_819,In_3856,In_1895);
and U820 (N_820,In_1222,In_1928);
nand U821 (N_821,In_866,In_3415);
xnor U822 (N_822,In_1202,In_2679);
nand U823 (N_823,In_2870,In_1343);
nor U824 (N_824,In_605,In_593);
or U825 (N_825,In_1028,In_1876);
and U826 (N_826,In_4519,In_4312);
nor U827 (N_827,In_4141,In_1889);
xnor U828 (N_828,In_3084,In_4074);
nand U829 (N_829,In_3952,In_4922);
and U830 (N_830,In_1953,In_3179);
and U831 (N_831,In_527,In_113);
or U832 (N_832,In_2353,In_3225);
and U833 (N_833,In_420,In_1499);
or U834 (N_834,In_1627,In_510);
xor U835 (N_835,In_4703,In_4209);
and U836 (N_836,In_440,In_4243);
and U837 (N_837,In_2804,In_3731);
and U838 (N_838,In_2597,In_1166);
or U839 (N_839,In_4897,In_1548);
nor U840 (N_840,In_4931,In_598);
nand U841 (N_841,In_315,In_4385);
nor U842 (N_842,In_4912,In_4066);
and U843 (N_843,In_2947,In_1554);
or U844 (N_844,In_1122,In_2263);
or U845 (N_845,In_4589,In_2193);
xor U846 (N_846,In_2209,In_11);
xor U847 (N_847,In_4594,In_922);
nand U848 (N_848,In_2693,In_1500);
nand U849 (N_849,In_3482,In_1607);
xor U850 (N_850,In_1744,In_327);
and U851 (N_851,In_2991,In_2707);
nand U852 (N_852,In_4578,In_4644);
nand U853 (N_853,In_235,In_2197);
nand U854 (N_854,In_2676,In_4969);
and U855 (N_855,In_3783,In_1127);
nor U856 (N_856,In_2699,In_476);
and U857 (N_857,In_2886,In_4335);
nor U858 (N_858,In_2596,In_1939);
nor U859 (N_859,In_160,In_2025);
nor U860 (N_860,In_2642,In_2687);
nand U861 (N_861,In_4245,In_155);
nor U862 (N_862,In_2616,In_2485);
and U863 (N_863,In_1145,In_2626);
xor U864 (N_864,In_2071,In_4175);
or U865 (N_865,In_1308,In_552);
or U866 (N_866,In_1065,In_4845);
nor U867 (N_867,In_1649,In_4707);
and U868 (N_868,In_4592,In_3272);
nor U869 (N_869,In_903,In_4617);
or U870 (N_870,In_1339,In_2066);
nand U871 (N_871,In_2549,In_4634);
nor U872 (N_872,In_1072,In_2235);
nor U873 (N_873,In_342,In_4689);
and U874 (N_874,In_2077,In_2432);
and U875 (N_875,In_4908,In_3169);
or U876 (N_876,In_495,In_4116);
or U877 (N_877,In_5,In_4085);
or U878 (N_878,In_4712,In_4927);
nor U879 (N_879,In_2464,In_2686);
nor U880 (N_880,In_499,In_3432);
or U881 (N_881,In_1648,In_3220);
and U882 (N_882,In_3015,In_541);
nor U883 (N_883,In_3657,In_3106);
and U884 (N_884,In_171,In_2013);
nand U885 (N_885,In_228,In_4287);
nor U886 (N_886,In_1162,In_4450);
nor U887 (N_887,In_2106,In_394);
nor U888 (N_888,In_2228,In_4949);
and U889 (N_889,In_3376,In_4300);
or U890 (N_890,In_609,In_2958);
or U891 (N_891,In_4193,In_4330);
nand U892 (N_892,In_3613,In_2952);
and U893 (N_893,In_4473,In_4522);
and U894 (N_894,In_1546,In_1828);
nor U895 (N_895,In_1571,In_2217);
and U896 (N_896,In_3125,In_625);
or U897 (N_897,In_1012,In_1079);
or U898 (N_898,In_1408,In_1205);
or U899 (N_899,In_3846,In_683);
xor U900 (N_900,In_496,In_2650);
nand U901 (N_901,In_4326,In_830);
nand U902 (N_902,In_2298,In_1773);
or U903 (N_903,In_1330,In_3786);
nor U904 (N_904,In_3083,In_3701);
nor U905 (N_905,In_960,In_4946);
and U906 (N_906,In_2020,In_954);
nor U907 (N_907,In_221,In_456);
or U908 (N_908,In_3016,In_3026);
and U909 (N_909,In_4379,In_2825);
nor U910 (N_910,In_1089,In_2884);
xor U911 (N_911,In_1825,In_4599);
xnor U912 (N_912,In_1301,In_3805);
nand U913 (N_913,In_4978,In_1719);
nor U914 (N_914,In_932,In_2939);
nand U915 (N_915,In_3065,In_4725);
nor U916 (N_916,In_2462,In_2279);
and U917 (N_917,In_4413,In_3612);
or U918 (N_918,In_1163,In_4673);
nor U919 (N_919,In_1470,In_4107);
xnor U920 (N_920,In_959,In_26);
nand U921 (N_921,In_2294,In_1963);
nor U922 (N_922,In_2606,In_1246);
or U923 (N_923,In_1125,In_1209);
and U924 (N_924,In_4575,In_1432);
or U925 (N_925,In_1359,In_3490);
nor U926 (N_926,In_3147,In_4183);
xnor U927 (N_927,In_2180,In_2437);
and U928 (N_928,In_4992,In_1838);
nor U929 (N_929,In_2811,In_2255);
nor U930 (N_930,In_1307,In_4964);
nand U931 (N_931,In_3346,In_4191);
xor U932 (N_932,In_858,In_3908);
nand U933 (N_933,In_1998,In_4958);
or U934 (N_934,In_4515,In_536);
and U935 (N_935,In_4148,In_447);
nor U936 (N_936,In_4104,In_4541);
xnor U937 (N_937,In_4047,In_2809);
or U938 (N_938,In_3362,In_1909);
nor U939 (N_939,In_1230,In_3837);
nor U940 (N_940,In_2571,In_1288);
nand U941 (N_941,In_3981,In_715);
nor U942 (N_942,In_1972,In_2214);
and U943 (N_943,In_2249,In_1355);
nand U944 (N_944,In_75,In_3306);
or U945 (N_945,In_4670,In_2062);
or U946 (N_946,In_2543,In_4751);
nand U947 (N_947,In_3560,In_3589);
nand U948 (N_948,In_2049,In_875);
nor U949 (N_949,In_3154,In_836);
nand U950 (N_950,In_3911,In_3568);
nor U951 (N_951,In_470,In_521);
or U952 (N_952,In_3123,In_1235);
or U953 (N_953,In_1946,In_4031);
nand U954 (N_954,In_2387,In_1629);
and U955 (N_955,In_2935,In_92);
nand U956 (N_956,In_1769,In_3344);
and U957 (N_957,In_1439,In_4609);
or U958 (N_958,In_772,In_1892);
and U959 (N_959,In_3207,In_3581);
xnor U960 (N_960,In_3077,In_933);
nor U961 (N_961,In_4309,In_3470);
nand U962 (N_962,In_1340,In_1224);
nand U963 (N_963,In_1107,In_909);
and U964 (N_964,In_635,In_1258);
nor U965 (N_965,In_1328,In_4355);
nor U966 (N_966,In_2183,In_2837);
or U967 (N_967,In_4772,In_1799);
and U968 (N_968,In_3690,In_2111);
xnor U969 (N_969,In_1390,In_240);
and U970 (N_970,In_4825,In_3694);
and U971 (N_971,In_4923,In_2359);
or U972 (N_972,In_3290,In_3532);
nor U973 (N_973,In_1049,In_2599);
nor U974 (N_974,In_3656,In_3733);
xnor U975 (N_975,In_3033,In_1691);
nor U976 (N_976,In_3677,In_2776);
and U977 (N_977,In_3525,In_2431);
nand U978 (N_978,In_2742,In_1411);
nand U979 (N_979,In_734,In_1206);
nand U980 (N_980,In_3153,In_3850);
and U981 (N_981,In_2469,In_3223);
nand U982 (N_982,In_1609,In_1720);
xnor U983 (N_983,In_2055,In_2850);
and U984 (N_984,In_4660,In_2863);
and U985 (N_985,In_4841,In_610);
nor U986 (N_986,In_3265,In_1839);
nor U987 (N_987,In_951,In_449);
xor U988 (N_988,In_3628,In_4878);
nand U989 (N_989,In_4749,In_3210);
nor U990 (N_990,In_3583,In_4021);
xor U991 (N_991,In_2902,In_1936);
nor U992 (N_992,In_3732,In_136);
and U993 (N_993,In_873,In_1306);
and U994 (N_994,In_2343,In_1880);
xnor U995 (N_995,In_1539,In_1840);
nor U996 (N_996,In_595,In_4648);
nand U997 (N_997,In_4614,In_4727);
and U998 (N_998,In_4898,In_914);
nand U999 (N_999,In_494,In_1754);
nor U1000 (N_1000,In_1514,In_2439);
nor U1001 (N_1001,In_2512,In_3969);
and U1002 (N_1002,In_4630,In_206);
nand U1003 (N_1003,In_1255,In_2061);
nand U1004 (N_1004,In_1321,In_2128);
xor U1005 (N_1005,In_4774,In_2080);
nand U1006 (N_1006,In_134,In_4204);
nor U1007 (N_1007,In_2338,In_1266);
or U1008 (N_1008,In_634,In_3110);
and U1009 (N_1009,In_3906,In_1389);
and U1010 (N_1010,In_1203,In_2167);
nand U1011 (N_1011,In_108,In_513);
or U1012 (N_1012,In_997,In_1265);
and U1013 (N_1013,In_2647,In_3496);
nand U1014 (N_1014,In_2323,In_3742);
or U1015 (N_1015,In_752,In_2487);
and U1016 (N_1016,In_832,In_1030);
or U1017 (N_1017,In_2454,In_4729);
or U1018 (N_1018,In_2505,In_364);
or U1019 (N_1019,In_4952,In_419);
nor U1020 (N_1020,In_3201,In_779);
nand U1021 (N_1021,In_4773,In_3451);
nand U1022 (N_1022,In_4460,In_1592);
nand U1023 (N_1023,In_3405,In_992);
and U1024 (N_1024,In_2847,In_700);
nor U1025 (N_1025,In_41,In_1319);
and U1026 (N_1026,In_4971,In_1393);
and U1027 (N_1027,In_2840,In_4622);
nor U1028 (N_1028,In_2317,In_3546);
nor U1029 (N_1029,In_2578,In_4829);
and U1030 (N_1030,In_3433,In_3205);
or U1031 (N_1031,In_973,In_2832);
or U1032 (N_1032,In_2638,In_1257);
and U1033 (N_1033,In_4806,In_1392);
or U1034 (N_1034,In_2914,In_4271);
and U1035 (N_1035,In_1759,In_3337);
nand U1036 (N_1036,In_4358,In_3661);
and U1037 (N_1037,In_3575,In_2920);
and U1038 (N_1038,In_2162,In_1660);
or U1039 (N_1039,In_1815,In_3307);
nand U1040 (N_1040,In_3185,In_414);
and U1041 (N_1041,In_153,In_1601);
or U1042 (N_1042,In_1779,In_2089);
nor U1043 (N_1043,In_239,In_3672);
nor U1044 (N_1044,In_1256,In_4615);
and U1045 (N_1045,In_2336,In_1426);
nor U1046 (N_1046,In_1919,In_2058);
nand U1047 (N_1047,In_1458,In_2592);
nor U1048 (N_1048,In_3759,In_3971);
and U1049 (N_1049,In_4152,In_3684);
nor U1050 (N_1050,In_895,In_107);
and U1051 (N_1051,In_3463,In_3291);
or U1052 (N_1052,In_2761,In_1282);
xnor U1053 (N_1053,In_4797,In_3926);
and U1054 (N_1054,In_1772,In_3804);
xnor U1055 (N_1055,In_2570,In_4651);
or U1056 (N_1056,In_2565,In_3852);
and U1057 (N_1057,In_3042,In_2544);
or U1058 (N_1058,In_3947,In_692);
nand U1059 (N_1059,In_1325,In_4192);
nand U1060 (N_1060,In_4536,In_1191);
and U1061 (N_1061,In_3596,In_223);
nor U1062 (N_1062,In_2903,In_2550);
nor U1063 (N_1063,In_4099,In_757);
and U1064 (N_1064,In_3222,In_378);
and U1065 (N_1065,In_4724,In_4064);
nand U1066 (N_1066,In_3094,In_3492);
nor U1067 (N_1067,In_2390,In_1298);
nor U1068 (N_1068,In_2985,In_1478);
and U1069 (N_1069,In_4343,In_3211);
or U1070 (N_1070,In_612,In_4757);
nand U1071 (N_1071,In_1196,In_52);
and U1072 (N_1072,In_3312,In_3057);
nand U1073 (N_1073,In_2054,In_1324);
nor U1074 (N_1074,In_896,In_4403);
nand U1075 (N_1075,In_465,In_2556);
nand U1076 (N_1076,In_3680,In_2149);
nand U1077 (N_1077,In_3688,In_3076);
nand U1078 (N_1078,In_2119,In_1798);
nor U1079 (N_1079,In_3961,In_767);
nor U1080 (N_1080,In_2577,In_2259);
and U1081 (N_1081,In_626,In_2702);
and U1082 (N_1082,In_1486,In_2404);
xnor U1083 (N_1083,In_2364,In_4491);
nor U1084 (N_1084,In_1421,In_3504);
or U1085 (N_1085,In_2881,In_1156);
and U1086 (N_1086,In_3558,In_3543);
and U1087 (N_1087,In_2152,In_0);
nor U1088 (N_1088,In_4940,In_3442);
nand U1089 (N_1089,In_2486,In_2371);
or U1090 (N_1090,In_4683,In_788);
nor U1091 (N_1091,In_3318,In_1207);
nor U1092 (N_1092,In_4100,In_1226);
xnor U1093 (N_1093,In_4215,In_1868);
xor U1094 (N_1094,In_4685,In_963);
nor U1095 (N_1095,In_279,In_3407);
nand U1096 (N_1096,In_769,In_4702);
nand U1097 (N_1097,In_4400,In_4827);
and U1098 (N_1098,In_2801,In_3757);
or U1099 (N_1099,In_3702,In_3571);
or U1100 (N_1100,In_1452,In_1093);
nor U1101 (N_1101,In_4072,In_4306);
and U1102 (N_1102,In_1420,In_3513);
and U1103 (N_1103,In_3336,In_2916);
nor U1104 (N_1104,In_251,In_2945);
nand U1105 (N_1105,In_4097,In_1978);
nor U1106 (N_1106,In_344,In_1900);
or U1107 (N_1107,In_3061,In_4078);
nor U1108 (N_1108,In_3020,In_3872);
nand U1109 (N_1109,In_617,In_2735);
nand U1110 (N_1110,In_2021,In_3654);
nor U1111 (N_1111,In_3461,In_2705);
or U1112 (N_1112,In_2311,In_253);
or U1113 (N_1113,In_2213,In_1777);
and U1114 (N_1114,In_2185,In_1182);
nand U1115 (N_1115,In_3032,In_3170);
nor U1116 (N_1116,In_3181,In_3390);
and U1117 (N_1117,In_1097,In_2402);
and U1118 (N_1118,In_1757,In_1593);
xnor U1119 (N_1119,In_4788,In_968);
nand U1120 (N_1120,In_1944,In_1341);
and U1121 (N_1121,In_3218,In_125);
or U1122 (N_1122,In_4577,In_1005);
and U1123 (N_1123,In_4548,In_4103);
nor U1124 (N_1124,In_2175,In_2664);
xnor U1125 (N_1125,In_2566,In_2981);
and U1126 (N_1126,In_3284,In_131);
nand U1127 (N_1127,In_2329,In_4526);
nand U1128 (N_1128,In_2785,In_615);
or U1129 (N_1129,In_12,In_1526);
and U1130 (N_1130,In_2654,In_68);
nor U1131 (N_1131,In_1204,In_318);
xnor U1132 (N_1132,In_1358,In_1523);
xor U1133 (N_1133,In_556,In_2508);
and U1134 (N_1134,In_705,In_432);
xor U1135 (N_1135,In_1487,In_2764);
and U1136 (N_1136,In_4873,In_2155);
or U1137 (N_1137,In_4801,In_4928);
nor U1138 (N_1138,In_2109,In_1704);
or U1139 (N_1139,In_4061,In_1818);
nand U1140 (N_1140,In_1685,In_3087);
nor U1141 (N_1141,In_254,In_193);
nor U1142 (N_1142,In_4282,In_2872);
nand U1143 (N_1143,In_1583,In_935);
nor U1144 (N_1144,In_3345,In_188);
nor U1145 (N_1145,In_3770,In_2007);
or U1146 (N_1146,In_2378,In_98);
or U1147 (N_1147,In_1988,In_4939);
or U1148 (N_1148,In_1619,In_2860);
or U1149 (N_1149,In_842,In_1185);
nor U1150 (N_1150,In_4933,In_4479);
xor U1151 (N_1151,In_3619,In_1563);
nor U1152 (N_1152,In_4274,In_3507);
and U1153 (N_1153,In_2755,In_3992);
or U1154 (N_1154,In_197,In_1817);
nand U1155 (N_1155,In_2527,In_1444);
xnor U1156 (N_1156,In_2949,In_553);
xor U1157 (N_1157,In_863,In_620);
and U1158 (N_1158,In_2100,In_986);
or U1159 (N_1159,In_3554,In_650);
or U1160 (N_1160,In_1017,In_1747);
nor U1161 (N_1161,In_1491,In_1335);
and U1162 (N_1162,In_82,In_853);
and U1163 (N_1163,In_328,In_4692);
and U1164 (N_1164,In_4081,In_2628);
or U1165 (N_1165,In_88,In_3340);
or U1166 (N_1166,In_2967,In_63);
and U1167 (N_1167,In_2492,In_4359);
nor U1168 (N_1168,In_4924,In_2953);
nand U1169 (N_1169,In_1933,In_4214);
and U1170 (N_1170,In_4987,In_1320);
or U1171 (N_1171,In_1422,In_2824);
and U1172 (N_1172,In_1118,In_2274);
nand U1173 (N_1173,In_4241,In_4697);
nor U1174 (N_1174,In_515,In_4647);
nor U1175 (N_1175,In_1616,In_354);
and U1176 (N_1176,In_3010,In_825);
nor U1177 (N_1177,In_809,In_2036);
or U1178 (N_1178,In_596,In_4415);
nor U1179 (N_1179,In_310,In_3974);
nor U1180 (N_1180,In_443,In_154);
or U1181 (N_1181,In_392,In_3097);
and U1182 (N_1182,In_3434,In_3615);
xnor U1183 (N_1183,In_1216,In_1819);
and U1184 (N_1184,In_2641,In_3954);
xnor U1185 (N_1185,In_4762,In_3052);
xor U1186 (N_1186,In_104,In_14);
and U1187 (N_1187,In_2682,In_435);
or U1188 (N_1188,In_2552,In_4399);
nand U1189 (N_1189,In_3929,In_2894);
nor U1190 (N_1190,In_586,In_1740);
nand U1191 (N_1191,In_219,In_4826);
nor U1192 (N_1192,In_1517,In_2190);
nor U1193 (N_1193,In_3685,In_3659);
nand U1194 (N_1194,In_3023,In_557);
xnor U1195 (N_1195,In_691,In_3314);
or U1196 (N_1196,In_1220,In_2195);
nor U1197 (N_1197,In_1021,In_3506);
nor U1198 (N_1198,In_1391,In_1864);
or U1199 (N_1199,In_2820,In_232);
nor U1200 (N_1200,In_1590,In_912);
nor U1201 (N_1201,In_2843,In_3905);
nand U1202 (N_1202,In_1561,In_1725);
nor U1203 (N_1203,In_4760,In_1714);
nor U1204 (N_1204,In_1263,In_4487);
or U1205 (N_1205,In_317,In_3454);
xnor U1206 (N_1206,In_2919,In_3630);
nor U1207 (N_1207,In_247,In_2086);
nor U1208 (N_1208,In_3343,In_4766);
xnor U1209 (N_1209,In_1999,In_3844);
nor U1210 (N_1210,In_4868,In_1669);
and U1211 (N_1211,In_4654,In_4573);
nand U1212 (N_1212,In_2888,In_4625);
and U1213 (N_1213,In_3068,In_1111);
xnor U1214 (N_1214,In_1337,In_3576);
and U1215 (N_1215,In_3922,In_1541);
nor U1216 (N_1216,In_2573,In_4555);
and U1217 (N_1217,In_2291,In_365);
nand U1218 (N_1218,In_2539,In_199);
and U1219 (N_1219,In_3260,In_2103);
xor U1220 (N_1220,In_1387,In_371);
nand U1221 (N_1221,In_633,In_2545);
and U1222 (N_1222,In_222,In_1940);
or U1223 (N_1223,In_4172,In_3338);
nand U1224 (N_1224,In_4848,In_3880);
nor U1225 (N_1225,In_1984,In_3189);
xor U1226 (N_1226,In_24,In_2315);
and U1227 (N_1227,In_3632,In_4737);
and U1228 (N_1228,In_181,In_3448);
nand U1229 (N_1229,In_775,In_3086);
nand U1230 (N_1230,In_3719,In_2653);
or U1231 (N_1231,In_2885,In_2085);
nor U1232 (N_1232,In_2159,In_644);
and U1233 (N_1233,In_2147,In_3278);
or U1234 (N_1234,In_4709,In_3939);
nor U1235 (N_1235,In_1628,In_4989);
nand U1236 (N_1236,In_3875,In_3914);
xor U1237 (N_1237,In_70,In_2064);
nor U1238 (N_1238,In_651,In_2714);
or U1239 (N_1239,In_802,In_3598);
nor U1240 (N_1240,In_359,In_4626);
and U1241 (N_1241,In_2515,In_822);
nand U1242 (N_1242,In_4591,In_574);
nor U1243 (N_1243,In_3079,In_3876);
nand U1244 (N_1244,In_1567,In_4658);
or U1245 (N_1245,In_1555,In_4836);
nand U1246 (N_1246,In_4823,In_1800);
nand U1247 (N_1247,In_3812,In_1574);
and U1248 (N_1248,In_159,In_297);
nand U1249 (N_1249,In_939,In_4619);
xnor U1250 (N_1250,In_2328,In_283);
nand U1251 (N_1251,In_4280,In_1903);
or U1252 (N_1252,In_4258,In_1467);
and U1253 (N_1253,In_1401,In_2019);
nor U1254 (N_1254,In_4769,In_666);
nand U1255 (N_1255,In_2504,In_2287);
nor U1256 (N_1256,In_987,In_761);
or U1257 (N_1257,In_2400,In_730);
nand U1258 (N_1258,In_4261,In_814);
xnor U1259 (N_1259,In_628,In_2398);
nand U1260 (N_1260,In_2153,In_673);
nand U1261 (N_1261,In_4851,In_372);
nor U1262 (N_1262,In_4249,In_3845);
and U1263 (N_1263,In_4256,In_4481);
xor U1264 (N_1264,In_1528,In_2014);
nand U1265 (N_1265,In_1178,In_4133);
nor U1266 (N_1266,In_1098,In_1064);
or U1267 (N_1267,In_1269,In_2376);
or U1268 (N_1268,In_1790,In_2132);
nor U1269 (N_1269,In_4179,In_2932);
nand U1270 (N_1270,In_1084,In_2484);
xnor U1271 (N_1271,In_4942,In_1821);
and U1272 (N_1272,In_1066,In_1835);
nor U1273 (N_1273,In_3790,In_4194);
and U1274 (N_1274,In_1680,In_4489);
or U1275 (N_1275,In_1460,In_4994);
or U1276 (N_1276,In_2002,In_4681);
nor U1277 (N_1277,In_2070,In_710);
or U1278 (N_1278,In_3266,In_4259);
nand U1279 (N_1279,In_1878,In_196);
or U1280 (N_1280,In_961,In_2576);
nor U1281 (N_1281,In_938,In_885);
nand U1282 (N_1282,In_2818,In_2352);
and U1283 (N_1283,In_4005,In_1025);
or U1284 (N_1284,In_488,In_3400);
nor U1285 (N_1285,In_638,In_4043);
nand U1286 (N_1286,In_4279,In_4019);
nand U1287 (N_1287,In_3486,In_4132);
nand U1288 (N_1288,In_3899,In_3557);
or U1289 (N_1289,In_976,In_2052);
or U1290 (N_1290,In_724,In_4899);
nor U1291 (N_1291,In_1060,In_1857);
nor U1292 (N_1292,In_1058,In_2059);
xor U1293 (N_1293,In_2964,In_175);
nor U1294 (N_1294,In_590,In_475);
nand U1295 (N_1295,In_1431,In_4357);
and U1296 (N_1296,In_646,In_4334);
and U1297 (N_1297,In_4346,In_3602);
and U1298 (N_1298,In_2874,In_2345);
or U1299 (N_1299,In_1508,In_233);
or U1300 (N_1300,In_4696,In_880);
or U1301 (N_1301,In_1170,In_2415);
or U1302 (N_1302,In_4252,In_3621);
nor U1303 (N_1303,In_3142,In_329);
and U1304 (N_1304,In_3136,In_2768);
nand U1305 (N_1305,In_1219,In_4554);
or U1306 (N_1306,In_2494,In_1816);
or U1307 (N_1307,In_3734,In_3968);
xor U1308 (N_1308,In_3945,In_3941);
nor U1309 (N_1309,In_4278,In_4372);
nor U1310 (N_1310,In_2470,In_4211);
or U1311 (N_1311,In_1322,In_1399);
and U1312 (N_1312,In_3862,In_2816);
nor U1313 (N_1313,In_3112,In_1041);
nand U1314 (N_1314,In_4435,In_4528);
nor U1315 (N_1315,In_2823,In_4865);
nor U1316 (N_1316,In_1456,In_2479);
nor U1317 (N_1317,In_1292,In_4720);
and U1318 (N_1318,In_4794,In_350);
xnor U1319 (N_1319,In_2176,In_546);
and U1320 (N_1320,In_4979,In_3885);
and U1321 (N_1321,In_3320,In_2083);
nand U1322 (N_1322,In_4077,In_2518);
and U1323 (N_1323,In_1862,In_2948);
nor U1324 (N_1324,In_34,In_1897);
nor U1325 (N_1325,In_1434,In_2452);
nand U1326 (N_1326,In_2891,In_4568);
and U1327 (N_1327,In_1874,In_2900);
and U1328 (N_1328,In_161,In_4604);
and U1329 (N_1329,In_2976,In_4963);
and U1330 (N_1330,In_4444,In_4205);
and U1331 (N_1331,In_804,In_3101);
nor U1332 (N_1332,In_4396,In_3391);
and U1333 (N_1333,In_4397,In_482);
and U1334 (N_1334,In_3419,In_806);
or U1335 (N_1335,In_178,In_1734);
nor U1336 (N_1336,In_2262,In_3477);
nor U1337 (N_1337,In_3606,In_4603);
and U1338 (N_1338,In_3237,In_2368);
xnor U1339 (N_1339,In_1398,In_1890);
nand U1340 (N_1340,In_4633,In_4549);
nor U1341 (N_1341,In_294,In_1270);
nor U1342 (N_1342,In_1904,In_2219);
nand U1343 (N_1343,In_3823,In_16);
or U1344 (N_1344,In_985,In_1727);
nand U1345 (N_1345,In_882,In_3566);
or U1346 (N_1346,In_2361,In_881);
nand U1347 (N_1347,In_3109,In_3963);
nand U1348 (N_1348,In_4970,In_2956);
or U1349 (N_1349,In_1001,In_580);
or U1350 (N_1350,In_1208,In_4879);
nand U1351 (N_1351,In_3360,In_4185);
xnor U1352 (N_1352,In_2581,In_277);
nand U1353 (N_1353,In_2724,In_64);
or U1354 (N_1354,In_1886,In_334);
and U1355 (N_1355,In_4296,In_1154);
nor U1356 (N_1356,In_1218,In_800);
nand U1357 (N_1357,In_411,In_215);
or U1358 (N_1358,In_1894,In_4468);
nand U1359 (N_1359,In_555,In_349);
or U1360 (N_1360,In_2652,In_4993);
and U1361 (N_1361,In_1507,In_3369);
and U1362 (N_1362,In_61,In_2034);
nor U1363 (N_1363,In_3967,In_2324);
nor U1364 (N_1364,In_1688,In_1276);
nor U1365 (N_1365,In_3034,In_600);
or U1366 (N_1366,In_2632,In_2851);
nand U1367 (N_1367,In_4715,In_3912);
and U1368 (N_1368,In_1681,In_2582);
or U1369 (N_1369,In_3163,In_3204);
or U1370 (N_1370,In_852,In_2468);
and U1371 (N_1371,In_425,In_4831);
or U1372 (N_1372,In_2251,In_701);
or U1373 (N_1373,In_4657,In_3011);
nor U1374 (N_1374,In_1673,In_3130);
xnor U1375 (N_1375,In_460,In_2443);
or U1376 (N_1376,In_1313,In_1366);
or U1377 (N_1377,In_3303,In_1347);
or U1378 (N_1378,In_671,In_2528);
and U1379 (N_1379,In_60,In_3012);
and U1380 (N_1380,In_321,In_1394);
nand U1381 (N_1381,In_3839,In_4586);
xnor U1382 (N_1382,In_930,In_1957);
or U1383 (N_1383,In_1280,In_1104);
nor U1384 (N_1384,In_1587,In_2342);
or U1385 (N_1385,In_4616,In_4288);
nor U1386 (N_1386,In_3847,In_698);
or U1387 (N_1387,In_4270,In_390);
and U1388 (N_1388,In_4311,In_4044);
and U1389 (N_1389,In_4471,In_2640);
nand U1390 (N_1390,In_3818,In_1142);
or U1391 (N_1391,In_2441,In_4167);
nand U1392 (N_1392,In_1436,In_1275);
or U1393 (N_1393,In_1611,In_2760);
nand U1394 (N_1394,In_765,In_2753);
and U1395 (N_1395,In_3003,In_1189);
or U1396 (N_1396,In_3221,In_763);
nor U1397 (N_1397,In_3605,In_3725);
or U1398 (N_1398,In_3476,In_4174);
nand U1399 (N_1399,In_1764,In_4344);
nand U1400 (N_1400,In_2438,In_1932);
nor U1401 (N_1401,In_4298,In_784);
nand U1402 (N_1402,In_4201,In_2181);
and U1403 (N_1403,In_2189,In_2188);
nor U1404 (N_1404,In_4291,In_927);
nor U1405 (N_1405,In_928,In_3241);
xnor U1406 (N_1406,In_3749,In_1700);
nor U1407 (N_1407,In_576,In_255);
or U1408 (N_1408,In_3206,In_652);
xnor U1409 (N_1409,In_1465,In_2168);
nor U1410 (N_1410,In_1659,In_2719);
or U1411 (N_1411,In_1213,In_597);
nand U1412 (N_1412,In_4383,In_2911);
and U1413 (N_1413,In_1760,In_4947);
and U1414 (N_1414,In_3505,In_1380);
nand U1415 (N_1415,In_1026,In_4532);
and U1416 (N_1416,In_3036,In_4543);
xnor U1417 (N_1417,In_4887,In_4684);
nand U1418 (N_1418,In_4905,In_4506);
nor U1419 (N_1419,In_3987,In_3599);
nand U1420 (N_1420,In_3363,In_1477);
nand U1421 (N_1421,In_1115,In_4004);
and U1422 (N_1422,In_3301,In_1351);
nor U1423 (N_1423,In_4700,In_58);
nor U1424 (N_1424,In_4483,In_3044);
and U1425 (N_1425,In_2227,In_2634);
nor U1426 (N_1426,In_4792,In_1232);
or U1427 (N_1427,In_2138,In_330);
and U1428 (N_1428,In_3639,In_1197);
and U1429 (N_1429,In_925,In_4424);
nand U1430 (N_1430,In_1608,In_697);
nand U1431 (N_1431,In_2033,In_3440);
nor U1432 (N_1432,In_993,In_1231);
or U1433 (N_1433,In_1599,In_2131);
nor U1434 (N_1434,In_3975,In_3397);
and U1435 (N_1435,In_815,In_1286);
and U1436 (N_1436,In_1331,In_2154);
xnor U1437 (N_1437,In_3801,In_3936);
or U1438 (N_1438,In_4283,In_478);
and U1439 (N_1439,In_4717,In_570);
nor U1440 (N_1440,In_51,In_33);
or U1441 (N_1441,In_3763,In_2095);
nor U1442 (N_1442,In_3691,In_3339);
or U1443 (N_1443,In_3965,In_702);
and U1444 (N_1444,In_1473,In_1803);
or U1445 (N_1445,In_217,In_3984);
nand U1446 (N_1446,In_129,In_2455);
nand U1447 (N_1447,In_1161,In_2115);
or U1448 (N_1448,In_4269,In_3066);
or U1449 (N_1449,In_2770,In_3863);
or U1450 (N_1450,In_2221,In_1241);
nor U1451 (N_1451,In_2211,In_3467);
nand U1452 (N_1452,In_551,In_1713);
and U1453 (N_1453,In_4034,In_4517);
nor U1454 (N_1454,In_1949,In_1634);
and U1455 (N_1455,In_2595,In_1615);
nor U1456 (N_1456,In_2306,In_3150);
and U1457 (N_1457,In_1403,In_3752);
nor U1458 (N_1458,In_1971,In_2148);
nor U1459 (N_1459,In_1124,In_4371);
and U1460 (N_1460,In_1492,In_4266);
or U1461 (N_1461,In_528,In_2199);
or U1462 (N_1462,In_4921,In_3214);
and U1463 (N_1463,In_2146,In_4014);
or U1464 (N_1464,In_4054,In_483);
and U1465 (N_1465,In_2384,In_3538);
or U1466 (N_1466,In_4547,In_1023);
xor U1467 (N_1467,In_1505,In_1385);
xnor U1468 (N_1468,In_915,In_258);
nand U1469 (N_1469,In_1896,In_723);
nor U1470 (N_1470,In_4929,In_3349);
xor U1471 (N_1471,In_4166,In_1378);
or U1472 (N_1472,In_2750,In_4694);
and U1473 (N_1473,In_4710,In_80);
or U1474 (N_1474,In_3972,In_3474);
xnor U1475 (N_1475,In_1731,In_3174);
nand U1476 (N_1476,In_111,In_1653);
or U1477 (N_1477,In_4406,In_2773);
and U1478 (N_1478,In_2172,In_1323);
nand U1479 (N_1479,In_4353,In_1525);
and U1480 (N_1480,In_2067,In_2270);
nand U1481 (N_1481,In_1522,In_1362);
xor U1482 (N_1482,In_1356,In_2129);
nor U1483 (N_1483,In_83,In_29);
and U1484 (N_1484,In_1873,In_1144);
or U1485 (N_1485,In_2955,In_2901);
nor U1486 (N_1486,In_4690,In_1223);
nor U1487 (N_1487,In_3053,In_4671);
or U1488 (N_1488,In_3446,In_4467);
or U1489 (N_1489,In_2476,In_1762);
xnor U1490 (N_1490,In_2187,In_4368);
nand U1491 (N_1491,In_1980,In_4394);
nor U1492 (N_1492,In_2943,In_39);
nor U1493 (N_1493,In_4608,In_2271);
xnor U1494 (N_1494,In_1309,In_744);
nor U1495 (N_1495,In_721,In_631);
xnor U1496 (N_1496,In_1074,In_4410);
nand U1497 (N_1497,In_2934,In_2889);
and U1498 (N_1498,In_409,In_3814);
and U1499 (N_1499,In_1253,In_4557);
and U1500 (N_1500,In_3215,In_4367);
xor U1501 (N_1501,In_35,In_4741);
and U1502 (N_1502,In_4203,In_4844);
nor U1503 (N_1503,In_2590,In_1654);
nand U1504 (N_1504,In_4656,In_2723);
and U1505 (N_1505,In_1923,In_3609);
nand U1506 (N_1506,In_4459,In_3305);
xor U1507 (N_1507,In_3744,In_1468);
and U1508 (N_1508,In_2672,In_3186);
or U1509 (N_1509,In_1136,In_2453);
nand U1510 (N_1510,In_2292,In_3779);
nand U1511 (N_1511,In_3674,In_280);
or U1512 (N_1512,In_2763,In_487);
or U1513 (N_1513,In_1618,In_4405);
nand U1514 (N_1514,In_805,In_716);
nor U1515 (N_1515,In_1914,In_1695);
or U1516 (N_1516,In_1990,In_2144);
nor U1517 (N_1517,In_272,In_787);
nor U1518 (N_1518,In_4920,In_1077);
nor U1519 (N_1519,In_3675,In_864);
nor U1520 (N_1520,In_1579,In_1155);
and U1521 (N_1521,In_571,In_1099);
nand U1522 (N_1522,In_1708,In_1905);
and U1523 (N_1523,In_1562,In_3904);
and U1524 (N_1524,In_190,In_509);
or U1525 (N_1525,In_2817,In_2267);
xnor U1526 (N_1526,In_834,In_1094);
nor U1527 (N_1527,In_1637,In_1960);
or U1528 (N_1528,In_3074,In_4990);
and U1529 (N_1529,In_4234,In_668);
and U1530 (N_1530,In_877,In_3627);
or U1531 (N_1531,In_1410,In_3696);
and U1532 (N_1532,In_4455,In_387);
nor U1533 (N_1533,In_1612,In_770);
and U1534 (N_1534,In_1488,In_636);
or U1535 (N_1535,In_3498,In_347);
and U1536 (N_1536,In_1251,In_1545);
or U1537 (N_1537,In_748,In_2137);
xnor U1538 (N_1538,In_2904,In_436);
nand U1539 (N_1539,In_4390,In_2554);
nand U1540 (N_1540,In_1139,In_139);
nand U1541 (N_1541,In_3572,In_2449);
nor U1542 (N_1542,In_1893,In_3964);
and U1543 (N_1543,In_1981,In_2551);
and U1544 (N_1544,In_412,In_1453);
xnor U1545 (N_1545,In_4349,In_1225);
and U1546 (N_1546,In_3807,In_2868);
or U1547 (N_1547,In_2677,In_4716);
nor U1548 (N_1548,In_4091,In_1610);
xor U1549 (N_1549,In_307,In_1802);
or U1550 (N_1550,In_819,In_1677);
and U1551 (N_1551,In_2610,In_396);
or U1552 (N_1552,In_4466,In_3500);
or U1553 (N_1553,In_3436,In_627);
xor U1554 (N_1554,In_2928,In_1445);
and U1555 (N_1555,In_4926,In_4811);
nor U1556 (N_1556,In_975,In_1625);
or U1557 (N_1557,In_3366,In_3250);
and U1558 (N_1558,In_2377,In_2299);
xor U1559 (N_1559,In_2426,In_1297);
nand U1560 (N_1560,In_3134,In_3289);
or U1561 (N_1561,In_1131,In_1419);
or U1562 (N_1562,In_2072,In_4022);
nand U1563 (N_1563,In_8,In_2930);
and U1564 (N_1564,In_340,In_1133);
or U1565 (N_1565,In_1888,In_3745);
and U1566 (N_1566,In_3636,In_3902);
and U1567 (N_1567,In_1056,In_1271);
nand U1568 (N_1568,In_2524,In_2990);
nor U1569 (N_1569,In_3861,In_908);
and U1570 (N_1570,In_4037,In_3269);
nor U1571 (N_1571,In_2655,In_522);
and U1572 (N_1572,In_733,In_2184);
nand U1573 (N_1573,In_3104,In_2564);
nor U1574 (N_1574,In_3256,In_1033);
or U1575 (N_1575,In_4783,In_3330);
nand U1576 (N_1576,In_3585,In_3956);
nor U1577 (N_1577,In_4301,In_2575);
or U1578 (N_1578,In_4909,In_2772);
nand U1579 (N_1579,In_245,In_888);
or U1580 (N_1580,In_4789,In_3009);
nor U1581 (N_1581,In_1472,In_567);
nor U1582 (N_1582,In_4202,In_4870);
or U1583 (N_1583,In_370,In_4364);
or U1584 (N_1584,In_1242,In_543);
and U1585 (N_1585,In_4944,In_4948);
or U1586 (N_1586,In_871,In_1464);
or U1587 (N_1587,In_3004,In_1997);
or U1588 (N_1588,In_2318,In_1109);
and U1589 (N_1589,In_4253,In_4039);
nand U1590 (N_1590,In_3176,In_2194);
or U1591 (N_1591,In_4962,In_2478);
nand U1592 (N_1592,In_273,In_2748);
and U1593 (N_1593,In_2038,In_3334);
or U1594 (N_1594,In_439,In_848);
nor U1595 (N_1595,In_2834,In_654);
and U1596 (N_1596,In_2743,In_4595);
and U1597 (N_1597,In_2333,In_399);
xor U1598 (N_1598,In_4916,In_4600);
nand U1599 (N_1599,In_2532,In_2670);
and U1600 (N_1600,In_2645,In_3797);
and U1601 (N_1601,In_811,In_1429);
and U1602 (N_1602,In_3209,In_2780);
nand U1603 (N_1603,In_2912,In_312);
and U1604 (N_1604,In_781,In_1632);
xnor U1605 (N_1605,In_3622,In_3938);
nor U1606 (N_1606,In_4484,In_962);
and U1607 (N_1607,In_2725,In_956);
nor U1608 (N_1608,In_1791,In_4911);
or U1609 (N_1609,In_647,In_4198);
or U1610 (N_1610,In_1929,In_2510);
nand U1611 (N_1611,In_4770,In_3070);
and U1612 (N_1612,In_1881,In_747);
and U1613 (N_1613,In_4469,In_3928);
and U1614 (N_1614,In_4495,In_1281);
xor U1615 (N_1615,In_1975,In_53);
nand U1616 (N_1616,In_4407,In_4508);
nor U1617 (N_1617,In_3820,In_735);
and U1618 (N_1618,In_73,In_4907);
nor U1619 (N_1619,In_1153,In_662);
nor U1620 (N_1620,In_4975,In_1955);
nand U1621 (N_1621,In_164,In_1884);
or U1622 (N_1622,In_3887,In_3287);
nand U1623 (N_1623,In_3953,In_2200);
or U1624 (N_1624,In_2534,In_4748);
nor U1625 (N_1625,In_4324,In_995);
nand U1626 (N_1626,In_707,In_2854);
nor U1627 (N_1627,In_4728,In_649);
nand U1628 (N_1628,In_2759,In_2697);
or U1629 (N_1629,In_718,In_3667);
xor U1630 (N_1630,In_3445,In_981);
nand U1631 (N_1631,In_2046,In_3288);
or U1632 (N_1632,In_2405,In_678);
nor U1633 (N_1633,In_1694,In_4582);
and U1634 (N_1634,In_3523,In_1513);
nor U1635 (N_1635,In_4365,In_2489);
and U1636 (N_1636,In_3896,In_3261);
or U1637 (N_1637,In_717,In_1238);
nor U1638 (N_1638,In_4570,In_680);
nor U1639 (N_1639,In_3487,In_1956);
nand U1640 (N_1640,In_177,In_1726);
or U1641 (N_1641,In_148,In_149);
and U1642 (N_1642,In_884,In_278);
nor U1643 (N_1643,In_2960,In_511);
xnor U1644 (N_1644,In_2747,In_2043);
xor U1645 (N_1645,In_1417,In_4485);
nand U1646 (N_1646,In_1054,In_603);
or U1647 (N_1647,In_1849,In_1532);
nand U1648 (N_1648,In_4169,In_2273);
or U1649 (N_1649,In_1349,In_862);
nor U1650 (N_1650,In_4115,In_4208);
nor U1651 (N_1651,In_1557,In_4759);
nor U1652 (N_1652,In_1316,In_292);
nand U1653 (N_1653,In_1733,In_3563);
and U1654 (N_1654,In_4027,In_119);
nand U1655 (N_1655,In_3859,In_558);
nor U1656 (N_1656,In_286,In_3604);
or U1657 (N_1657,In_582,In_4318);
nor U1658 (N_1658,In_3851,In_1743);
or U1659 (N_1659,In_4451,In_1303);
or U1660 (N_1660,In_3541,In_1622);
or U1661 (N_1661,In_4503,In_624);
and U1662 (N_1662,In_2314,In_759);
and U1663 (N_1663,In_1483,In_2799);
and U1664 (N_1664,In_851,In_3321);
xnor U1665 (N_1665,In_4507,In_4742);
nor U1666 (N_1666,In_3155,In_579);
or U1667 (N_1667,In_282,In_4053);
nor U1668 (N_1668,In_1687,In_3501);
xor U1669 (N_1669,In_2157,In_3048);
or U1670 (N_1670,In_1650,In_1368);
nand U1671 (N_1671,In_1121,In_1036);
and U1672 (N_1672,In_4030,In_3593);
nand U1673 (N_1673,In_3075,In_727);
xnor U1674 (N_1674,In_3535,In_3216);
and U1675 (N_1675,In_3923,In_489);
or U1676 (N_1676,In_4938,In_21);
nand U1677 (N_1677,In_1006,In_268);
nor U1678 (N_1678,In_913,In_2970);
nand U1679 (N_1679,In_1334,In_1763);
nand U1680 (N_1680,In_4117,In_4816);
nor U1681 (N_1681,In_203,In_1845);
or U1682 (N_1682,In_2663,In_4490);
or U1683 (N_1683,In_4581,In_3275);
nor U1684 (N_1684,In_2746,In_1437);
xnor U1685 (N_1685,In_1192,In_2140);
and U1686 (N_1686,In_2407,In_3489);
and U1687 (N_1687,In_1116,In_906);
or U1688 (N_1688,In_2658,In_1781);
and U1689 (N_1689,In_1784,In_1885);
nor U1690 (N_1690,In_3528,In_3234);
nand U1691 (N_1691,In_4935,In_1462);
and U1692 (N_1692,In_4662,In_3081);
nand U1693 (N_1693,In_4576,In_1299);
nand U1694 (N_1694,In_4013,In_602);
nand U1695 (N_1695,In_2092,In_2738);
nor U1696 (N_1696,In_1388,In_685);
nand U1697 (N_1697,In_3873,In_1381);
nor U1698 (N_1698,In_1742,In_2347);
and U1699 (N_1699,In_65,In_4574);
nand U1700 (N_1700,In_1277,In_4289);
nor U1701 (N_1701,In_2608,In_934);
and U1702 (N_1702,In_290,In_323);
and U1703 (N_1703,In_892,In_3782);
and U1704 (N_1704,In_505,In_3460);
nand U1705 (N_1705,In_1261,In_1506);
or U1706 (N_1706,In_72,In_4977);
nand U1707 (N_1707,In_868,In_2516);
nor U1708 (N_1708,In_1037,In_3165);
nand U1709 (N_1709,In_3518,In_335);
xor U1710 (N_1710,In_2436,In_2848);
and U1711 (N_1711,In_3919,In_4461);
nand U1712 (N_1712,In_3796,In_4239);
and U1713 (N_1713,In_431,In_2356);
and U1714 (N_1714,In_3229,In_1509);
or U1715 (N_1715,In_1214,In_2908);
and U1716 (N_1716,In_2247,In_3254);
xor U1717 (N_1717,In_1544,In_2704);
or U1718 (N_1718,In_1002,In_1014);
nand U1719 (N_1719,In_2203,In_4688);
nor U1720 (N_1720,In_3761,In_1038);
nor U1721 (N_1721,In_415,In_3);
nor U1722 (N_1722,In_1134,In_1010);
nand U1723 (N_1723,In_1771,In_2122);
nor U1724 (N_1724,In_2413,In_4677);
xnor U1725 (N_1725,In_1510,In_2540);
xor U1726 (N_1726,In_4659,In_656);
or U1727 (N_1727,In_870,In_4231);
and U1728 (N_1728,In_4052,In_4212);
nand U1729 (N_1729,In_4853,In_2698);
nand U1730 (N_1730,In_4950,In_3341);
and U1731 (N_1731,In_2409,In_1120);
nand U1732 (N_1732,In_4620,In_1697);
and U1733 (N_1733,In_1570,In_2475);
and U1734 (N_1734,In_4747,In_714);
nand U1735 (N_1735,In_4598,In_1503);
xnor U1736 (N_1736,In_304,In_4220);
nor U1737 (N_1737,In_13,In_3587);
xor U1738 (N_1738,In_751,In_3297);
nor U1739 (N_1739,In_1938,In_3418);
nor U1740 (N_1740,In_4474,In_2056);
xor U1741 (N_1741,In_785,In_4308);
or U1742 (N_1742,In_4527,In_1383);
and U1743 (N_1743,In_3834,In_4389);
xor U1744 (N_1744,In_1179,In_2098);
and U1745 (N_1745,In_4505,In_706);
nand U1746 (N_1746,In_4010,In_969);
or U1747 (N_1747,In_271,In_1228);
xor U1748 (N_1748,In_4925,In_2666);
nand U1749 (N_1749,In_952,In_3526);
xnor U1750 (N_1750,In_4734,In_2560);
nand U1751 (N_1751,In_84,In_1416);
xor U1752 (N_1752,In_1176,In_2150);
or U1753 (N_1753,In_2457,In_320);
nand U1754 (N_1754,In_1789,In_1088);
and U1755 (N_1755,In_4369,In_2865);
nor U1756 (N_1756,In_362,In_2458);
or U1757 (N_1757,In_2481,In_244);
and U1758 (N_1758,In_2240,In_3648);
and U1759 (N_1759,In_4795,In_946);
or U1760 (N_1760,In_4653,In_1785);
and U1761 (N_1761,In_4857,In_123);
or U1762 (N_1762,In_3027,In_1861);
nand U1763 (N_1763,In_2703,In_492);
nand U1764 (N_1764,In_1496,In_4242);
or U1765 (N_1765,In_3005,In_4839);
xor U1766 (N_1766,In_1068,In_4106);
and U1767 (N_1767,In_1386,In_4153);
or U1768 (N_1768,In_3756,In_1834);
and U1769 (N_1769,In_741,In_1675);
or U1770 (N_1770,In_2048,In_2787);
nand U1771 (N_1771,In_4889,In_966);
nand U1772 (N_1772,In_4663,In_2344);
xnor U1773 (N_1773,In_1234,In_4189);
nand U1774 (N_1774,In_835,In_4882);
xnor U1775 (N_1775,In_428,In_2756);
nand U1776 (N_1776,In_1924,In_3799);
or U1777 (N_1777,In_23,In_3119);
and U1778 (N_1778,In_3721,In_2786);
or U1779 (N_1779,In_2337,In_648);
or U1780 (N_1780,In_549,In_1441);
or U1781 (N_1781,In_2226,In_2957);
or U1782 (N_1782,In_2630,In_4961);
nor U1783 (N_1783,In_3769,In_4959);
nand U1784 (N_1784,In_270,In_1723);
nand U1785 (N_1785,In_3456,In_3751);
nor U1786 (N_1786,In_3634,In_3586);
or U1787 (N_1787,In_1586,In_397);
nand U1788 (N_1788,In_4058,In_182);
xnor U1789 (N_1789,In_2910,In_1352);
nand U1790 (N_1790,In_3755,In_950);
and U1791 (N_1791,In_398,In_486);
nor U1792 (N_1792,In_4815,In_2587);
or U1793 (N_1793,In_1438,In_1604);
or U1794 (N_1794,In_4809,In_1418);
and U1795 (N_1795,In_2421,In_1879);
nand U1796 (N_1796,In_3663,In_424);
or U1797 (N_1797,In_141,In_753);
nand U1798 (N_1798,In_4796,In_1148);
and U1799 (N_1799,In_3948,In_4743);
nand U1800 (N_1800,In_4051,In_3798);
xnor U1801 (N_1801,In_3724,In_573);
or U1802 (N_1802,In_1062,In_820);
or U1803 (N_1803,In_4284,In_2326);
and U1804 (N_1804,In_238,In_4856);
or U1805 (N_1805,In_308,In_179);
nand U1806 (N_1806,In_55,In_2265);
xor U1807 (N_1807,In_1626,In_4917);
and U1808 (N_1808,In_1201,In_4793);
and U1809 (N_1809,In_1296,In_2079);
and U1810 (N_1810,In_3177,In_3037);
or U1811 (N_1811,In_446,In_4226);
nor U1812 (N_1812,In_3736,In_4808);
or U1813 (N_1813,In_1229,In_1572);
and U1814 (N_1814,In_3900,In_865);
nor U1815 (N_1815,In_4476,In_1912);
nor U1816 (N_1816,In_2688,In_4292);
nand U1817 (N_1817,In_250,In_2026);
and U1818 (N_1818,In_3894,In_4161);
or U1819 (N_1819,In_2030,In_337);
and U1820 (N_1820,In_794,In_1540);
and U1821 (N_1821,In_2726,In_3372);
and U1822 (N_1822,In_3510,In_4919);
or U1823 (N_1823,In_1083,In_1081);
nor U1824 (N_1824,In_3711,In_4219);
and U1825 (N_1825,In_1175,In_3480);
nand U1826 (N_1826,In_2503,In_1907);
xnor U1827 (N_1827,In_3556,In_3521);
nor U1828 (N_1828,In_4218,In_3458);
or U1829 (N_1829,In_3378,In_2237);
nand U1830 (N_1830,In_295,In_1128);
nand U1831 (N_1831,In_1699,In_2656);
nor U1832 (N_1832,In_4432,In_798);
nor U1833 (N_1833,In_3115,In_1530);
nor U1834 (N_1834,In_429,In_3356);
or U1835 (N_1835,In_3857,In_1872);
xor U1836 (N_1836,In_1413,In_786);
nor U1837 (N_1837,In_4627,In_1542);
or U1838 (N_1838,In_1243,In_1451);
or U1839 (N_1839,In_2450,In_410);
nor U1840 (N_1840,In_1715,In_4199);
nor U1841 (N_1841,In_3988,In_1254);
and U1842 (N_1842,In_2940,In_479);
nor U1843 (N_1843,In_4158,In_1565);
nand U1844 (N_1844,In_972,In_2558);
nor U1845 (N_1845,In_4597,In_2223);
nand U1846 (N_1846,In_1193,In_3323);
nor U1847 (N_1847,In_1015,In_231);
nand U1848 (N_1848,In_2143,In_2588);
or U1849 (N_1849,In_4529,In_4046);
nor U1850 (N_1850,In_2998,In_4361);
and U1851 (N_1851,In_2730,In_3516);
or U1852 (N_1852,In_1718,In_48);
or U1853 (N_1853,In_890,In_3188);
xnor U1854 (N_1854,In_4638,In_1745);
or U1855 (N_1855,In_2207,In_4779);
nand U1856 (N_1856,In_1404,In_689);
nor U1857 (N_1857,In_506,In_1373);
nor U1858 (N_1858,In_38,In_4516);
nand U1859 (N_1859,In_3640,In_62);
nor U1860 (N_1860,In_3921,In_3853);
or U1861 (N_1861,In_3389,In_2812);
nor U1862 (N_1862,In_3028,In_4112);
or U1863 (N_1863,In_3246,In_4988);
xnor U1864 (N_1864,In_2493,In_3652);
or U1865 (N_1865,In_808,In_3383);
nor U1866 (N_1866,In_4534,In_4337);
xor U1867 (N_1867,In_117,In_1346);
nor U1868 (N_1868,In_264,In_3402);
nand U1869 (N_1869,In_201,In_2636);
or U1870 (N_1870,In_4126,In_353);
or U1871 (N_1871,In_746,In_355);
or U1872 (N_1872,In_1529,In_3379);
nand U1873 (N_1873,In_2613,In_2631);
nor U1874 (N_1874,In_1985,In_2685);
nor U1875 (N_1875,In_3315,In_93);
and U1876 (N_1876,In_1961,In_3520);
and U1877 (N_1877,In_3662,In_403);
nor U1878 (N_1878,In_1813,In_452);
nand U1879 (N_1879,In_1942,In_2965);
or U1880 (N_1880,In_4838,In_3191);
or U1881 (N_1881,In_4500,In_4903);
xnor U1882 (N_1882,In_3727,In_3898);
nand U1883 (N_1883,In_4332,In_4035);
nor U1884 (N_1884,In_1027,In_322);
nand U1885 (N_1885,In_2514,In_3983);
or U1886 (N_1886,In_4631,In_3625);
nand U1887 (N_1887,In_4342,In_696);
and U1888 (N_1888,In_3673,In_4695);
and U1889 (N_1889,In_3443,In_1405);
and U1890 (N_1890,In_964,In_3821);
and U1891 (N_1891,In_67,In_4163);
or U1892 (N_1892,In_899,In_2406);
or U1893 (N_1893,In_4798,In_1063);
or U1894 (N_1894,In_4101,In_3118);
nand U1895 (N_1895,In_2533,In_4427);
nand U1896 (N_1896,In_4462,In_2615);
nand U1897 (N_1897,In_4340,In_4012);
or U1898 (N_1898,In_4867,In_4611);
or U1899 (N_1899,In_1117,In_540);
xor U1900 (N_1900,In_2068,In_2506);
nand U1901 (N_1901,In_4159,In_3633);
xnor U1902 (N_1902,In_4409,In_3013);
nand U1903 (N_1903,In_1995,In_1428);
nor U1904 (N_1904,In_3071,In_2815);
or U1905 (N_1905,In_4055,In_4446);
and U1906 (N_1906,In_1767,In_3979);
xor U1907 (N_1907,In_3319,In_4629);
or U1908 (N_1908,In_472,In_3631);
nor U1909 (N_1909,In_2522,In_2798);
nor U1910 (N_1910,In_4628,In_3295);
nand U1911 (N_1911,In_1008,In_1497);
or U1912 (N_1912,In_3243,In_764);
and U1913 (N_1913,In_591,In_2695);
nor U1914 (N_1914,In_3380,In_2810);
xnor U1915 (N_1915,In_142,In_3382);
xor U1916 (N_1916,In_2151,In_2261);
and U1917 (N_1917,In_2320,In_2272);
and U1918 (N_1918,In_3708,In_3311);
and U1919 (N_1919,In_4079,In_2739);
and U1920 (N_1920,In_2258,In_1221);
or U1921 (N_1921,In_144,In_1147);
and U1922 (N_1922,In_2202,In_4238);
nor U1923 (N_1923,In_4164,In_25);
nor U1924 (N_1924,In_375,In_351);
and U1925 (N_1925,In_1290,In_3198);
nand U1926 (N_1926,In_3836,In_955);
and U1927 (N_1927,In_4000,In_3439);
nand U1928 (N_1928,In_3854,In_2266);
xor U1929 (N_1929,In_2112,In_889);
xor U1930 (N_1930,In_3137,In_3178);
or U1931 (N_1931,In_2041,In_1967);
and U1932 (N_1932,In_2737,In_4652);
xnor U1933 (N_1933,In_828,In_4565);
and U1934 (N_1934,In_2110,In_2627);
or U1935 (N_1935,In_2120,In_345);
xor U1936 (N_1936,In_1795,In_2108);
nand U1937 (N_1937,In_2803,In_4197);
nand U1938 (N_1938,In_4472,In_3073);
nand U1939 (N_1939,In_4736,In_3473);
or U1940 (N_1940,In_3040,In_158);
xnor U1941 (N_1941,In_1709,In_2639);
xnor U1942 (N_1942,In_1061,In_3864);
and U1943 (N_1943,In_1046,In_893);
nor U1944 (N_1944,In_4965,In_2530);
or U1945 (N_1945,In_3014,In_3925);
nor U1946 (N_1946,In_2305,In_202);
or U1947 (N_1947,In_1620,In_4740);
or U1948 (N_1948,In_4967,In_750);
and U1949 (N_1949,In_4071,In_1177);
nor U1950 (N_1950,In_1706,In_4676);
nor U1951 (N_1951,In_4596,In_572);
nand U1952 (N_1952,In_2445,In_1843);
nand U1953 (N_1953,In_637,In_4294);
and U1954 (N_1954,In_1870,In_1582);
nor U1955 (N_1955,In_1076,In_2210);
or U1956 (N_1956,In_4184,In_818);
and U1957 (N_1957,In_1640,In_2694);
or U1958 (N_1958,In_3056,In_4998);
nand U1959 (N_1959,In_2133,In_4567);
nor U1960 (N_1960,In_4803,In_3277);
nand U1961 (N_1961,In_4521,In_1279);
or U1962 (N_1962,In_4240,In_4976);
or U1963 (N_1963,In_2836,In_101);
nand U1964 (N_1964,In_4,In_3626);
or U1965 (N_1965,In_2562,In_948);
and U1966 (N_1966,In_1621,In_1515);
xnor U1967 (N_1967,In_1925,In_2883);
nor U1968 (N_1968,In_2355,In_2373);
nor U1969 (N_1969,In_4610,In_406);
and U1970 (N_1970,In_3117,In_1761);
nor U1971 (N_1971,In_1245,In_4008);
or U1972 (N_1972,In_4454,In_2513);
xnor U1973 (N_1973,In_2101,In_3282);
xnor U1974 (N_1974,In_621,In_920);
nor U1975 (N_1975,In_2488,In_578);
nor U1976 (N_1976,In_629,In_3800);
nand U1977 (N_1977,In_1644,In_305);
and U1978 (N_1978,In_4790,In_3051);
nor U1979 (N_1979,In_1728,In_1829);
nor U1980 (N_1980,In_4714,In_4233);
and U1981 (N_1981,In_947,In_2665);
or U1982 (N_1982,In_3668,In_4960);
nor U1983 (N_1983,In_3698,In_28);
nor U1984 (N_1984,In_2088,In_2087);
and U1985 (N_1985,In_4551,In_2936);
and U1986 (N_1986,In_4672,In_331);
nor U1987 (N_1987,In_4537,In_166);
nand U1988 (N_1988,In_2607,In_1809);
nor U1989 (N_1989,In_4321,In_4504);
or U1990 (N_1990,In_4075,In_560);
nor U1991 (N_1991,In_10,In_4285);
and U1992 (N_1992,In_1755,In_2680);
nor U1993 (N_1993,In_4738,In_2623);
nand U1994 (N_1994,In_3224,In_1780);
and U1995 (N_1995,In_1382,In_817);
nor U1996 (N_1996,In_225,In_3934);
xor U1997 (N_1997,In_1252,In_469);
nor U1998 (N_1998,In_1239,In_4062);
xnor U1999 (N_1999,In_2192,In_352);
and U2000 (N_2000,In_466,In_120);
or U2001 (N_2001,In_3107,In_4315);
and U2002 (N_2002,In_712,In_1174);
nand U2003 (N_2003,In_4862,In_2142);
nand U2004 (N_2004,In_530,In_514);
nor U2005 (N_2005,In_623,In_1770);
nor U2006 (N_2006,In_474,In_3868);
and U2007 (N_2007,In_4863,In_688);
or U2008 (N_2008,In_3064,In_2963);
and U2009 (N_2009,In_1797,In_777);
or U2010 (N_2010,In_40,In_3855);
nand U2011 (N_2011,In_2915,In_1576);
nor U2012 (N_2012,In_275,In_2502);
and U2013 (N_2013,In_43,In_1705);
and U2014 (N_2014,In_4441,In_3120);
xnor U2015 (N_2015,In_2993,In_3102);
nand U2016 (N_2016,In_3093,In_4754);
or U2017 (N_2017,In_2117,In_773);
nor U2018 (N_2018,In_3421,In_4566);
or U2019 (N_2019,In_1645,In_684);
xor U2020 (N_2020,In_2350,In_59);
nand U2021 (N_2021,In_1812,In_3331);
nor U2022 (N_2022,In_2950,In_4020);
or U2023 (N_2023,In_2433,In_3399);
and U2024 (N_2024,In_3687,In_2536);
and U2025 (N_2025,In_15,In_4699);
nand U2026 (N_2026,In_1701,In_4718);
nor U2027 (N_2027,In_4200,In_4953);
nand U2028 (N_2028,In_451,In_266);
nand U2029 (N_2029,In_4584,In_1663);
nand U2030 (N_2030,In_2010,In_91);
nand U2031 (N_2031,In_4373,In_4834);
nor U2032 (N_2032,In_978,In_4666);
or U2033 (N_2033,In_1463,In_3714);
nand U2034 (N_2034,In_2774,In_1948);
and U2035 (N_2035,In_1521,In_2541);
nand U2036 (N_2036,In_2561,In_3580);
xnor U2037 (N_2037,In_1113,In_4830);
nor U2038 (N_2038,In_243,In_2031);
xor U2039 (N_2039,In_3193,In_112);
or U2040 (N_2040,In_2859,In_1594);
and U2041 (N_2041,In_661,In_1376);
or U2042 (N_2042,In_1498,In_4090);
nor U2043 (N_2043,In_719,In_3140);
xor U2044 (N_2044,In_2215,In_361);
nor U2045 (N_2045,In_2954,In_165);
nor U2046 (N_2046,In_4538,In_3754);
nor U2047 (N_2047,In_1977,In_74);
nor U2048 (N_2048,In_3664,In_2275);
and U2049 (N_2049,In_534,In_126);
and U2050 (N_2050,In_3577,In_1922);
and U2051 (N_2051,In_559,In_4855);
nand U2052 (N_2052,In_749,In_1987);
nand U2053 (N_2053,In_2871,In_1227);
nand U2054 (N_2054,In_4711,In_176);
or U2055 (N_2055,In_4267,In_1051);
or U2056 (N_2056,In_1931,In_2045);
and U2057 (N_2057,In_3249,In_1181);
or U2058 (N_2058,In_2913,In_3039);
nor U2059 (N_2059,In_2875,In_3469);
nand U2060 (N_2060,In_1751,In_887);
and U2061 (N_2061,In_4182,In_1564);
and U2062 (N_2062,In_1160,In_622);
or U2063 (N_2063,In_151,In_4885);
or U2064 (N_2064,In_923,In_3388);
nand U2065 (N_2065,In_3531,In_1146);
nor U2066 (N_2066,In_1674,In_336);
or U2067 (N_2067,In_4745,In_3300);
or U2068 (N_2068,In_388,In_3244);
and U2069 (N_2069,In_3326,In_1024);
or U2070 (N_2070,In_3203,In_1566);
and U2071 (N_2071,In_3466,In_4006);
and U2072 (N_2072,In_2880,In_4331);
nor U2073 (N_2073,In_4533,In_4387);
or U2074 (N_2074,In_4080,In_3549);
nand U2075 (N_2075,In_4602,In_2105);
xnor U2076 (N_2076,In_2234,In_3335);
nand U2077 (N_2077,In_1149,In_3175);
or U2078 (N_2078,In_2191,In_2862);
nor U2079 (N_2079,In_4771,In_3704);
or U2080 (N_2080,In_2348,In_4299);
and U2081 (N_2081,In_3392,In_4874);
nand U2082 (N_2082,In_657,In_2684);
nor U2083 (N_2083,In_4561,In_66);
or U2084 (N_2084,In_1291,In_3353);
nor U2085 (N_2085,In_1485,In_517);
nor U2086 (N_2086,In_1667,In_3310);
and U2087 (N_2087,In_3707,In_2389);
nand U2088 (N_2088,In_3208,In_4154);
and U2089 (N_2089,In_1283,In_3091);
or U2090 (N_2090,In_1087,In_3354);
and U2091 (N_2091,In_4168,In_2231);
xor U2092 (N_2092,In_1671,In_2789);
or U2093 (N_2093,In_2861,In_4800);
or U2094 (N_2094,In_4746,In_2091);
or U2095 (N_2095,In_4520,In_2975);
or U2096 (N_2096,In_667,In_2099);
nand U2097 (N_2097,In_640,In_4572);
or U2098 (N_2098,In_2419,In_1504);
nor U2099 (N_2099,In_2257,In_1822);
nand U2100 (N_2100,In_4111,In_936);
nor U2101 (N_2101,In_1183,In_3703);
and U2102 (N_2102,In_4263,In_2831);
nor U2103 (N_2103,In_1090,In_801);
or U2104 (N_2104,In_3930,In_3920);
or U2105 (N_2105,In_2392,In_1326);
nor U2106 (N_2106,In_2208,In_2220);
and U2107 (N_2107,In_2757,In_4945);
and U2108 (N_2108,In_358,In_2805);
and U2109 (N_2109,In_2979,In_611);
nor U2110 (N_2110,In_2741,In_725);
or U2111 (N_2111,In_4350,In_3258);
nor U2112 (N_2112,In_4837,In_1329);
and U2113 (N_2113,In_4463,In_1945);
or U2114 (N_2114,In_3143,In_4854);
and U2115 (N_2115,In_2256,In_1004);
and U2116 (N_2116,In_564,In_2819);
nand U2117 (N_2117,In_3294,In_1856);
nor U2118 (N_2118,In_4178,In_1906);
and U2119 (N_2119,In_1986,In_535);
nand U2120 (N_2120,In_4750,In_4149);
and U2121 (N_2121,In_1958,In_4139);
nor U2122 (N_2122,In_4247,In_301);
or U2123 (N_2123,In_2073,In_1357);
nor U2124 (N_2124,In_4866,In_3826);
nand U2125 (N_2125,In_1137,In_2977);
and U2126 (N_2126,In_3429,In_690);
or U2127 (N_2127,In_2179,In_4902);
nor U2128 (N_2128,In_1549,In_3635);
nor U2129 (N_2129,In_4430,In_2917);
nor U2130 (N_2130,In_448,In_791);
and U2131 (N_2131,In_1414,In_3058);
nor U2132 (N_2132,In_693,In_1595);
nand U2133 (N_2133,In_3697,In_1310);
and U2134 (N_2134,In_1793,In_538);
nor U2135 (N_2135,In_919,In_316);
xor U2136 (N_2136,In_417,In_191);
nor U2137 (N_2137,In_3374,In_4421);
and U2138 (N_2138,In_1345,In_4428);
nand U2139 (N_2139,In_3423,In_1842);
and U2140 (N_2140,In_3713,In_2733);
and U2141 (N_2141,In_2078,In_2614);
or U2142 (N_2142,In_4391,In_1511);
or U2143 (N_2143,In_3874,In_86);
xor U2144 (N_2144,In_293,In_3462);
or U2145 (N_2145,In_3999,In_3357);
nor U2146 (N_2146,In_4655,In_1057);
and U2147 (N_2147,In_2727,In_1820);
nand U2148 (N_2148,In_3565,In_220);
or U2149 (N_2149,In_2385,In_2096);
nand U2150 (N_2150,In_3406,In_2360);
xor U2151 (N_2151,In_183,In_1187);
nor U2152 (N_2152,In_1338,In_2526);
nand U2153 (N_2153,In_1670,In_4333);
or U2154 (N_2154,In_2435,In_3219);
nor U2155 (N_2155,In_3403,In_4735);
nor U2156 (N_2156,In_4327,In_3710);
nand U2157 (N_2157,In_4539,In_2800);
nand U2158 (N_2158,In_4420,In_4127);
nor U2159 (N_2159,In_3890,In_4057);
nand U2160 (N_2160,In_1883,In_3472);
nand U2161 (N_2161,In_3351,In_1657);
and U2162 (N_2162,In_1918,In_3931);
and U2163 (N_2163,In_2548,In_3268);
and U2164 (N_2164,In_3252,In_400);
nand U2165 (N_2165,In_1159,In_1396);
nand U2166 (N_2166,In_3452,In_699);
nor U2167 (N_2167,In_2233,In_762);
nand U2168 (N_2168,In_3348,In_2396);
nand U2169 (N_2169,In_1602,In_4828);
nor U2170 (N_2170,In_4986,In_900);
and U2171 (N_2171,In_1643,In_4763);
nor U2172 (N_2172,In_309,In_4366);
or U2173 (N_2173,In_1738,In_1141);
and U2174 (N_2174,In_2683,In_1729);
and U2175 (N_2175,In_3059,In_2093);
nand U2176 (N_2176,In_2712,In_3768);
xor U2177 (N_2177,In_3450,In_3285);
and U2178 (N_2178,In_313,In_1167);
nor U2179 (N_2179,In_708,In_1029);
nor U2180 (N_2180,In_3441,In_2307);
nand U2181 (N_2181,In_4386,In_3517);
nand U2182 (N_2182,In_2224,In_533);
xnor U2183 (N_2183,In_803,In_2728);
and U2184 (N_2184,In_3991,In_2178);
nor U2185 (N_2185,In_1210,In_498);
and U2186 (N_2186,In_2777,In_776);
xor U2187 (N_2187,In_1964,In_4784);
nor U2188 (N_2188,In_4966,In_3514);
nor U2189 (N_2189,In_4888,In_1851);
nand U2190 (N_2190,In_2341,In_2381);
xor U2191 (N_2191,In_4497,In_1577);
nor U2192 (N_2192,In_4880,In_642);
and U2193 (N_2193,In_1796,In_4402);
or U2194 (N_2194,In_1071,In_4569);
nand U2195 (N_2195,In_236,In_3248);
nand U2196 (N_2196,In_3665,In_2929);
nand U2197 (N_2197,In_2878,In_4954);
and U2198 (N_2198,In_490,In_497);
xor U2199 (N_2199,In_422,In_3878);
nand U2200 (N_2200,In_3022,In_2999);
and U2201 (N_2201,In_3877,In_2491);
nor U2202 (N_2202,In_3444,In_778);
and U2203 (N_2203,In_3660,In_47);
and U2204 (N_2204,In_4316,In_4151);
nand U2205 (N_2205,In_2160,In_3913);
nor U2206 (N_2206,In_4996,In_4563);
nand U2207 (N_2207,In_2978,In_3509);
nor U2208 (N_2208,In_1552,In_287);
nand U2209 (N_2209,In_3428,In_3879);
xnor U2210 (N_2210,In_3966,In_2316);
and U2211 (N_2211,In_2873,In_4580);
nor U2212 (N_2212,In_2201,In_1807);
or U2213 (N_2213,In_248,In_3099);
or U2214 (N_2214,In_2731,In_4915);
and U2215 (N_2215,In_2678,In_373);
and U2216 (N_2216,In_4216,In_3603);
xor U2217 (N_2217,In_2580,In_2537);
and U2218 (N_2218,In_4765,In_1898);
nor U2219 (N_2219,In_146,In_2793);
nand U2220 (N_2220,In_3114,In_3228);
and U2221 (N_2221,In_150,In_4144);
nor U2222 (N_2222,In_2285,In_1850);
and U2223 (N_2223,In_2771,In_3182);
and U2224 (N_2224,In_2354,In_4374);
or U2225 (N_2225,In_4290,In_3748);
or U2226 (N_2226,In_1684,In_2060);
or U2227 (N_2227,In_4585,In_2158);
or U2228 (N_2228,In_4820,In_1788);
or U2229 (N_2229,In_4119,In_3491);
or U2230 (N_2230,In_4128,In_1534);
nor U2231 (N_2231,In_3511,In_2141);
and U2232 (N_2232,In_869,In_4093);
or U2233 (N_2233,In_970,In_2281);
nor U2234 (N_2234,In_2116,In_1247);
or U2235 (N_2235,In_3730,In_2039);
nor U2236 (N_2236,In_1047,In_1927);
and U2237 (N_2237,In_3638,In_2637);
or U2238 (N_2238,In_2842,In_4941);
nand U2239 (N_2239,In_2662,In_462);
or U2240 (N_2240,In_3162,In_4860);
or U2241 (N_2241,In_1293,In_2358);
nor U2242 (N_2242,In_3958,In_4425);
and U2243 (N_2243,In_659,In_1311);
xnor U2244 (N_2244,In_4345,In_4705);
xnor U2245 (N_2245,In_3689,In_4980);
nor U2246 (N_2246,In_377,In_2309);
nand U2247 (N_2247,In_4412,In_4448);
nand U2248 (N_2248,In_3281,In_2444);
nor U2249 (N_2249,In_4140,In_1123);
nand U2250 (N_2250,In_4180,In_3173);
nand U2251 (N_2251,In_3737,In_2206);
nor U2252 (N_2252,In_1516,In_3515);
nor U2253 (N_2253,In_2418,In_4295);
and U2254 (N_2254,In_2017,In_1641);
xor U2255 (N_2255,In_4913,In_2557);
nand U2256 (N_2256,In_3989,In_3164);
and U2257 (N_2257,In_156,In_660);
and U2258 (N_2258,In_2681,In_3431);
nor U2259 (N_2259,In_1930,In_3002);
nand U2260 (N_2260,In_4254,In_1461);
and U2261 (N_2261,In_4621,In_943);
or U2262 (N_2262,In_4323,In_1400);
nor U2263 (N_2263,In_581,In_3280);
or U2264 (N_2264,In_4129,In_1424);
or U2265 (N_2265,In_4886,In_3601);
nand U2266 (N_2266,In_1129,In_3085);
or U2267 (N_2267,In_4036,In_4804);
nand U2268 (N_2268,In_3438,In_4142);
nor U2269 (N_2269,In_2669,In_2618);
and U2270 (N_2270,In_2846,In_2821);
nand U2271 (N_2271,In_3607,In_2252);
nand U2272 (N_2272,In_4664,In_4314);
nor U2273 (N_2273,In_2461,In_2047);
nor U2274 (N_2274,In_1794,In_4478);
or U2275 (N_2275,In_878,In_1332);
nor U2276 (N_2276,In_1732,In_931);
nand U2277 (N_2277,In_4893,In_114);
xnor U2278 (N_2278,In_2420,In_2024);
nor U2279 (N_2279,In_1244,In_812);
or U2280 (N_2280,In_4228,In_3495);
nor U2281 (N_2281,In_4733,In_100);
or U2282 (N_2282,In_3146,In_1011);
or U2283 (N_2283,In_737,In_4250);
nor U2284 (N_2284,In_1364,In_1085);
or U2285 (N_2285,In_2845,In_3588);
and U2286 (N_2286,In_1568,In_2959);
nor U2287 (N_2287,In_1284,In_172);
nand U2288 (N_2288,In_2718,In_3226);
nor U2289 (N_2289,In_1722,In_3584);
xor U2290 (N_2290,In_1976,In_2807);
and U2291 (N_2291,In_1765,In_1415);
nand U2292 (N_2292,In_1739,In_458);
and U2293 (N_2293,In_3427,In_821);
nand U2294 (N_2294,In_810,In_3567);
or U2295 (N_2295,In_4583,In_4038);
nand U2296 (N_2296,In_2379,In_444);
nand U2297 (N_2297,In_4524,In_1295);
nand U2298 (N_2298,In_1966,In_4641);
nor U2299 (N_2299,In_376,In_686);
nor U2300 (N_2300,In_1580,In_1866);
or U2301 (N_2301,In_682,In_2907);
and U2302 (N_2302,In_3886,In_152);
xor U2303 (N_2303,In_3247,In_1920);
nor U2304 (N_2304,In_886,In_4698);
and U2305 (N_2305,In_4170,In_106);
and U2306 (N_2306,In_1490,In_1353);
or U2307 (N_2307,In_3122,In_607);
nor U2308 (N_2308,In_4678,In_2864);
or U2309 (N_2309,In_2982,In_4082);
nand U2310 (N_2310,In_1287,In_3771);
and U2311 (N_2311,In_3322,In_3766);
and U2312 (N_2312,In_237,In_346);
and U2313 (N_2313,In_1591,In_3190);
nor U2314 (N_2314,In_897,In_1481);
nand U2315 (N_2315,In_1138,In_299);
and U2316 (N_2316,In_4195,In_3935);
or U2317 (N_2317,In_1721,In_984);
xor U2318 (N_2318,In_393,In_2423);
nor U2319 (N_2319,In_989,In_4639);
or U2320 (N_2320,In_4040,In_1996);
and U2321 (N_2321,In_2668,In_4257);
and U2322 (N_2322,In_709,In_608);
nor U2323 (N_2323,In_138,In_2244);
xor U2324 (N_2324,In_4590,In_544);
and U2325 (N_2325,In_2611,In_4805);
nor U2326 (N_2326,In_2740,In_4060);
nor U2327 (N_2327,In_1752,In_3784);
or U2328 (N_2328,In_2205,In_3540);
nor U2329 (N_2329,In_94,In_3430);
xnor U2330 (N_2330,In_4739,In_4131);
nor U2331 (N_2331,In_81,In_4761);
xnor U2332 (N_2332,In_520,In_2983);
nor U2333 (N_2333,In_121,In_3238);
nor U2334 (N_2334,In_1476,In_4981);
nor U2335 (N_2335,In_4408,In_2890);
nand U2336 (N_2336,In_4713,In_3840);
nand U2337 (N_2337,In_3471,In_4162);
xnor U2338 (N_2338,In_3151,In_849);
nand U2339 (N_2339,In_4445,In_4875);
and U2340 (N_2340,In_3271,In_2887);
nor U2341 (N_2341,In_3918,In_2855);
or U2342 (N_2342,In_421,In_2716);
or U2343 (N_2343,In_3192,In_1489);
nand U2344 (N_2344,In_4995,In_502);
xnor U2345 (N_2345,In_563,In_3367);
nand U2346 (N_2346,In_4564,In_916);
nor U2347 (N_2347,In_1855,In_3651);
nor U2348 (N_2348,In_575,In_4173);
nor U2349 (N_2349,In_4276,In_1035);
nand U2350 (N_2350,In_3180,In_1180);
and U2351 (N_2351,In_1073,In_9);
or U2352 (N_2352,In_1446,In_3658);
or U2353 (N_2353,In_4275,In_4934);
nor U2354 (N_2354,In_2646,In_1573);
nand U2355 (N_2355,In_3485,In_1703);
nor U2356 (N_2356,In_416,In_1766);
nand U2357 (N_2357,In_1100,In_77);
nand U2358 (N_2358,In_4339,In_3653);
or U2359 (N_2359,In_2525,In_137);
nand U2360 (N_2360,In_4286,In_4752);
xor U2361 (N_2361,In_827,In_288);
nand U2362 (N_2362,In_2892,In_227);
nand U2363 (N_2363,In_3128,In_3377);
or U2364 (N_2364,In_713,In_2174);
nand U2365 (N_2365,In_2300,In_3891);
or U2366 (N_2366,In_1157,In_732);
xor U2367 (N_2367,In_1537,In_872);
or U2368 (N_2368,In_1524,In_384);
nor U2369 (N_2369,In_1348,In_789);
and U2370 (N_2370,In_3328,In_3195);
and U2371 (N_2371,In_2877,In_1448);
and U2372 (N_2372,In_2456,In_3316);
and U2373 (N_2373,In_2782,In_924);
or U2374 (N_2374,In_3937,In_4447);
and U2375 (N_2375,In_4114,In_1067);
nor U2376 (N_2376,In_442,In_4310);
or U2377 (N_2377,In_3129,In_4686);
and U2378 (N_2378,In_2473,In_796);
nor U2379 (N_2379,In_2063,In_306);
nor U2380 (N_2380,In_3562,In_1934);
xnor U2381 (N_2381,In_3655,In_790);
and U2382 (N_2382,In_2711,In_740);
or U2383 (N_2383,In_1853,In_3973);
or U2384 (N_2384,In_2649,In_4032);
and U2385 (N_2385,In_1951,In_4687);
nor U2386 (N_2386,In_4273,In_4135);
nor U2387 (N_2387,In_4098,In_2946);
and U2388 (N_2388,In_2517,In_974);
nand U2389 (N_2389,In_658,In_3716);
nand U2390 (N_2390,In_3544,In_3832);
or U2391 (N_2391,In_187,In_1312);
nor U2392 (N_2392,In_3332,In_1811);
and U2393 (N_2393,In_1639,In_4842);
nor U2394 (N_2394,In_2276,In_1792);
and U2395 (N_2395,In_1965,In_3883);
nor U2396 (N_2396,In_252,In_4160);
nand U2397 (N_2397,In_2605,In_2905);
and U2398 (N_2398,In_4791,In_937);
or U2399 (N_2399,In_4118,In_4731);
nand U2400 (N_2400,In_4511,In_2822);
and U2401 (N_2401,In_3995,In_4509);
nand U2402 (N_2402,In_4222,In_4635);
or U2403 (N_2403,In_2973,In_3808);
nor U2404 (N_2404,In_2362,In_4121);
and U2405 (N_2405,In_1042,In_1215);
nand U2406 (N_2406,In_124,In_3738);
and U2407 (N_2407,In_360,In_3375);
nand U2408 (N_2408,In_3740,In_1867);
and U2409 (N_2409,In_385,In_583);
or U2410 (N_2410,In_2752,In_4411);
and U2411 (N_2411,In_2542,In_2941);
and U2412 (N_2412,In_4883,In_4553);
xnor U2413 (N_2413,In_4456,In_2118);
nor U2414 (N_2414,In_2844,In_566);
or U2415 (N_2415,In_1032,In_1787);
or U2416 (N_2416,In_1363,In_4417);
and U2417 (N_2417,In_742,In_2795);
nor U2418 (N_2418,In_1103,In_4307);
nor U2419 (N_2419,In_133,In_2778);
and U2420 (N_2420,In_4381,In_405);
nor U2421 (N_2421,In_4530,In_3273);
or U2422 (N_2422,In_2500,In_1412);
and U2423 (N_2423,In_1019,In_1315);
xor U2424 (N_2424,In_2242,In_3642);
nand U2425 (N_2425,In_994,In_4571);
or U2426 (N_2426,In_2312,In_3943);
and U2427 (N_2427,In_3132,In_1165);
nor U2428 (N_2428,In_4246,In_2042);
nand U2429 (N_2429,In_4914,In_3949);
xor U2430 (N_2430,In_4016,In_4475);
and U2431 (N_2431,In_4480,In_1808);
and U2432 (N_2432,In_226,In_3133);
or U2433 (N_2433,In_4512,In_4562);
nand U2434 (N_2434,In_675,In_2003);
nand U2435 (N_2435,In_813,In_4559);
nand U2436 (N_2436,In_2308,In_2230);
nand U2437 (N_2437,In_453,In_2053);
nand U2438 (N_2438,In_508,In_3368);
nand U2439 (N_2439,In_1935,In_4846);
nor U2440 (N_2440,In_4338,In_167);
and U2441 (N_2441,In_2604,In_1646);
or U2442 (N_2442,In_2791,In_2035);
nand U2443 (N_2443,In_2962,In_433);
nor U2444 (N_2444,In_4088,In_1558);
or U2445 (N_2445,In_891,In_588);
or U2446 (N_2446,In_859,In_85);
or U2447 (N_2447,In_2924,In_3699);
or U2448 (N_2448,In_4388,In_3187);
xnor U2449 (N_2449,In_4002,In_4492);
and U2450 (N_2450,In_4322,In_3830);
and U2451 (N_2451,In_4320,In_3152);
xnor U2452 (N_2452,In_755,In_2869);
or U2453 (N_2453,In_2022,In_2293);
or U2454 (N_2454,In_4224,In_4637);
nand U2455 (N_2455,In_1259,In_3426);
nor U2456 (N_2456,In_3903,In_366);
and U2457 (N_2457,In_2156,In_523);
or U2458 (N_2458,In_4380,In_4632);
or U2459 (N_2459,In_2896,In_1877);
nand U2460 (N_2460,In_1108,In_768);
nor U2461 (N_2461,In_170,In_3666);
and U2462 (N_2462,In_982,In_2509);
nor U2463 (N_2463,In_3610,In_493);
or U2464 (N_2464,In_3789,In_3990);
and U2465 (N_2465,In_184,In_2380);
nand U2466 (N_2466,In_3693,In_2286);
nand U2467 (N_2467,In_2987,In_4419);
or U2468 (N_2468,In_2164,In_3774);
and U2469 (N_2469,In_655,In_1344);
nand U2470 (N_2470,In_3158,In_991);
and U2471 (N_2471,In_2357,In_1569);
or U2472 (N_2472,In_4464,In_4587);
nor U2473 (N_2473,In_4753,In_568);
nand U2474 (N_2474,In_1034,In_2425);
nor U2475 (N_2475,In_3764,In_3025);
nor U2476 (N_2476,In_4488,In_2297);
and U2477 (N_2477,In_1518,In_4347);
or U2478 (N_2478,In_4433,In_4213);
or U2479 (N_2479,In_1,In_2849);
nor U2480 (N_2480,In_4661,In_1804);
or U2481 (N_2481,In_2758,In_1119);
or U2482 (N_2482,In_743,In_720);
nand U2483 (N_2483,In_2988,In_4601);
nand U2484 (N_2484,In_4138,In_3359);
and U2485 (N_2485,In_2721,In_461);
nand U2486 (N_2486,In_4056,In_192);
nand U2487 (N_2487,In_2909,In_4084);
and U2488 (N_2488,In_3750,In_4593);
nor U2489 (N_2489,In_1336,In_3692);
or U2490 (N_2490,In_996,In_4145);
or U2491 (N_2491,In_2327,In_3449);
and U2492 (N_2492,In_2004,In_4852);
and U2493 (N_2493,In_1262,In_2754);
or U2494 (N_2494,In_3547,In_4157);
nand U2495 (N_2495,In_2082,In_2986);
or U2496 (N_2496,In_169,In_1600);
nor U2497 (N_2497,In_427,In_677);
nand U2498 (N_2498,In_4732,In_2296);
nand U2499 (N_2499,In_3417,In_4109);
nand U2500 (N_2500,In_132,In_4145);
nand U2501 (N_2501,In_1842,In_4921);
nor U2502 (N_2502,In_122,In_4019);
xor U2503 (N_2503,In_1371,In_4889);
nand U2504 (N_2504,In_1358,In_1492);
or U2505 (N_2505,In_4610,In_1601);
xnor U2506 (N_2506,In_2421,In_2423);
or U2507 (N_2507,In_766,In_3805);
and U2508 (N_2508,In_1152,In_288);
and U2509 (N_2509,In_4215,In_3068);
nor U2510 (N_2510,In_2757,In_1649);
nor U2511 (N_2511,In_2848,In_3957);
xnor U2512 (N_2512,In_859,In_3157);
nor U2513 (N_2513,In_2409,In_4448);
nor U2514 (N_2514,In_3322,In_4692);
and U2515 (N_2515,In_3865,In_3193);
nor U2516 (N_2516,In_3711,In_1199);
and U2517 (N_2517,In_1943,In_4174);
and U2518 (N_2518,In_2643,In_2677);
and U2519 (N_2519,In_3541,In_2040);
nor U2520 (N_2520,In_2769,In_2632);
nand U2521 (N_2521,In_1835,In_3240);
nor U2522 (N_2522,In_3830,In_4699);
and U2523 (N_2523,In_1987,In_1831);
and U2524 (N_2524,In_4832,In_4159);
nor U2525 (N_2525,In_1501,In_4077);
and U2526 (N_2526,In_4135,In_3227);
nor U2527 (N_2527,In_2673,In_3406);
and U2528 (N_2528,In_4812,In_3075);
nor U2529 (N_2529,In_1366,In_3697);
and U2530 (N_2530,In_2816,In_4005);
nor U2531 (N_2531,In_3451,In_2333);
or U2532 (N_2532,In_4875,In_1234);
and U2533 (N_2533,In_1622,In_4642);
xor U2534 (N_2534,In_2287,In_419);
nand U2535 (N_2535,In_4138,In_1264);
or U2536 (N_2536,In_203,In_1997);
and U2537 (N_2537,In_2742,In_1768);
nand U2538 (N_2538,In_1758,In_1389);
nand U2539 (N_2539,In_2991,In_2705);
nand U2540 (N_2540,In_1770,In_3362);
nor U2541 (N_2541,In_1477,In_2365);
and U2542 (N_2542,In_4322,In_630);
xor U2543 (N_2543,In_3236,In_2205);
and U2544 (N_2544,In_1894,In_3582);
or U2545 (N_2545,In_2410,In_448);
and U2546 (N_2546,In_4571,In_1428);
or U2547 (N_2547,In_941,In_1711);
nand U2548 (N_2548,In_672,In_4259);
and U2549 (N_2549,In_2687,In_4766);
xnor U2550 (N_2550,In_4776,In_658);
nand U2551 (N_2551,In_3187,In_2010);
and U2552 (N_2552,In_38,In_3271);
xnor U2553 (N_2553,In_988,In_1928);
or U2554 (N_2554,In_3959,In_1112);
nand U2555 (N_2555,In_4419,In_2329);
nor U2556 (N_2556,In_4304,In_3105);
nor U2557 (N_2557,In_2789,In_4376);
nor U2558 (N_2558,In_2120,In_1454);
nor U2559 (N_2559,In_1204,In_3834);
or U2560 (N_2560,In_4499,In_196);
nor U2561 (N_2561,In_3615,In_2357);
nor U2562 (N_2562,In_2998,In_2079);
nand U2563 (N_2563,In_2429,In_4084);
nand U2564 (N_2564,In_2315,In_3256);
and U2565 (N_2565,In_3950,In_4689);
and U2566 (N_2566,In_4211,In_422);
nand U2567 (N_2567,In_1421,In_2797);
and U2568 (N_2568,In_3205,In_1437);
nand U2569 (N_2569,In_2976,In_2009);
nor U2570 (N_2570,In_1278,In_2489);
and U2571 (N_2571,In_3612,In_11);
or U2572 (N_2572,In_468,In_544);
nand U2573 (N_2573,In_562,In_981);
nand U2574 (N_2574,In_4570,In_4852);
and U2575 (N_2575,In_3112,In_3298);
and U2576 (N_2576,In_1014,In_1542);
nand U2577 (N_2577,In_4695,In_326);
nand U2578 (N_2578,In_1484,In_1458);
nor U2579 (N_2579,In_1093,In_3779);
or U2580 (N_2580,In_2705,In_3474);
nand U2581 (N_2581,In_2211,In_1559);
and U2582 (N_2582,In_4097,In_3715);
nor U2583 (N_2583,In_1358,In_1035);
nand U2584 (N_2584,In_1363,In_4853);
xor U2585 (N_2585,In_4431,In_1334);
or U2586 (N_2586,In_652,In_3332);
nor U2587 (N_2587,In_2589,In_3367);
nand U2588 (N_2588,In_2526,In_841);
or U2589 (N_2589,In_3666,In_3755);
nor U2590 (N_2590,In_1714,In_3468);
nor U2591 (N_2591,In_4183,In_4385);
nor U2592 (N_2592,In_7,In_1984);
or U2593 (N_2593,In_1802,In_4473);
and U2594 (N_2594,In_4528,In_2418);
xor U2595 (N_2595,In_2176,In_497);
nor U2596 (N_2596,In_3872,In_1252);
and U2597 (N_2597,In_4329,In_4081);
and U2598 (N_2598,In_768,In_4780);
or U2599 (N_2599,In_1014,In_4429);
or U2600 (N_2600,In_2797,In_3958);
or U2601 (N_2601,In_870,In_1288);
nor U2602 (N_2602,In_4654,In_3618);
and U2603 (N_2603,In_2587,In_1027);
and U2604 (N_2604,In_2460,In_2948);
and U2605 (N_2605,In_2404,In_3417);
xnor U2606 (N_2606,In_1096,In_3660);
or U2607 (N_2607,In_2106,In_3155);
nor U2608 (N_2608,In_3632,In_295);
nor U2609 (N_2609,In_3092,In_2951);
or U2610 (N_2610,In_2408,In_2834);
or U2611 (N_2611,In_2091,In_342);
nand U2612 (N_2612,In_4040,In_2474);
nand U2613 (N_2613,In_402,In_1469);
xor U2614 (N_2614,In_695,In_2183);
or U2615 (N_2615,In_3802,In_4662);
nand U2616 (N_2616,In_268,In_1809);
nand U2617 (N_2617,In_2802,In_3420);
and U2618 (N_2618,In_2746,In_3111);
and U2619 (N_2619,In_2430,In_2992);
xnor U2620 (N_2620,In_1958,In_2797);
and U2621 (N_2621,In_773,In_1488);
and U2622 (N_2622,In_1746,In_891);
or U2623 (N_2623,In_907,In_977);
or U2624 (N_2624,In_505,In_4244);
or U2625 (N_2625,In_56,In_2310);
and U2626 (N_2626,In_3710,In_920);
or U2627 (N_2627,In_1935,In_2941);
or U2628 (N_2628,In_3386,In_2668);
and U2629 (N_2629,In_4397,In_2714);
or U2630 (N_2630,In_1591,In_4041);
or U2631 (N_2631,In_3476,In_974);
or U2632 (N_2632,In_3854,In_3688);
nor U2633 (N_2633,In_3346,In_158);
and U2634 (N_2634,In_4306,In_2752);
xnor U2635 (N_2635,In_2038,In_4924);
or U2636 (N_2636,In_1166,In_1661);
or U2637 (N_2637,In_3456,In_640);
and U2638 (N_2638,In_2266,In_1532);
or U2639 (N_2639,In_1235,In_479);
nand U2640 (N_2640,In_3037,In_3403);
xor U2641 (N_2641,In_2517,In_357);
nand U2642 (N_2642,In_2381,In_26);
and U2643 (N_2643,In_2263,In_2286);
or U2644 (N_2644,In_1982,In_140);
and U2645 (N_2645,In_1374,In_853);
nand U2646 (N_2646,In_4585,In_1014);
or U2647 (N_2647,In_2785,In_4468);
xnor U2648 (N_2648,In_3678,In_3947);
or U2649 (N_2649,In_1004,In_432);
xor U2650 (N_2650,In_3248,In_3102);
nor U2651 (N_2651,In_1064,In_2906);
or U2652 (N_2652,In_1211,In_1184);
nor U2653 (N_2653,In_2449,In_1585);
or U2654 (N_2654,In_991,In_599);
nor U2655 (N_2655,In_2090,In_3459);
or U2656 (N_2656,In_4923,In_2270);
or U2657 (N_2657,In_3792,In_230);
nand U2658 (N_2658,In_576,In_1121);
nand U2659 (N_2659,In_470,In_3992);
nand U2660 (N_2660,In_1510,In_2430);
and U2661 (N_2661,In_3337,In_3850);
nand U2662 (N_2662,In_3535,In_627);
and U2663 (N_2663,In_4944,In_3940);
xor U2664 (N_2664,In_873,In_4249);
nor U2665 (N_2665,In_4768,In_978);
nor U2666 (N_2666,In_4852,In_4079);
nor U2667 (N_2667,In_317,In_366);
nand U2668 (N_2668,In_1607,In_3158);
or U2669 (N_2669,In_1686,In_4533);
and U2670 (N_2670,In_1207,In_1873);
or U2671 (N_2671,In_4241,In_3250);
xor U2672 (N_2672,In_1289,In_1008);
and U2673 (N_2673,In_2889,In_3416);
nor U2674 (N_2674,In_1476,In_1240);
nor U2675 (N_2675,In_2791,In_1889);
or U2676 (N_2676,In_4363,In_4196);
or U2677 (N_2677,In_2007,In_1297);
nor U2678 (N_2678,In_2456,In_3138);
nor U2679 (N_2679,In_2617,In_765);
nor U2680 (N_2680,In_4117,In_4576);
nand U2681 (N_2681,In_1504,In_4196);
and U2682 (N_2682,In_3220,In_3630);
and U2683 (N_2683,In_2442,In_209);
and U2684 (N_2684,In_2403,In_1487);
nand U2685 (N_2685,In_1863,In_2759);
xor U2686 (N_2686,In_1235,In_2998);
or U2687 (N_2687,In_4522,In_3616);
nand U2688 (N_2688,In_1665,In_2731);
nand U2689 (N_2689,In_2473,In_3655);
or U2690 (N_2690,In_4341,In_3455);
nor U2691 (N_2691,In_4466,In_4514);
nor U2692 (N_2692,In_2025,In_4101);
nor U2693 (N_2693,In_2999,In_2305);
nor U2694 (N_2694,In_3743,In_3630);
or U2695 (N_2695,In_4593,In_1872);
and U2696 (N_2696,In_4403,In_2960);
nor U2697 (N_2697,In_3177,In_1773);
nand U2698 (N_2698,In_310,In_1637);
nand U2699 (N_2699,In_1158,In_2949);
nand U2700 (N_2700,In_1651,In_3231);
and U2701 (N_2701,In_3185,In_1391);
or U2702 (N_2702,In_2660,In_4650);
xnor U2703 (N_2703,In_3415,In_2911);
nand U2704 (N_2704,In_294,In_933);
nor U2705 (N_2705,In_1535,In_1812);
xor U2706 (N_2706,In_3363,In_3271);
xor U2707 (N_2707,In_3624,In_4587);
nor U2708 (N_2708,In_4153,In_1010);
nand U2709 (N_2709,In_4121,In_1672);
nand U2710 (N_2710,In_2733,In_3387);
xor U2711 (N_2711,In_3292,In_3171);
xor U2712 (N_2712,In_1986,In_3852);
nor U2713 (N_2713,In_1129,In_1833);
xnor U2714 (N_2714,In_3981,In_3818);
or U2715 (N_2715,In_1918,In_2443);
nand U2716 (N_2716,In_629,In_795);
nor U2717 (N_2717,In_4266,In_4077);
nand U2718 (N_2718,In_2801,In_1569);
nor U2719 (N_2719,In_856,In_3883);
nand U2720 (N_2720,In_4039,In_1998);
nor U2721 (N_2721,In_4605,In_2993);
nor U2722 (N_2722,In_1488,In_4044);
and U2723 (N_2723,In_4759,In_882);
or U2724 (N_2724,In_2080,In_3114);
and U2725 (N_2725,In_2084,In_756);
nor U2726 (N_2726,In_3098,In_819);
nor U2727 (N_2727,In_3374,In_3159);
or U2728 (N_2728,In_3237,In_107);
and U2729 (N_2729,In_2492,In_4390);
nand U2730 (N_2730,In_2155,In_1239);
nand U2731 (N_2731,In_3484,In_957);
and U2732 (N_2732,In_3437,In_1500);
nand U2733 (N_2733,In_1460,In_2445);
nand U2734 (N_2734,In_2040,In_785);
and U2735 (N_2735,In_3504,In_1853);
or U2736 (N_2736,In_3726,In_4427);
or U2737 (N_2737,In_578,In_1013);
xnor U2738 (N_2738,In_1821,In_4713);
and U2739 (N_2739,In_1540,In_4234);
or U2740 (N_2740,In_2661,In_3541);
or U2741 (N_2741,In_275,In_1008);
or U2742 (N_2742,In_468,In_4272);
xnor U2743 (N_2743,In_280,In_4537);
and U2744 (N_2744,In_3142,In_3394);
and U2745 (N_2745,In_183,In_2212);
nor U2746 (N_2746,In_3265,In_3891);
and U2747 (N_2747,In_3811,In_3184);
nand U2748 (N_2748,In_3574,In_1008);
or U2749 (N_2749,In_2384,In_4929);
nor U2750 (N_2750,In_758,In_1443);
xnor U2751 (N_2751,In_1273,In_4644);
nand U2752 (N_2752,In_2760,In_1603);
nand U2753 (N_2753,In_4476,In_2882);
xor U2754 (N_2754,In_2642,In_737);
or U2755 (N_2755,In_3168,In_1123);
nor U2756 (N_2756,In_4511,In_3215);
nand U2757 (N_2757,In_3982,In_4020);
nand U2758 (N_2758,In_2795,In_3363);
nand U2759 (N_2759,In_819,In_3110);
nor U2760 (N_2760,In_3791,In_277);
xor U2761 (N_2761,In_4148,In_2032);
and U2762 (N_2762,In_2849,In_2452);
or U2763 (N_2763,In_3387,In_121);
nand U2764 (N_2764,In_3139,In_3342);
nand U2765 (N_2765,In_2378,In_92);
xor U2766 (N_2766,In_2252,In_4024);
and U2767 (N_2767,In_4843,In_4942);
xor U2768 (N_2768,In_2625,In_1123);
or U2769 (N_2769,In_1613,In_4518);
nand U2770 (N_2770,In_2927,In_1648);
xnor U2771 (N_2771,In_850,In_1044);
and U2772 (N_2772,In_4558,In_2869);
or U2773 (N_2773,In_3480,In_2243);
or U2774 (N_2774,In_3823,In_2556);
xnor U2775 (N_2775,In_491,In_968);
nor U2776 (N_2776,In_2406,In_1556);
and U2777 (N_2777,In_2139,In_1834);
nor U2778 (N_2778,In_1646,In_1420);
nand U2779 (N_2779,In_712,In_1740);
or U2780 (N_2780,In_4541,In_284);
and U2781 (N_2781,In_696,In_496);
or U2782 (N_2782,In_3776,In_1289);
or U2783 (N_2783,In_3604,In_1336);
nor U2784 (N_2784,In_2754,In_3645);
nand U2785 (N_2785,In_3842,In_4258);
xor U2786 (N_2786,In_1153,In_1214);
and U2787 (N_2787,In_2032,In_2051);
nand U2788 (N_2788,In_4647,In_2155);
and U2789 (N_2789,In_1916,In_757);
or U2790 (N_2790,In_196,In_206);
nor U2791 (N_2791,In_1715,In_2019);
and U2792 (N_2792,In_721,In_3947);
nor U2793 (N_2793,In_1662,In_4128);
nand U2794 (N_2794,In_3100,In_2558);
nand U2795 (N_2795,In_1921,In_3486);
and U2796 (N_2796,In_4218,In_4824);
and U2797 (N_2797,In_1549,In_1438);
nand U2798 (N_2798,In_2438,In_3568);
nor U2799 (N_2799,In_4072,In_3031);
and U2800 (N_2800,In_2742,In_3833);
and U2801 (N_2801,In_1020,In_1650);
and U2802 (N_2802,In_4908,In_4617);
and U2803 (N_2803,In_3119,In_3445);
nor U2804 (N_2804,In_3561,In_2594);
or U2805 (N_2805,In_960,In_4689);
xnor U2806 (N_2806,In_3255,In_4485);
xnor U2807 (N_2807,In_1477,In_3392);
nor U2808 (N_2808,In_642,In_1508);
nand U2809 (N_2809,In_2680,In_4312);
and U2810 (N_2810,In_2282,In_698);
nand U2811 (N_2811,In_4326,In_629);
nor U2812 (N_2812,In_993,In_3841);
nor U2813 (N_2813,In_4014,In_2430);
nand U2814 (N_2814,In_1608,In_3369);
and U2815 (N_2815,In_516,In_2933);
nor U2816 (N_2816,In_3124,In_204);
or U2817 (N_2817,In_1383,In_321);
or U2818 (N_2818,In_1120,In_2402);
nor U2819 (N_2819,In_4912,In_2286);
and U2820 (N_2820,In_2770,In_3698);
nor U2821 (N_2821,In_2374,In_1125);
xor U2822 (N_2822,In_3757,In_2947);
or U2823 (N_2823,In_4932,In_1908);
xnor U2824 (N_2824,In_2468,In_711);
xor U2825 (N_2825,In_4748,In_2927);
nor U2826 (N_2826,In_3852,In_4337);
nand U2827 (N_2827,In_553,In_1746);
nand U2828 (N_2828,In_2947,In_3457);
or U2829 (N_2829,In_2731,In_3239);
xnor U2830 (N_2830,In_1289,In_1530);
and U2831 (N_2831,In_4113,In_4879);
nor U2832 (N_2832,In_2949,In_4350);
and U2833 (N_2833,In_189,In_1812);
or U2834 (N_2834,In_846,In_79);
and U2835 (N_2835,In_50,In_276);
nand U2836 (N_2836,In_556,In_3615);
or U2837 (N_2837,In_4893,In_2814);
or U2838 (N_2838,In_3010,In_3424);
and U2839 (N_2839,In_461,In_464);
nand U2840 (N_2840,In_4741,In_1967);
nor U2841 (N_2841,In_1951,In_1758);
or U2842 (N_2842,In_152,In_2514);
or U2843 (N_2843,In_366,In_3255);
nand U2844 (N_2844,In_3187,In_3563);
nor U2845 (N_2845,In_4563,In_498);
and U2846 (N_2846,In_2768,In_4698);
xnor U2847 (N_2847,In_3233,In_2467);
nand U2848 (N_2848,In_2882,In_2829);
nor U2849 (N_2849,In_97,In_4902);
or U2850 (N_2850,In_3492,In_1283);
and U2851 (N_2851,In_3285,In_3386);
xnor U2852 (N_2852,In_2546,In_4733);
nand U2853 (N_2853,In_3533,In_4241);
and U2854 (N_2854,In_2585,In_4660);
and U2855 (N_2855,In_3619,In_408);
or U2856 (N_2856,In_4219,In_2867);
or U2857 (N_2857,In_4204,In_3924);
nor U2858 (N_2858,In_4057,In_124);
nor U2859 (N_2859,In_4959,In_1696);
or U2860 (N_2860,In_28,In_3780);
nand U2861 (N_2861,In_2418,In_3158);
nor U2862 (N_2862,In_4767,In_3685);
or U2863 (N_2863,In_4162,In_4017);
or U2864 (N_2864,In_2974,In_244);
or U2865 (N_2865,In_4484,In_3039);
nand U2866 (N_2866,In_1689,In_1723);
nand U2867 (N_2867,In_4497,In_3437);
and U2868 (N_2868,In_868,In_4479);
and U2869 (N_2869,In_4417,In_366);
and U2870 (N_2870,In_3018,In_3348);
nand U2871 (N_2871,In_1740,In_1367);
xor U2872 (N_2872,In_3794,In_4979);
nand U2873 (N_2873,In_1498,In_4957);
or U2874 (N_2874,In_2276,In_1568);
nand U2875 (N_2875,In_1064,In_4006);
or U2876 (N_2876,In_4098,In_2827);
or U2877 (N_2877,In_213,In_3181);
nand U2878 (N_2878,In_16,In_848);
xor U2879 (N_2879,In_540,In_3795);
xor U2880 (N_2880,In_596,In_159);
and U2881 (N_2881,In_1728,In_2539);
nand U2882 (N_2882,In_2401,In_3746);
or U2883 (N_2883,In_796,In_4161);
and U2884 (N_2884,In_1971,In_1966);
nand U2885 (N_2885,In_4107,In_2606);
and U2886 (N_2886,In_1164,In_448);
nor U2887 (N_2887,In_3607,In_3466);
or U2888 (N_2888,In_4303,In_485);
nor U2889 (N_2889,In_3579,In_757);
nor U2890 (N_2890,In_263,In_2016);
nor U2891 (N_2891,In_1670,In_1510);
nor U2892 (N_2892,In_1581,In_4836);
nor U2893 (N_2893,In_132,In_726);
or U2894 (N_2894,In_966,In_4625);
nand U2895 (N_2895,In_3332,In_4791);
and U2896 (N_2896,In_3601,In_2600);
or U2897 (N_2897,In_258,In_3287);
nand U2898 (N_2898,In_2059,In_1826);
nand U2899 (N_2899,In_805,In_1045);
and U2900 (N_2900,In_2971,In_4514);
or U2901 (N_2901,In_3738,In_3431);
nand U2902 (N_2902,In_861,In_4649);
and U2903 (N_2903,In_2257,In_4402);
and U2904 (N_2904,In_1357,In_155);
and U2905 (N_2905,In_1305,In_3967);
or U2906 (N_2906,In_1666,In_2060);
nor U2907 (N_2907,In_4273,In_2837);
and U2908 (N_2908,In_2429,In_2879);
or U2909 (N_2909,In_1018,In_2939);
nand U2910 (N_2910,In_200,In_4055);
or U2911 (N_2911,In_39,In_459);
and U2912 (N_2912,In_2129,In_1234);
nor U2913 (N_2913,In_3642,In_4652);
or U2914 (N_2914,In_1755,In_1843);
nor U2915 (N_2915,In_1035,In_2916);
nand U2916 (N_2916,In_3204,In_1135);
nor U2917 (N_2917,In_4890,In_172);
and U2918 (N_2918,In_2026,In_333);
nor U2919 (N_2919,In_836,In_4280);
nor U2920 (N_2920,In_3007,In_3159);
nor U2921 (N_2921,In_4720,In_4234);
or U2922 (N_2922,In_1245,In_1397);
and U2923 (N_2923,In_2819,In_1100);
and U2924 (N_2924,In_1460,In_168);
nand U2925 (N_2925,In_3968,In_1301);
nor U2926 (N_2926,In_3214,In_4486);
nand U2927 (N_2927,In_3579,In_195);
nor U2928 (N_2928,In_1251,In_2431);
and U2929 (N_2929,In_4637,In_504);
or U2930 (N_2930,In_2104,In_4327);
and U2931 (N_2931,In_1339,In_3052);
and U2932 (N_2932,In_2550,In_3774);
or U2933 (N_2933,In_310,In_3343);
and U2934 (N_2934,In_3860,In_4876);
nor U2935 (N_2935,In_4009,In_4538);
or U2936 (N_2936,In_405,In_3867);
or U2937 (N_2937,In_2617,In_3894);
and U2938 (N_2938,In_621,In_1951);
nor U2939 (N_2939,In_1855,In_927);
nand U2940 (N_2940,In_1222,In_4838);
and U2941 (N_2941,In_3813,In_1629);
or U2942 (N_2942,In_2637,In_2939);
nor U2943 (N_2943,In_3017,In_2840);
and U2944 (N_2944,In_946,In_3553);
nor U2945 (N_2945,In_2605,In_1228);
nor U2946 (N_2946,In_467,In_2254);
and U2947 (N_2947,In_2721,In_4420);
and U2948 (N_2948,In_2835,In_1786);
nor U2949 (N_2949,In_1353,In_2458);
and U2950 (N_2950,In_1859,In_4122);
nor U2951 (N_2951,In_1640,In_3583);
nand U2952 (N_2952,In_598,In_1956);
and U2953 (N_2953,In_934,In_1356);
and U2954 (N_2954,In_2173,In_3940);
and U2955 (N_2955,In_3886,In_4680);
nor U2956 (N_2956,In_2678,In_4587);
nand U2957 (N_2957,In_4445,In_3497);
or U2958 (N_2958,In_3482,In_2550);
and U2959 (N_2959,In_1732,In_3225);
xnor U2960 (N_2960,In_3200,In_1689);
and U2961 (N_2961,In_3302,In_1917);
nand U2962 (N_2962,In_2440,In_3751);
or U2963 (N_2963,In_4270,In_3173);
nor U2964 (N_2964,In_1650,In_1987);
and U2965 (N_2965,In_891,In_1855);
and U2966 (N_2966,In_2582,In_3768);
nor U2967 (N_2967,In_2108,In_804);
and U2968 (N_2968,In_4627,In_281);
or U2969 (N_2969,In_4124,In_2882);
nor U2970 (N_2970,In_4192,In_4034);
xor U2971 (N_2971,In_4597,In_4833);
nor U2972 (N_2972,In_809,In_4077);
or U2973 (N_2973,In_4198,In_3259);
nor U2974 (N_2974,In_4292,In_2324);
or U2975 (N_2975,In_4998,In_3826);
and U2976 (N_2976,In_2860,In_4699);
or U2977 (N_2977,In_4874,In_225);
nand U2978 (N_2978,In_2848,In_2853);
nand U2979 (N_2979,In_841,In_2032);
nor U2980 (N_2980,In_3126,In_3526);
nor U2981 (N_2981,In_1530,In_3575);
nor U2982 (N_2982,In_3791,In_4395);
nand U2983 (N_2983,In_2134,In_766);
and U2984 (N_2984,In_3906,In_57);
and U2985 (N_2985,In_1265,In_1694);
or U2986 (N_2986,In_137,In_1892);
nand U2987 (N_2987,In_4070,In_2806);
and U2988 (N_2988,In_2602,In_2468);
xnor U2989 (N_2989,In_3303,In_202);
or U2990 (N_2990,In_2490,In_282);
or U2991 (N_2991,In_1832,In_4125);
or U2992 (N_2992,In_2101,In_712);
or U2993 (N_2993,In_3128,In_4327);
nand U2994 (N_2994,In_2980,In_794);
nor U2995 (N_2995,In_432,In_2321);
xnor U2996 (N_2996,In_3511,In_1962);
or U2997 (N_2997,In_1238,In_3581);
nand U2998 (N_2998,In_44,In_4796);
or U2999 (N_2999,In_4832,In_4765);
or U3000 (N_3000,In_1512,In_4689);
nand U3001 (N_3001,In_56,In_4070);
nor U3002 (N_3002,In_3275,In_1638);
nor U3003 (N_3003,In_2995,In_2030);
nand U3004 (N_3004,In_4059,In_2532);
or U3005 (N_3005,In_3566,In_39);
and U3006 (N_3006,In_418,In_4210);
xnor U3007 (N_3007,In_1531,In_1950);
nor U3008 (N_3008,In_1735,In_4864);
nand U3009 (N_3009,In_4959,In_3726);
nor U3010 (N_3010,In_2424,In_3457);
nand U3011 (N_3011,In_1277,In_3172);
xor U3012 (N_3012,In_660,In_4319);
nand U3013 (N_3013,In_827,In_1179);
or U3014 (N_3014,In_1480,In_2337);
or U3015 (N_3015,In_2823,In_3117);
xnor U3016 (N_3016,In_4196,In_2814);
or U3017 (N_3017,In_2256,In_278);
nor U3018 (N_3018,In_2532,In_3707);
or U3019 (N_3019,In_800,In_3098);
nor U3020 (N_3020,In_4223,In_646);
and U3021 (N_3021,In_2695,In_4058);
nor U3022 (N_3022,In_3114,In_1701);
and U3023 (N_3023,In_1460,In_2075);
nor U3024 (N_3024,In_2771,In_4275);
or U3025 (N_3025,In_964,In_2892);
xnor U3026 (N_3026,In_3073,In_3645);
and U3027 (N_3027,In_4306,In_3647);
nand U3028 (N_3028,In_3203,In_1392);
nor U3029 (N_3029,In_2788,In_4499);
nand U3030 (N_3030,In_1063,In_955);
or U3031 (N_3031,In_4672,In_4627);
xor U3032 (N_3032,In_2826,In_4245);
nor U3033 (N_3033,In_2953,In_2702);
nor U3034 (N_3034,In_862,In_2255);
nand U3035 (N_3035,In_196,In_3671);
nor U3036 (N_3036,In_3679,In_3612);
nor U3037 (N_3037,In_1433,In_4193);
and U3038 (N_3038,In_3283,In_2467);
xnor U3039 (N_3039,In_2826,In_870);
and U3040 (N_3040,In_857,In_3139);
xnor U3041 (N_3041,In_2503,In_3612);
and U3042 (N_3042,In_567,In_808);
nor U3043 (N_3043,In_457,In_4093);
or U3044 (N_3044,In_1513,In_3792);
nor U3045 (N_3045,In_4015,In_1842);
nor U3046 (N_3046,In_4766,In_2266);
nor U3047 (N_3047,In_2224,In_2211);
xnor U3048 (N_3048,In_1579,In_2463);
or U3049 (N_3049,In_2272,In_1649);
or U3050 (N_3050,In_2715,In_3259);
and U3051 (N_3051,In_3256,In_511);
and U3052 (N_3052,In_3817,In_3925);
nand U3053 (N_3053,In_1713,In_2191);
and U3054 (N_3054,In_1090,In_1039);
nor U3055 (N_3055,In_2383,In_4900);
and U3056 (N_3056,In_742,In_2247);
nor U3057 (N_3057,In_4263,In_4439);
nor U3058 (N_3058,In_51,In_4439);
and U3059 (N_3059,In_4227,In_2611);
nand U3060 (N_3060,In_2901,In_3108);
nor U3061 (N_3061,In_4056,In_106);
nand U3062 (N_3062,In_4214,In_243);
or U3063 (N_3063,In_1631,In_3407);
nor U3064 (N_3064,In_775,In_3501);
nor U3065 (N_3065,In_3280,In_2909);
or U3066 (N_3066,In_328,In_3345);
or U3067 (N_3067,In_3358,In_2505);
nand U3068 (N_3068,In_3772,In_2595);
and U3069 (N_3069,In_2478,In_4890);
or U3070 (N_3070,In_2820,In_3458);
nand U3071 (N_3071,In_1932,In_346);
or U3072 (N_3072,In_1396,In_3605);
nor U3073 (N_3073,In_3109,In_3859);
nor U3074 (N_3074,In_420,In_2668);
nand U3075 (N_3075,In_873,In_3497);
or U3076 (N_3076,In_3885,In_457);
xnor U3077 (N_3077,In_1299,In_3829);
nor U3078 (N_3078,In_3692,In_1225);
or U3079 (N_3079,In_25,In_2122);
xor U3080 (N_3080,In_2242,In_395);
nor U3081 (N_3081,In_3811,In_776);
and U3082 (N_3082,In_3222,In_939);
and U3083 (N_3083,In_1160,In_3559);
or U3084 (N_3084,In_3261,In_3901);
nor U3085 (N_3085,In_3270,In_2739);
and U3086 (N_3086,In_4748,In_4195);
or U3087 (N_3087,In_448,In_3755);
or U3088 (N_3088,In_438,In_3605);
nand U3089 (N_3089,In_2929,In_1066);
or U3090 (N_3090,In_4209,In_333);
nor U3091 (N_3091,In_2497,In_4703);
or U3092 (N_3092,In_2136,In_2486);
and U3093 (N_3093,In_4581,In_453);
nand U3094 (N_3094,In_4897,In_2775);
and U3095 (N_3095,In_419,In_4224);
nor U3096 (N_3096,In_1649,In_143);
and U3097 (N_3097,In_4280,In_3973);
xor U3098 (N_3098,In_899,In_24);
nand U3099 (N_3099,In_2626,In_2655);
xor U3100 (N_3100,In_756,In_4789);
nor U3101 (N_3101,In_3848,In_505);
or U3102 (N_3102,In_4290,In_323);
and U3103 (N_3103,In_3183,In_2184);
or U3104 (N_3104,In_1204,In_1103);
and U3105 (N_3105,In_368,In_3112);
or U3106 (N_3106,In_4733,In_2011);
nand U3107 (N_3107,In_4117,In_1058);
xnor U3108 (N_3108,In_1321,In_4367);
and U3109 (N_3109,In_4544,In_2668);
nand U3110 (N_3110,In_4857,In_4846);
nand U3111 (N_3111,In_99,In_416);
or U3112 (N_3112,In_3443,In_4853);
and U3113 (N_3113,In_2156,In_2210);
or U3114 (N_3114,In_1862,In_4204);
xnor U3115 (N_3115,In_1811,In_514);
nand U3116 (N_3116,In_4589,In_3198);
or U3117 (N_3117,In_1685,In_2955);
and U3118 (N_3118,In_3776,In_1928);
xnor U3119 (N_3119,In_2678,In_397);
nor U3120 (N_3120,In_4236,In_1047);
xnor U3121 (N_3121,In_3852,In_2272);
or U3122 (N_3122,In_2784,In_632);
nor U3123 (N_3123,In_594,In_830);
or U3124 (N_3124,In_1789,In_634);
and U3125 (N_3125,In_2144,In_3651);
or U3126 (N_3126,In_3412,In_346);
nor U3127 (N_3127,In_443,In_706);
nor U3128 (N_3128,In_1796,In_2647);
nand U3129 (N_3129,In_3708,In_1975);
nand U3130 (N_3130,In_3981,In_1964);
nor U3131 (N_3131,In_3576,In_1968);
nand U3132 (N_3132,In_3284,In_4440);
and U3133 (N_3133,In_1553,In_2680);
or U3134 (N_3134,In_1571,In_1226);
xnor U3135 (N_3135,In_4140,In_4111);
nand U3136 (N_3136,In_3114,In_1458);
and U3137 (N_3137,In_1353,In_2910);
or U3138 (N_3138,In_1700,In_2012);
and U3139 (N_3139,In_2383,In_4315);
or U3140 (N_3140,In_2477,In_1069);
nor U3141 (N_3141,In_1733,In_4065);
and U3142 (N_3142,In_344,In_3919);
or U3143 (N_3143,In_361,In_1598);
and U3144 (N_3144,In_1445,In_3257);
nand U3145 (N_3145,In_2907,In_4325);
or U3146 (N_3146,In_4544,In_3249);
and U3147 (N_3147,In_2076,In_2182);
and U3148 (N_3148,In_3686,In_771);
or U3149 (N_3149,In_4643,In_1482);
nand U3150 (N_3150,In_3384,In_1218);
xor U3151 (N_3151,In_4101,In_3626);
xor U3152 (N_3152,In_906,In_134);
or U3153 (N_3153,In_1040,In_3310);
nor U3154 (N_3154,In_3842,In_182);
nor U3155 (N_3155,In_2359,In_4129);
and U3156 (N_3156,In_2028,In_578);
nand U3157 (N_3157,In_2538,In_4313);
nand U3158 (N_3158,In_4213,In_3362);
xor U3159 (N_3159,In_150,In_1964);
nor U3160 (N_3160,In_1561,In_2687);
nor U3161 (N_3161,In_1955,In_1235);
nor U3162 (N_3162,In_876,In_4050);
nand U3163 (N_3163,In_2885,In_1671);
nand U3164 (N_3164,In_2021,In_1361);
nand U3165 (N_3165,In_831,In_2132);
xnor U3166 (N_3166,In_4760,In_319);
nor U3167 (N_3167,In_1055,In_4213);
nor U3168 (N_3168,In_780,In_382);
nand U3169 (N_3169,In_690,In_4853);
or U3170 (N_3170,In_126,In_4653);
and U3171 (N_3171,In_3705,In_529);
or U3172 (N_3172,In_17,In_3251);
nor U3173 (N_3173,In_3065,In_3128);
nor U3174 (N_3174,In_2849,In_1311);
nor U3175 (N_3175,In_4665,In_1534);
nor U3176 (N_3176,In_3102,In_450);
nand U3177 (N_3177,In_792,In_653);
nand U3178 (N_3178,In_943,In_737);
and U3179 (N_3179,In_1456,In_3107);
nor U3180 (N_3180,In_2910,In_82);
nand U3181 (N_3181,In_3928,In_4862);
or U3182 (N_3182,In_3628,In_4433);
nor U3183 (N_3183,In_3950,In_3535);
and U3184 (N_3184,In_4385,In_4994);
xor U3185 (N_3185,In_231,In_4342);
and U3186 (N_3186,In_2695,In_2626);
and U3187 (N_3187,In_1903,In_395);
nand U3188 (N_3188,In_2442,In_2832);
and U3189 (N_3189,In_4409,In_4988);
nand U3190 (N_3190,In_2020,In_4192);
and U3191 (N_3191,In_3640,In_478);
and U3192 (N_3192,In_3290,In_3809);
or U3193 (N_3193,In_1036,In_2670);
and U3194 (N_3194,In_4001,In_1996);
nand U3195 (N_3195,In_2143,In_401);
nor U3196 (N_3196,In_1129,In_1585);
or U3197 (N_3197,In_150,In_4301);
nand U3198 (N_3198,In_2708,In_877);
and U3199 (N_3199,In_1321,In_3837);
or U3200 (N_3200,In_832,In_1350);
nand U3201 (N_3201,In_4176,In_1630);
or U3202 (N_3202,In_4849,In_2169);
xor U3203 (N_3203,In_1099,In_4742);
nor U3204 (N_3204,In_4904,In_3918);
nand U3205 (N_3205,In_375,In_989);
or U3206 (N_3206,In_3450,In_2247);
nand U3207 (N_3207,In_381,In_3156);
nor U3208 (N_3208,In_4267,In_1524);
nor U3209 (N_3209,In_4994,In_1559);
nand U3210 (N_3210,In_4505,In_2202);
nor U3211 (N_3211,In_2740,In_3106);
nor U3212 (N_3212,In_3411,In_1672);
and U3213 (N_3213,In_1464,In_4318);
xor U3214 (N_3214,In_3088,In_4078);
nor U3215 (N_3215,In_3242,In_2764);
xor U3216 (N_3216,In_2343,In_2991);
nand U3217 (N_3217,In_1258,In_3338);
xor U3218 (N_3218,In_2520,In_3044);
nand U3219 (N_3219,In_3327,In_4834);
nand U3220 (N_3220,In_1431,In_694);
nor U3221 (N_3221,In_1404,In_1849);
or U3222 (N_3222,In_2751,In_3827);
or U3223 (N_3223,In_4549,In_11);
nor U3224 (N_3224,In_1463,In_681);
nor U3225 (N_3225,In_3207,In_2299);
nor U3226 (N_3226,In_201,In_2096);
and U3227 (N_3227,In_4187,In_3280);
xnor U3228 (N_3228,In_2661,In_4379);
nand U3229 (N_3229,In_223,In_258);
nor U3230 (N_3230,In_4697,In_210);
nand U3231 (N_3231,In_2659,In_1521);
nor U3232 (N_3232,In_834,In_1951);
nor U3233 (N_3233,In_4521,In_3852);
nor U3234 (N_3234,In_4816,In_4601);
and U3235 (N_3235,In_1038,In_4511);
nand U3236 (N_3236,In_4701,In_1340);
nor U3237 (N_3237,In_2216,In_2255);
nand U3238 (N_3238,In_1083,In_4464);
nand U3239 (N_3239,In_390,In_875);
xor U3240 (N_3240,In_4351,In_1435);
nand U3241 (N_3241,In_2661,In_3510);
nand U3242 (N_3242,In_2851,In_395);
nand U3243 (N_3243,In_2227,In_2762);
and U3244 (N_3244,In_685,In_4869);
or U3245 (N_3245,In_3243,In_2485);
nand U3246 (N_3246,In_4256,In_3780);
and U3247 (N_3247,In_4931,In_259);
nor U3248 (N_3248,In_2698,In_3065);
and U3249 (N_3249,In_2400,In_745);
nand U3250 (N_3250,In_188,In_1801);
and U3251 (N_3251,In_3607,In_3043);
and U3252 (N_3252,In_2160,In_3461);
nand U3253 (N_3253,In_3936,In_2739);
and U3254 (N_3254,In_4188,In_1426);
xor U3255 (N_3255,In_1379,In_254);
nand U3256 (N_3256,In_2605,In_236);
or U3257 (N_3257,In_688,In_819);
and U3258 (N_3258,In_4360,In_3521);
nor U3259 (N_3259,In_4277,In_2904);
and U3260 (N_3260,In_476,In_253);
nand U3261 (N_3261,In_4369,In_3576);
and U3262 (N_3262,In_1221,In_137);
nand U3263 (N_3263,In_2699,In_254);
nand U3264 (N_3264,In_1813,In_1878);
nor U3265 (N_3265,In_3918,In_3523);
xor U3266 (N_3266,In_342,In_3154);
nand U3267 (N_3267,In_3676,In_2816);
nand U3268 (N_3268,In_52,In_1489);
xnor U3269 (N_3269,In_1421,In_2276);
and U3270 (N_3270,In_2997,In_4868);
and U3271 (N_3271,In_3968,In_3551);
nor U3272 (N_3272,In_1560,In_3791);
and U3273 (N_3273,In_3501,In_326);
nand U3274 (N_3274,In_4192,In_3283);
and U3275 (N_3275,In_4814,In_513);
nor U3276 (N_3276,In_717,In_1328);
nand U3277 (N_3277,In_4675,In_45);
and U3278 (N_3278,In_4846,In_593);
xor U3279 (N_3279,In_3646,In_1600);
or U3280 (N_3280,In_3434,In_494);
nor U3281 (N_3281,In_3062,In_69);
nor U3282 (N_3282,In_4578,In_1523);
and U3283 (N_3283,In_338,In_3481);
nand U3284 (N_3284,In_2660,In_3504);
nand U3285 (N_3285,In_650,In_1670);
nor U3286 (N_3286,In_1963,In_3266);
xor U3287 (N_3287,In_2572,In_4369);
and U3288 (N_3288,In_4093,In_4936);
or U3289 (N_3289,In_340,In_4042);
nor U3290 (N_3290,In_4576,In_3234);
nand U3291 (N_3291,In_4037,In_2703);
nor U3292 (N_3292,In_2495,In_2743);
and U3293 (N_3293,In_3394,In_3882);
and U3294 (N_3294,In_2667,In_9);
and U3295 (N_3295,In_603,In_2301);
and U3296 (N_3296,In_1116,In_3508);
nor U3297 (N_3297,In_3140,In_3363);
and U3298 (N_3298,In_1713,In_3666);
and U3299 (N_3299,In_1198,In_4933);
nand U3300 (N_3300,In_3351,In_4134);
nand U3301 (N_3301,In_4448,In_1806);
and U3302 (N_3302,In_4488,In_3329);
nand U3303 (N_3303,In_3770,In_1678);
and U3304 (N_3304,In_1017,In_4318);
nor U3305 (N_3305,In_2262,In_4919);
xor U3306 (N_3306,In_2737,In_3849);
nor U3307 (N_3307,In_4702,In_3508);
nand U3308 (N_3308,In_213,In_1778);
and U3309 (N_3309,In_2422,In_3809);
and U3310 (N_3310,In_992,In_92);
or U3311 (N_3311,In_4771,In_3016);
and U3312 (N_3312,In_1774,In_760);
xor U3313 (N_3313,In_867,In_3969);
nor U3314 (N_3314,In_2915,In_1487);
and U3315 (N_3315,In_616,In_481);
and U3316 (N_3316,In_4924,In_4729);
nor U3317 (N_3317,In_167,In_589);
xor U3318 (N_3318,In_1108,In_1654);
or U3319 (N_3319,In_2695,In_4356);
nand U3320 (N_3320,In_3414,In_3081);
or U3321 (N_3321,In_4780,In_3403);
xor U3322 (N_3322,In_1171,In_4097);
and U3323 (N_3323,In_1872,In_1311);
and U3324 (N_3324,In_1255,In_1138);
or U3325 (N_3325,In_2755,In_3702);
or U3326 (N_3326,In_4774,In_1294);
nand U3327 (N_3327,In_4306,In_1650);
nand U3328 (N_3328,In_3490,In_1252);
and U3329 (N_3329,In_4057,In_2260);
and U3330 (N_3330,In_1323,In_3519);
nor U3331 (N_3331,In_495,In_1715);
nor U3332 (N_3332,In_1847,In_816);
nand U3333 (N_3333,In_1033,In_4053);
xnor U3334 (N_3334,In_2992,In_374);
nor U3335 (N_3335,In_2049,In_4484);
nand U3336 (N_3336,In_1664,In_184);
and U3337 (N_3337,In_3580,In_740);
xor U3338 (N_3338,In_4895,In_4333);
and U3339 (N_3339,In_4787,In_337);
and U3340 (N_3340,In_4633,In_2731);
xnor U3341 (N_3341,In_3143,In_3821);
and U3342 (N_3342,In_1962,In_1499);
or U3343 (N_3343,In_1055,In_4257);
nor U3344 (N_3344,In_2916,In_343);
xor U3345 (N_3345,In_1138,In_1925);
nor U3346 (N_3346,In_2053,In_97);
nor U3347 (N_3347,In_1921,In_2425);
or U3348 (N_3348,In_3874,In_2864);
xor U3349 (N_3349,In_4688,In_3245);
and U3350 (N_3350,In_3070,In_4410);
xor U3351 (N_3351,In_2641,In_4407);
nor U3352 (N_3352,In_3657,In_4992);
nand U3353 (N_3353,In_4860,In_1204);
or U3354 (N_3354,In_2380,In_2944);
nand U3355 (N_3355,In_1361,In_4914);
nand U3356 (N_3356,In_3174,In_2576);
nand U3357 (N_3357,In_4183,In_4808);
nor U3358 (N_3358,In_1503,In_2184);
nor U3359 (N_3359,In_2922,In_570);
or U3360 (N_3360,In_983,In_3688);
or U3361 (N_3361,In_3313,In_3926);
or U3362 (N_3362,In_1745,In_3307);
or U3363 (N_3363,In_1008,In_1276);
and U3364 (N_3364,In_2581,In_4860);
or U3365 (N_3365,In_3379,In_4574);
nor U3366 (N_3366,In_2569,In_357);
or U3367 (N_3367,In_4881,In_263);
nand U3368 (N_3368,In_2526,In_3857);
nor U3369 (N_3369,In_71,In_1730);
and U3370 (N_3370,In_4701,In_1004);
nor U3371 (N_3371,In_536,In_3685);
nand U3372 (N_3372,In_1169,In_471);
and U3373 (N_3373,In_3275,In_4108);
nor U3374 (N_3374,In_2592,In_290);
nor U3375 (N_3375,In_2216,In_1114);
or U3376 (N_3376,In_1668,In_3461);
nand U3377 (N_3377,In_478,In_3358);
nor U3378 (N_3378,In_4561,In_2992);
xnor U3379 (N_3379,In_2011,In_3174);
nor U3380 (N_3380,In_1328,In_2999);
nor U3381 (N_3381,In_3899,In_3438);
or U3382 (N_3382,In_1218,In_1515);
nand U3383 (N_3383,In_819,In_2423);
nand U3384 (N_3384,In_2184,In_3490);
nor U3385 (N_3385,In_4776,In_2177);
or U3386 (N_3386,In_3986,In_870);
nor U3387 (N_3387,In_1456,In_3393);
and U3388 (N_3388,In_2804,In_3323);
nand U3389 (N_3389,In_1680,In_3285);
or U3390 (N_3390,In_4770,In_286);
xnor U3391 (N_3391,In_969,In_4446);
nand U3392 (N_3392,In_3056,In_4094);
xor U3393 (N_3393,In_2664,In_2705);
nor U3394 (N_3394,In_1000,In_587);
nor U3395 (N_3395,In_1877,In_2673);
xnor U3396 (N_3396,In_2618,In_384);
nor U3397 (N_3397,In_425,In_1448);
nor U3398 (N_3398,In_3527,In_1168);
nand U3399 (N_3399,In_2303,In_1374);
nor U3400 (N_3400,In_2438,In_3511);
or U3401 (N_3401,In_3510,In_4353);
or U3402 (N_3402,In_3243,In_2047);
or U3403 (N_3403,In_314,In_4906);
nor U3404 (N_3404,In_2799,In_3861);
nand U3405 (N_3405,In_2160,In_4783);
or U3406 (N_3406,In_4687,In_1872);
xnor U3407 (N_3407,In_4693,In_2788);
and U3408 (N_3408,In_803,In_2621);
or U3409 (N_3409,In_2269,In_3188);
and U3410 (N_3410,In_2747,In_1508);
nand U3411 (N_3411,In_2447,In_1777);
xnor U3412 (N_3412,In_4002,In_36);
nand U3413 (N_3413,In_418,In_4369);
and U3414 (N_3414,In_1181,In_1288);
xor U3415 (N_3415,In_1168,In_4641);
nand U3416 (N_3416,In_930,In_862);
and U3417 (N_3417,In_328,In_4180);
nand U3418 (N_3418,In_1743,In_244);
nand U3419 (N_3419,In_721,In_3215);
xnor U3420 (N_3420,In_496,In_4876);
nor U3421 (N_3421,In_2317,In_247);
and U3422 (N_3422,In_4862,In_1236);
xnor U3423 (N_3423,In_1803,In_1355);
or U3424 (N_3424,In_1993,In_4563);
xnor U3425 (N_3425,In_4200,In_3114);
and U3426 (N_3426,In_2212,In_2447);
nand U3427 (N_3427,In_4751,In_3310);
nor U3428 (N_3428,In_1672,In_2312);
or U3429 (N_3429,In_1712,In_1345);
nand U3430 (N_3430,In_3953,In_430);
nand U3431 (N_3431,In_2607,In_3720);
and U3432 (N_3432,In_93,In_351);
or U3433 (N_3433,In_4804,In_4281);
nand U3434 (N_3434,In_2641,In_3011);
or U3435 (N_3435,In_1594,In_3210);
nand U3436 (N_3436,In_1061,In_1525);
nor U3437 (N_3437,In_2543,In_3404);
nand U3438 (N_3438,In_2605,In_1604);
or U3439 (N_3439,In_4640,In_2850);
nor U3440 (N_3440,In_2825,In_4105);
nand U3441 (N_3441,In_4866,In_1383);
or U3442 (N_3442,In_2364,In_3988);
nor U3443 (N_3443,In_2532,In_4236);
and U3444 (N_3444,In_838,In_4771);
nand U3445 (N_3445,In_687,In_2302);
nand U3446 (N_3446,In_3999,In_2246);
or U3447 (N_3447,In_4043,In_3147);
nor U3448 (N_3448,In_2747,In_3827);
nor U3449 (N_3449,In_1165,In_416);
nand U3450 (N_3450,In_1755,In_3584);
or U3451 (N_3451,In_1040,In_4409);
nand U3452 (N_3452,In_1476,In_1892);
and U3453 (N_3453,In_3610,In_588);
nand U3454 (N_3454,In_2574,In_2925);
and U3455 (N_3455,In_1103,In_2003);
and U3456 (N_3456,In_4151,In_4300);
or U3457 (N_3457,In_2176,In_2625);
and U3458 (N_3458,In_4493,In_4962);
nor U3459 (N_3459,In_340,In_4884);
or U3460 (N_3460,In_1006,In_3882);
and U3461 (N_3461,In_54,In_3432);
nor U3462 (N_3462,In_1477,In_147);
nand U3463 (N_3463,In_4188,In_2704);
nor U3464 (N_3464,In_443,In_2223);
or U3465 (N_3465,In_3248,In_4223);
or U3466 (N_3466,In_2322,In_1090);
or U3467 (N_3467,In_4336,In_2322);
or U3468 (N_3468,In_1884,In_458);
or U3469 (N_3469,In_3580,In_660);
and U3470 (N_3470,In_4990,In_4758);
xor U3471 (N_3471,In_2493,In_4296);
xnor U3472 (N_3472,In_261,In_2690);
or U3473 (N_3473,In_4871,In_2757);
and U3474 (N_3474,In_3700,In_1765);
and U3475 (N_3475,In_453,In_1151);
and U3476 (N_3476,In_2354,In_2993);
and U3477 (N_3477,In_2330,In_1162);
nor U3478 (N_3478,In_4586,In_1653);
xnor U3479 (N_3479,In_277,In_3505);
and U3480 (N_3480,In_1356,In_1754);
or U3481 (N_3481,In_2090,In_1495);
and U3482 (N_3482,In_4711,In_4523);
and U3483 (N_3483,In_4611,In_927);
xnor U3484 (N_3484,In_2316,In_3159);
nor U3485 (N_3485,In_1057,In_3225);
xor U3486 (N_3486,In_4118,In_2450);
nand U3487 (N_3487,In_3802,In_3671);
xnor U3488 (N_3488,In_2119,In_2350);
nand U3489 (N_3489,In_2447,In_3117);
nand U3490 (N_3490,In_4683,In_1995);
nand U3491 (N_3491,In_3065,In_4176);
nand U3492 (N_3492,In_4705,In_3935);
nand U3493 (N_3493,In_2294,In_3325);
nor U3494 (N_3494,In_10,In_4561);
and U3495 (N_3495,In_4293,In_2692);
or U3496 (N_3496,In_1785,In_2327);
and U3497 (N_3497,In_1869,In_577);
or U3498 (N_3498,In_2363,In_3941);
and U3499 (N_3499,In_4622,In_1317);
nor U3500 (N_3500,In_1052,In_3827);
xor U3501 (N_3501,In_370,In_4229);
xor U3502 (N_3502,In_3016,In_3974);
nand U3503 (N_3503,In_3110,In_3768);
xnor U3504 (N_3504,In_2758,In_3042);
or U3505 (N_3505,In_3930,In_2466);
nor U3506 (N_3506,In_1922,In_4429);
or U3507 (N_3507,In_1073,In_1485);
xnor U3508 (N_3508,In_461,In_4537);
or U3509 (N_3509,In_2317,In_2193);
nand U3510 (N_3510,In_4496,In_320);
nor U3511 (N_3511,In_3793,In_1831);
or U3512 (N_3512,In_2793,In_2622);
and U3513 (N_3513,In_385,In_705);
xor U3514 (N_3514,In_1884,In_4557);
nand U3515 (N_3515,In_563,In_1293);
nor U3516 (N_3516,In_3150,In_1081);
or U3517 (N_3517,In_600,In_2013);
nand U3518 (N_3518,In_657,In_2764);
nor U3519 (N_3519,In_1374,In_691);
xor U3520 (N_3520,In_746,In_382);
nor U3521 (N_3521,In_4105,In_4199);
nor U3522 (N_3522,In_1651,In_717);
nor U3523 (N_3523,In_2045,In_411);
or U3524 (N_3524,In_285,In_1174);
or U3525 (N_3525,In_877,In_2713);
nor U3526 (N_3526,In_1916,In_2919);
and U3527 (N_3527,In_3125,In_3558);
or U3528 (N_3528,In_913,In_263);
nor U3529 (N_3529,In_309,In_4023);
and U3530 (N_3530,In_942,In_678);
or U3531 (N_3531,In_4078,In_4966);
nor U3532 (N_3532,In_3434,In_2056);
nand U3533 (N_3533,In_1504,In_1739);
nor U3534 (N_3534,In_862,In_4466);
nand U3535 (N_3535,In_3519,In_1395);
or U3536 (N_3536,In_2314,In_4135);
and U3537 (N_3537,In_3419,In_2129);
and U3538 (N_3538,In_3186,In_3558);
nand U3539 (N_3539,In_159,In_1738);
nor U3540 (N_3540,In_3028,In_1688);
or U3541 (N_3541,In_4467,In_3486);
or U3542 (N_3542,In_1311,In_698);
nand U3543 (N_3543,In_727,In_1528);
nor U3544 (N_3544,In_1553,In_4241);
nand U3545 (N_3545,In_976,In_2795);
nor U3546 (N_3546,In_3353,In_2520);
and U3547 (N_3547,In_1121,In_2146);
or U3548 (N_3548,In_531,In_2031);
or U3549 (N_3549,In_4017,In_1492);
or U3550 (N_3550,In_2146,In_1516);
or U3551 (N_3551,In_2556,In_4079);
nor U3552 (N_3552,In_4099,In_4274);
and U3553 (N_3553,In_4652,In_473);
nor U3554 (N_3554,In_91,In_4853);
xor U3555 (N_3555,In_2955,In_2739);
nor U3556 (N_3556,In_4585,In_3328);
and U3557 (N_3557,In_4072,In_4006);
nor U3558 (N_3558,In_1607,In_2345);
xnor U3559 (N_3559,In_4099,In_2722);
xor U3560 (N_3560,In_2360,In_4337);
and U3561 (N_3561,In_3728,In_4751);
nand U3562 (N_3562,In_3568,In_145);
and U3563 (N_3563,In_340,In_3083);
xnor U3564 (N_3564,In_3138,In_3123);
nor U3565 (N_3565,In_962,In_2167);
and U3566 (N_3566,In_1147,In_2637);
or U3567 (N_3567,In_374,In_37);
nor U3568 (N_3568,In_4293,In_2905);
or U3569 (N_3569,In_3649,In_1554);
and U3570 (N_3570,In_4609,In_3174);
nor U3571 (N_3571,In_4807,In_4500);
or U3572 (N_3572,In_1517,In_2369);
nor U3573 (N_3573,In_586,In_2788);
and U3574 (N_3574,In_770,In_861);
nand U3575 (N_3575,In_1242,In_1811);
or U3576 (N_3576,In_2476,In_4941);
nor U3577 (N_3577,In_3335,In_3603);
and U3578 (N_3578,In_3070,In_4653);
nor U3579 (N_3579,In_4172,In_4037);
nor U3580 (N_3580,In_1601,In_4508);
nor U3581 (N_3581,In_1099,In_3207);
nand U3582 (N_3582,In_4228,In_4790);
nor U3583 (N_3583,In_2712,In_1305);
nor U3584 (N_3584,In_2864,In_829);
nand U3585 (N_3585,In_2620,In_3181);
or U3586 (N_3586,In_1188,In_3199);
and U3587 (N_3587,In_2790,In_3057);
nand U3588 (N_3588,In_2971,In_4941);
nor U3589 (N_3589,In_1852,In_2189);
and U3590 (N_3590,In_1879,In_1288);
nand U3591 (N_3591,In_2604,In_1379);
and U3592 (N_3592,In_3911,In_1077);
or U3593 (N_3593,In_2163,In_4536);
nor U3594 (N_3594,In_357,In_380);
or U3595 (N_3595,In_4125,In_4530);
nor U3596 (N_3596,In_669,In_4226);
xnor U3597 (N_3597,In_2585,In_496);
or U3598 (N_3598,In_2718,In_3024);
or U3599 (N_3599,In_3602,In_3010);
xor U3600 (N_3600,In_3980,In_1836);
and U3601 (N_3601,In_46,In_4629);
nand U3602 (N_3602,In_3752,In_1221);
and U3603 (N_3603,In_430,In_705);
and U3604 (N_3604,In_3958,In_3729);
or U3605 (N_3605,In_3652,In_789);
or U3606 (N_3606,In_4080,In_3234);
or U3607 (N_3607,In_1163,In_4528);
and U3608 (N_3608,In_643,In_2481);
xor U3609 (N_3609,In_3416,In_466);
and U3610 (N_3610,In_2655,In_3819);
or U3611 (N_3611,In_2756,In_814);
and U3612 (N_3612,In_3789,In_2438);
nand U3613 (N_3613,In_3104,In_2116);
nor U3614 (N_3614,In_50,In_3566);
nand U3615 (N_3615,In_754,In_3547);
and U3616 (N_3616,In_3710,In_4314);
nor U3617 (N_3617,In_894,In_705);
xor U3618 (N_3618,In_2385,In_3623);
nor U3619 (N_3619,In_3322,In_2178);
and U3620 (N_3620,In_1922,In_2114);
xnor U3621 (N_3621,In_3976,In_4555);
or U3622 (N_3622,In_4033,In_3035);
and U3623 (N_3623,In_4879,In_1785);
and U3624 (N_3624,In_4064,In_2806);
xor U3625 (N_3625,In_995,In_4542);
or U3626 (N_3626,In_3526,In_4908);
xnor U3627 (N_3627,In_2156,In_525);
or U3628 (N_3628,In_2715,In_1631);
or U3629 (N_3629,In_2041,In_4943);
nand U3630 (N_3630,In_535,In_3328);
or U3631 (N_3631,In_3369,In_1116);
or U3632 (N_3632,In_4274,In_4724);
nand U3633 (N_3633,In_249,In_4284);
or U3634 (N_3634,In_651,In_3288);
nand U3635 (N_3635,In_1304,In_743);
or U3636 (N_3636,In_4576,In_2992);
xor U3637 (N_3637,In_3736,In_2136);
nand U3638 (N_3638,In_4727,In_1855);
and U3639 (N_3639,In_935,In_3108);
nand U3640 (N_3640,In_2323,In_3445);
and U3641 (N_3641,In_406,In_2872);
nand U3642 (N_3642,In_1818,In_3462);
or U3643 (N_3643,In_3580,In_1860);
nor U3644 (N_3644,In_3378,In_689);
nand U3645 (N_3645,In_3602,In_733);
and U3646 (N_3646,In_711,In_2753);
nand U3647 (N_3647,In_3824,In_2511);
nor U3648 (N_3648,In_4563,In_3750);
or U3649 (N_3649,In_3374,In_2604);
nand U3650 (N_3650,In_1898,In_3989);
or U3651 (N_3651,In_64,In_4925);
and U3652 (N_3652,In_2658,In_4177);
nor U3653 (N_3653,In_204,In_2316);
or U3654 (N_3654,In_3890,In_4374);
nand U3655 (N_3655,In_3427,In_4303);
and U3656 (N_3656,In_1349,In_3425);
and U3657 (N_3657,In_3148,In_1702);
or U3658 (N_3658,In_201,In_1417);
and U3659 (N_3659,In_619,In_1483);
nand U3660 (N_3660,In_2834,In_1906);
nand U3661 (N_3661,In_1860,In_4295);
nand U3662 (N_3662,In_2982,In_4152);
and U3663 (N_3663,In_4406,In_1609);
nand U3664 (N_3664,In_2739,In_1058);
nand U3665 (N_3665,In_2650,In_1898);
nand U3666 (N_3666,In_898,In_2372);
nand U3667 (N_3667,In_1276,In_4312);
or U3668 (N_3668,In_4131,In_1866);
nor U3669 (N_3669,In_3075,In_4605);
or U3670 (N_3670,In_2305,In_2973);
or U3671 (N_3671,In_669,In_3416);
nand U3672 (N_3672,In_2575,In_3444);
nor U3673 (N_3673,In_1254,In_415);
nand U3674 (N_3674,In_122,In_1188);
xor U3675 (N_3675,In_3125,In_4592);
nand U3676 (N_3676,In_3434,In_4406);
or U3677 (N_3677,In_4883,In_1799);
nor U3678 (N_3678,In_1436,In_528);
nor U3679 (N_3679,In_1911,In_4182);
nand U3680 (N_3680,In_3189,In_4267);
nand U3681 (N_3681,In_4116,In_954);
or U3682 (N_3682,In_4451,In_2955);
and U3683 (N_3683,In_534,In_3910);
nor U3684 (N_3684,In_2200,In_4676);
xnor U3685 (N_3685,In_3414,In_4330);
and U3686 (N_3686,In_4804,In_2195);
nand U3687 (N_3687,In_3709,In_3029);
or U3688 (N_3688,In_4314,In_4025);
or U3689 (N_3689,In_1316,In_100);
nor U3690 (N_3690,In_2063,In_502);
or U3691 (N_3691,In_817,In_2175);
and U3692 (N_3692,In_3643,In_4138);
nor U3693 (N_3693,In_4053,In_661);
and U3694 (N_3694,In_4464,In_2292);
and U3695 (N_3695,In_1847,In_4648);
nor U3696 (N_3696,In_3903,In_934);
nand U3697 (N_3697,In_2797,In_2293);
nand U3698 (N_3698,In_1363,In_1693);
or U3699 (N_3699,In_428,In_4705);
nand U3700 (N_3700,In_4221,In_4207);
or U3701 (N_3701,In_2450,In_604);
nor U3702 (N_3702,In_4727,In_3108);
nand U3703 (N_3703,In_2123,In_3631);
nor U3704 (N_3704,In_4248,In_1620);
nor U3705 (N_3705,In_3510,In_4708);
and U3706 (N_3706,In_567,In_4659);
and U3707 (N_3707,In_137,In_4497);
nor U3708 (N_3708,In_1010,In_2555);
or U3709 (N_3709,In_746,In_948);
or U3710 (N_3710,In_192,In_3794);
nor U3711 (N_3711,In_3732,In_1653);
nand U3712 (N_3712,In_4270,In_249);
nor U3713 (N_3713,In_3512,In_1691);
xor U3714 (N_3714,In_4819,In_2837);
xnor U3715 (N_3715,In_1813,In_4358);
nor U3716 (N_3716,In_3483,In_1739);
nand U3717 (N_3717,In_2248,In_3532);
and U3718 (N_3718,In_2490,In_3445);
and U3719 (N_3719,In_245,In_240);
nand U3720 (N_3720,In_3490,In_736);
or U3721 (N_3721,In_931,In_1408);
and U3722 (N_3722,In_673,In_4507);
or U3723 (N_3723,In_3178,In_2744);
nor U3724 (N_3724,In_1278,In_1374);
nand U3725 (N_3725,In_782,In_1344);
or U3726 (N_3726,In_4972,In_3359);
and U3727 (N_3727,In_424,In_3626);
or U3728 (N_3728,In_4486,In_3525);
and U3729 (N_3729,In_1699,In_2883);
nor U3730 (N_3730,In_1475,In_1687);
and U3731 (N_3731,In_607,In_4103);
or U3732 (N_3732,In_3816,In_3958);
xor U3733 (N_3733,In_3631,In_3679);
nand U3734 (N_3734,In_978,In_263);
nand U3735 (N_3735,In_4164,In_3941);
or U3736 (N_3736,In_4085,In_4278);
nor U3737 (N_3737,In_3674,In_2571);
or U3738 (N_3738,In_4501,In_2903);
and U3739 (N_3739,In_3912,In_4809);
xor U3740 (N_3740,In_3570,In_511);
and U3741 (N_3741,In_156,In_2681);
nor U3742 (N_3742,In_694,In_520);
nand U3743 (N_3743,In_4366,In_1051);
nand U3744 (N_3744,In_1657,In_1994);
nor U3745 (N_3745,In_3303,In_4973);
and U3746 (N_3746,In_4204,In_4208);
nor U3747 (N_3747,In_1293,In_1574);
nand U3748 (N_3748,In_42,In_2571);
and U3749 (N_3749,In_2673,In_1035);
and U3750 (N_3750,In_63,In_3719);
xor U3751 (N_3751,In_808,In_3589);
nor U3752 (N_3752,In_1842,In_2242);
or U3753 (N_3753,In_2643,In_3218);
nor U3754 (N_3754,In_2425,In_2212);
and U3755 (N_3755,In_4430,In_3773);
nand U3756 (N_3756,In_3427,In_1494);
nor U3757 (N_3757,In_2188,In_2677);
nor U3758 (N_3758,In_2579,In_65);
nand U3759 (N_3759,In_621,In_2380);
and U3760 (N_3760,In_2585,In_3458);
nand U3761 (N_3761,In_1463,In_394);
or U3762 (N_3762,In_1892,In_1646);
xnor U3763 (N_3763,In_1997,In_3554);
or U3764 (N_3764,In_2294,In_1316);
nor U3765 (N_3765,In_3116,In_2606);
or U3766 (N_3766,In_885,In_1611);
nor U3767 (N_3767,In_2210,In_401);
or U3768 (N_3768,In_160,In_4613);
nor U3769 (N_3769,In_2660,In_1415);
or U3770 (N_3770,In_4814,In_4890);
xnor U3771 (N_3771,In_436,In_2339);
nand U3772 (N_3772,In_2082,In_4517);
and U3773 (N_3773,In_2656,In_1285);
or U3774 (N_3774,In_4623,In_1565);
nand U3775 (N_3775,In_3518,In_4933);
nor U3776 (N_3776,In_196,In_954);
xnor U3777 (N_3777,In_3947,In_424);
nor U3778 (N_3778,In_1905,In_2070);
or U3779 (N_3779,In_4334,In_722);
nor U3780 (N_3780,In_4347,In_4660);
or U3781 (N_3781,In_2713,In_1983);
nor U3782 (N_3782,In_2704,In_3869);
or U3783 (N_3783,In_4670,In_3533);
nor U3784 (N_3784,In_3375,In_3446);
and U3785 (N_3785,In_4663,In_1496);
nand U3786 (N_3786,In_4046,In_3861);
nand U3787 (N_3787,In_205,In_2775);
xor U3788 (N_3788,In_4109,In_3997);
and U3789 (N_3789,In_2140,In_2383);
nor U3790 (N_3790,In_905,In_4573);
or U3791 (N_3791,In_1589,In_4579);
and U3792 (N_3792,In_2068,In_335);
nor U3793 (N_3793,In_3083,In_3362);
nor U3794 (N_3794,In_1807,In_4520);
nand U3795 (N_3795,In_1284,In_710);
and U3796 (N_3796,In_1965,In_2486);
and U3797 (N_3797,In_178,In_2890);
or U3798 (N_3798,In_4553,In_3557);
nand U3799 (N_3799,In_1378,In_2208);
and U3800 (N_3800,In_2328,In_2921);
nor U3801 (N_3801,In_3017,In_1666);
nor U3802 (N_3802,In_4203,In_950);
and U3803 (N_3803,In_4130,In_1585);
nor U3804 (N_3804,In_4584,In_1064);
nor U3805 (N_3805,In_3604,In_3961);
or U3806 (N_3806,In_260,In_941);
nor U3807 (N_3807,In_2223,In_197);
nand U3808 (N_3808,In_4546,In_4286);
and U3809 (N_3809,In_2836,In_2474);
nor U3810 (N_3810,In_4614,In_911);
xor U3811 (N_3811,In_2027,In_776);
and U3812 (N_3812,In_2455,In_3786);
nand U3813 (N_3813,In_435,In_1206);
nand U3814 (N_3814,In_93,In_2053);
nand U3815 (N_3815,In_1346,In_2665);
or U3816 (N_3816,In_220,In_4809);
or U3817 (N_3817,In_3460,In_2012);
and U3818 (N_3818,In_635,In_3704);
nand U3819 (N_3819,In_3200,In_39);
nand U3820 (N_3820,In_293,In_2141);
nor U3821 (N_3821,In_4296,In_2273);
or U3822 (N_3822,In_124,In_4647);
xnor U3823 (N_3823,In_1143,In_2045);
nand U3824 (N_3824,In_2103,In_752);
nand U3825 (N_3825,In_2646,In_2450);
and U3826 (N_3826,In_465,In_852);
and U3827 (N_3827,In_275,In_2592);
and U3828 (N_3828,In_1557,In_1016);
and U3829 (N_3829,In_2534,In_3964);
nor U3830 (N_3830,In_3522,In_3364);
and U3831 (N_3831,In_3500,In_560);
nand U3832 (N_3832,In_190,In_2859);
xor U3833 (N_3833,In_25,In_1418);
or U3834 (N_3834,In_4538,In_1344);
and U3835 (N_3835,In_1352,In_1905);
nor U3836 (N_3836,In_1400,In_3274);
nor U3837 (N_3837,In_465,In_3029);
nand U3838 (N_3838,In_3214,In_4061);
nor U3839 (N_3839,In_597,In_3275);
and U3840 (N_3840,In_4448,In_2826);
xnor U3841 (N_3841,In_477,In_1564);
nor U3842 (N_3842,In_3288,In_4492);
nor U3843 (N_3843,In_3544,In_516);
nor U3844 (N_3844,In_3919,In_3794);
nor U3845 (N_3845,In_4181,In_990);
nand U3846 (N_3846,In_2086,In_209);
or U3847 (N_3847,In_2882,In_4754);
nand U3848 (N_3848,In_2154,In_611);
and U3849 (N_3849,In_4165,In_1204);
xnor U3850 (N_3850,In_1669,In_3492);
nand U3851 (N_3851,In_1916,In_1266);
nand U3852 (N_3852,In_4736,In_3491);
nor U3853 (N_3853,In_205,In_3766);
or U3854 (N_3854,In_718,In_2636);
nand U3855 (N_3855,In_2371,In_715);
nand U3856 (N_3856,In_1376,In_1314);
or U3857 (N_3857,In_4770,In_4054);
nor U3858 (N_3858,In_4444,In_698);
or U3859 (N_3859,In_4672,In_4781);
or U3860 (N_3860,In_1377,In_36);
nor U3861 (N_3861,In_4611,In_1078);
or U3862 (N_3862,In_2239,In_358);
nor U3863 (N_3863,In_4398,In_590);
and U3864 (N_3864,In_904,In_3912);
or U3865 (N_3865,In_2067,In_720);
and U3866 (N_3866,In_4533,In_4038);
or U3867 (N_3867,In_3235,In_2807);
nand U3868 (N_3868,In_3870,In_567);
xor U3869 (N_3869,In_1846,In_4422);
nand U3870 (N_3870,In_916,In_2054);
nor U3871 (N_3871,In_2997,In_1490);
or U3872 (N_3872,In_4403,In_3945);
nor U3873 (N_3873,In_4369,In_842);
and U3874 (N_3874,In_4583,In_2149);
or U3875 (N_3875,In_183,In_1612);
xor U3876 (N_3876,In_1244,In_1344);
xnor U3877 (N_3877,In_3663,In_475);
or U3878 (N_3878,In_2265,In_1036);
nor U3879 (N_3879,In_995,In_172);
and U3880 (N_3880,In_247,In_3672);
nand U3881 (N_3881,In_2270,In_3660);
xnor U3882 (N_3882,In_1564,In_750);
or U3883 (N_3883,In_648,In_731);
and U3884 (N_3884,In_2839,In_3616);
and U3885 (N_3885,In_1008,In_2134);
nand U3886 (N_3886,In_1501,In_1255);
nand U3887 (N_3887,In_4345,In_629);
xor U3888 (N_3888,In_4004,In_3158);
nor U3889 (N_3889,In_4772,In_847);
nand U3890 (N_3890,In_3488,In_2542);
or U3891 (N_3891,In_4373,In_1345);
nor U3892 (N_3892,In_3351,In_4294);
nor U3893 (N_3893,In_3162,In_957);
or U3894 (N_3894,In_2158,In_362);
xnor U3895 (N_3895,In_816,In_4889);
or U3896 (N_3896,In_1705,In_289);
nor U3897 (N_3897,In_3088,In_3096);
nor U3898 (N_3898,In_1481,In_2754);
nand U3899 (N_3899,In_4360,In_2791);
nor U3900 (N_3900,In_3887,In_3766);
nand U3901 (N_3901,In_855,In_971);
nand U3902 (N_3902,In_2238,In_3274);
nand U3903 (N_3903,In_3662,In_2038);
xnor U3904 (N_3904,In_2372,In_2727);
nand U3905 (N_3905,In_2437,In_2506);
nand U3906 (N_3906,In_1259,In_1594);
and U3907 (N_3907,In_703,In_2021);
nand U3908 (N_3908,In_4931,In_2458);
xor U3909 (N_3909,In_2390,In_518);
and U3910 (N_3910,In_3605,In_3724);
nand U3911 (N_3911,In_4857,In_2438);
nand U3912 (N_3912,In_4340,In_104);
xnor U3913 (N_3913,In_4035,In_2958);
nand U3914 (N_3914,In_1006,In_2295);
and U3915 (N_3915,In_638,In_2310);
nor U3916 (N_3916,In_4665,In_549);
or U3917 (N_3917,In_3611,In_1502);
or U3918 (N_3918,In_1722,In_4834);
nand U3919 (N_3919,In_2747,In_808);
nor U3920 (N_3920,In_4695,In_216);
nand U3921 (N_3921,In_1379,In_882);
and U3922 (N_3922,In_2463,In_2526);
or U3923 (N_3923,In_3830,In_226);
nor U3924 (N_3924,In_705,In_3144);
nand U3925 (N_3925,In_2189,In_2062);
and U3926 (N_3926,In_2675,In_2904);
and U3927 (N_3927,In_1680,In_4942);
and U3928 (N_3928,In_3422,In_4117);
nor U3929 (N_3929,In_1241,In_784);
nor U3930 (N_3930,In_1269,In_1996);
nand U3931 (N_3931,In_4668,In_4009);
or U3932 (N_3932,In_2292,In_4140);
and U3933 (N_3933,In_3940,In_2747);
nand U3934 (N_3934,In_508,In_3109);
or U3935 (N_3935,In_3826,In_1470);
or U3936 (N_3936,In_4294,In_2033);
xnor U3937 (N_3937,In_4161,In_825);
nor U3938 (N_3938,In_593,In_1222);
nor U3939 (N_3939,In_4814,In_451);
xnor U3940 (N_3940,In_23,In_3736);
nand U3941 (N_3941,In_4519,In_465);
nand U3942 (N_3942,In_380,In_2759);
nand U3943 (N_3943,In_166,In_3866);
nor U3944 (N_3944,In_14,In_4317);
nand U3945 (N_3945,In_580,In_4101);
nor U3946 (N_3946,In_4794,In_786);
or U3947 (N_3947,In_2495,In_2841);
nand U3948 (N_3948,In_20,In_2375);
or U3949 (N_3949,In_4512,In_2087);
or U3950 (N_3950,In_98,In_1303);
and U3951 (N_3951,In_410,In_897);
xnor U3952 (N_3952,In_4005,In_3959);
or U3953 (N_3953,In_564,In_4247);
and U3954 (N_3954,In_3639,In_4524);
nor U3955 (N_3955,In_1271,In_828);
or U3956 (N_3956,In_3172,In_1699);
nand U3957 (N_3957,In_1560,In_3767);
nand U3958 (N_3958,In_4348,In_803);
nand U3959 (N_3959,In_559,In_259);
nand U3960 (N_3960,In_1095,In_3225);
nor U3961 (N_3961,In_440,In_2715);
nand U3962 (N_3962,In_2932,In_4715);
nor U3963 (N_3963,In_2503,In_4914);
or U3964 (N_3964,In_1984,In_1055);
or U3965 (N_3965,In_7,In_3624);
nor U3966 (N_3966,In_333,In_3132);
nor U3967 (N_3967,In_2631,In_935);
nor U3968 (N_3968,In_768,In_2384);
and U3969 (N_3969,In_1468,In_1816);
nor U3970 (N_3970,In_892,In_151);
or U3971 (N_3971,In_684,In_3703);
and U3972 (N_3972,In_1683,In_4725);
and U3973 (N_3973,In_2227,In_1065);
or U3974 (N_3974,In_1118,In_520);
nand U3975 (N_3975,In_1153,In_3749);
nor U3976 (N_3976,In_531,In_240);
or U3977 (N_3977,In_4270,In_3507);
nand U3978 (N_3978,In_4048,In_696);
and U3979 (N_3979,In_3493,In_3754);
nand U3980 (N_3980,In_2852,In_1119);
nor U3981 (N_3981,In_1670,In_4439);
and U3982 (N_3982,In_3703,In_3422);
and U3983 (N_3983,In_4765,In_862);
or U3984 (N_3984,In_65,In_843);
or U3985 (N_3985,In_1722,In_3027);
xor U3986 (N_3986,In_121,In_2703);
xor U3987 (N_3987,In_4871,In_2065);
nor U3988 (N_3988,In_2910,In_4182);
or U3989 (N_3989,In_4025,In_740);
and U3990 (N_3990,In_596,In_4941);
or U3991 (N_3991,In_2500,In_2746);
nor U3992 (N_3992,In_1452,In_904);
and U3993 (N_3993,In_310,In_4107);
nand U3994 (N_3994,In_2060,In_2385);
and U3995 (N_3995,In_3817,In_1370);
nor U3996 (N_3996,In_4684,In_4901);
and U3997 (N_3997,In_4746,In_3209);
and U3998 (N_3998,In_731,In_3465);
nand U3999 (N_3999,In_3008,In_2536);
nand U4000 (N_4000,In_4369,In_478);
or U4001 (N_4001,In_3418,In_2896);
and U4002 (N_4002,In_274,In_4385);
nand U4003 (N_4003,In_1974,In_4943);
or U4004 (N_4004,In_2624,In_4476);
and U4005 (N_4005,In_168,In_1618);
nor U4006 (N_4006,In_2212,In_701);
and U4007 (N_4007,In_303,In_3074);
or U4008 (N_4008,In_1037,In_4287);
nand U4009 (N_4009,In_2080,In_3094);
nand U4010 (N_4010,In_4255,In_4413);
nand U4011 (N_4011,In_485,In_2423);
or U4012 (N_4012,In_460,In_360);
and U4013 (N_4013,In_1844,In_3136);
nor U4014 (N_4014,In_2075,In_4063);
xor U4015 (N_4015,In_4899,In_2953);
and U4016 (N_4016,In_3934,In_4281);
or U4017 (N_4017,In_3568,In_336);
or U4018 (N_4018,In_3572,In_4118);
nand U4019 (N_4019,In_602,In_3010);
or U4020 (N_4020,In_4829,In_4556);
and U4021 (N_4021,In_3157,In_3434);
nand U4022 (N_4022,In_3145,In_4989);
nor U4023 (N_4023,In_3449,In_1039);
or U4024 (N_4024,In_2397,In_3994);
and U4025 (N_4025,In_1114,In_2259);
nand U4026 (N_4026,In_3885,In_3253);
nand U4027 (N_4027,In_95,In_1379);
and U4028 (N_4028,In_1759,In_1074);
or U4029 (N_4029,In_1764,In_591);
nor U4030 (N_4030,In_4567,In_1162);
xnor U4031 (N_4031,In_4587,In_4687);
and U4032 (N_4032,In_620,In_4273);
or U4033 (N_4033,In_3793,In_2658);
and U4034 (N_4034,In_3825,In_4136);
or U4035 (N_4035,In_317,In_4470);
or U4036 (N_4036,In_1921,In_2652);
nand U4037 (N_4037,In_3931,In_3139);
nor U4038 (N_4038,In_4462,In_3862);
and U4039 (N_4039,In_2077,In_4712);
nand U4040 (N_4040,In_2791,In_690);
nand U4041 (N_4041,In_4001,In_579);
or U4042 (N_4042,In_3287,In_2146);
and U4043 (N_4043,In_1251,In_580);
or U4044 (N_4044,In_1871,In_2012);
nor U4045 (N_4045,In_1482,In_4846);
nand U4046 (N_4046,In_3139,In_1977);
nand U4047 (N_4047,In_4737,In_2961);
nand U4048 (N_4048,In_2598,In_1119);
nor U4049 (N_4049,In_2775,In_571);
or U4050 (N_4050,In_854,In_4456);
xor U4051 (N_4051,In_931,In_1927);
and U4052 (N_4052,In_268,In_3085);
or U4053 (N_4053,In_2493,In_4980);
and U4054 (N_4054,In_1087,In_2432);
and U4055 (N_4055,In_339,In_1357);
nor U4056 (N_4056,In_1837,In_712);
nor U4057 (N_4057,In_4173,In_3260);
and U4058 (N_4058,In_1300,In_3619);
nor U4059 (N_4059,In_82,In_1272);
nor U4060 (N_4060,In_4254,In_4675);
and U4061 (N_4061,In_281,In_3442);
nand U4062 (N_4062,In_1509,In_4805);
nor U4063 (N_4063,In_1087,In_160);
or U4064 (N_4064,In_321,In_11);
xnor U4065 (N_4065,In_331,In_2440);
or U4066 (N_4066,In_1561,In_4491);
nor U4067 (N_4067,In_3882,In_1130);
and U4068 (N_4068,In_3551,In_4137);
or U4069 (N_4069,In_4372,In_4353);
or U4070 (N_4070,In_217,In_1097);
and U4071 (N_4071,In_1752,In_4722);
or U4072 (N_4072,In_2734,In_2016);
nor U4073 (N_4073,In_2876,In_1063);
nand U4074 (N_4074,In_1798,In_4100);
xnor U4075 (N_4075,In_4884,In_4729);
nor U4076 (N_4076,In_4368,In_2302);
or U4077 (N_4077,In_3945,In_2640);
xor U4078 (N_4078,In_4684,In_1698);
nand U4079 (N_4079,In_2176,In_2152);
and U4080 (N_4080,In_3443,In_949);
nor U4081 (N_4081,In_212,In_3189);
nor U4082 (N_4082,In_1968,In_278);
nor U4083 (N_4083,In_1658,In_475);
nor U4084 (N_4084,In_4221,In_2142);
and U4085 (N_4085,In_18,In_2136);
and U4086 (N_4086,In_3854,In_468);
xor U4087 (N_4087,In_4870,In_3185);
and U4088 (N_4088,In_3237,In_3965);
and U4089 (N_4089,In_2994,In_4953);
nor U4090 (N_4090,In_4044,In_3234);
nand U4091 (N_4091,In_428,In_4220);
or U4092 (N_4092,In_2532,In_2458);
nor U4093 (N_4093,In_4092,In_825);
xnor U4094 (N_4094,In_585,In_4662);
or U4095 (N_4095,In_830,In_2648);
xor U4096 (N_4096,In_3633,In_3127);
nor U4097 (N_4097,In_2642,In_3400);
nor U4098 (N_4098,In_1046,In_4727);
nor U4099 (N_4099,In_1661,In_4221);
nand U4100 (N_4100,In_1886,In_724);
nor U4101 (N_4101,In_4233,In_2635);
or U4102 (N_4102,In_3486,In_2012);
nand U4103 (N_4103,In_887,In_3355);
nand U4104 (N_4104,In_4549,In_4097);
nor U4105 (N_4105,In_2133,In_4959);
and U4106 (N_4106,In_4494,In_4124);
xnor U4107 (N_4107,In_242,In_3254);
nor U4108 (N_4108,In_403,In_978);
xnor U4109 (N_4109,In_468,In_3957);
or U4110 (N_4110,In_1413,In_3389);
and U4111 (N_4111,In_4271,In_1913);
nand U4112 (N_4112,In_1553,In_4780);
nor U4113 (N_4113,In_510,In_3623);
nand U4114 (N_4114,In_2064,In_1085);
nor U4115 (N_4115,In_840,In_4463);
nand U4116 (N_4116,In_1424,In_3897);
and U4117 (N_4117,In_2660,In_718);
and U4118 (N_4118,In_1096,In_4011);
nor U4119 (N_4119,In_4062,In_1802);
or U4120 (N_4120,In_4885,In_4718);
xnor U4121 (N_4121,In_1320,In_4028);
nor U4122 (N_4122,In_4606,In_3440);
or U4123 (N_4123,In_1942,In_3836);
nor U4124 (N_4124,In_3929,In_3335);
and U4125 (N_4125,In_2580,In_1128);
nor U4126 (N_4126,In_1694,In_1610);
nor U4127 (N_4127,In_1261,In_2061);
nand U4128 (N_4128,In_1139,In_4200);
or U4129 (N_4129,In_542,In_2532);
and U4130 (N_4130,In_4206,In_4412);
or U4131 (N_4131,In_1789,In_4667);
nand U4132 (N_4132,In_4764,In_1873);
nand U4133 (N_4133,In_679,In_3961);
nand U4134 (N_4134,In_3075,In_4840);
nor U4135 (N_4135,In_1901,In_4069);
xnor U4136 (N_4136,In_2087,In_357);
nand U4137 (N_4137,In_3230,In_3619);
or U4138 (N_4138,In_2528,In_2498);
nor U4139 (N_4139,In_4048,In_2011);
or U4140 (N_4140,In_3566,In_1174);
and U4141 (N_4141,In_4309,In_2846);
nor U4142 (N_4142,In_4587,In_2160);
or U4143 (N_4143,In_1545,In_1207);
xnor U4144 (N_4144,In_2720,In_224);
nand U4145 (N_4145,In_2515,In_129);
or U4146 (N_4146,In_4498,In_443);
and U4147 (N_4147,In_360,In_296);
and U4148 (N_4148,In_1867,In_1641);
nor U4149 (N_4149,In_2823,In_162);
xor U4150 (N_4150,In_3359,In_3809);
xor U4151 (N_4151,In_4752,In_4672);
xor U4152 (N_4152,In_463,In_2185);
nand U4153 (N_4153,In_881,In_4604);
and U4154 (N_4154,In_1670,In_4918);
and U4155 (N_4155,In_4221,In_762);
and U4156 (N_4156,In_2857,In_1803);
nand U4157 (N_4157,In_982,In_3116);
and U4158 (N_4158,In_3256,In_1168);
nand U4159 (N_4159,In_4612,In_1180);
or U4160 (N_4160,In_1810,In_144);
nor U4161 (N_4161,In_4039,In_3307);
nand U4162 (N_4162,In_3412,In_4875);
xor U4163 (N_4163,In_841,In_2145);
nand U4164 (N_4164,In_4510,In_4363);
nand U4165 (N_4165,In_4136,In_1903);
nand U4166 (N_4166,In_641,In_3224);
xor U4167 (N_4167,In_3464,In_4348);
nand U4168 (N_4168,In_2521,In_3362);
and U4169 (N_4169,In_3593,In_77);
and U4170 (N_4170,In_3998,In_2882);
nor U4171 (N_4171,In_2510,In_4830);
or U4172 (N_4172,In_3421,In_223);
or U4173 (N_4173,In_4510,In_4643);
or U4174 (N_4174,In_887,In_4540);
and U4175 (N_4175,In_1257,In_4404);
and U4176 (N_4176,In_3111,In_2837);
nand U4177 (N_4177,In_2169,In_691);
nand U4178 (N_4178,In_4001,In_1002);
or U4179 (N_4179,In_3452,In_1874);
and U4180 (N_4180,In_868,In_382);
nand U4181 (N_4181,In_4667,In_3677);
nand U4182 (N_4182,In_3871,In_375);
nor U4183 (N_4183,In_2000,In_4915);
and U4184 (N_4184,In_3748,In_4370);
nand U4185 (N_4185,In_1663,In_3156);
nand U4186 (N_4186,In_4716,In_739);
nand U4187 (N_4187,In_4227,In_3738);
nand U4188 (N_4188,In_3747,In_4878);
and U4189 (N_4189,In_3566,In_4756);
or U4190 (N_4190,In_2557,In_1389);
xnor U4191 (N_4191,In_3698,In_578);
nor U4192 (N_4192,In_4332,In_4405);
or U4193 (N_4193,In_1660,In_257);
and U4194 (N_4194,In_3439,In_1569);
and U4195 (N_4195,In_123,In_1965);
and U4196 (N_4196,In_2730,In_3434);
nand U4197 (N_4197,In_1471,In_1670);
xor U4198 (N_4198,In_150,In_4527);
and U4199 (N_4199,In_3353,In_4438);
and U4200 (N_4200,In_2956,In_4425);
nor U4201 (N_4201,In_4101,In_3245);
xor U4202 (N_4202,In_4413,In_1115);
nand U4203 (N_4203,In_1893,In_3145);
or U4204 (N_4204,In_742,In_1798);
nor U4205 (N_4205,In_561,In_2907);
or U4206 (N_4206,In_3939,In_745);
and U4207 (N_4207,In_3195,In_2417);
and U4208 (N_4208,In_4090,In_4452);
xor U4209 (N_4209,In_2732,In_2560);
xor U4210 (N_4210,In_3867,In_4891);
and U4211 (N_4211,In_1451,In_4259);
nor U4212 (N_4212,In_4134,In_137);
nor U4213 (N_4213,In_2492,In_1808);
nand U4214 (N_4214,In_3138,In_4104);
or U4215 (N_4215,In_1335,In_1711);
or U4216 (N_4216,In_4441,In_4486);
or U4217 (N_4217,In_1922,In_3997);
or U4218 (N_4218,In_2128,In_2897);
and U4219 (N_4219,In_940,In_517);
xnor U4220 (N_4220,In_4785,In_4015);
and U4221 (N_4221,In_4281,In_1741);
and U4222 (N_4222,In_2014,In_4890);
or U4223 (N_4223,In_4427,In_1850);
or U4224 (N_4224,In_3650,In_144);
nor U4225 (N_4225,In_1889,In_4354);
and U4226 (N_4226,In_4578,In_2825);
or U4227 (N_4227,In_1873,In_844);
nand U4228 (N_4228,In_2438,In_4983);
nand U4229 (N_4229,In_4491,In_1260);
nand U4230 (N_4230,In_4111,In_4300);
xnor U4231 (N_4231,In_2661,In_3994);
or U4232 (N_4232,In_1136,In_3321);
nor U4233 (N_4233,In_2732,In_4436);
and U4234 (N_4234,In_3263,In_2269);
or U4235 (N_4235,In_923,In_4556);
nor U4236 (N_4236,In_4021,In_4649);
nand U4237 (N_4237,In_4197,In_626);
nand U4238 (N_4238,In_3812,In_3118);
and U4239 (N_4239,In_4341,In_1477);
nor U4240 (N_4240,In_1729,In_4096);
nand U4241 (N_4241,In_3380,In_928);
and U4242 (N_4242,In_1729,In_2155);
and U4243 (N_4243,In_3262,In_2726);
nor U4244 (N_4244,In_1522,In_2930);
and U4245 (N_4245,In_3860,In_3197);
xor U4246 (N_4246,In_461,In_2320);
xnor U4247 (N_4247,In_2885,In_771);
nand U4248 (N_4248,In_4625,In_1398);
nor U4249 (N_4249,In_442,In_1142);
and U4250 (N_4250,In_3128,In_3346);
or U4251 (N_4251,In_4728,In_4916);
and U4252 (N_4252,In_2543,In_3432);
nor U4253 (N_4253,In_2080,In_918);
nand U4254 (N_4254,In_416,In_3098);
or U4255 (N_4255,In_2073,In_1137);
nand U4256 (N_4256,In_4436,In_4783);
nand U4257 (N_4257,In_3909,In_3663);
and U4258 (N_4258,In_1452,In_4776);
nand U4259 (N_4259,In_1125,In_303);
nor U4260 (N_4260,In_3695,In_995);
or U4261 (N_4261,In_3281,In_1948);
nor U4262 (N_4262,In_3232,In_4480);
or U4263 (N_4263,In_391,In_2635);
and U4264 (N_4264,In_4584,In_3690);
nor U4265 (N_4265,In_248,In_4984);
or U4266 (N_4266,In_1137,In_4860);
nand U4267 (N_4267,In_4473,In_3930);
nand U4268 (N_4268,In_1616,In_24);
nor U4269 (N_4269,In_3050,In_2561);
xnor U4270 (N_4270,In_2108,In_702);
or U4271 (N_4271,In_3016,In_3299);
nor U4272 (N_4272,In_4909,In_3251);
and U4273 (N_4273,In_1695,In_1053);
xnor U4274 (N_4274,In_300,In_283);
nor U4275 (N_4275,In_4566,In_413);
and U4276 (N_4276,In_2244,In_2532);
nand U4277 (N_4277,In_3822,In_1956);
nand U4278 (N_4278,In_4202,In_63);
or U4279 (N_4279,In_4611,In_2737);
nand U4280 (N_4280,In_1832,In_2326);
nand U4281 (N_4281,In_1956,In_452);
nand U4282 (N_4282,In_1597,In_341);
and U4283 (N_4283,In_2167,In_1135);
or U4284 (N_4284,In_2951,In_3891);
nor U4285 (N_4285,In_4662,In_4726);
and U4286 (N_4286,In_1678,In_4117);
xor U4287 (N_4287,In_1775,In_3951);
and U4288 (N_4288,In_4056,In_3349);
or U4289 (N_4289,In_789,In_4599);
xor U4290 (N_4290,In_2212,In_71);
or U4291 (N_4291,In_3839,In_4476);
nand U4292 (N_4292,In_1941,In_4167);
or U4293 (N_4293,In_1841,In_3967);
nand U4294 (N_4294,In_294,In_1352);
nor U4295 (N_4295,In_2600,In_1608);
nor U4296 (N_4296,In_3692,In_1860);
nor U4297 (N_4297,In_3243,In_445);
nand U4298 (N_4298,In_1301,In_3092);
or U4299 (N_4299,In_1841,In_3265);
nand U4300 (N_4300,In_4810,In_1930);
nor U4301 (N_4301,In_4566,In_3507);
or U4302 (N_4302,In_1199,In_3021);
and U4303 (N_4303,In_2781,In_4724);
or U4304 (N_4304,In_2718,In_3665);
nor U4305 (N_4305,In_3804,In_4620);
nand U4306 (N_4306,In_3409,In_3381);
and U4307 (N_4307,In_49,In_1363);
or U4308 (N_4308,In_3750,In_2896);
xor U4309 (N_4309,In_3535,In_3983);
or U4310 (N_4310,In_2627,In_3981);
nand U4311 (N_4311,In_3259,In_3375);
and U4312 (N_4312,In_732,In_1220);
or U4313 (N_4313,In_4246,In_4142);
and U4314 (N_4314,In_1626,In_4904);
nor U4315 (N_4315,In_4912,In_806);
and U4316 (N_4316,In_4378,In_10);
nand U4317 (N_4317,In_3530,In_770);
and U4318 (N_4318,In_3813,In_2533);
or U4319 (N_4319,In_1908,In_1620);
nand U4320 (N_4320,In_2169,In_3251);
nor U4321 (N_4321,In_3392,In_856);
xor U4322 (N_4322,In_2420,In_4676);
and U4323 (N_4323,In_4728,In_2757);
xnor U4324 (N_4324,In_3185,In_2655);
and U4325 (N_4325,In_1498,In_2887);
xor U4326 (N_4326,In_2140,In_616);
nand U4327 (N_4327,In_2973,In_58);
or U4328 (N_4328,In_2605,In_4995);
nand U4329 (N_4329,In_713,In_3843);
xnor U4330 (N_4330,In_16,In_2497);
or U4331 (N_4331,In_3664,In_3286);
nand U4332 (N_4332,In_4499,In_4472);
or U4333 (N_4333,In_1930,In_3374);
nand U4334 (N_4334,In_41,In_4503);
and U4335 (N_4335,In_4332,In_4494);
nor U4336 (N_4336,In_1002,In_2558);
xnor U4337 (N_4337,In_4681,In_2885);
nand U4338 (N_4338,In_3200,In_1511);
and U4339 (N_4339,In_4342,In_3495);
or U4340 (N_4340,In_1669,In_4353);
nand U4341 (N_4341,In_3726,In_4765);
nand U4342 (N_4342,In_518,In_4909);
nand U4343 (N_4343,In_4503,In_3132);
nand U4344 (N_4344,In_2006,In_571);
nand U4345 (N_4345,In_3539,In_2526);
nand U4346 (N_4346,In_4915,In_2344);
or U4347 (N_4347,In_849,In_3714);
xnor U4348 (N_4348,In_2044,In_2030);
nand U4349 (N_4349,In_2897,In_1156);
nand U4350 (N_4350,In_3232,In_3788);
nor U4351 (N_4351,In_344,In_2527);
nand U4352 (N_4352,In_3886,In_744);
or U4353 (N_4353,In_3782,In_1199);
nor U4354 (N_4354,In_1532,In_250);
nand U4355 (N_4355,In_2984,In_4594);
and U4356 (N_4356,In_1896,In_4872);
xor U4357 (N_4357,In_4135,In_4101);
or U4358 (N_4358,In_1000,In_3182);
nor U4359 (N_4359,In_3490,In_969);
xor U4360 (N_4360,In_33,In_4740);
and U4361 (N_4361,In_187,In_431);
nand U4362 (N_4362,In_4766,In_2471);
xnor U4363 (N_4363,In_552,In_4686);
and U4364 (N_4364,In_3080,In_2940);
nor U4365 (N_4365,In_3134,In_3676);
nor U4366 (N_4366,In_3949,In_1574);
nor U4367 (N_4367,In_3674,In_1972);
and U4368 (N_4368,In_3303,In_1723);
or U4369 (N_4369,In_3133,In_3590);
or U4370 (N_4370,In_4723,In_676);
and U4371 (N_4371,In_1936,In_1545);
xor U4372 (N_4372,In_4066,In_2556);
nor U4373 (N_4373,In_509,In_3378);
nor U4374 (N_4374,In_1897,In_487);
or U4375 (N_4375,In_190,In_1086);
nand U4376 (N_4376,In_812,In_1655);
or U4377 (N_4377,In_3837,In_3041);
nor U4378 (N_4378,In_1807,In_2135);
or U4379 (N_4379,In_1250,In_2577);
nor U4380 (N_4380,In_2491,In_2012);
or U4381 (N_4381,In_1225,In_1203);
or U4382 (N_4382,In_2630,In_3936);
nand U4383 (N_4383,In_4975,In_1544);
nor U4384 (N_4384,In_2381,In_932);
nand U4385 (N_4385,In_1466,In_2510);
or U4386 (N_4386,In_3175,In_4275);
and U4387 (N_4387,In_3320,In_4624);
nand U4388 (N_4388,In_1384,In_1979);
nand U4389 (N_4389,In_4298,In_3315);
nand U4390 (N_4390,In_3508,In_1140);
nand U4391 (N_4391,In_2112,In_1487);
nor U4392 (N_4392,In_3951,In_2500);
and U4393 (N_4393,In_1498,In_890);
nand U4394 (N_4394,In_3500,In_4443);
and U4395 (N_4395,In_4991,In_4417);
and U4396 (N_4396,In_1190,In_162);
and U4397 (N_4397,In_3840,In_4084);
and U4398 (N_4398,In_4506,In_499);
and U4399 (N_4399,In_191,In_1612);
nor U4400 (N_4400,In_2424,In_1346);
nand U4401 (N_4401,In_921,In_4319);
xor U4402 (N_4402,In_4800,In_1118);
nand U4403 (N_4403,In_3735,In_4932);
and U4404 (N_4404,In_2180,In_943);
nand U4405 (N_4405,In_4008,In_3398);
nor U4406 (N_4406,In_1577,In_4333);
or U4407 (N_4407,In_1165,In_206);
nor U4408 (N_4408,In_1833,In_4992);
nor U4409 (N_4409,In_1651,In_277);
nand U4410 (N_4410,In_1386,In_2545);
and U4411 (N_4411,In_184,In_4649);
or U4412 (N_4412,In_3792,In_3912);
or U4413 (N_4413,In_1615,In_2402);
nand U4414 (N_4414,In_2169,In_2161);
nand U4415 (N_4415,In_4702,In_2086);
and U4416 (N_4416,In_4907,In_4278);
or U4417 (N_4417,In_3652,In_2129);
nand U4418 (N_4418,In_634,In_4101);
nor U4419 (N_4419,In_566,In_289);
nand U4420 (N_4420,In_3161,In_196);
nand U4421 (N_4421,In_3055,In_982);
and U4422 (N_4422,In_1441,In_3135);
xor U4423 (N_4423,In_3792,In_4663);
nand U4424 (N_4424,In_394,In_2062);
xnor U4425 (N_4425,In_179,In_3957);
nor U4426 (N_4426,In_2624,In_1287);
and U4427 (N_4427,In_904,In_2329);
nor U4428 (N_4428,In_1431,In_1155);
or U4429 (N_4429,In_3612,In_608);
or U4430 (N_4430,In_3010,In_3334);
nand U4431 (N_4431,In_3910,In_4384);
and U4432 (N_4432,In_572,In_215);
xnor U4433 (N_4433,In_3532,In_2493);
nor U4434 (N_4434,In_2797,In_163);
nor U4435 (N_4435,In_1544,In_940);
nor U4436 (N_4436,In_3897,In_1715);
and U4437 (N_4437,In_3216,In_3805);
and U4438 (N_4438,In_4344,In_1377);
and U4439 (N_4439,In_2595,In_4218);
nor U4440 (N_4440,In_3199,In_1054);
nor U4441 (N_4441,In_1708,In_4554);
or U4442 (N_4442,In_3887,In_4935);
and U4443 (N_4443,In_4653,In_628);
and U4444 (N_4444,In_864,In_121);
and U4445 (N_4445,In_3509,In_618);
xnor U4446 (N_4446,In_912,In_384);
nor U4447 (N_4447,In_831,In_775);
nor U4448 (N_4448,In_823,In_3931);
and U4449 (N_4449,In_3054,In_543);
nor U4450 (N_4450,In_3222,In_3183);
or U4451 (N_4451,In_634,In_4382);
nand U4452 (N_4452,In_1344,In_366);
nor U4453 (N_4453,In_4723,In_2489);
and U4454 (N_4454,In_2970,In_3544);
or U4455 (N_4455,In_1604,In_4194);
nand U4456 (N_4456,In_3571,In_4105);
or U4457 (N_4457,In_4150,In_3846);
nand U4458 (N_4458,In_1849,In_2779);
nand U4459 (N_4459,In_762,In_909);
nor U4460 (N_4460,In_753,In_4113);
nand U4461 (N_4461,In_506,In_2813);
and U4462 (N_4462,In_1824,In_3860);
and U4463 (N_4463,In_1037,In_295);
nor U4464 (N_4464,In_1722,In_1545);
nand U4465 (N_4465,In_734,In_2164);
and U4466 (N_4466,In_2362,In_940);
and U4467 (N_4467,In_3701,In_868);
or U4468 (N_4468,In_856,In_2409);
nand U4469 (N_4469,In_4270,In_4901);
nand U4470 (N_4470,In_4705,In_1334);
nor U4471 (N_4471,In_779,In_2100);
or U4472 (N_4472,In_2666,In_4619);
and U4473 (N_4473,In_3210,In_229);
nand U4474 (N_4474,In_2265,In_995);
or U4475 (N_4475,In_4400,In_4470);
or U4476 (N_4476,In_2361,In_87);
nor U4477 (N_4477,In_3430,In_3869);
xnor U4478 (N_4478,In_111,In_2249);
nand U4479 (N_4479,In_4169,In_300);
or U4480 (N_4480,In_2890,In_3590);
nor U4481 (N_4481,In_4326,In_1468);
nor U4482 (N_4482,In_3264,In_2060);
and U4483 (N_4483,In_4058,In_4492);
and U4484 (N_4484,In_3953,In_1647);
nand U4485 (N_4485,In_3841,In_1306);
nand U4486 (N_4486,In_187,In_3772);
nand U4487 (N_4487,In_3941,In_1639);
xor U4488 (N_4488,In_2947,In_1310);
nand U4489 (N_4489,In_753,In_546);
or U4490 (N_4490,In_4004,In_314);
nor U4491 (N_4491,In_2843,In_3405);
nor U4492 (N_4492,In_4124,In_1405);
and U4493 (N_4493,In_4620,In_2522);
nand U4494 (N_4494,In_2336,In_1159);
and U4495 (N_4495,In_2273,In_1856);
nand U4496 (N_4496,In_3978,In_2540);
nor U4497 (N_4497,In_2923,In_1469);
nor U4498 (N_4498,In_3380,In_1468);
or U4499 (N_4499,In_159,In_2610);
or U4500 (N_4500,In_3624,In_3356);
nor U4501 (N_4501,In_1813,In_3133);
and U4502 (N_4502,In_4157,In_2826);
nand U4503 (N_4503,In_4069,In_4729);
and U4504 (N_4504,In_1782,In_247);
and U4505 (N_4505,In_3352,In_4132);
nor U4506 (N_4506,In_960,In_3333);
and U4507 (N_4507,In_4592,In_4213);
nand U4508 (N_4508,In_1394,In_182);
nand U4509 (N_4509,In_1689,In_3324);
and U4510 (N_4510,In_178,In_4590);
nor U4511 (N_4511,In_3451,In_4088);
nor U4512 (N_4512,In_3376,In_1889);
nand U4513 (N_4513,In_4011,In_2887);
xor U4514 (N_4514,In_349,In_87);
nor U4515 (N_4515,In_2966,In_3077);
xor U4516 (N_4516,In_31,In_1917);
nor U4517 (N_4517,In_519,In_113);
nor U4518 (N_4518,In_4315,In_3909);
or U4519 (N_4519,In_2513,In_907);
nor U4520 (N_4520,In_3837,In_18);
xor U4521 (N_4521,In_3890,In_3744);
or U4522 (N_4522,In_2160,In_1998);
and U4523 (N_4523,In_2930,In_2721);
or U4524 (N_4524,In_753,In_2277);
xor U4525 (N_4525,In_1110,In_1190);
xnor U4526 (N_4526,In_4806,In_3180);
or U4527 (N_4527,In_1485,In_1641);
or U4528 (N_4528,In_4264,In_1831);
and U4529 (N_4529,In_1156,In_4598);
nand U4530 (N_4530,In_1178,In_4107);
or U4531 (N_4531,In_2906,In_2128);
xor U4532 (N_4532,In_2058,In_853);
nand U4533 (N_4533,In_4011,In_2895);
nand U4534 (N_4534,In_803,In_2230);
and U4535 (N_4535,In_4923,In_2389);
nand U4536 (N_4536,In_2690,In_1752);
or U4537 (N_4537,In_257,In_568);
nand U4538 (N_4538,In_4853,In_2061);
or U4539 (N_4539,In_4901,In_4931);
and U4540 (N_4540,In_1497,In_186);
and U4541 (N_4541,In_2551,In_4287);
or U4542 (N_4542,In_3926,In_661);
nand U4543 (N_4543,In_1383,In_3156);
nor U4544 (N_4544,In_4909,In_2339);
and U4545 (N_4545,In_2029,In_2000);
and U4546 (N_4546,In_2190,In_192);
and U4547 (N_4547,In_236,In_1635);
and U4548 (N_4548,In_1069,In_2568);
xor U4549 (N_4549,In_4384,In_4032);
nor U4550 (N_4550,In_2821,In_132);
and U4551 (N_4551,In_4578,In_1521);
or U4552 (N_4552,In_3223,In_4196);
xor U4553 (N_4553,In_413,In_3732);
or U4554 (N_4554,In_4566,In_4848);
and U4555 (N_4555,In_3902,In_1594);
xor U4556 (N_4556,In_3896,In_2296);
xnor U4557 (N_4557,In_4137,In_3738);
nor U4558 (N_4558,In_3272,In_3357);
nand U4559 (N_4559,In_2740,In_1305);
nand U4560 (N_4560,In_3171,In_2596);
nand U4561 (N_4561,In_4685,In_806);
xnor U4562 (N_4562,In_549,In_1443);
nor U4563 (N_4563,In_4602,In_2384);
nor U4564 (N_4564,In_327,In_2493);
xnor U4565 (N_4565,In_3293,In_3180);
nand U4566 (N_4566,In_4893,In_1117);
and U4567 (N_4567,In_4110,In_3672);
nor U4568 (N_4568,In_1618,In_3894);
or U4569 (N_4569,In_4365,In_1791);
nand U4570 (N_4570,In_1953,In_3147);
nand U4571 (N_4571,In_4192,In_2646);
nor U4572 (N_4572,In_1437,In_2041);
and U4573 (N_4573,In_2935,In_2920);
nor U4574 (N_4574,In_4773,In_3);
or U4575 (N_4575,In_3414,In_3649);
nor U4576 (N_4576,In_2196,In_3890);
and U4577 (N_4577,In_3701,In_2938);
nand U4578 (N_4578,In_4278,In_3133);
nor U4579 (N_4579,In_1309,In_4792);
or U4580 (N_4580,In_3128,In_472);
and U4581 (N_4581,In_1461,In_1818);
nand U4582 (N_4582,In_3281,In_3006);
nor U4583 (N_4583,In_1081,In_2684);
nor U4584 (N_4584,In_604,In_3925);
nand U4585 (N_4585,In_4244,In_499);
and U4586 (N_4586,In_3886,In_4627);
and U4587 (N_4587,In_2369,In_1296);
and U4588 (N_4588,In_2953,In_3647);
nand U4589 (N_4589,In_1404,In_4561);
or U4590 (N_4590,In_3822,In_3307);
nand U4591 (N_4591,In_499,In_2289);
nand U4592 (N_4592,In_3231,In_118);
nor U4593 (N_4593,In_4914,In_972);
nand U4594 (N_4594,In_524,In_2217);
xor U4595 (N_4595,In_1096,In_2899);
xor U4596 (N_4596,In_3448,In_2893);
or U4597 (N_4597,In_4096,In_4130);
nand U4598 (N_4598,In_638,In_1713);
xnor U4599 (N_4599,In_4035,In_2572);
nor U4600 (N_4600,In_400,In_770);
and U4601 (N_4601,In_4857,In_4391);
or U4602 (N_4602,In_28,In_3910);
nand U4603 (N_4603,In_3502,In_1057);
or U4604 (N_4604,In_3787,In_1813);
and U4605 (N_4605,In_1500,In_2244);
xnor U4606 (N_4606,In_1762,In_2524);
nand U4607 (N_4607,In_3016,In_1131);
nor U4608 (N_4608,In_3028,In_77);
nor U4609 (N_4609,In_2342,In_2599);
or U4610 (N_4610,In_4766,In_460);
nand U4611 (N_4611,In_1274,In_988);
and U4612 (N_4612,In_4767,In_4301);
or U4613 (N_4613,In_3221,In_643);
nor U4614 (N_4614,In_1815,In_3460);
or U4615 (N_4615,In_1519,In_4823);
and U4616 (N_4616,In_2795,In_1342);
nand U4617 (N_4617,In_668,In_3459);
and U4618 (N_4618,In_3867,In_3866);
nor U4619 (N_4619,In_926,In_454);
nor U4620 (N_4620,In_2561,In_4962);
or U4621 (N_4621,In_3606,In_991);
or U4622 (N_4622,In_2433,In_782);
and U4623 (N_4623,In_3522,In_3028);
nand U4624 (N_4624,In_3780,In_1679);
nor U4625 (N_4625,In_468,In_3337);
nand U4626 (N_4626,In_973,In_1486);
nor U4627 (N_4627,In_2098,In_4818);
and U4628 (N_4628,In_1979,In_4399);
xor U4629 (N_4629,In_3157,In_339);
or U4630 (N_4630,In_2221,In_860);
nor U4631 (N_4631,In_3730,In_2031);
nor U4632 (N_4632,In_2252,In_4589);
nand U4633 (N_4633,In_4726,In_4274);
or U4634 (N_4634,In_4649,In_3843);
or U4635 (N_4635,In_3695,In_3032);
or U4636 (N_4636,In_3752,In_211);
or U4637 (N_4637,In_1720,In_3440);
nand U4638 (N_4638,In_1870,In_4791);
nor U4639 (N_4639,In_243,In_508);
xor U4640 (N_4640,In_218,In_1834);
nor U4641 (N_4641,In_1199,In_771);
nand U4642 (N_4642,In_2293,In_3645);
xor U4643 (N_4643,In_576,In_1634);
and U4644 (N_4644,In_871,In_2147);
nand U4645 (N_4645,In_3628,In_1114);
and U4646 (N_4646,In_1813,In_35);
nand U4647 (N_4647,In_718,In_4923);
nand U4648 (N_4648,In_1690,In_4386);
nor U4649 (N_4649,In_2507,In_3642);
or U4650 (N_4650,In_992,In_10);
nor U4651 (N_4651,In_3485,In_2738);
xnor U4652 (N_4652,In_2897,In_2153);
nand U4653 (N_4653,In_4108,In_4922);
or U4654 (N_4654,In_214,In_4899);
or U4655 (N_4655,In_930,In_4089);
and U4656 (N_4656,In_2271,In_1246);
and U4657 (N_4657,In_2582,In_134);
or U4658 (N_4658,In_2299,In_301);
or U4659 (N_4659,In_1200,In_2354);
nor U4660 (N_4660,In_2444,In_4497);
xor U4661 (N_4661,In_183,In_1391);
or U4662 (N_4662,In_4362,In_4516);
nand U4663 (N_4663,In_628,In_1005);
nand U4664 (N_4664,In_2375,In_2560);
nor U4665 (N_4665,In_3140,In_4190);
nor U4666 (N_4666,In_2134,In_4388);
and U4667 (N_4667,In_2501,In_4364);
nand U4668 (N_4668,In_2555,In_3855);
and U4669 (N_4669,In_1402,In_1898);
nor U4670 (N_4670,In_4091,In_3085);
nor U4671 (N_4671,In_2790,In_3771);
or U4672 (N_4672,In_3717,In_454);
nor U4673 (N_4673,In_3232,In_3185);
nand U4674 (N_4674,In_1585,In_2800);
and U4675 (N_4675,In_3376,In_4084);
nand U4676 (N_4676,In_525,In_3083);
nor U4677 (N_4677,In_3916,In_4024);
and U4678 (N_4678,In_1428,In_4729);
nor U4679 (N_4679,In_4134,In_3844);
and U4680 (N_4680,In_1125,In_4104);
and U4681 (N_4681,In_1626,In_4738);
nor U4682 (N_4682,In_2253,In_630);
xor U4683 (N_4683,In_2170,In_1250);
or U4684 (N_4684,In_4257,In_3927);
or U4685 (N_4685,In_4237,In_943);
nor U4686 (N_4686,In_2501,In_430);
and U4687 (N_4687,In_375,In_3222);
nor U4688 (N_4688,In_938,In_3773);
nand U4689 (N_4689,In_3181,In_1235);
nand U4690 (N_4690,In_3174,In_4712);
nand U4691 (N_4691,In_80,In_4615);
nor U4692 (N_4692,In_1208,In_4542);
nor U4693 (N_4693,In_4184,In_1878);
and U4694 (N_4694,In_1909,In_1558);
or U4695 (N_4695,In_1004,In_927);
or U4696 (N_4696,In_3782,In_1076);
and U4697 (N_4697,In_4965,In_1889);
nor U4698 (N_4698,In_1885,In_3517);
and U4699 (N_4699,In_2520,In_516);
or U4700 (N_4700,In_3982,In_3962);
and U4701 (N_4701,In_3562,In_1781);
or U4702 (N_4702,In_3940,In_508);
and U4703 (N_4703,In_2129,In_928);
and U4704 (N_4704,In_4557,In_1706);
nand U4705 (N_4705,In_2305,In_2992);
nand U4706 (N_4706,In_3133,In_2025);
nor U4707 (N_4707,In_2988,In_3883);
and U4708 (N_4708,In_4887,In_4123);
or U4709 (N_4709,In_4135,In_4822);
nand U4710 (N_4710,In_1948,In_4135);
nand U4711 (N_4711,In_910,In_694);
or U4712 (N_4712,In_3352,In_2785);
and U4713 (N_4713,In_2907,In_174);
and U4714 (N_4714,In_3956,In_63);
or U4715 (N_4715,In_1785,In_1294);
nor U4716 (N_4716,In_4301,In_174);
or U4717 (N_4717,In_3126,In_4984);
nand U4718 (N_4718,In_2612,In_4731);
nand U4719 (N_4719,In_4062,In_773);
and U4720 (N_4720,In_2425,In_3825);
nand U4721 (N_4721,In_333,In_3190);
nand U4722 (N_4722,In_1846,In_3999);
nor U4723 (N_4723,In_1660,In_4682);
or U4724 (N_4724,In_1893,In_3464);
or U4725 (N_4725,In_2320,In_1326);
and U4726 (N_4726,In_2924,In_4216);
nor U4727 (N_4727,In_2731,In_3754);
nand U4728 (N_4728,In_86,In_3430);
and U4729 (N_4729,In_2724,In_2829);
and U4730 (N_4730,In_2189,In_3636);
or U4731 (N_4731,In_497,In_2270);
xnor U4732 (N_4732,In_1816,In_399);
nor U4733 (N_4733,In_4849,In_843);
and U4734 (N_4734,In_4671,In_4873);
nand U4735 (N_4735,In_2335,In_3882);
and U4736 (N_4736,In_4972,In_97);
nor U4737 (N_4737,In_2222,In_642);
nor U4738 (N_4738,In_269,In_2949);
nor U4739 (N_4739,In_1368,In_533);
nand U4740 (N_4740,In_1058,In_178);
and U4741 (N_4741,In_4563,In_2490);
or U4742 (N_4742,In_3452,In_2677);
and U4743 (N_4743,In_2499,In_3346);
or U4744 (N_4744,In_2371,In_2106);
xor U4745 (N_4745,In_2004,In_182);
nor U4746 (N_4746,In_826,In_3485);
and U4747 (N_4747,In_3251,In_625);
or U4748 (N_4748,In_1262,In_3345);
nand U4749 (N_4749,In_3279,In_1539);
nor U4750 (N_4750,In_4652,In_578);
nor U4751 (N_4751,In_2811,In_3288);
or U4752 (N_4752,In_1689,In_2049);
nand U4753 (N_4753,In_4591,In_1432);
nor U4754 (N_4754,In_3696,In_1166);
or U4755 (N_4755,In_3955,In_3893);
nor U4756 (N_4756,In_331,In_2576);
and U4757 (N_4757,In_646,In_1804);
nor U4758 (N_4758,In_1253,In_2015);
nor U4759 (N_4759,In_465,In_3519);
and U4760 (N_4760,In_1199,In_1544);
nand U4761 (N_4761,In_3659,In_4825);
nor U4762 (N_4762,In_2568,In_1184);
or U4763 (N_4763,In_3058,In_1805);
nand U4764 (N_4764,In_3208,In_3155);
or U4765 (N_4765,In_3331,In_3596);
nand U4766 (N_4766,In_4429,In_305);
nand U4767 (N_4767,In_3492,In_1364);
nor U4768 (N_4768,In_1809,In_4841);
nand U4769 (N_4769,In_4722,In_4694);
nand U4770 (N_4770,In_1871,In_2963);
xnor U4771 (N_4771,In_3914,In_865);
nor U4772 (N_4772,In_4345,In_3463);
and U4773 (N_4773,In_2483,In_4782);
and U4774 (N_4774,In_4635,In_4707);
xnor U4775 (N_4775,In_3871,In_3381);
nand U4776 (N_4776,In_4329,In_591);
nand U4777 (N_4777,In_514,In_4182);
nor U4778 (N_4778,In_19,In_4290);
nand U4779 (N_4779,In_690,In_1842);
nand U4780 (N_4780,In_1701,In_964);
nand U4781 (N_4781,In_603,In_1311);
or U4782 (N_4782,In_2064,In_1977);
or U4783 (N_4783,In_3411,In_3111);
nor U4784 (N_4784,In_68,In_3473);
and U4785 (N_4785,In_605,In_3003);
or U4786 (N_4786,In_1536,In_4335);
nand U4787 (N_4787,In_4325,In_3532);
nand U4788 (N_4788,In_3834,In_1631);
nand U4789 (N_4789,In_671,In_3856);
or U4790 (N_4790,In_3095,In_4825);
nand U4791 (N_4791,In_4657,In_981);
nor U4792 (N_4792,In_3045,In_98);
nand U4793 (N_4793,In_4201,In_1846);
and U4794 (N_4794,In_3839,In_3009);
nand U4795 (N_4795,In_2005,In_4622);
nand U4796 (N_4796,In_4765,In_638);
and U4797 (N_4797,In_1672,In_1202);
or U4798 (N_4798,In_3371,In_1195);
nor U4799 (N_4799,In_1460,In_3311);
or U4800 (N_4800,In_30,In_3363);
nor U4801 (N_4801,In_3633,In_3309);
nand U4802 (N_4802,In_4872,In_114);
or U4803 (N_4803,In_3469,In_846);
nand U4804 (N_4804,In_3494,In_2861);
nor U4805 (N_4805,In_1822,In_2602);
xor U4806 (N_4806,In_221,In_1006);
and U4807 (N_4807,In_4788,In_1384);
nor U4808 (N_4808,In_2936,In_1160);
or U4809 (N_4809,In_415,In_4376);
nand U4810 (N_4810,In_678,In_309);
xor U4811 (N_4811,In_700,In_3367);
nand U4812 (N_4812,In_2340,In_4758);
or U4813 (N_4813,In_839,In_2444);
nor U4814 (N_4814,In_3424,In_2130);
and U4815 (N_4815,In_3756,In_3168);
xnor U4816 (N_4816,In_4329,In_689);
nand U4817 (N_4817,In_2213,In_3387);
nor U4818 (N_4818,In_2923,In_1977);
nor U4819 (N_4819,In_2062,In_2797);
nand U4820 (N_4820,In_1649,In_4074);
nor U4821 (N_4821,In_1009,In_601);
xor U4822 (N_4822,In_2150,In_2878);
nand U4823 (N_4823,In_687,In_1273);
nor U4824 (N_4824,In_1325,In_2132);
or U4825 (N_4825,In_1146,In_2506);
nor U4826 (N_4826,In_961,In_1465);
nand U4827 (N_4827,In_2649,In_249);
nor U4828 (N_4828,In_4476,In_3627);
nand U4829 (N_4829,In_3058,In_4869);
or U4830 (N_4830,In_951,In_4755);
or U4831 (N_4831,In_2230,In_1042);
and U4832 (N_4832,In_4516,In_2246);
nor U4833 (N_4833,In_4042,In_3363);
nor U4834 (N_4834,In_4137,In_2722);
or U4835 (N_4835,In_1373,In_878);
and U4836 (N_4836,In_2352,In_3539);
nand U4837 (N_4837,In_1478,In_3299);
nor U4838 (N_4838,In_368,In_4509);
and U4839 (N_4839,In_4068,In_453);
and U4840 (N_4840,In_3462,In_3713);
nand U4841 (N_4841,In_3867,In_3138);
nor U4842 (N_4842,In_71,In_358);
nor U4843 (N_4843,In_2410,In_3789);
xnor U4844 (N_4844,In_2408,In_2111);
and U4845 (N_4845,In_4939,In_2455);
nor U4846 (N_4846,In_4810,In_3969);
nand U4847 (N_4847,In_3914,In_491);
and U4848 (N_4848,In_993,In_1509);
or U4849 (N_4849,In_2507,In_2575);
nand U4850 (N_4850,In_1786,In_161);
xnor U4851 (N_4851,In_4344,In_1468);
nor U4852 (N_4852,In_4601,In_1448);
or U4853 (N_4853,In_1242,In_928);
nor U4854 (N_4854,In_570,In_4064);
and U4855 (N_4855,In_907,In_1773);
nor U4856 (N_4856,In_4583,In_682);
nor U4857 (N_4857,In_4965,In_4732);
or U4858 (N_4858,In_1100,In_1778);
nor U4859 (N_4859,In_989,In_1190);
nor U4860 (N_4860,In_1253,In_2576);
xnor U4861 (N_4861,In_633,In_4257);
nor U4862 (N_4862,In_4467,In_4038);
nor U4863 (N_4863,In_1761,In_2417);
nand U4864 (N_4864,In_1087,In_688);
nor U4865 (N_4865,In_2250,In_648);
and U4866 (N_4866,In_3571,In_3164);
nor U4867 (N_4867,In_1147,In_2526);
and U4868 (N_4868,In_2870,In_1838);
nor U4869 (N_4869,In_2370,In_2954);
nor U4870 (N_4870,In_2391,In_4600);
xnor U4871 (N_4871,In_2436,In_3016);
or U4872 (N_4872,In_1390,In_2377);
xnor U4873 (N_4873,In_1692,In_227);
nor U4874 (N_4874,In_2086,In_1937);
and U4875 (N_4875,In_2858,In_3429);
nor U4876 (N_4876,In_3215,In_3318);
nor U4877 (N_4877,In_2609,In_1491);
and U4878 (N_4878,In_4769,In_3219);
nor U4879 (N_4879,In_893,In_4020);
and U4880 (N_4880,In_2508,In_2325);
or U4881 (N_4881,In_4871,In_3206);
or U4882 (N_4882,In_877,In_684);
nor U4883 (N_4883,In_2642,In_4862);
and U4884 (N_4884,In_4176,In_4673);
and U4885 (N_4885,In_4173,In_4121);
nor U4886 (N_4886,In_4994,In_257);
and U4887 (N_4887,In_2610,In_564);
nor U4888 (N_4888,In_4872,In_3474);
xor U4889 (N_4889,In_3870,In_1452);
or U4890 (N_4890,In_674,In_4542);
nand U4891 (N_4891,In_2328,In_3315);
nand U4892 (N_4892,In_387,In_1460);
or U4893 (N_4893,In_4318,In_2242);
and U4894 (N_4894,In_1303,In_999);
xor U4895 (N_4895,In_1229,In_2205);
and U4896 (N_4896,In_4622,In_3516);
or U4897 (N_4897,In_3290,In_2680);
nand U4898 (N_4898,In_2479,In_2149);
or U4899 (N_4899,In_3859,In_2919);
and U4900 (N_4900,In_2117,In_117);
xnor U4901 (N_4901,In_3036,In_1490);
nand U4902 (N_4902,In_1204,In_1420);
nand U4903 (N_4903,In_4109,In_2146);
and U4904 (N_4904,In_2676,In_4503);
xnor U4905 (N_4905,In_3009,In_1090);
nor U4906 (N_4906,In_1090,In_4242);
and U4907 (N_4907,In_4934,In_558);
xnor U4908 (N_4908,In_2539,In_1575);
or U4909 (N_4909,In_3568,In_596);
and U4910 (N_4910,In_97,In_1287);
nor U4911 (N_4911,In_3038,In_1163);
xnor U4912 (N_4912,In_2833,In_1483);
nor U4913 (N_4913,In_2497,In_1587);
or U4914 (N_4914,In_2190,In_1422);
xor U4915 (N_4915,In_781,In_1125);
or U4916 (N_4916,In_2612,In_3274);
nand U4917 (N_4917,In_741,In_2640);
or U4918 (N_4918,In_2987,In_2211);
and U4919 (N_4919,In_1908,In_2407);
and U4920 (N_4920,In_2102,In_2109);
or U4921 (N_4921,In_2157,In_3562);
nor U4922 (N_4922,In_2010,In_1943);
and U4923 (N_4923,In_393,In_2210);
or U4924 (N_4924,In_2912,In_3785);
xor U4925 (N_4925,In_1565,In_793);
or U4926 (N_4926,In_2589,In_1824);
nand U4927 (N_4927,In_1678,In_2433);
xor U4928 (N_4928,In_991,In_3769);
nand U4929 (N_4929,In_2864,In_2105);
xor U4930 (N_4930,In_415,In_534);
nor U4931 (N_4931,In_963,In_596);
xor U4932 (N_4932,In_2815,In_2581);
nand U4933 (N_4933,In_1411,In_3925);
or U4934 (N_4934,In_4472,In_804);
or U4935 (N_4935,In_2024,In_1219);
or U4936 (N_4936,In_3910,In_1851);
nor U4937 (N_4937,In_4116,In_1395);
nor U4938 (N_4938,In_610,In_1231);
and U4939 (N_4939,In_4039,In_929);
nand U4940 (N_4940,In_3331,In_3433);
nand U4941 (N_4941,In_826,In_4123);
nand U4942 (N_4942,In_2358,In_3404);
xnor U4943 (N_4943,In_1311,In_3887);
xor U4944 (N_4944,In_2069,In_4533);
or U4945 (N_4945,In_3954,In_3988);
or U4946 (N_4946,In_1195,In_168);
nand U4947 (N_4947,In_4089,In_834);
nand U4948 (N_4948,In_855,In_2555);
nor U4949 (N_4949,In_2313,In_3302);
or U4950 (N_4950,In_3474,In_551);
and U4951 (N_4951,In_3971,In_2904);
and U4952 (N_4952,In_4522,In_4932);
or U4953 (N_4953,In_4254,In_1579);
and U4954 (N_4954,In_4204,In_4766);
or U4955 (N_4955,In_4500,In_2423);
and U4956 (N_4956,In_4025,In_2546);
or U4957 (N_4957,In_2340,In_420);
and U4958 (N_4958,In_4997,In_362);
or U4959 (N_4959,In_4759,In_216);
nand U4960 (N_4960,In_2986,In_857);
or U4961 (N_4961,In_1949,In_4242);
nand U4962 (N_4962,In_1083,In_2213);
xnor U4963 (N_4963,In_41,In_482);
nor U4964 (N_4964,In_1377,In_1061);
nor U4965 (N_4965,In_3595,In_4589);
and U4966 (N_4966,In_2881,In_3848);
nand U4967 (N_4967,In_626,In_739);
xor U4968 (N_4968,In_3615,In_1156);
or U4969 (N_4969,In_4701,In_2222);
or U4970 (N_4970,In_2181,In_1555);
or U4971 (N_4971,In_4073,In_975);
and U4972 (N_4972,In_707,In_2834);
and U4973 (N_4973,In_2444,In_4255);
or U4974 (N_4974,In_3963,In_3086);
nand U4975 (N_4975,In_4178,In_2873);
or U4976 (N_4976,In_4865,In_1906);
nor U4977 (N_4977,In_675,In_1723);
nor U4978 (N_4978,In_1148,In_234);
and U4979 (N_4979,In_2710,In_300);
nand U4980 (N_4980,In_2937,In_3339);
or U4981 (N_4981,In_1006,In_4398);
or U4982 (N_4982,In_307,In_2748);
and U4983 (N_4983,In_221,In_2701);
nor U4984 (N_4984,In_3929,In_3008);
nor U4985 (N_4985,In_2357,In_2726);
nand U4986 (N_4986,In_22,In_2963);
or U4987 (N_4987,In_2737,In_2389);
xor U4988 (N_4988,In_3393,In_3126);
or U4989 (N_4989,In_92,In_2420);
or U4990 (N_4990,In_742,In_3357);
and U4991 (N_4991,In_1142,In_4092);
xnor U4992 (N_4992,In_778,In_3569);
or U4993 (N_4993,In_2469,In_4664);
or U4994 (N_4994,In_3685,In_2179);
nand U4995 (N_4995,In_3830,In_3460);
nor U4996 (N_4996,In_3470,In_834);
nor U4997 (N_4997,In_4110,In_4639);
or U4998 (N_4998,In_3677,In_2092);
and U4999 (N_4999,In_439,In_3624);
nand U5000 (N_5000,In_413,In_4331);
or U5001 (N_5001,In_240,In_2901);
or U5002 (N_5002,In_1431,In_3208);
nand U5003 (N_5003,In_3462,In_3823);
and U5004 (N_5004,In_3965,In_968);
or U5005 (N_5005,In_3045,In_4313);
nand U5006 (N_5006,In_672,In_2413);
nor U5007 (N_5007,In_329,In_3389);
or U5008 (N_5008,In_1290,In_4609);
or U5009 (N_5009,In_4009,In_2883);
or U5010 (N_5010,In_1908,In_3540);
xnor U5011 (N_5011,In_1303,In_3135);
nand U5012 (N_5012,In_2168,In_1493);
or U5013 (N_5013,In_4315,In_608);
or U5014 (N_5014,In_4359,In_369);
and U5015 (N_5015,In_1316,In_1282);
or U5016 (N_5016,In_2436,In_1738);
or U5017 (N_5017,In_886,In_3130);
and U5018 (N_5018,In_4887,In_1258);
and U5019 (N_5019,In_1086,In_2789);
nor U5020 (N_5020,In_970,In_1494);
and U5021 (N_5021,In_1460,In_3194);
nand U5022 (N_5022,In_3755,In_4995);
xor U5023 (N_5023,In_757,In_1991);
xor U5024 (N_5024,In_1747,In_1382);
nand U5025 (N_5025,In_63,In_4326);
nor U5026 (N_5026,In_4530,In_1348);
or U5027 (N_5027,In_2424,In_4072);
or U5028 (N_5028,In_1723,In_2058);
nor U5029 (N_5029,In_926,In_3899);
nor U5030 (N_5030,In_2270,In_2803);
and U5031 (N_5031,In_1451,In_4791);
nor U5032 (N_5032,In_3957,In_4319);
nand U5033 (N_5033,In_4558,In_4511);
nand U5034 (N_5034,In_4122,In_4234);
and U5035 (N_5035,In_484,In_3359);
or U5036 (N_5036,In_668,In_3812);
nor U5037 (N_5037,In_4682,In_2341);
nand U5038 (N_5038,In_129,In_1993);
and U5039 (N_5039,In_555,In_1822);
or U5040 (N_5040,In_3175,In_1077);
nor U5041 (N_5041,In_410,In_2250);
nor U5042 (N_5042,In_1261,In_4075);
and U5043 (N_5043,In_172,In_4063);
and U5044 (N_5044,In_3409,In_3681);
nand U5045 (N_5045,In_446,In_3224);
or U5046 (N_5046,In_1685,In_3725);
xnor U5047 (N_5047,In_2391,In_1617);
and U5048 (N_5048,In_731,In_4210);
or U5049 (N_5049,In_3163,In_4092);
and U5050 (N_5050,In_4320,In_1510);
or U5051 (N_5051,In_1605,In_1449);
nor U5052 (N_5052,In_840,In_2601);
nor U5053 (N_5053,In_882,In_474);
and U5054 (N_5054,In_1838,In_950);
or U5055 (N_5055,In_3037,In_1980);
xnor U5056 (N_5056,In_2481,In_4995);
nor U5057 (N_5057,In_2367,In_3743);
nor U5058 (N_5058,In_168,In_2824);
nor U5059 (N_5059,In_443,In_3233);
and U5060 (N_5060,In_1113,In_2955);
and U5061 (N_5061,In_2781,In_1803);
and U5062 (N_5062,In_3820,In_2523);
or U5063 (N_5063,In_2700,In_2034);
or U5064 (N_5064,In_2712,In_1273);
or U5065 (N_5065,In_310,In_3692);
nand U5066 (N_5066,In_4209,In_1236);
and U5067 (N_5067,In_1049,In_1134);
nand U5068 (N_5068,In_981,In_2094);
and U5069 (N_5069,In_2880,In_1061);
nand U5070 (N_5070,In_1294,In_3939);
nor U5071 (N_5071,In_879,In_3219);
xnor U5072 (N_5072,In_853,In_51);
nor U5073 (N_5073,In_366,In_2459);
and U5074 (N_5074,In_1895,In_1985);
and U5075 (N_5075,In_1262,In_1280);
and U5076 (N_5076,In_1636,In_4941);
nand U5077 (N_5077,In_4836,In_4791);
or U5078 (N_5078,In_3878,In_3909);
xor U5079 (N_5079,In_2847,In_777);
or U5080 (N_5080,In_3519,In_2987);
and U5081 (N_5081,In_4885,In_1687);
xor U5082 (N_5082,In_2517,In_4731);
nand U5083 (N_5083,In_2473,In_1523);
nand U5084 (N_5084,In_781,In_35);
nand U5085 (N_5085,In_4483,In_812);
nand U5086 (N_5086,In_1930,In_418);
and U5087 (N_5087,In_1887,In_215);
and U5088 (N_5088,In_4499,In_1278);
nor U5089 (N_5089,In_4630,In_581);
nor U5090 (N_5090,In_4066,In_3484);
and U5091 (N_5091,In_3069,In_3338);
nand U5092 (N_5092,In_2027,In_1526);
nand U5093 (N_5093,In_506,In_458);
nor U5094 (N_5094,In_3352,In_3510);
nand U5095 (N_5095,In_99,In_2575);
nor U5096 (N_5096,In_3716,In_3347);
xnor U5097 (N_5097,In_2596,In_4966);
nand U5098 (N_5098,In_4348,In_1454);
xor U5099 (N_5099,In_1214,In_2035);
and U5100 (N_5100,In_1598,In_1188);
nand U5101 (N_5101,In_4123,In_101);
nand U5102 (N_5102,In_4259,In_4105);
nand U5103 (N_5103,In_3748,In_583);
and U5104 (N_5104,In_2021,In_462);
nand U5105 (N_5105,In_3508,In_3331);
xor U5106 (N_5106,In_4379,In_4080);
or U5107 (N_5107,In_1514,In_4644);
and U5108 (N_5108,In_2431,In_2921);
and U5109 (N_5109,In_464,In_4445);
and U5110 (N_5110,In_941,In_228);
or U5111 (N_5111,In_1412,In_2589);
nor U5112 (N_5112,In_43,In_3194);
xnor U5113 (N_5113,In_442,In_4847);
and U5114 (N_5114,In_3820,In_721);
or U5115 (N_5115,In_2465,In_904);
nand U5116 (N_5116,In_2937,In_1333);
or U5117 (N_5117,In_3795,In_3822);
nand U5118 (N_5118,In_1057,In_2196);
nand U5119 (N_5119,In_3348,In_2182);
nor U5120 (N_5120,In_1885,In_2320);
nand U5121 (N_5121,In_1781,In_757);
nor U5122 (N_5122,In_2412,In_4686);
xor U5123 (N_5123,In_3849,In_1430);
and U5124 (N_5124,In_1894,In_977);
nor U5125 (N_5125,In_111,In_4116);
nand U5126 (N_5126,In_3895,In_4973);
nor U5127 (N_5127,In_3589,In_3700);
or U5128 (N_5128,In_1559,In_3906);
nand U5129 (N_5129,In_1314,In_2494);
xnor U5130 (N_5130,In_1345,In_1505);
and U5131 (N_5131,In_1028,In_2435);
nand U5132 (N_5132,In_2825,In_4571);
and U5133 (N_5133,In_841,In_4046);
xnor U5134 (N_5134,In_1063,In_4911);
and U5135 (N_5135,In_4253,In_4750);
nor U5136 (N_5136,In_688,In_1901);
nor U5137 (N_5137,In_2314,In_1564);
nor U5138 (N_5138,In_3457,In_4010);
and U5139 (N_5139,In_3991,In_847);
and U5140 (N_5140,In_1509,In_3555);
nor U5141 (N_5141,In_212,In_1228);
and U5142 (N_5142,In_2589,In_957);
nor U5143 (N_5143,In_2732,In_135);
nor U5144 (N_5144,In_507,In_2383);
nor U5145 (N_5145,In_713,In_288);
or U5146 (N_5146,In_3996,In_958);
xnor U5147 (N_5147,In_1799,In_3053);
nand U5148 (N_5148,In_3608,In_2090);
and U5149 (N_5149,In_266,In_4869);
and U5150 (N_5150,In_470,In_890);
nand U5151 (N_5151,In_1636,In_3794);
xnor U5152 (N_5152,In_2936,In_1867);
nor U5153 (N_5153,In_83,In_112);
and U5154 (N_5154,In_1459,In_855);
nand U5155 (N_5155,In_1541,In_3848);
nand U5156 (N_5156,In_1123,In_3148);
and U5157 (N_5157,In_1564,In_4546);
and U5158 (N_5158,In_3228,In_2301);
and U5159 (N_5159,In_2601,In_2245);
xnor U5160 (N_5160,In_1263,In_3429);
or U5161 (N_5161,In_1979,In_2456);
or U5162 (N_5162,In_4195,In_365);
and U5163 (N_5163,In_2828,In_2288);
and U5164 (N_5164,In_1222,In_3132);
nand U5165 (N_5165,In_1413,In_3426);
and U5166 (N_5166,In_1170,In_1154);
xor U5167 (N_5167,In_538,In_344);
or U5168 (N_5168,In_45,In_4552);
and U5169 (N_5169,In_1553,In_1362);
nor U5170 (N_5170,In_3541,In_4472);
and U5171 (N_5171,In_814,In_271);
and U5172 (N_5172,In_2678,In_662);
or U5173 (N_5173,In_2060,In_641);
nand U5174 (N_5174,In_207,In_1475);
nand U5175 (N_5175,In_3911,In_1578);
nand U5176 (N_5176,In_2033,In_1232);
xor U5177 (N_5177,In_3148,In_3949);
nand U5178 (N_5178,In_3954,In_3870);
xnor U5179 (N_5179,In_637,In_96);
nor U5180 (N_5180,In_297,In_924);
xnor U5181 (N_5181,In_4000,In_2867);
nand U5182 (N_5182,In_3291,In_3855);
nor U5183 (N_5183,In_904,In_977);
and U5184 (N_5184,In_3698,In_1225);
nand U5185 (N_5185,In_1203,In_2131);
and U5186 (N_5186,In_2373,In_806);
and U5187 (N_5187,In_2460,In_2451);
nor U5188 (N_5188,In_1172,In_405);
nor U5189 (N_5189,In_1422,In_2589);
xnor U5190 (N_5190,In_1177,In_4674);
xnor U5191 (N_5191,In_3054,In_385);
nor U5192 (N_5192,In_4414,In_653);
nand U5193 (N_5193,In_2557,In_4426);
and U5194 (N_5194,In_3047,In_312);
and U5195 (N_5195,In_3461,In_3300);
nand U5196 (N_5196,In_2959,In_2046);
nand U5197 (N_5197,In_2282,In_4286);
nor U5198 (N_5198,In_1324,In_1995);
and U5199 (N_5199,In_1256,In_1473);
or U5200 (N_5200,In_459,In_4429);
xor U5201 (N_5201,In_1637,In_3067);
and U5202 (N_5202,In_991,In_3946);
nor U5203 (N_5203,In_3739,In_1280);
nor U5204 (N_5204,In_1031,In_3839);
or U5205 (N_5205,In_3075,In_2069);
nand U5206 (N_5206,In_1599,In_4572);
or U5207 (N_5207,In_3019,In_4684);
or U5208 (N_5208,In_844,In_2476);
nor U5209 (N_5209,In_402,In_3196);
nand U5210 (N_5210,In_894,In_1878);
nand U5211 (N_5211,In_4428,In_3874);
nor U5212 (N_5212,In_4300,In_3691);
xnor U5213 (N_5213,In_2912,In_4417);
and U5214 (N_5214,In_4003,In_3855);
nand U5215 (N_5215,In_570,In_1161);
or U5216 (N_5216,In_1640,In_2027);
nand U5217 (N_5217,In_1243,In_1563);
or U5218 (N_5218,In_4346,In_3023);
nand U5219 (N_5219,In_1795,In_1402);
or U5220 (N_5220,In_3097,In_2258);
and U5221 (N_5221,In_990,In_4365);
nor U5222 (N_5222,In_4604,In_3370);
nand U5223 (N_5223,In_4458,In_2783);
xnor U5224 (N_5224,In_534,In_3308);
nand U5225 (N_5225,In_1236,In_2632);
or U5226 (N_5226,In_4121,In_894);
nand U5227 (N_5227,In_2207,In_1305);
nor U5228 (N_5228,In_1547,In_780);
nor U5229 (N_5229,In_2152,In_3452);
and U5230 (N_5230,In_3246,In_1517);
and U5231 (N_5231,In_2983,In_4801);
and U5232 (N_5232,In_4822,In_2892);
nor U5233 (N_5233,In_820,In_2129);
and U5234 (N_5234,In_1129,In_1912);
or U5235 (N_5235,In_4592,In_1148);
nand U5236 (N_5236,In_4567,In_2215);
and U5237 (N_5237,In_1421,In_968);
nor U5238 (N_5238,In_738,In_2468);
nand U5239 (N_5239,In_1571,In_1835);
or U5240 (N_5240,In_3994,In_909);
or U5241 (N_5241,In_3738,In_2773);
nand U5242 (N_5242,In_3170,In_1139);
nand U5243 (N_5243,In_1164,In_2547);
nor U5244 (N_5244,In_2672,In_2454);
and U5245 (N_5245,In_2679,In_2223);
or U5246 (N_5246,In_4012,In_375);
nor U5247 (N_5247,In_1633,In_3938);
or U5248 (N_5248,In_4304,In_3000);
or U5249 (N_5249,In_4859,In_4660);
nand U5250 (N_5250,In_1146,In_518);
nand U5251 (N_5251,In_4199,In_2696);
or U5252 (N_5252,In_3508,In_1541);
nand U5253 (N_5253,In_4865,In_4933);
nand U5254 (N_5254,In_1848,In_4854);
nor U5255 (N_5255,In_2081,In_1845);
and U5256 (N_5256,In_2781,In_106);
nand U5257 (N_5257,In_1847,In_2066);
nand U5258 (N_5258,In_2387,In_572);
nand U5259 (N_5259,In_3920,In_3671);
nand U5260 (N_5260,In_316,In_723);
nor U5261 (N_5261,In_589,In_4293);
or U5262 (N_5262,In_2558,In_1558);
and U5263 (N_5263,In_2330,In_3328);
nand U5264 (N_5264,In_2321,In_3126);
nand U5265 (N_5265,In_2285,In_901);
nor U5266 (N_5266,In_3871,In_183);
nand U5267 (N_5267,In_3911,In_307);
nand U5268 (N_5268,In_2855,In_3589);
nand U5269 (N_5269,In_2809,In_1397);
and U5270 (N_5270,In_1174,In_1287);
nand U5271 (N_5271,In_4740,In_858);
xnor U5272 (N_5272,In_1688,In_2406);
or U5273 (N_5273,In_8,In_365);
or U5274 (N_5274,In_43,In_845);
and U5275 (N_5275,In_1485,In_3304);
or U5276 (N_5276,In_1120,In_4646);
or U5277 (N_5277,In_3489,In_3540);
nand U5278 (N_5278,In_1479,In_2123);
or U5279 (N_5279,In_2635,In_3194);
xnor U5280 (N_5280,In_2598,In_320);
nand U5281 (N_5281,In_3113,In_4770);
and U5282 (N_5282,In_2608,In_4389);
and U5283 (N_5283,In_2263,In_2515);
nand U5284 (N_5284,In_2456,In_3785);
xnor U5285 (N_5285,In_2114,In_3108);
and U5286 (N_5286,In_3793,In_3457);
nor U5287 (N_5287,In_1819,In_2273);
nand U5288 (N_5288,In_1122,In_4554);
nor U5289 (N_5289,In_4015,In_4617);
or U5290 (N_5290,In_1530,In_3635);
nor U5291 (N_5291,In_516,In_1348);
or U5292 (N_5292,In_1930,In_3351);
and U5293 (N_5293,In_4871,In_1856);
nor U5294 (N_5294,In_2524,In_377);
nor U5295 (N_5295,In_4183,In_1413);
and U5296 (N_5296,In_4456,In_888);
xnor U5297 (N_5297,In_1519,In_2801);
nand U5298 (N_5298,In_2444,In_4803);
nor U5299 (N_5299,In_139,In_3211);
nand U5300 (N_5300,In_3896,In_519);
and U5301 (N_5301,In_649,In_480);
nor U5302 (N_5302,In_197,In_4416);
nand U5303 (N_5303,In_1204,In_1644);
nand U5304 (N_5304,In_562,In_2620);
nor U5305 (N_5305,In_4763,In_1099);
nor U5306 (N_5306,In_2428,In_4856);
nor U5307 (N_5307,In_4774,In_2867);
or U5308 (N_5308,In_4563,In_968);
and U5309 (N_5309,In_296,In_1569);
nand U5310 (N_5310,In_1190,In_1952);
xnor U5311 (N_5311,In_2742,In_2384);
nor U5312 (N_5312,In_337,In_1425);
and U5313 (N_5313,In_1040,In_647);
or U5314 (N_5314,In_2833,In_4217);
nand U5315 (N_5315,In_4228,In_1301);
xnor U5316 (N_5316,In_3375,In_1527);
nor U5317 (N_5317,In_173,In_2211);
and U5318 (N_5318,In_4316,In_315);
xor U5319 (N_5319,In_3331,In_2815);
nand U5320 (N_5320,In_1767,In_3624);
nor U5321 (N_5321,In_1372,In_4086);
or U5322 (N_5322,In_1545,In_4218);
nor U5323 (N_5323,In_3970,In_347);
or U5324 (N_5324,In_3082,In_1541);
nor U5325 (N_5325,In_53,In_3557);
nand U5326 (N_5326,In_2671,In_3274);
or U5327 (N_5327,In_4855,In_1758);
nor U5328 (N_5328,In_3979,In_3989);
and U5329 (N_5329,In_4861,In_4864);
nor U5330 (N_5330,In_1906,In_740);
and U5331 (N_5331,In_3024,In_2070);
and U5332 (N_5332,In_4908,In_3990);
or U5333 (N_5333,In_799,In_4599);
nand U5334 (N_5334,In_4592,In_3377);
xor U5335 (N_5335,In_3486,In_4914);
xor U5336 (N_5336,In_580,In_1454);
or U5337 (N_5337,In_4789,In_855);
and U5338 (N_5338,In_1642,In_3065);
and U5339 (N_5339,In_4679,In_14);
and U5340 (N_5340,In_2746,In_935);
or U5341 (N_5341,In_1150,In_4792);
nor U5342 (N_5342,In_4275,In_1835);
and U5343 (N_5343,In_4246,In_889);
and U5344 (N_5344,In_3584,In_4090);
and U5345 (N_5345,In_2649,In_4298);
xnor U5346 (N_5346,In_588,In_1692);
nand U5347 (N_5347,In_2455,In_2105);
xor U5348 (N_5348,In_1643,In_3082);
nand U5349 (N_5349,In_1009,In_2212);
and U5350 (N_5350,In_433,In_4213);
or U5351 (N_5351,In_4651,In_3577);
or U5352 (N_5352,In_313,In_2929);
and U5353 (N_5353,In_4868,In_2691);
nand U5354 (N_5354,In_1025,In_2279);
or U5355 (N_5355,In_3978,In_4281);
nor U5356 (N_5356,In_1770,In_3356);
and U5357 (N_5357,In_3783,In_1415);
nand U5358 (N_5358,In_4363,In_2636);
or U5359 (N_5359,In_3987,In_1839);
and U5360 (N_5360,In_4716,In_3209);
nor U5361 (N_5361,In_4934,In_2564);
and U5362 (N_5362,In_3393,In_2839);
or U5363 (N_5363,In_3376,In_2606);
nor U5364 (N_5364,In_3168,In_722);
and U5365 (N_5365,In_1452,In_1783);
nand U5366 (N_5366,In_1787,In_2180);
nor U5367 (N_5367,In_2144,In_3292);
nor U5368 (N_5368,In_2947,In_2074);
nor U5369 (N_5369,In_3108,In_2093);
nand U5370 (N_5370,In_1295,In_3786);
and U5371 (N_5371,In_159,In_2143);
nand U5372 (N_5372,In_3634,In_4979);
xor U5373 (N_5373,In_4017,In_3505);
nand U5374 (N_5374,In_2071,In_3180);
and U5375 (N_5375,In_2344,In_3921);
and U5376 (N_5376,In_733,In_1890);
xor U5377 (N_5377,In_2982,In_3960);
or U5378 (N_5378,In_3886,In_4673);
and U5379 (N_5379,In_3710,In_2167);
nor U5380 (N_5380,In_1709,In_1807);
nand U5381 (N_5381,In_4398,In_4708);
or U5382 (N_5382,In_1517,In_4890);
nor U5383 (N_5383,In_3975,In_42);
nand U5384 (N_5384,In_3877,In_48);
and U5385 (N_5385,In_687,In_2006);
nand U5386 (N_5386,In_4334,In_4747);
or U5387 (N_5387,In_1356,In_1446);
nor U5388 (N_5388,In_1092,In_2716);
and U5389 (N_5389,In_3393,In_3634);
or U5390 (N_5390,In_896,In_853);
or U5391 (N_5391,In_2998,In_2242);
nand U5392 (N_5392,In_570,In_92);
nor U5393 (N_5393,In_3514,In_1416);
and U5394 (N_5394,In_758,In_2009);
or U5395 (N_5395,In_3438,In_3011);
xor U5396 (N_5396,In_4395,In_1698);
or U5397 (N_5397,In_4150,In_2017);
nor U5398 (N_5398,In_31,In_2505);
and U5399 (N_5399,In_2262,In_3270);
and U5400 (N_5400,In_2743,In_3530);
and U5401 (N_5401,In_1454,In_4134);
nand U5402 (N_5402,In_2823,In_2061);
or U5403 (N_5403,In_339,In_3113);
nor U5404 (N_5404,In_2111,In_3260);
nor U5405 (N_5405,In_3305,In_1028);
xor U5406 (N_5406,In_2545,In_2921);
nor U5407 (N_5407,In_3993,In_641);
xnor U5408 (N_5408,In_4223,In_1736);
xnor U5409 (N_5409,In_2665,In_2704);
or U5410 (N_5410,In_4119,In_2356);
nor U5411 (N_5411,In_181,In_2852);
xnor U5412 (N_5412,In_462,In_3560);
and U5413 (N_5413,In_1186,In_2713);
or U5414 (N_5414,In_3259,In_3684);
nor U5415 (N_5415,In_1951,In_3964);
or U5416 (N_5416,In_4415,In_3183);
xnor U5417 (N_5417,In_3596,In_3564);
and U5418 (N_5418,In_562,In_1358);
nor U5419 (N_5419,In_3614,In_2646);
and U5420 (N_5420,In_3384,In_4164);
or U5421 (N_5421,In_1973,In_3705);
and U5422 (N_5422,In_1467,In_2456);
or U5423 (N_5423,In_4931,In_1491);
and U5424 (N_5424,In_2620,In_2107);
and U5425 (N_5425,In_4844,In_3865);
nand U5426 (N_5426,In_1595,In_4198);
nor U5427 (N_5427,In_4194,In_4500);
nor U5428 (N_5428,In_3487,In_97);
and U5429 (N_5429,In_2239,In_3178);
or U5430 (N_5430,In_4715,In_2367);
nand U5431 (N_5431,In_1596,In_1524);
nand U5432 (N_5432,In_4604,In_30);
and U5433 (N_5433,In_3918,In_2389);
xnor U5434 (N_5434,In_2926,In_3215);
and U5435 (N_5435,In_3941,In_3080);
nand U5436 (N_5436,In_1751,In_4231);
nand U5437 (N_5437,In_1506,In_3147);
nor U5438 (N_5438,In_424,In_2655);
nor U5439 (N_5439,In_412,In_4091);
nand U5440 (N_5440,In_2665,In_3457);
and U5441 (N_5441,In_2934,In_347);
or U5442 (N_5442,In_1455,In_4020);
nor U5443 (N_5443,In_3646,In_4890);
or U5444 (N_5444,In_1514,In_3780);
nand U5445 (N_5445,In_381,In_1970);
xor U5446 (N_5446,In_617,In_4733);
and U5447 (N_5447,In_3549,In_2200);
nand U5448 (N_5448,In_1511,In_232);
or U5449 (N_5449,In_18,In_4915);
nor U5450 (N_5450,In_671,In_2894);
nor U5451 (N_5451,In_2068,In_552);
nor U5452 (N_5452,In_1414,In_3271);
and U5453 (N_5453,In_3549,In_1420);
nor U5454 (N_5454,In_2743,In_3876);
nor U5455 (N_5455,In_4902,In_2504);
or U5456 (N_5456,In_119,In_2054);
or U5457 (N_5457,In_4105,In_3678);
and U5458 (N_5458,In_917,In_4695);
and U5459 (N_5459,In_1057,In_2062);
or U5460 (N_5460,In_1531,In_699);
nor U5461 (N_5461,In_3264,In_2195);
or U5462 (N_5462,In_4227,In_4239);
nor U5463 (N_5463,In_1559,In_4749);
nand U5464 (N_5464,In_2984,In_608);
nand U5465 (N_5465,In_4193,In_2074);
or U5466 (N_5466,In_1055,In_379);
or U5467 (N_5467,In_4786,In_1332);
and U5468 (N_5468,In_2658,In_4239);
or U5469 (N_5469,In_431,In_931);
nand U5470 (N_5470,In_510,In_773);
and U5471 (N_5471,In_4388,In_140);
or U5472 (N_5472,In_2757,In_1493);
nand U5473 (N_5473,In_1180,In_1637);
nand U5474 (N_5474,In_4796,In_2321);
nor U5475 (N_5475,In_1283,In_3740);
and U5476 (N_5476,In_340,In_813);
and U5477 (N_5477,In_2004,In_3831);
nand U5478 (N_5478,In_4497,In_4012);
or U5479 (N_5479,In_85,In_561);
nor U5480 (N_5480,In_273,In_4028);
and U5481 (N_5481,In_2203,In_1659);
nand U5482 (N_5482,In_4742,In_867);
nand U5483 (N_5483,In_1319,In_1962);
or U5484 (N_5484,In_135,In_4203);
nand U5485 (N_5485,In_3013,In_2251);
nand U5486 (N_5486,In_2812,In_677);
or U5487 (N_5487,In_842,In_2863);
nor U5488 (N_5488,In_1671,In_4307);
nor U5489 (N_5489,In_1096,In_3648);
nand U5490 (N_5490,In_358,In_4501);
and U5491 (N_5491,In_1743,In_722);
nor U5492 (N_5492,In_2192,In_2620);
nor U5493 (N_5493,In_681,In_4696);
nand U5494 (N_5494,In_4293,In_37);
and U5495 (N_5495,In_4409,In_1281);
and U5496 (N_5496,In_1122,In_3484);
or U5497 (N_5497,In_3111,In_871);
xor U5498 (N_5498,In_3968,In_4751);
and U5499 (N_5499,In_386,In_287);
or U5500 (N_5500,In_387,In_4253);
or U5501 (N_5501,In_1409,In_4243);
xnor U5502 (N_5502,In_3426,In_243);
and U5503 (N_5503,In_1895,In_1412);
and U5504 (N_5504,In_3178,In_2063);
or U5505 (N_5505,In_1037,In_3343);
nand U5506 (N_5506,In_2771,In_1664);
xnor U5507 (N_5507,In_3063,In_2783);
or U5508 (N_5508,In_4363,In_1010);
nand U5509 (N_5509,In_1999,In_3006);
or U5510 (N_5510,In_3961,In_3702);
nand U5511 (N_5511,In_66,In_3035);
nor U5512 (N_5512,In_2685,In_3137);
and U5513 (N_5513,In_1989,In_2853);
xnor U5514 (N_5514,In_2114,In_3953);
nor U5515 (N_5515,In_3147,In_728);
nor U5516 (N_5516,In_1909,In_504);
nand U5517 (N_5517,In_4831,In_2580);
nand U5518 (N_5518,In_3909,In_4106);
and U5519 (N_5519,In_1642,In_696);
nor U5520 (N_5520,In_2752,In_4367);
nand U5521 (N_5521,In_4837,In_2279);
xnor U5522 (N_5522,In_3753,In_227);
or U5523 (N_5523,In_4841,In_4092);
nand U5524 (N_5524,In_812,In_2491);
nand U5525 (N_5525,In_4879,In_3599);
xnor U5526 (N_5526,In_4613,In_4540);
or U5527 (N_5527,In_63,In_2059);
or U5528 (N_5528,In_2697,In_734);
or U5529 (N_5529,In_858,In_527);
nand U5530 (N_5530,In_1159,In_4779);
and U5531 (N_5531,In_1747,In_122);
nand U5532 (N_5532,In_4929,In_4453);
nand U5533 (N_5533,In_3315,In_759);
nand U5534 (N_5534,In_3338,In_1547);
or U5535 (N_5535,In_3234,In_2083);
xnor U5536 (N_5536,In_4283,In_3116);
nor U5537 (N_5537,In_1471,In_4313);
xnor U5538 (N_5538,In_2278,In_4815);
nand U5539 (N_5539,In_592,In_3026);
or U5540 (N_5540,In_2624,In_4587);
nand U5541 (N_5541,In_2387,In_3120);
xnor U5542 (N_5542,In_4443,In_2491);
xor U5543 (N_5543,In_3622,In_3245);
and U5544 (N_5544,In_4082,In_787);
nor U5545 (N_5545,In_976,In_4641);
or U5546 (N_5546,In_4773,In_936);
nor U5547 (N_5547,In_2031,In_4463);
nor U5548 (N_5548,In_4875,In_4336);
nor U5549 (N_5549,In_3491,In_193);
xor U5550 (N_5550,In_1606,In_157);
nand U5551 (N_5551,In_189,In_495);
nand U5552 (N_5552,In_2639,In_868);
nor U5553 (N_5553,In_1320,In_985);
and U5554 (N_5554,In_618,In_560);
nand U5555 (N_5555,In_1241,In_109);
and U5556 (N_5556,In_4110,In_3731);
nor U5557 (N_5557,In_401,In_3805);
nand U5558 (N_5558,In_1518,In_2743);
and U5559 (N_5559,In_3429,In_3285);
xnor U5560 (N_5560,In_4064,In_2486);
xor U5561 (N_5561,In_1271,In_2663);
nand U5562 (N_5562,In_4646,In_4911);
nand U5563 (N_5563,In_1715,In_3144);
nor U5564 (N_5564,In_1840,In_607);
or U5565 (N_5565,In_3390,In_3861);
and U5566 (N_5566,In_1073,In_332);
nand U5567 (N_5567,In_4831,In_599);
nand U5568 (N_5568,In_3454,In_744);
and U5569 (N_5569,In_3835,In_528);
nor U5570 (N_5570,In_3764,In_2673);
nor U5571 (N_5571,In_2291,In_2474);
xnor U5572 (N_5572,In_3669,In_3331);
or U5573 (N_5573,In_1631,In_4506);
nor U5574 (N_5574,In_4279,In_4221);
nand U5575 (N_5575,In_6,In_2317);
nor U5576 (N_5576,In_3003,In_3332);
or U5577 (N_5577,In_1579,In_3202);
nand U5578 (N_5578,In_2016,In_1623);
and U5579 (N_5579,In_4977,In_2964);
nor U5580 (N_5580,In_61,In_4181);
nor U5581 (N_5581,In_697,In_2385);
nand U5582 (N_5582,In_1936,In_3145);
nor U5583 (N_5583,In_3581,In_1652);
nor U5584 (N_5584,In_3370,In_1928);
nor U5585 (N_5585,In_2940,In_3159);
nor U5586 (N_5586,In_1674,In_161);
nand U5587 (N_5587,In_666,In_4655);
nor U5588 (N_5588,In_4535,In_3526);
nand U5589 (N_5589,In_3239,In_4440);
or U5590 (N_5590,In_4991,In_1975);
or U5591 (N_5591,In_2943,In_1232);
or U5592 (N_5592,In_3957,In_2941);
nor U5593 (N_5593,In_985,In_2251);
nand U5594 (N_5594,In_3065,In_3301);
xor U5595 (N_5595,In_918,In_2072);
nor U5596 (N_5596,In_4695,In_2380);
nor U5597 (N_5597,In_4971,In_4122);
nor U5598 (N_5598,In_4303,In_4166);
and U5599 (N_5599,In_4699,In_1465);
and U5600 (N_5600,In_2085,In_1131);
or U5601 (N_5601,In_1289,In_2077);
nand U5602 (N_5602,In_927,In_2905);
or U5603 (N_5603,In_4048,In_2765);
or U5604 (N_5604,In_4233,In_4327);
xor U5605 (N_5605,In_1230,In_1584);
or U5606 (N_5606,In_152,In_1508);
xnor U5607 (N_5607,In_4548,In_133);
and U5608 (N_5608,In_1281,In_4950);
nor U5609 (N_5609,In_3224,In_3601);
and U5610 (N_5610,In_1940,In_1339);
or U5611 (N_5611,In_4471,In_3697);
and U5612 (N_5612,In_3467,In_1256);
and U5613 (N_5613,In_1502,In_3985);
and U5614 (N_5614,In_4187,In_2748);
or U5615 (N_5615,In_3509,In_3655);
or U5616 (N_5616,In_3515,In_2841);
and U5617 (N_5617,In_513,In_2852);
or U5618 (N_5618,In_632,In_1792);
nand U5619 (N_5619,In_1456,In_2317);
and U5620 (N_5620,In_1208,In_931);
and U5621 (N_5621,In_985,In_4165);
and U5622 (N_5622,In_4235,In_4895);
nor U5623 (N_5623,In_4804,In_567);
nor U5624 (N_5624,In_4183,In_3509);
and U5625 (N_5625,In_3641,In_4257);
nand U5626 (N_5626,In_2705,In_3522);
nor U5627 (N_5627,In_1409,In_2555);
xnor U5628 (N_5628,In_2087,In_2157);
nor U5629 (N_5629,In_3814,In_942);
or U5630 (N_5630,In_396,In_4389);
or U5631 (N_5631,In_4025,In_2650);
and U5632 (N_5632,In_4236,In_4740);
and U5633 (N_5633,In_3736,In_71);
nand U5634 (N_5634,In_3974,In_4824);
nor U5635 (N_5635,In_823,In_3072);
nand U5636 (N_5636,In_3938,In_1365);
nand U5637 (N_5637,In_2538,In_3833);
or U5638 (N_5638,In_1936,In_343);
nor U5639 (N_5639,In_2723,In_2305);
or U5640 (N_5640,In_1768,In_4955);
or U5641 (N_5641,In_859,In_256);
xnor U5642 (N_5642,In_3550,In_3976);
or U5643 (N_5643,In_1675,In_1800);
nand U5644 (N_5644,In_1484,In_4487);
or U5645 (N_5645,In_4107,In_3053);
or U5646 (N_5646,In_3607,In_4867);
and U5647 (N_5647,In_3393,In_86);
xnor U5648 (N_5648,In_755,In_2332);
or U5649 (N_5649,In_838,In_3397);
or U5650 (N_5650,In_2649,In_3740);
and U5651 (N_5651,In_2847,In_1842);
and U5652 (N_5652,In_1076,In_3909);
nand U5653 (N_5653,In_4235,In_3557);
or U5654 (N_5654,In_4205,In_2140);
or U5655 (N_5655,In_1127,In_1179);
or U5656 (N_5656,In_2724,In_1515);
nand U5657 (N_5657,In_4519,In_4167);
nand U5658 (N_5658,In_986,In_4851);
and U5659 (N_5659,In_3884,In_3152);
and U5660 (N_5660,In_4291,In_4017);
and U5661 (N_5661,In_2380,In_394);
and U5662 (N_5662,In_1849,In_1754);
nor U5663 (N_5663,In_3383,In_4473);
nor U5664 (N_5664,In_1684,In_2486);
and U5665 (N_5665,In_1657,In_4331);
and U5666 (N_5666,In_1224,In_1138);
and U5667 (N_5667,In_1541,In_4986);
nor U5668 (N_5668,In_1025,In_2641);
and U5669 (N_5669,In_562,In_4100);
nor U5670 (N_5670,In_4610,In_79);
and U5671 (N_5671,In_2664,In_2704);
and U5672 (N_5672,In_1332,In_3861);
nand U5673 (N_5673,In_623,In_442);
and U5674 (N_5674,In_3223,In_3898);
or U5675 (N_5675,In_4992,In_993);
nor U5676 (N_5676,In_2422,In_3837);
and U5677 (N_5677,In_4841,In_330);
or U5678 (N_5678,In_3701,In_3834);
nand U5679 (N_5679,In_3233,In_3234);
nor U5680 (N_5680,In_2933,In_570);
and U5681 (N_5681,In_3224,In_1761);
or U5682 (N_5682,In_3276,In_1704);
and U5683 (N_5683,In_1251,In_1073);
nor U5684 (N_5684,In_3681,In_346);
nor U5685 (N_5685,In_1954,In_3039);
nand U5686 (N_5686,In_780,In_1063);
nand U5687 (N_5687,In_3491,In_3381);
or U5688 (N_5688,In_2322,In_2705);
nand U5689 (N_5689,In_4948,In_4641);
nor U5690 (N_5690,In_4166,In_2694);
nand U5691 (N_5691,In_1854,In_4678);
nand U5692 (N_5692,In_961,In_2316);
nand U5693 (N_5693,In_2977,In_3540);
nand U5694 (N_5694,In_84,In_3670);
nand U5695 (N_5695,In_786,In_4657);
and U5696 (N_5696,In_1612,In_2147);
xor U5697 (N_5697,In_2234,In_4495);
and U5698 (N_5698,In_76,In_4661);
xnor U5699 (N_5699,In_2977,In_1658);
nor U5700 (N_5700,In_3541,In_738);
or U5701 (N_5701,In_3040,In_3704);
and U5702 (N_5702,In_633,In_2986);
nand U5703 (N_5703,In_1682,In_2202);
xor U5704 (N_5704,In_3225,In_3196);
nand U5705 (N_5705,In_1552,In_4514);
or U5706 (N_5706,In_722,In_1524);
and U5707 (N_5707,In_4045,In_173);
xnor U5708 (N_5708,In_3795,In_2938);
nor U5709 (N_5709,In_2400,In_4114);
and U5710 (N_5710,In_1151,In_1272);
nor U5711 (N_5711,In_2229,In_2077);
and U5712 (N_5712,In_842,In_4518);
nand U5713 (N_5713,In_1270,In_1116);
nor U5714 (N_5714,In_2672,In_1304);
xor U5715 (N_5715,In_204,In_4950);
and U5716 (N_5716,In_4749,In_1025);
nand U5717 (N_5717,In_1165,In_447);
nand U5718 (N_5718,In_3760,In_672);
nor U5719 (N_5719,In_3466,In_1919);
nand U5720 (N_5720,In_4697,In_183);
nand U5721 (N_5721,In_1627,In_2063);
nand U5722 (N_5722,In_4813,In_310);
nand U5723 (N_5723,In_3494,In_4772);
and U5724 (N_5724,In_3802,In_1723);
and U5725 (N_5725,In_1737,In_1923);
or U5726 (N_5726,In_1139,In_692);
or U5727 (N_5727,In_3543,In_215);
nor U5728 (N_5728,In_593,In_3053);
nor U5729 (N_5729,In_4644,In_4770);
xor U5730 (N_5730,In_317,In_2350);
or U5731 (N_5731,In_4800,In_3281);
nand U5732 (N_5732,In_4641,In_2282);
and U5733 (N_5733,In_2655,In_626);
and U5734 (N_5734,In_2940,In_2636);
or U5735 (N_5735,In_2164,In_2033);
or U5736 (N_5736,In_327,In_4426);
nor U5737 (N_5737,In_1995,In_1436);
xnor U5738 (N_5738,In_4776,In_3626);
or U5739 (N_5739,In_2985,In_231);
or U5740 (N_5740,In_4227,In_950);
or U5741 (N_5741,In_607,In_2077);
and U5742 (N_5742,In_2483,In_51);
xor U5743 (N_5743,In_3535,In_1036);
nand U5744 (N_5744,In_2742,In_1821);
nand U5745 (N_5745,In_1185,In_4946);
nor U5746 (N_5746,In_4124,In_489);
nor U5747 (N_5747,In_3799,In_3774);
nor U5748 (N_5748,In_3026,In_926);
nand U5749 (N_5749,In_2139,In_2449);
nor U5750 (N_5750,In_4069,In_1962);
or U5751 (N_5751,In_1990,In_1164);
nor U5752 (N_5752,In_693,In_3177);
nand U5753 (N_5753,In_2522,In_2225);
xor U5754 (N_5754,In_4766,In_2911);
nand U5755 (N_5755,In_134,In_2738);
xnor U5756 (N_5756,In_2672,In_4126);
nor U5757 (N_5757,In_258,In_3822);
nand U5758 (N_5758,In_839,In_2027);
nor U5759 (N_5759,In_905,In_4545);
nor U5760 (N_5760,In_4960,In_648);
nor U5761 (N_5761,In_1118,In_4997);
and U5762 (N_5762,In_3374,In_2717);
or U5763 (N_5763,In_616,In_3993);
or U5764 (N_5764,In_4105,In_1514);
xnor U5765 (N_5765,In_3685,In_4708);
and U5766 (N_5766,In_2725,In_2720);
or U5767 (N_5767,In_59,In_3785);
nand U5768 (N_5768,In_2732,In_2179);
nand U5769 (N_5769,In_695,In_36);
or U5770 (N_5770,In_3286,In_4546);
or U5771 (N_5771,In_1530,In_3571);
and U5772 (N_5772,In_904,In_1384);
nor U5773 (N_5773,In_4112,In_4104);
nor U5774 (N_5774,In_4621,In_3757);
xnor U5775 (N_5775,In_4185,In_3906);
or U5776 (N_5776,In_1095,In_1491);
nand U5777 (N_5777,In_2065,In_279);
and U5778 (N_5778,In_1848,In_3666);
xnor U5779 (N_5779,In_3914,In_739);
nand U5780 (N_5780,In_981,In_1133);
xnor U5781 (N_5781,In_570,In_836);
nand U5782 (N_5782,In_4553,In_4124);
nand U5783 (N_5783,In_230,In_2465);
and U5784 (N_5784,In_350,In_1976);
xnor U5785 (N_5785,In_3649,In_4977);
and U5786 (N_5786,In_15,In_1227);
and U5787 (N_5787,In_4600,In_3886);
nor U5788 (N_5788,In_3742,In_1014);
nor U5789 (N_5789,In_337,In_4035);
nand U5790 (N_5790,In_1780,In_3608);
xnor U5791 (N_5791,In_3863,In_789);
nor U5792 (N_5792,In_2136,In_2361);
or U5793 (N_5793,In_731,In_1692);
nor U5794 (N_5794,In_2965,In_1214);
and U5795 (N_5795,In_974,In_1652);
xnor U5796 (N_5796,In_2682,In_2117);
and U5797 (N_5797,In_17,In_1586);
nand U5798 (N_5798,In_2094,In_2355);
nor U5799 (N_5799,In_3923,In_3720);
and U5800 (N_5800,In_2766,In_3952);
nand U5801 (N_5801,In_3668,In_149);
nand U5802 (N_5802,In_3482,In_1522);
nand U5803 (N_5803,In_895,In_4442);
and U5804 (N_5804,In_2167,In_252);
or U5805 (N_5805,In_4611,In_1473);
nand U5806 (N_5806,In_2720,In_2452);
and U5807 (N_5807,In_2015,In_3964);
or U5808 (N_5808,In_398,In_4934);
and U5809 (N_5809,In_4363,In_3949);
nor U5810 (N_5810,In_4026,In_570);
or U5811 (N_5811,In_1919,In_4623);
xor U5812 (N_5812,In_4749,In_1082);
or U5813 (N_5813,In_4311,In_686);
or U5814 (N_5814,In_2897,In_4616);
or U5815 (N_5815,In_3482,In_4753);
or U5816 (N_5816,In_1580,In_636);
nand U5817 (N_5817,In_4048,In_3634);
and U5818 (N_5818,In_2520,In_1205);
or U5819 (N_5819,In_2630,In_2496);
and U5820 (N_5820,In_3673,In_1900);
or U5821 (N_5821,In_3178,In_1756);
and U5822 (N_5822,In_2379,In_1312);
nand U5823 (N_5823,In_4698,In_4561);
or U5824 (N_5824,In_1724,In_3088);
and U5825 (N_5825,In_3461,In_55);
or U5826 (N_5826,In_3062,In_2975);
xnor U5827 (N_5827,In_924,In_2412);
or U5828 (N_5828,In_976,In_3296);
and U5829 (N_5829,In_4328,In_1855);
xnor U5830 (N_5830,In_1794,In_1243);
nor U5831 (N_5831,In_3010,In_3537);
or U5832 (N_5832,In_2025,In_2059);
nor U5833 (N_5833,In_217,In_4070);
xnor U5834 (N_5834,In_2175,In_4837);
nor U5835 (N_5835,In_2289,In_1117);
nand U5836 (N_5836,In_4429,In_1241);
or U5837 (N_5837,In_3050,In_4763);
nand U5838 (N_5838,In_4741,In_1867);
nand U5839 (N_5839,In_657,In_328);
nor U5840 (N_5840,In_1762,In_1798);
or U5841 (N_5841,In_1106,In_2443);
nand U5842 (N_5842,In_1261,In_66);
or U5843 (N_5843,In_1744,In_3494);
or U5844 (N_5844,In_4735,In_3131);
or U5845 (N_5845,In_4105,In_3036);
and U5846 (N_5846,In_2703,In_2849);
and U5847 (N_5847,In_372,In_4868);
nand U5848 (N_5848,In_2695,In_3440);
and U5849 (N_5849,In_3310,In_2136);
xnor U5850 (N_5850,In_2416,In_1607);
nor U5851 (N_5851,In_4735,In_2501);
xor U5852 (N_5852,In_2486,In_839);
and U5853 (N_5853,In_2469,In_4543);
nor U5854 (N_5854,In_1576,In_4747);
nor U5855 (N_5855,In_186,In_672);
or U5856 (N_5856,In_3612,In_1647);
nand U5857 (N_5857,In_4116,In_3455);
or U5858 (N_5858,In_624,In_3635);
nand U5859 (N_5859,In_3002,In_2858);
nor U5860 (N_5860,In_4005,In_111);
nor U5861 (N_5861,In_47,In_4419);
and U5862 (N_5862,In_3845,In_163);
and U5863 (N_5863,In_1664,In_3588);
and U5864 (N_5864,In_3133,In_4433);
nor U5865 (N_5865,In_208,In_4720);
nand U5866 (N_5866,In_3896,In_2066);
xnor U5867 (N_5867,In_1910,In_1971);
xnor U5868 (N_5868,In_1836,In_4313);
nor U5869 (N_5869,In_4904,In_4613);
or U5870 (N_5870,In_793,In_2974);
or U5871 (N_5871,In_1883,In_579);
nor U5872 (N_5872,In_2637,In_3099);
and U5873 (N_5873,In_2930,In_4706);
or U5874 (N_5874,In_1644,In_2612);
nor U5875 (N_5875,In_1870,In_1906);
and U5876 (N_5876,In_1598,In_1465);
or U5877 (N_5877,In_125,In_118);
nor U5878 (N_5878,In_711,In_2383);
nand U5879 (N_5879,In_155,In_4419);
or U5880 (N_5880,In_1762,In_3452);
xor U5881 (N_5881,In_1280,In_1693);
or U5882 (N_5882,In_3449,In_1273);
nor U5883 (N_5883,In_2122,In_1072);
and U5884 (N_5884,In_2037,In_3258);
or U5885 (N_5885,In_3925,In_4122);
xor U5886 (N_5886,In_4244,In_4665);
or U5887 (N_5887,In_742,In_4390);
or U5888 (N_5888,In_1321,In_3442);
nor U5889 (N_5889,In_4462,In_2078);
xor U5890 (N_5890,In_937,In_2600);
nand U5891 (N_5891,In_263,In_3209);
and U5892 (N_5892,In_711,In_1474);
nor U5893 (N_5893,In_4574,In_3410);
nand U5894 (N_5894,In_1389,In_1177);
or U5895 (N_5895,In_1323,In_4378);
and U5896 (N_5896,In_1482,In_2063);
and U5897 (N_5897,In_3970,In_3226);
and U5898 (N_5898,In_3409,In_3454);
nor U5899 (N_5899,In_668,In_4823);
xor U5900 (N_5900,In_3180,In_1650);
nor U5901 (N_5901,In_156,In_1909);
and U5902 (N_5902,In_3698,In_3582);
nor U5903 (N_5903,In_1042,In_3054);
nor U5904 (N_5904,In_4314,In_76);
or U5905 (N_5905,In_4790,In_2889);
xor U5906 (N_5906,In_1616,In_1590);
or U5907 (N_5907,In_610,In_4107);
or U5908 (N_5908,In_4598,In_4993);
and U5909 (N_5909,In_2042,In_3077);
and U5910 (N_5910,In_26,In_1877);
nand U5911 (N_5911,In_2100,In_3991);
xor U5912 (N_5912,In_4560,In_2101);
xor U5913 (N_5913,In_1825,In_3460);
and U5914 (N_5914,In_1808,In_1025);
and U5915 (N_5915,In_2959,In_811);
nand U5916 (N_5916,In_2106,In_3854);
nor U5917 (N_5917,In_3975,In_3957);
nor U5918 (N_5918,In_1370,In_1899);
and U5919 (N_5919,In_623,In_4086);
or U5920 (N_5920,In_2464,In_1031);
xnor U5921 (N_5921,In_2377,In_4929);
or U5922 (N_5922,In_4249,In_1191);
or U5923 (N_5923,In_4371,In_3814);
nor U5924 (N_5924,In_3130,In_2662);
or U5925 (N_5925,In_1941,In_2592);
nand U5926 (N_5926,In_100,In_4275);
xor U5927 (N_5927,In_4074,In_3288);
or U5928 (N_5928,In_2763,In_1860);
and U5929 (N_5929,In_4707,In_1831);
and U5930 (N_5930,In_1696,In_478);
nor U5931 (N_5931,In_3613,In_2717);
nor U5932 (N_5932,In_3038,In_1950);
or U5933 (N_5933,In_1348,In_19);
and U5934 (N_5934,In_1502,In_3474);
nand U5935 (N_5935,In_2189,In_2900);
and U5936 (N_5936,In_4948,In_3866);
and U5937 (N_5937,In_4691,In_1664);
and U5938 (N_5938,In_3784,In_4187);
nor U5939 (N_5939,In_1428,In_3479);
nor U5940 (N_5940,In_1621,In_1316);
nand U5941 (N_5941,In_2111,In_1764);
or U5942 (N_5942,In_1827,In_1672);
nor U5943 (N_5943,In_4288,In_2527);
or U5944 (N_5944,In_4635,In_3971);
and U5945 (N_5945,In_4085,In_4144);
or U5946 (N_5946,In_3205,In_3338);
nand U5947 (N_5947,In_4574,In_4093);
nor U5948 (N_5948,In_1102,In_3706);
xor U5949 (N_5949,In_994,In_3297);
nand U5950 (N_5950,In_2634,In_4332);
and U5951 (N_5951,In_4445,In_1265);
nand U5952 (N_5952,In_1615,In_4607);
or U5953 (N_5953,In_2905,In_1579);
nand U5954 (N_5954,In_662,In_1097);
or U5955 (N_5955,In_4579,In_1196);
xor U5956 (N_5956,In_670,In_3006);
nand U5957 (N_5957,In_1806,In_2159);
and U5958 (N_5958,In_1064,In_4563);
nand U5959 (N_5959,In_2794,In_4921);
nor U5960 (N_5960,In_1484,In_2743);
or U5961 (N_5961,In_1805,In_217);
and U5962 (N_5962,In_3975,In_1545);
and U5963 (N_5963,In_1048,In_3801);
and U5964 (N_5964,In_4877,In_3005);
xor U5965 (N_5965,In_1220,In_3841);
nor U5966 (N_5966,In_3632,In_2861);
and U5967 (N_5967,In_298,In_3372);
nand U5968 (N_5968,In_765,In_2901);
and U5969 (N_5969,In_4491,In_1962);
and U5970 (N_5970,In_3902,In_1021);
nand U5971 (N_5971,In_2405,In_4117);
and U5972 (N_5972,In_3614,In_2387);
nor U5973 (N_5973,In_1571,In_2105);
or U5974 (N_5974,In_1150,In_3246);
nor U5975 (N_5975,In_2493,In_1527);
xnor U5976 (N_5976,In_2612,In_2829);
or U5977 (N_5977,In_3753,In_2158);
nor U5978 (N_5978,In_711,In_3321);
nor U5979 (N_5979,In_1103,In_1741);
or U5980 (N_5980,In_484,In_332);
and U5981 (N_5981,In_3644,In_2600);
and U5982 (N_5982,In_2807,In_2692);
nand U5983 (N_5983,In_789,In_461);
nor U5984 (N_5984,In_978,In_3696);
nand U5985 (N_5985,In_250,In_1506);
xor U5986 (N_5986,In_4784,In_2041);
xnor U5987 (N_5987,In_1929,In_2115);
and U5988 (N_5988,In_2572,In_1133);
nor U5989 (N_5989,In_1300,In_3171);
or U5990 (N_5990,In_4132,In_2984);
and U5991 (N_5991,In_1372,In_16);
xor U5992 (N_5992,In_4140,In_1262);
or U5993 (N_5993,In_2687,In_811);
nand U5994 (N_5994,In_3988,In_2202);
and U5995 (N_5995,In_1761,In_4305);
or U5996 (N_5996,In_2988,In_748);
or U5997 (N_5997,In_3442,In_2744);
and U5998 (N_5998,In_4611,In_1216);
nor U5999 (N_5999,In_3192,In_3067);
xnor U6000 (N_6000,In_1957,In_351);
and U6001 (N_6001,In_4789,In_2539);
nand U6002 (N_6002,In_750,In_4943);
and U6003 (N_6003,In_1117,In_3006);
or U6004 (N_6004,In_3728,In_2526);
nor U6005 (N_6005,In_643,In_820);
or U6006 (N_6006,In_1305,In_4769);
and U6007 (N_6007,In_1081,In_3023);
xor U6008 (N_6008,In_2942,In_628);
nor U6009 (N_6009,In_4356,In_1153);
nor U6010 (N_6010,In_1498,In_58);
nor U6011 (N_6011,In_454,In_1188);
nor U6012 (N_6012,In_4277,In_41);
nor U6013 (N_6013,In_2315,In_3673);
or U6014 (N_6014,In_4364,In_1135);
nor U6015 (N_6015,In_4663,In_4033);
and U6016 (N_6016,In_1071,In_1560);
xnor U6017 (N_6017,In_3850,In_3809);
and U6018 (N_6018,In_22,In_4102);
nor U6019 (N_6019,In_3222,In_2748);
nor U6020 (N_6020,In_4293,In_1120);
nor U6021 (N_6021,In_713,In_3778);
nand U6022 (N_6022,In_2885,In_4329);
nor U6023 (N_6023,In_1891,In_942);
or U6024 (N_6024,In_1188,In_3524);
nand U6025 (N_6025,In_908,In_1945);
and U6026 (N_6026,In_2665,In_3252);
nand U6027 (N_6027,In_1921,In_3761);
nand U6028 (N_6028,In_3076,In_3250);
and U6029 (N_6029,In_4404,In_546);
xor U6030 (N_6030,In_3142,In_3858);
nand U6031 (N_6031,In_4940,In_977);
or U6032 (N_6032,In_1976,In_1320);
and U6033 (N_6033,In_2007,In_762);
nand U6034 (N_6034,In_1934,In_939);
and U6035 (N_6035,In_4492,In_2981);
and U6036 (N_6036,In_2370,In_4779);
and U6037 (N_6037,In_2693,In_3435);
nand U6038 (N_6038,In_4956,In_3001);
and U6039 (N_6039,In_755,In_1835);
xnor U6040 (N_6040,In_2747,In_2576);
nand U6041 (N_6041,In_4452,In_975);
or U6042 (N_6042,In_139,In_2119);
and U6043 (N_6043,In_2505,In_4852);
or U6044 (N_6044,In_849,In_3248);
xor U6045 (N_6045,In_1232,In_4745);
or U6046 (N_6046,In_2550,In_1584);
nand U6047 (N_6047,In_1757,In_4385);
and U6048 (N_6048,In_2424,In_2756);
nor U6049 (N_6049,In_2992,In_370);
nor U6050 (N_6050,In_190,In_1362);
nand U6051 (N_6051,In_1490,In_4441);
or U6052 (N_6052,In_1136,In_583);
nand U6053 (N_6053,In_741,In_1762);
xnor U6054 (N_6054,In_1931,In_2558);
or U6055 (N_6055,In_4644,In_948);
nor U6056 (N_6056,In_4158,In_229);
nand U6057 (N_6057,In_2356,In_3403);
and U6058 (N_6058,In_4951,In_4770);
xor U6059 (N_6059,In_4055,In_319);
and U6060 (N_6060,In_4925,In_2885);
or U6061 (N_6061,In_2542,In_2987);
nor U6062 (N_6062,In_3853,In_3207);
and U6063 (N_6063,In_4862,In_3492);
and U6064 (N_6064,In_4990,In_231);
nand U6065 (N_6065,In_891,In_3528);
nand U6066 (N_6066,In_125,In_4537);
nor U6067 (N_6067,In_3333,In_2840);
nand U6068 (N_6068,In_4861,In_4001);
nand U6069 (N_6069,In_3521,In_3477);
and U6070 (N_6070,In_2788,In_2085);
or U6071 (N_6071,In_1688,In_2613);
or U6072 (N_6072,In_3447,In_198);
or U6073 (N_6073,In_4745,In_2339);
nor U6074 (N_6074,In_2954,In_2329);
nand U6075 (N_6075,In_180,In_1438);
nor U6076 (N_6076,In_4933,In_3549);
or U6077 (N_6077,In_938,In_2246);
and U6078 (N_6078,In_1930,In_1358);
and U6079 (N_6079,In_1099,In_3290);
or U6080 (N_6080,In_2667,In_885);
xnor U6081 (N_6081,In_3921,In_866);
or U6082 (N_6082,In_3830,In_1032);
and U6083 (N_6083,In_312,In_4868);
nand U6084 (N_6084,In_236,In_2621);
nand U6085 (N_6085,In_4775,In_1861);
or U6086 (N_6086,In_884,In_166);
or U6087 (N_6087,In_4960,In_231);
nand U6088 (N_6088,In_882,In_3279);
nor U6089 (N_6089,In_3957,In_3061);
nand U6090 (N_6090,In_2336,In_667);
and U6091 (N_6091,In_701,In_1350);
nor U6092 (N_6092,In_4279,In_1523);
and U6093 (N_6093,In_3622,In_317);
xor U6094 (N_6094,In_2850,In_999);
nor U6095 (N_6095,In_3686,In_592);
nand U6096 (N_6096,In_288,In_3832);
nand U6097 (N_6097,In_1799,In_1101);
nor U6098 (N_6098,In_4167,In_305);
and U6099 (N_6099,In_4427,In_817);
nor U6100 (N_6100,In_120,In_4976);
xor U6101 (N_6101,In_505,In_918);
and U6102 (N_6102,In_2327,In_3325);
nand U6103 (N_6103,In_4383,In_4869);
xnor U6104 (N_6104,In_838,In_2046);
xor U6105 (N_6105,In_1287,In_2102);
and U6106 (N_6106,In_1755,In_249);
or U6107 (N_6107,In_4784,In_737);
or U6108 (N_6108,In_3980,In_1368);
nor U6109 (N_6109,In_4883,In_3314);
nor U6110 (N_6110,In_1909,In_2634);
nand U6111 (N_6111,In_1895,In_3794);
nor U6112 (N_6112,In_889,In_1919);
or U6113 (N_6113,In_1676,In_1471);
or U6114 (N_6114,In_1890,In_2682);
nand U6115 (N_6115,In_2562,In_1767);
xnor U6116 (N_6116,In_753,In_801);
or U6117 (N_6117,In_4024,In_2093);
xor U6118 (N_6118,In_192,In_4610);
nand U6119 (N_6119,In_3537,In_2867);
and U6120 (N_6120,In_957,In_2366);
and U6121 (N_6121,In_2347,In_2539);
or U6122 (N_6122,In_1586,In_2711);
nor U6123 (N_6123,In_2658,In_633);
nor U6124 (N_6124,In_2881,In_754);
or U6125 (N_6125,In_3334,In_1064);
and U6126 (N_6126,In_2753,In_1049);
nor U6127 (N_6127,In_2611,In_3403);
xor U6128 (N_6128,In_3843,In_4313);
and U6129 (N_6129,In_134,In_857);
nand U6130 (N_6130,In_2049,In_3675);
nand U6131 (N_6131,In_3566,In_4183);
or U6132 (N_6132,In_3081,In_1648);
nand U6133 (N_6133,In_4369,In_1726);
nand U6134 (N_6134,In_191,In_684);
nor U6135 (N_6135,In_1648,In_3975);
nand U6136 (N_6136,In_1218,In_524);
and U6137 (N_6137,In_858,In_4574);
or U6138 (N_6138,In_3594,In_2706);
nand U6139 (N_6139,In_4507,In_1701);
and U6140 (N_6140,In_1096,In_3408);
or U6141 (N_6141,In_3837,In_362);
xor U6142 (N_6142,In_3932,In_1237);
xnor U6143 (N_6143,In_4280,In_4777);
nand U6144 (N_6144,In_680,In_4223);
nand U6145 (N_6145,In_2216,In_4123);
nand U6146 (N_6146,In_4509,In_1133);
nand U6147 (N_6147,In_4125,In_127);
and U6148 (N_6148,In_3309,In_4261);
nor U6149 (N_6149,In_95,In_1836);
and U6150 (N_6150,In_3778,In_1542);
nand U6151 (N_6151,In_629,In_3928);
and U6152 (N_6152,In_3325,In_3572);
and U6153 (N_6153,In_3008,In_1182);
nand U6154 (N_6154,In_190,In_2535);
and U6155 (N_6155,In_2692,In_2296);
nor U6156 (N_6156,In_1036,In_643);
and U6157 (N_6157,In_4415,In_1513);
and U6158 (N_6158,In_2725,In_2987);
and U6159 (N_6159,In_1539,In_3829);
and U6160 (N_6160,In_1200,In_422);
nor U6161 (N_6161,In_3786,In_1725);
nor U6162 (N_6162,In_1529,In_518);
nand U6163 (N_6163,In_1273,In_1288);
or U6164 (N_6164,In_1390,In_779);
xor U6165 (N_6165,In_4607,In_2703);
and U6166 (N_6166,In_654,In_1558);
nor U6167 (N_6167,In_4682,In_2051);
nor U6168 (N_6168,In_1199,In_1826);
xor U6169 (N_6169,In_1113,In_2578);
and U6170 (N_6170,In_2532,In_4324);
or U6171 (N_6171,In_137,In_3110);
nor U6172 (N_6172,In_2401,In_68);
xnor U6173 (N_6173,In_3181,In_4053);
nand U6174 (N_6174,In_4455,In_1008);
nor U6175 (N_6175,In_529,In_734);
nor U6176 (N_6176,In_4431,In_105);
or U6177 (N_6177,In_3843,In_4096);
nor U6178 (N_6178,In_4945,In_2049);
nor U6179 (N_6179,In_2643,In_4878);
or U6180 (N_6180,In_2312,In_204);
xnor U6181 (N_6181,In_2872,In_230);
and U6182 (N_6182,In_2438,In_647);
or U6183 (N_6183,In_2610,In_1824);
nand U6184 (N_6184,In_2100,In_4360);
or U6185 (N_6185,In_1614,In_2076);
and U6186 (N_6186,In_857,In_849);
xnor U6187 (N_6187,In_2117,In_2445);
xnor U6188 (N_6188,In_1529,In_2642);
nor U6189 (N_6189,In_1680,In_2653);
nor U6190 (N_6190,In_4440,In_3746);
nor U6191 (N_6191,In_2851,In_504);
or U6192 (N_6192,In_1678,In_3340);
nor U6193 (N_6193,In_3523,In_2868);
and U6194 (N_6194,In_3988,In_1048);
and U6195 (N_6195,In_14,In_2794);
or U6196 (N_6196,In_2317,In_2357);
and U6197 (N_6197,In_3386,In_3489);
and U6198 (N_6198,In_4075,In_4970);
or U6199 (N_6199,In_1832,In_3682);
and U6200 (N_6200,In_2097,In_1470);
nor U6201 (N_6201,In_4675,In_3538);
and U6202 (N_6202,In_2327,In_2132);
nand U6203 (N_6203,In_2085,In_123);
or U6204 (N_6204,In_2276,In_4663);
and U6205 (N_6205,In_3635,In_2050);
or U6206 (N_6206,In_1890,In_3364);
nor U6207 (N_6207,In_4686,In_1634);
or U6208 (N_6208,In_2960,In_926);
nor U6209 (N_6209,In_1681,In_3651);
xor U6210 (N_6210,In_3976,In_584);
nor U6211 (N_6211,In_4899,In_2552);
nand U6212 (N_6212,In_759,In_3355);
nor U6213 (N_6213,In_793,In_2779);
nand U6214 (N_6214,In_1443,In_1306);
nand U6215 (N_6215,In_89,In_2535);
or U6216 (N_6216,In_4017,In_246);
or U6217 (N_6217,In_3000,In_83);
nand U6218 (N_6218,In_663,In_3991);
nand U6219 (N_6219,In_1088,In_1181);
nor U6220 (N_6220,In_2765,In_2388);
and U6221 (N_6221,In_2871,In_3151);
or U6222 (N_6222,In_1295,In_1618);
nand U6223 (N_6223,In_1905,In_1187);
nand U6224 (N_6224,In_1283,In_3016);
or U6225 (N_6225,In_2912,In_1015);
or U6226 (N_6226,In_862,In_4493);
and U6227 (N_6227,In_3288,In_3728);
or U6228 (N_6228,In_769,In_4723);
nor U6229 (N_6229,In_1344,In_764);
nor U6230 (N_6230,In_1372,In_1696);
nand U6231 (N_6231,In_2495,In_3010);
or U6232 (N_6232,In_1001,In_3567);
nor U6233 (N_6233,In_4859,In_2442);
nand U6234 (N_6234,In_1640,In_1955);
or U6235 (N_6235,In_2765,In_977);
nand U6236 (N_6236,In_3572,In_1303);
and U6237 (N_6237,In_186,In_1476);
and U6238 (N_6238,In_4293,In_1496);
and U6239 (N_6239,In_3879,In_4997);
and U6240 (N_6240,In_2068,In_1835);
and U6241 (N_6241,In_700,In_242);
xor U6242 (N_6242,In_4272,In_1300);
nand U6243 (N_6243,In_4789,In_1617);
nand U6244 (N_6244,In_4616,In_3541);
xnor U6245 (N_6245,In_2381,In_1574);
nand U6246 (N_6246,In_4890,In_4417);
nand U6247 (N_6247,In_1429,In_3502);
nor U6248 (N_6248,In_4513,In_1083);
and U6249 (N_6249,In_719,In_890);
and U6250 (N_6250,In_1166,In_3511);
and U6251 (N_6251,In_2688,In_4109);
nor U6252 (N_6252,In_2557,In_3227);
and U6253 (N_6253,In_1632,In_1751);
nand U6254 (N_6254,In_372,In_3787);
nand U6255 (N_6255,In_2298,In_3721);
and U6256 (N_6256,In_2179,In_2948);
nor U6257 (N_6257,In_992,In_2015);
nor U6258 (N_6258,In_3041,In_3580);
nor U6259 (N_6259,In_2704,In_3090);
and U6260 (N_6260,In_2709,In_3208);
nor U6261 (N_6261,In_2279,In_189);
or U6262 (N_6262,In_4906,In_3962);
and U6263 (N_6263,In_3839,In_2126);
or U6264 (N_6264,In_3561,In_3715);
nand U6265 (N_6265,In_2766,In_3149);
xor U6266 (N_6266,In_3938,In_3789);
and U6267 (N_6267,In_4097,In_3856);
or U6268 (N_6268,In_1858,In_3943);
nand U6269 (N_6269,In_1171,In_153);
nor U6270 (N_6270,In_3757,In_1689);
nor U6271 (N_6271,In_1416,In_4760);
xnor U6272 (N_6272,In_189,In_4950);
and U6273 (N_6273,In_2560,In_2482);
and U6274 (N_6274,In_3024,In_3629);
nor U6275 (N_6275,In_2704,In_3137);
and U6276 (N_6276,In_1812,In_3262);
or U6277 (N_6277,In_3008,In_427);
and U6278 (N_6278,In_2610,In_1915);
nor U6279 (N_6279,In_563,In_2587);
xnor U6280 (N_6280,In_2730,In_2888);
nand U6281 (N_6281,In_1239,In_2033);
nand U6282 (N_6282,In_4679,In_2750);
nand U6283 (N_6283,In_297,In_2810);
nand U6284 (N_6284,In_1590,In_3250);
nand U6285 (N_6285,In_1402,In_146);
and U6286 (N_6286,In_3555,In_3451);
nor U6287 (N_6287,In_4233,In_4406);
nand U6288 (N_6288,In_1397,In_4541);
xnor U6289 (N_6289,In_1067,In_26);
or U6290 (N_6290,In_2678,In_4549);
or U6291 (N_6291,In_786,In_3275);
or U6292 (N_6292,In_584,In_2045);
and U6293 (N_6293,In_4592,In_2220);
or U6294 (N_6294,In_4829,In_2448);
or U6295 (N_6295,In_4165,In_399);
and U6296 (N_6296,In_980,In_698);
nand U6297 (N_6297,In_1824,In_4414);
and U6298 (N_6298,In_3256,In_721);
xor U6299 (N_6299,In_263,In_4167);
xor U6300 (N_6300,In_10,In_3141);
nand U6301 (N_6301,In_3913,In_1599);
and U6302 (N_6302,In_3004,In_702);
or U6303 (N_6303,In_1836,In_3534);
nand U6304 (N_6304,In_4108,In_399);
nor U6305 (N_6305,In_1705,In_1242);
nand U6306 (N_6306,In_704,In_3493);
nor U6307 (N_6307,In_2178,In_847);
nand U6308 (N_6308,In_3970,In_3872);
xor U6309 (N_6309,In_4837,In_3873);
xor U6310 (N_6310,In_796,In_4647);
and U6311 (N_6311,In_1464,In_2277);
and U6312 (N_6312,In_4398,In_1682);
nor U6313 (N_6313,In_3975,In_2491);
nand U6314 (N_6314,In_2625,In_561);
and U6315 (N_6315,In_621,In_3202);
nor U6316 (N_6316,In_3225,In_4591);
or U6317 (N_6317,In_1776,In_4475);
and U6318 (N_6318,In_3147,In_2783);
nand U6319 (N_6319,In_487,In_4129);
nand U6320 (N_6320,In_1637,In_4843);
and U6321 (N_6321,In_4553,In_4421);
xor U6322 (N_6322,In_1573,In_2291);
and U6323 (N_6323,In_1290,In_3649);
nand U6324 (N_6324,In_3651,In_126);
and U6325 (N_6325,In_2866,In_530);
and U6326 (N_6326,In_1952,In_2357);
and U6327 (N_6327,In_3640,In_4003);
and U6328 (N_6328,In_4188,In_2078);
nand U6329 (N_6329,In_895,In_4196);
and U6330 (N_6330,In_3149,In_3469);
nor U6331 (N_6331,In_3385,In_2838);
nand U6332 (N_6332,In_4417,In_1536);
xnor U6333 (N_6333,In_4027,In_2992);
nor U6334 (N_6334,In_1662,In_3541);
xor U6335 (N_6335,In_602,In_4466);
and U6336 (N_6336,In_2173,In_3773);
or U6337 (N_6337,In_2220,In_3061);
nand U6338 (N_6338,In_2585,In_2226);
and U6339 (N_6339,In_2899,In_1377);
nor U6340 (N_6340,In_4563,In_3793);
nor U6341 (N_6341,In_923,In_1164);
or U6342 (N_6342,In_1187,In_3260);
and U6343 (N_6343,In_3448,In_1262);
or U6344 (N_6344,In_3483,In_658);
nand U6345 (N_6345,In_4670,In_1359);
nand U6346 (N_6346,In_2536,In_38);
and U6347 (N_6347,In_118,In_1355);
nand U6348 (N_6348,In_4401,In_3773);
nor U6349 (N_6349,In_4152,In_3836);
or U6350 (N_6350,In_4783,In_1978);
nand U6351 (N_6351,In_592,In_3506);
nor U6352 (N_6352,In_1574,In_3118);
nand U6353 (N_6353,In_3875,In_4013);
nor U6354 (N_6354,In_2749,In_1451);
and U6355 (N_6355,In_3228,In_1427);
or U6356 (N_6356,In_2740,In_4432);
xnor U6357 (N_6357,In_1395,In_4782);
nor U6358 (N_6358,In_4903,In_1404);
or U6359 (N_6359,In_4169,In_3403);
and U6360 (N_6360,In_1751,In_1315);
nor U6361 (N_6361,In_2998,In_4728);
or U6362 (N_6362,In_3052,In_3416);
nand U6363 (N_6363,In_4615,In_771);
nor U6364 (N_6364,In_615,In_2325);
and U6365 (N_6365,In_2976,In_1048);
and U6366 (N_6366,In_1006,In_4115);
xnor U6367 (N_6367,In_4058,In_4293);
nand U6368 (N_6368,In_733,In_1390);
nor U6369 (N_6369,In_654,In_225);
or U6370 (N_6370,In_2723,In_4076);
nand U6371 (N_6371,In_4575,In_2075);
nand U6372 (N_6372,In_4644,In_3378);
and U6373 (N_6373,In_520,In_4717);
and U6374 (N_6374,In_629,In_649);
and U6375 (N_6375,In_4624,In_743);
xnor U6376 (N_6376,In_2629,In_4228);
nor U6377 (N_6377,In_2864,In_2573);
nor U6378 (N_6378,In_504,In_464);
nand U6379 (N_6379,In_934,In_4685);
or U6380 (N_6380,In_4657,In_3409);
or U6381 (N_6381,In_4850,In_2592);
nor U6382 (N_6382,In_4312,In_726);
or U6383 (N_6383,In_3725,In_2731);
nor U6384 (N_6384,In_1301,In_1549);
or U6385 (N_6385,In_3243,In_2984);
nand U6386 (N_6386,In_3597,In_4981);
or U6387 (N_6387,In_264,In_3649);
and U6388 (N_6388,In_1385,In_3639);
or U6389 (N_6389,In_4687,In_3160);
or U6390 (N_6390,In_1528,In_3077);
nor U6391 (N_6391,In_2907,In_1823);
or U6392 (N_6392,In_1355,In_709);
nand U6393 (N_6393,In_1472,In_1255);
and U6394 (N_6394,In_3087,In_4941);
and U6395 (N_6395,In_599,In_3154);
and U6396 (N_6396,In_3608,In_1865);
or U6397 (N_6397,In_3964,In_51);
or U6398 (N_6398,In_748,In_3854);
nand U6399 (N_6399,In_4330,In_3897);
nor U6400 (N_6400,In_1214,In_544);
and U6401 (N_6401,In_2006,In_4714);
xor U6402 (N_6402,In_3415,In_2521);
nand U6403 (N_6403,In_4730,In_3995);
and U6404 (N_6404,In_1881,In_1762);
nor U6405 (N_6405,In_2314,In_3770);
nand U6406 (N_6406,In_2878,In_2907);
or U6407 (N_6407,In_1866,In_3949);
nor U6408 (N_6408,In_3823,In_2521);
nand U6409 (N_6409,In_511,In_2657);
nand U6410 (N_6410,In_4181,In_3540);
or U6411 (N_6411,In_1554,In_58);
and U6412 (N_6412,In_2275,In_2513);
nor U6413 (N_6413,In_567,In_1799);
nand U6414 (N_6414,In_3626,In_780);
nand U6415 (N_6415,In_4744,In_3921);
nor U6416 (N_6416,In_226,In_2192);
nand U6417 (N_6417,In_2293,In_2653);
nor U6418 (N_6418,In_3336,In_1619);
xnor U6419 (N_6419,In_2157,In_1006);
xnor U6420 (N_6420,In_537,In_4567);
nor U6421 (N_6421,In_1945,In_1317);
nor U6422 (N_6422,In_2546,In_1016);
and U6423 (N_6423,In_2752,In_4968);
nor U6424 (N_6424,In_4331,In_1178);
and U6425 (N_6425,In_4415,In_4903);
or U6426 (N_6426,In_26,In_1942);
or U6427 (N_6427,In_2422,In_3777);
xnor U6428 (N_6428,In_1067,In_2002);
and U6429 (N_6429,In_4246,In_65);
and U6430 (N_6430,In_3515,In_2943);
xnor U6431 (N_6431,In_4995,In_2347);
and U6432 (N_6432,In_3144,In_290);
and U6433 (N_6433,In_4164,In_4629);
and U6434 (N_6434,In_1326,In_3460);
xnor U6435 (N_6435,In_1225,In_3589);
nand U6436 (N_6436,In_4089,In_2726);
nand U6437 (N_6437,In_2532,In_4034);
and U6438 (N_6438,In_878,In_417);
nor U6439 (N_6439,In_1515,In_2858);
nor U6440 (N_6440,In_3662,In_4826);
or U6441 (N_6441,In_2283,In_4389);
and U6442 (N_6442,In_4532,In_1823);
and U6443 (N_6443,In_534,In_3309);
nand U6444 (N_6444,In_3507,In_4999);
and U6445 (N_6445,In_1529,In_3757);
or U6446 (N_6446,In_998,In_1964);
nand U6447 (N_6447,In_4757,In_3769);
nor U6448 (N_6448,In_2521,In_3681);
nand U6449 (N_6449,In_4885,In_1312);
and U6450 (N_6450,In_2636,In_4957);
nor U6451 (N_6451,In_2826,In_562);
nand U6452 (N_6452,In_2454,In_1861);
or U6453 (N_6453,In_4808,In_1866);
xor U6454 (N_6454,In_1190,In_4933);
or U6455 (N_6455,In_2809,In_4020);
nor U6456 (N_6456,In_1284,In_1311);
and U6457 (N_6457,In_3315,In_325);
and U6458 (N_6458,In_374,In_2348);
and U6459 (N_6459,In_4224,In_3829);
xor U6460 (N_6460,In_535,In_2080);
and U6461 (N_6461,In_1360,In_4630);
nor U6462 (N_6462,In_2971,In_2327);
and U6463 (N_6463,In_2907,In_238);
nand U6464 (N_6464,In_2003,In_4044);
or U6465 (N_6465,In_4909,In_4491);
xor U6466 (N_6466,In_1646,In_2886);
nand U6467 (N_6467,In_4838,In_4695);
and U6468 (N_6468,In_4914,In_2883);
nor U6469 (N_6469,In_4245,In_3585);
or U6470 (N_6470,In_4007,In_3572);
and U6471 (N_6471,In_879,In_1138);
nand U6472 (N_6472,In_1355,In_784);
and U6473 (N_6473,In_771,In_115);
or U6474 (N_6474,In_1218,In_3638);
and U6475 (N_6475,In_2499,In_4001);
or U6476 (N_6476,In_4312,In_1219);
or U6477 (N_6477,In_2182,In_4255);
and U6478 (N_6478,In_3451,In_4807);
and U6479 (N_6479,In_3848,In_183);
nor U6480 (N_6480,In_216,In_2849);
nor U6481 (N_6481,In_4611,In_3432);
nand U6482 (N_6482,In_1683,In_2969);
nand U6483 (N_6483,In_1930,In_1544);
nor U6484 (N_6484,In_2858,In_2384);
nor U6485 (N_6485,In_516,In_2458);
and U6486 (N_6486,In_2719,In_4160);
nor U6487 (N_6487,In_3449,In_3386);
nand U6488 (N_6488,In_3032,In_3796);
or U6489 (N_6489,In_3517,In_3248);
nor U6490 (N_6490,In_3119,In_2028);
nor U6491 (N_6491,In_720,In_4404);
or U6492 (N_6492,In_1510,In_3333);
xor U6493 (N_6493,In_3299,In_354);
and U6494 (N_6494,In_3832,In_1324);
xor U6495 (N_6495,In_905,In_3997);
or U6496 (N_6496,In_3662,In_1573);
nor U6497 (N_6497,In_2788,In_4942);
and U6498 (N_6498,In_956,In_173);
or U6499 (N_6499,In_1034,In_4478);
or U6500 (N_6500,In_4881,In_893);
xor U6501 (N_6501,In_95,In_1883);
or U6502 (N_6502,In_2884,In_1837);
and U6503 (N_6503,In_107,In_139);
nor U6504 (N_6504,In_1783,In_5);
nand U6505 (N_6505,In_3565,In_4362);
nor U6506 (N_6506,In_4723,In_2332);
nor U6507 (N_6507,In_1279,In_2177);
xnor U6508 (N_6508,In_1194,In_2305);
nand U6509 (N_6509,In_4572,In_429);
and U6510 (N_6510,In_334,In_2248);
xnor U6511 (N_6511,In_3592,In_4463);
and U6512 (N_6512,In_3186,In_2216);
nor U6513 (N_6513,In_4972,In_1357);
nor U6514 (N_6514,In_1093,In_1724);
and U6515 (N_6515,In_701,In_400);
and U6516 (N_6516,In_4565,In_1424);
nor U6517 (N_6517,In_1509,In_4395);
nor U6518 (N_6518,In_3649,In_4566);
xor U6519 (N_6519,In_769,In_2990);
and U6520 (N_6520,In_2107,In_4434);
nand U6521 (N_6521,In_4138,In_2814);
nand U6522 (N_6522,In_86,In_2547);
nand U6523 (N_6523,In_4076,In_3269);
or U6524 (N_6524,In_386,In_3657);
nand U6525 (N_6525,In_4988,In_1277);
nor U6526 (N_6526,In_2275,In_3695);
nand U6527 (N_6527,In_2849,In_1661);
and U6528 (N_6528,In_4113,In_3756);
or U6529 (N_6529,In_1230,In_3350);
nand U6530 (N_6530,In_3835,In_2943);
nand U6531 (N_6531,In_1089,In_3);
nor U6532 (N_6532,In_3193,In_3833);
and U6533 (N_6533,In_4977,In_3235);
or U6534 (N_6534,In_4098,In_2455);
nor U6535 (N_6535,In_1358,In_2097);
nand U6536 (N_6536,In_2870,In_71);
nand U6537 (N_6537,In_574,In_2308);
nor U6538 (N_6538,In_3514,In_855);
nand U6539 (N_6539,In_3779,In_3170);
or U6540 (N_6540,In_3794,In_4028);
xnor U6541 (N_6541,In_1907,In_2536);
or U6542 (N_6542,In_376,In_4374);
xnor U6543 (N_6543,In_4192,In_2967);
nand U6544 (N_6544,In_68,In_4189);
or U6545 (N_6545,In_1825,In_3730);
or U6546 (N_6546,In_2099,In_3787);
nor U6547 (N_6547,In_3512,In_350);
xor U6548 (N_6548,In_3633,In_2670);
nor U6549 (N_6549,In_664,In_3419);
and U6550 (N_6550,In_2887,In_4718);
nand U6551 (N_6551,In_2250,In_944);
xor U6552 (N_6552,In_438,In_3368);
and U6553 (N_6553,In_141,In_4485);
or U6554 (N_6554,In_4462,In_2343);
and U6555 (N_6555,In_3562,In_2910);
nand U6556 (N_6556,In_2109,In_3177);
xor U6557 (N_6557,In_3763,In_525);
xnor U6558 (N_6558,In_3099,In_1135);
nand U6559 (N_6559,In_3776,In_3189);
nor U6560 (N_6560,In_4192,In_2920);
xnor U6561 (N_6561,In_4325,In_1676);
xor U6562 (N_6562,In_408,In_2219);
and U6563 (N_6563,In_3474,In_2502);
nor U6564 (N_6564,In_802,In_3190);
xnor U6565 (N_6565,In_1460,In_4935);
nor U6566 (N_6566,In_3810,In_3911);
or U6567 (N_6567,In_4408,In_4091);
nand U6568 (N_6568,In_372,In_4535);
and U6569 (N_6569,In_4254,In_4405);
and U6570 (N_6570,In_1648,In_2065);
nor U6571 (N_6571,In_1228,In_4049);
nand U6572 (N_6572,In_1175,In_4548);
nor U6573 (N_6573,In_1897,In_4471);
and U6574 (N_6574,In_1486,In_3202);
nor U6575 (N_6575,In_1810,In_321);
and U6576 (N_6576,In_968,In_1068);
and U6577 (N_6577,In_4264,In_4363);
nand U6578 (N_6578,In_2060,In_2308);
nor U6579 (N_6579,In_1605,In_3499);
nand U6580 (N_6580,In_2701,In_2063);
nand U6581 (N_6581,In_1440,In_4067);
nor U6582 (N_6582,In_1578,In_1683);
nor U6583 (N_6583,In_819,In_493);
xnor U6584 (N_6584,In_1349,In_4541);
or U6585 (N_6585,In_382,In_3504);
nor U6586 (N_6586,In_3986,In_2567);
nor U6587 (N_6587,In_1164,In_1586);
and U6588 (N_6588,In_1971,In_4350);
and U6589 (N_6589,In_438,In_1640);
and U6590 (N_6590,In_775,In_4475);
and U6591 (N_6591,In_2783,In_4945);
xor U6592 (N_6592,In_3645,In_2991);
or U6593 (N_6593,In_2400,In_4568);
or U6594 (N_6594,In_990,In_2805);
and U6595 (N_6595,In_3392,In_4525);
nor U6596 (N_6596,In_1656,In_1192);
xor U6597 (N_6597,In_985,In_2570);
and U6598 (N_6598,In_2626,In_1969);
nor U6599 (N_6599,In_2138,In_4945);
nor U6600 (N_6600,In_1357,In_4923);
or U6601 (N_6601,In_1937,In_1542);
nor U6602 (N_6602,In_4266,In_1708);
nor U6603 (N_6603,In_2240,In_1555);
nor U6604 (N_6604,In_1159,In_734);
or U6605 (N_6605,In_2325,In_3779);
and U6606 (N_6606,In_3551,In_1601);
or U6607 (N_6607,In_1039,In_4251);
and U6608 (N_6608,In_146,In_1966);
nand U6609 (N_6609,In_2396,In_828);
nand U6610 (N_6610,In_1314,In_2821);
or U6611 (N_6611,In_575,In_4228);
nand U6612 (N_6612,In_2705,In_4536);
nor U6613 (N_6613,In_3561,In_1800);
nor U6614 (N_6614,In_4907,In_454);
and U6615 (N_6615,In_962,In_3772);
nand U6616 (N_6616,In_898,In_3331);
nor U6617 (N_6617,In_2749,In_2659);
nor U6618 (N_6618,In_4890,In_3040);
and U6619 (N_6619,In_4804,In_1008);
nand U6620 (N_6620,In_1032,In_359);
xnor U6621 (N_6621,In_2792,In_138);
or U6622 (N_6622,In_3773,In_4465);
or U6623 (N_6623,In_4636,In_3007);
and U6624 (N_6624,In_3452,In_2375);
nand U6625 (N_6625,In_969,In_4283);
and U6626 (N_6626,In_1583,In_1057);
or U6627 (N_6627,In_1605,In_4035);
xnor U6628 (N_6628,In_394,In_356);
xor U6629 (N_6629,In_851,In_1183);
or U6630 (N_6630,In_4369,In_865);
xnor U6631 (N_6631,In_2023,In_4531);
or U6632 (N_6632,In_1720,In_960);
or U6633 (N_6633,In_3704,In_1273);
nor U6634 (N_6634,In_3982,In_1913);
nor U6635 (N_6635,In_1773,In_1591);
and U6636 (N_6636,In_2306,In_4805);
xor U6637 (N_6637,In_4716,In_2415);
or U6638 (N_6638,In_1848,In_731);
and U6639 (N_6639,In_2067,In_3255);
nor U6640 (N_6640,In_2607,In_3672);
and U6641 (N_6641,In_1107,In_2234);
or U6642 (N_6642,In_1927,In_3824);
nor U6643 (N_6643,In_237,In_1891);
and U6644 (N_6644,In_370,In_2881);
and U6645 (N_6645,In_1226,In_3618);
nor U6646 (N_6646,In_2180,In_293);
and U6647 (N_6647,In_2886,In_3541);
nand U6648 (N_6648,In_2576,In_3800);
xor U6649 (N_6649,In_626,In_960);
nor U6650 (N_6650,In_413,In_746);
xor U6651 (N_6651,In_3860,In_863);
or U6652 (N_6652,In_4394,In_3616);
and U6653 (N_6653,In_2460,In_3588);
or U6654 (N_6654,In_3109,In_2943);
or U6655 (N_6655,In_4483,In_3163);
nand U6656 (N_6656,In_3337,In_3875);
nand U6657 (N_6657,In_2075,In_4672);
and U6658 (N_6658,In_1894,In_425);
and U6659 (N_6659,In_3947,In_3655);
nor U6660 (N_6660,In_1389,In_2333);
nor U6661 (N_6661,In_1993,In_3924);
and U6662 (N_6662,In_4750,In_524);
and U6663 (N_6663,In_868,In_4384);
or U6664 (N_6664,In_1819,In_1981);
and U6665 (N_6665,In_1477,In_1344);
xnor U6666 (N_6666,In_3380,In_3315);
nor U6667 (N_6667,In_2291,In_159);
nand U6668 (N_6668,In_4313,In_4948);
or U6669 (N_6669,In_3470,In_2723);
or U6670 (N_6670,In_3068,In_2236);
xor U6671 (N_6671,In_2187,In_24);
nor U6672 (N_6672,In_900,In_1684);
nand U6673 (N_6673,In_974,In_3961);
nand U6674 (N_6674,In_3404,In_4263);
or U6675 (N_6675,In_345,In_81);
or U6676 (N_6676,In_2193,In_3245);
or U6677 (N_6677,In_3693,In_1049);
and U6678 (N_6678,In_2388,In_3793);
and U6679 (N_6679,In_1084,In_3937);
or U6680 (N_6680,In_1178,In_3147);
nand U6681 (N_6681,In_3975,In_2705);
nor U6682 (N_6682,In_1638,In_4875);
nand U6683 (N_6683,In_1573,In_796);
nor U6684 (N_6684,In_132,In_2218);
or U6685 (N_6685,In_2454,In_2308);
xor U6686 (N_6686,In_3323,In_2801);
xor U6687 (N_6687,In_1107,In_924);
nand U6688 (N_6688,In_2698,In_1750);
nor U6689 (N_6689,In_1817,In_3340);
nand U6690 (N_6690,In_946,In_3103);
and U6691 (N_6691,In_2966,In_1836);
nor U6692 (N_6692,In_535,In_66);
nand U6693 (N_6693,In_598,In_2470);
nor U6694 (N_6694,In_681,In_4069);
nand U6695 (N_6695,In_2290,In_4871);
nand U6696 (N_6696,In_86,In_1246);
or U6697 (N_6697,In_276,In_3771);
and U6698 (N_6698,In_4018,In_2730);
and U6699 (N_6699,In_1986,In_3615);
and U6700 (N_6700,In_969,In_63);
and U6701 (N_6701,In_3289,In_995);
and U6702 (N_6702,In_2169,In_2342);
nor U6703 (N_6703,In_3487,In_2218);
or U6704 (N_6704,In_2393,In_4605);
or U6705 (N_6705,In_1279,In_2519);
nor U6706 (N_6706,In_1565,In_3420);
or U6707 (N_6707,In_2652,In_2990);
nor U6708 (N_6708,In_412,In_2449);
and U6709 (N_6709,In_4386,In_3582);
nor U6710 (N_6710,In_4579,In_909);
nor U6711 (N_6711,In_1499,In_1124);
nor U6712 (N_6712,In_3587,In_4530);
or U6713 (N_6713,In_2661,In_1654);
nand U6714 (N_6714,In_1747,In_372);
nand U6715 (N_6715,In_234,In_389);
nand U6716 (N_6716,In_3394,In_1554);
nand U6717 (N_6717,In_4088,In_858);
or U6718 (N_6718,In_2356,In_2468);
nand U6719 (N_6719,In_2500,In_961);
nand U6720 (N_6720,In_2711,In_2015);
nor U6721 (N_6721,In_2327,In_1345);
xor U6722 (N_6722,In_2217,In_2923);
nor U6723 (N_6723,In_3997,In_4787);
and U6724 (N_6724,In_3342,In_2699);
nor U6725 (N_6725,In_3037,In_3624);
or U6726 (N_6726,In_1212,In_1180);
nor U6727 (N_6727,In_4531,In_3032);
or U6728 (N_6728,In_2513,In_3040);
nor U6729 (N_6729,In_735,In_574);
nand U6730 (N_6730,In_1384,In_4625);
or U6731 (N_6731,In_1037,In_2149);
or U6732 (N_6732,In_1963,In_3268);
or U6733 (N_6733,In_3702,In_573);
and U6734 (N_6734,In_444,In_1752);
nor U6735 (N_6735,In_4914,In_717);
xnor U6736 (N_6736,In_245,In_4441);
nor U6737 (N_6737,In_2194,In_3609);
and U6738 (N_6738,In_1383,In_665);
xnor U6739 (N_6739,In_3295,In_1970);
or U6740 (N_6740,In_2115,In_2371);
nor U6741 (N_6741,In_17,In_1964);
and U6742 (N_6742,In_4341,In_4607);
nor U6743 (N_6743,In_92,In_3150);
or U6744 (N_6744,In_168,In_26);
nor U6745 (N_6745,In_1926,In_1962);
xor U6746 (N_6746,In_2992,In_4601);
or U6747 (N_6747,In_1813,In_3962);
nand U6748 (N_6748,In_4464,In_3231);
xnor U6749 (N_6749,In_1066,In_4504);
nand U6750 (N_6750,In_4217,In_2328);
or U6751 (N_6751,In_1839,In_952);
nor U6752 (N_6752,In_1505,In_1720);
nor U6753 (N_6753,In_4787,In_230);
and U6754 (N_6754,In_646,In_2074);
and U6755 (N_6755,In_2745,In_2593);
nand U6756 (N_6756,In_2218,In_2264);
and U6757 (N_6757,In_4002,In_3383);
or U6758 (N_6758,In_1324,In_79);
and U6759 (N_6759,In_138,In_4128);
or U6760 (N_6760,In_4645,In_4069);
nand U6761 (N_6761,In_1169,In_4133);
and U6762 (N_6762,In_435,In_3860);
nand U6763 (N_6763,In_4862,In_2257);
nor U6764 (N_6764,In_724,In_1058);
or U6765 (N_6765,In_3642,In_3026);
nor U6766 (N_6766,In_3595,In_531);
and U6767 (N_6767,In_4786,In_1124);
and U6768 (N_6768,In_2336,In_3122);
nor U6769 (N_6769,In_3244,In_3251);
nor U6770 (N_6770,In_2389,In_953);
nand U6771 (N_6771,In_3095,In_3463);
xor U6772 (N_6772,In_4764,In_3683);
nor U6773 (N_6773,In_3560,In_3910);
or U6774 (N_6774,In_3839,In_2997);
nand U6775 (N_6775,In_2605,In_1394);
or U6776 (N_6776,In_4175,In_4737);
nor U6777 (N_6777,In_3145,In_4740);
or U6778 (N_6778,In_2385,In_790);
nor U6779 (N_6779,In_146,In_3027);
or U6780 (N_6780,In_112,In_1872);
and U6781 (N_6781,In_2494,In_4439);
and U6782 (N_6782,In_1568,In_3033);
and U6783 (N_6783,In_1272,In_3434);
xor U6784 (N_6784,In_959,In_1703);
nand U6785 (N_6785,In_3353,In_2794);
and U6786 (N_6786,In_4820,In_4689);
or U6787 (N_6787,In_2345,In_4048);
nor U6788 (N_6788,In_3789,In_1929);
nor U6789 (N_6789,In_1534,In_2986);
or U6790 (N_6790,In_2064,In_1027);
nand U6791 (N_6791,In_3711,In_4754);
nand U6792 (N_6792,In_1075,In_2803);
nand U6793 (N_6793,In_2968,In_23);
xor U6794 (N_6794,In_2696,In_660);
nand U6795 (N_6795,In_121,In_1805);
or U6796 (N_6796,In_2851,In_4609);
nor U6797 (N_6797,In_126,In_1066);
or U6798 (N_6798,In_528,In_2706);
nor U6799 (N_6799,In_4228,In_1073);
or U6800 (N_6800,In_1896,In_2050);
and U6801 (N_6801,In_1705,In_2531);
xor U6802 (N_6802,In_1941,In_4512);
and U6803 (N_6803,In_1644,In_2568);
and U6804 (N_6804,In_1860,In_3941);
nand U6805 (N_6805,In_2810,In_3613);
nor U6806 (N_6806,In_4361,In_2655);
and U6807 (N_6807,In_1342,In_1441);
xor U6808 (N_6808,In_91,In_353);
nor U6809 (N_6809,In_4292,In_3434);
or U6810 (N_6810,In_2280,In_2419);
or U6811 (N_6811,In_4967,In_1247);
nor U6812 (N_6812,In_4934,In_488);
xor U6813 (N_6813,In_1688,In_3162);
or U6814 (N_6814,In_395,In_996);
nand U6815 (N_6815,In_4603,In_4286);
or U6816 (N_6816,In_2034,In_4478);
and U6817 (N_6817,In_1095,In_4179);
nand U6818 (N_6818,In_267,In_1443);
nand U6819 (N_6819,In_2074,In_116);
or U6820 (N_6820,In_17,In_566);
or U6821 (N_6821,In_3358,In_1885);
nand U6822 (N_6822,In_1320,In_3301);
or U6823 (N_6823,In_2294,In_2428);
nand U6824 (N_6824,In_2957,In_270);
and U6825 (N_6825,In_739,In_2512);
or U6826 (N_6826,In_2735,In_3813);
xor U6827 (N_6827,In_4868,In_2635);
nand U6828 (N_6828,In_107,In_2045);
or U6829 (N_6829,In_2368,In_1451);
nand U6830 (N_6830,In_3695,In_1492);
nand U6831 (N_6831,In_223,In_3807);
and U6832 (N_6832,In_874,In_1940);
xor U6833 (N_6833,In_3069,In_1713);
xnor U6834 (N_6834,In_4206,In_2702);
or U6835 (N_6835,In_4365,In_46);
or U6836 (N_6836,In_710,In_317);
xnor U6837 (N_6837,In_4122,In_3320);
nand U6838 (N_6838,In_2540,In_2959);
or U6839 (N_6839,In_4717,In_4920);
or U6840 (N_6840,In_1909,In_2862);
or U6841 (N_6841,In_1845,In_1713);
and U6842 (N_6842,In_3572,In_1959);
xor U6843 (N_6843,In_2365,In_2664);
nand U6844 (N_6844,In_970,In_1246);
and U6845 (N_6845,In_282,In_3191);
xor U6846 (N_6846,In_889,In_191);
or U6847 (N_6847,In_2273,In_2462);
and U6848 (N_6848,In_3376,In_4360);
nor U6849 (N_6849,In_3849,In_862);
nor U6850 (N_6850,In_2509,In_2995);
xnor U6851 (N_6851,In_4811,In_4161);
and U6852 (N_6852,In_3660,In_592);
nand U6853 (N_6853,In_4740,In_671);
or U6854 (N_6854,In_4440,In_4732);
xnor U6855 (N_6855,In_3449,In_1388);
nor U6856 (N_6856,In_3562,In_2052);
or U6857 (N_6857,In_1049,In_1523);
and U6858 (N_6858,In_4394,In_1945);
and U6859 (N_6859,In_1783,In_2998);
or U6860 (N_6860,In_1934,In_161);
or U6861 (N_6861,In_1551,In_105);
xor U6862 (N_6862,In_2385,In_1552);
or U6863 (N_6863,In_4688,In_4740);
or U6864 (N_6864,In_2019,In_4353);
nand U6865 (N_6865,In_3647,In_3619);
or U6866 (N_6866,In_1283,In_2017);
and U6867 (N_6867,In_663,In_4284);
nand U6868 (N_6868,In_4242,In_4406);
nor U6869 (N_6869,In_3995,In_227);
xnor U6870 (N_6870,In_4516,In_4835);
and U6871 (N_6871,In_2854,In_1124);
nand U6872 (N_6872,In_1390,In_2813);
nand U6873 (N_6873,In_2893,In_3763);
nor U6874 (N_6874,In_1529,In_4386);
nor U6875 (N_6875,In_4927,In_2460);
or U6876 (N_6876,In_1469,In_2033);
or U6877 (N_6877,In_4561,In_4995);
and U6878 (N_6878,In_3904,In_2670);
xor U6879 (N_6879,In_3468,In_4726);
nor U6880 (N_6880,In_1798,In_1305);
or U6881 (N_6881,In_3606,In_965);
or U6882 (N_6882,In_4825,In_3284);
xor U6883 (N_6883,In_1064,In_1673);
and U6884 (N_6884,In_1023,In_3376);
nand U6885 (N_6885,In_2633,In_2285);
nand U6886 (N_6886,In_4244,In_1739);
and U6887 (N_6887,In_1783,In_3434);
or U6888 (N_6888,In_2852,In_3679);
nor U6889 (N_6889,In_272,In_4352);
and U6890 (N_6890,In_3210,In_2392);
or U6891 (N_6891,In_618,In_4606);
and U6892 (N_6892,In_2004,In_270);
xor U6893 (N_6893,In_3511,In_3637);
xnor U6894 (N_6894,In_2379,In_2838);
or U6895 (N_6895,In_520,In_2762);
nand U6896 (N_6896,In_1126,In_1471);
and U6897 (N_6897,In_4830,In_1200);
nand U6898 (N_6898,In_50,In_481);
or U6899 (N_6899,In_511,In_3870);
or U6900 (N_6900,In_1868,In_4716);
and U6901 (N_6901,In_3492,In_1038);
or U6902 (N_6902,In_4281,In_4800);
or U6903 (N_6903,In_4674,In_4367);
nand U6904 (N_6904,In_2709,In_1227);
nor U6905 (N_6905,In_1074,In_3860);
or U6906 (N_6906,In_1722,In_3679);
nor U6907 (N_6907,In_4221,In_1282);
and U6908 (N_6908,In_604,In_901);
nor U6909 (N_6909,In_3190,In_4922);
nor U6910 (N_6910,In_4322,In_3601);
and U6911 (N_6911,In_3158,In_3977);
nand U6912 (N_6912,In_4213,In_2516);
nor U6913 (N_6913,In_2805,In_3663);
nand U6914 (N_6914,In_2955,In_2291);
nand U6915 (N_6915,In_2119,In_2480);
or U6916 (N_6916,In_2168,In_446);
or U6917 (N_6917,In_781,In_2392);
nand U6918 (N_6918,In_1994,In_2678);
or U6919 (N_6919,In_2397,In_1429);
or U6920 (N_6920,In_1198,In_2442);
nor U6921 (N_6921,In_4950,In_2411);
and U6922 (N_6922,In_1172,In_941);
and U6923 (N_6923,In_4774,In_4702);
and U6924 (N_6924,In_468,In_3632);
or U6925 (N_6925,In_3689,In_1129);
nor U6926 (N_6926,In_3845,In_3055);
or U6927 (N_6927,In_857,In_3084);
xor U6928 (N_6928,In_1859,In_2105);
and U6929 (N_6929,In_1842,In_4207);
xor U6930 (N_6930,In_1014,In_1627);
nand U6931 (N_6931,In_2472,In_517);
or U6932 (N_6932,In_2616,In_1960);
nor U6933 (N_6933,In_314,In_2507);
nor U6934 (N_6934,In_4500,In_4988);
and U6935 (N_6935,In_3682,In_4385);
and U6936 (N_6936,In_2511,In_2683);
or U6937 (N_6937,In_1269,In_817);
xnor U6938 (N_6938,In_3966,In_1093);
and U6939 (N_6939,In_3834,In_1168);
nor U6940 (N_6940,In_4885,In_4912);
nand U6941 (N_6941,In_234,In_3124);
nor U6942 (N_6942,In_4396,In_3687);
nor U6943 (N_6943,In_3663,In_1713);
nand U6944 (N_6944,In_2045,In_398);
and U6945 (N_6945,In_308,In_990);
or U6946 (N_6946,In_3416,In_3011);
nand U6947 (N_6947,In_3060,In_3801);
or U6948 (N_6948,In_4757,In_2487);
xor U6949 (N_6949,In_453,In_4178);
or U6950 (N_6950,In_3743,In_2757);
and U6951 (N_6951,In_1217,In_4319);
or U6952 (N_6952,In_3708,In_434);
nor U6953 (N_6953,In_2217,In_4852);
and U6954 (N_6954,In_3110,In_3646);
and U6955 (N_6955,In_157,In_4711);
nand U6956 (N_6956,In_4034,In_3183);
or U6957 (N_6957,In_4969,In_997);
xnor U6958 (N_6958,In_1503,In_2704);
nor U6959 (N_6959,In_3857,In_1319);
nor U6960 (N_6960,In_2033,In_4979);
and U6961 (N_6961,In_2520,In_1422);
and U6962 (N_6962,In_2261,In_3187);
xor U6963 (N_6963,In_3829,In_3272);
and U6964 (N_6964,In_2934,In_2813);
and U6965 (N_6965,In_959,In_2259);
nand U6966 (N_6966,In_4377,In_1948);
xor U6967 (N_6967,In_3229,In_98);
nor U6968 (N_6968,In_4042,In_3353);
nor U6969 (N_6969,In_634,In_2394);
or U6970 (N_6970,In_4002,In_4011);
or U6971 (N_6971,In_2325,In_1729);
or U6972 (N_6972,In_3551,In_164);
nand U6973 (N_6973,In_3706,In_2901);
nor U6974 (N_6974,In_1733,In_278);
or U6975 (N_6975,In_4828,In_380);
nor U6976 (N_6976,In_2241,In_646);
and U6977 (N_6977,In_4957,In_4183);
and U6978 (N_6978,In_2848,In_823);
nor U6979 (N_6979,In_3790,In_3302);
and U6980 (N_6980,In_3828,In_1356);
nand U6981 (N_6981,In_4837,In_1235);
nor U6982 (N_6982,In_4099,In_4811);
nand U6983 (N_6983,In_6,In_704);
or U6984 (N_6984,In_2245,In_1003);
or U6985 (N_6985,In_4973,In_3832);
nor U6986 (N_6986,In_2000,In_267);
and U6987 (N_6987,In_3811,In_1662);
nor U6988 (N_6988,In_3381,In_4625);
or U6989 (N_6989,In_909,In_3775);
nand U6990 (N_6990,In_4331,In_4497);
or U6991 (N_6991,In_3521,In_4335);
nand U6992 (N_6992,In_1788,In_3960);
xnor U6993 (N_6993,In_4661,In_3136);
nand U6994 (N_6994,In_1152,In_2491);
nand U6995 (N_6995,In_3812,In_2174);
nand U6996 (N_6996,In_1136,In_977);
or U6997 (N_6997,In_2776,In_4312);
and U6998 (N_6998,In_3920,In_4880);
and U6999 (N_6999,In_125,In_1392);
xor U7000 (N_7000,In_2224,In_924);
or U7001 (N_7001,In_2076,In_4724);
nor U7002 (N_7002,In_3530,In_785);
or U7003 (N_7003,In_3889,In_3199);
xor U7004 (N_7004,In_2239,In_3595);
and U7005 (N_7005,In_1852,In_2295);
or U7006 (N_7006,In_2516,In_614);
nand U7007 (N_7007,In_3757,In_1309);
and U7008 (N_7008,In_77,In_4983);
and U7009 (N_7009,In_2726,In_4700);
nand U7010 (N_7010,In_2877,In_1476);
and U7011 (N_7011,In_415,In_834);
nand U7012 (N_7012,In_3550,In_3319);
and U7013 (N_7013,In_3766,In_4577);
xnor U7014 (N_7014,In_4797,In_4302);
or U7015 (N_7015,In_876,In_3928);
nor U7016 (N_7016,In_2876,In_1530);
and U7017 (N_7017,In_3032,In_1638);
and U7018 (N_7018,In_3879,In_416);
xnor U7019 (N_7019,In_559,In_2760);
nor U7020 (N_7020,In_4851,In_523);
nand U7021 (N_7021,In_1,In_593);
and U7022 (N_7022,In_2879,In_1149);
and U7023 (N_7023,In_3225,In_1207);
nor U7024 (N_7024,In_2650,In_3136);
nand U7025 (N_7025,In_4115,In_3160);
nand U7026 (N_7026,In_2407,In_2765);
nor U7027 (N_7027,In_1101,In_158);
nand U7028 (N_7028,In_4141,In_640);
nand U7029 (N_7029,In_4187,In_620);
or U7030 (N_7030,In_2871,In_4553);
nor U7031 (N_7031,In_3315,In_3083);
nor U7032 (N_7032,In_2842,In_364);
nand U7033 (N_7033,In_2710,In_4207);
and U7034 (N_7034,In_4399,In_3757);
nor U7035 (N_7035,In_2859,In_4849);
nor U7036 (N_7036,In_415,In_2876);
nand U7037 (N_7037,In_467,In_3094);
and U7038 (N_7038,In_3847,In_4937);
nand U7039 (N_7039,In_1498,In_3064);
nor U7040 (N_7040,In_1757,In_1726);
nand U7041 (N_7041,In_3673,In_2850);
and U7042 (N_7042,In_2845,In_2109);
and U7043 (N_7043,In_4709,In_2338);
nand U7044 (N_7044,In_4536,In_135);
or U7045 (N_7045,In_786,In_2527);
or U7046 (N_7046,In_2718,In_505);
and U7047 (N_7047,In_1267,In_4875);
xnor U7048 (N_7048,In_1907,In_2346);
nor U7049 (N_7049,In_3593,In_2210);
or U7050 (N_7050,In_4390,In_2460);
xnor U7051 (N_7051,In_4058,In_4402);
or U7052 (N_7052,In_514,In_728);
nor U7053 (N_7053,In_2562,In_1062);
nand U7054 (N_7054,In_888,In_2913);
nand U7055 (N_7055,In_4259,In_3265);
and U7056 (N_7056,In_637,In_3406);
nor U7057 (N_7057,In_347,In_3250);
nor U7058 (N_7058,In_51,In_3363);
nor U7059 (N_7059,In_1679,In_2170);
nand U7060 (N_7060,In_172,In_201);
nand U7061 (N_7061,In_608,In_1145);
or U7062 (N_7062,In_4102,In_3890);
or U7063 (N_7063,In_1305,In_3567);
or U7064 (N_7064,In_2197,In_3548);
nand U7065 (N_7065,In_1556,In_1218);
xor U7066 (N_7066,In_229,In_298);
nand U7067 (N_7067,In_2904,In_1183);
or U7068 (N_7068,In_3338,In_4546);
nand U7069 (N_7069,In_3308,In_4441);
nor U7070 (N_7070,In_673,In_2654);
nand U7071 (N_7071,In_4212,In_475);
nand U7072 (N_7072,In_1324,In_2028);
and U7073 (N_7073,In_1434,In_65);
nor U7074 (N_7074,In_903,In_3764);
xor U7075 (N_7075,In_4723,In_289);
or U7076 (N_7076,In_3856,In_4973);
and U7077 (N_7077,In_1943,In_2507);
or U7078 (N_7078,In_3082,In_3838);
and U7079 (N_7079,In_4227,In_3375);
nand U7080 (N_7080,In_169,In_2060);
nand U7081 (N_7081,In_370,In_330);
nand U7082 (N_7082,In_3263,In_1095);
nor U7083 (N_7083,In_1548,In_2057);
nand U7084 (N_7084,In_3736,In_4616);
xnor U7085 (N_7085,In_1196,In_4720);
nor U7086 (N_7086,In_4548,In_2393);
or U7087 (N_7087,In_2923,In_2255);
nand U7088 (N_7088,In_232,In_671);
or U7089 (N_7089,In_1469,In_2307);
or U7090 (N_7090,In_4968,In_1517);
and U7091 (N_7091,In_3200,In_4560);
nor U7092 (N_7092,In_2505,In_1649);
or U7093 (N_7093,In_997,In_312);
or U7094 (N_7094,In_3068,In_1579);
nand U7095 (N_7095,In_2795,In_1112);
nand U7096 (N_7096,In_3298,In_3737);
and U7097 (N_7097,In_4486,In_4054);
nand U7098 (N_7098,In_3298,In_4074);
or U7099 (N_7099,In_3476,In_3767);
or U7100 (N_7100,In_1514,In_409);
nand U7101 (N_7101,In_1427,In_2899);
or U7102 (N_7102,In_3791,In_3251);
nand U7103 (N_7103,In_4098,In_3786);
or U7104 (N_7104,In_4707,In_3811);
or U7105 (N_7105,In_3812,In_897);
nand U7106 (N_7106,In_38,In_3031);
or U7107 (N_7107,In_512,In_351);
nand U7108 (N_7108,In_3225,In_1076);
nor U7109 (N_7109,In_3007,In_4059);
nand U7110 (N_7110,In_4175,In_2631);
xnor U7111 (N_7111,In_1091,In_3797);
xnor U7112 (N_7112,In_3323,In_2963);
or U7113 (N_7113,In_2850,In_3904);
nand U7114 (N_7114,In_268,In_4247);
nand U7115 (N_7115,In_4974,In_3709);
nand U7116 (N_7116,In_1101,In_2320);
and U7117 (N_7117,In_2232,In_1483);
nor U7118 (N_7118,In_3402,In_2298);
or U7119 (N_7119,In_4891,In_591);
nor U7120 (N_7120,In_1463,In_4254);
nand U7121 (N_7121,In_1395,In_3962);
nand U7122 (N_7122,In_130,In_3367);
nor U7123 (N_7123,In_4554,In_2209);
or U7124 (N_7124,In_4303,In_1774);
and U7125 (N_7125,In_1207,In_4625);
or U7126 (N_7126,In_2481,In_3917);
and U7127 (N_7127,In_2352,In_913);
and U7128 (N_7128,In_475,In_2957);
xnor U7129 (N_7129,In_3366,In_422);
nor U7130 (N_7130,In_2227,In_487);
xnor U7131 (N_7131,In_3070,In_531);
nand U7132 (N_7132,In_1138,In_1665);
xor U7133 (N_7133,In_755,In_3679);
nand U7134 (N_7134,In_3482,In_2664);
xnor U7135 (N_7135,In_3478,In_3329);
or U7136 (N_7136,In_757,In_1860);
and U7137 (N_7137,In_3687,In_2948);
and U7138 (N_7138,In_3775,In_1722);
and U7139 (N_7139,In_4651,In_2220);
nand U7140 (N_7140,In_2974,In_4365);
nand U7141 (N_7141,In_1969,In_2233);
nor U7142 (N_7142,In_1540,In_27);
xor U7143 (N_7143,In_1487,In_1513);
nand U7144 (N_7144,In_984,In_2581);
and U7145 (N_7145,In_701,In_1638);
xnor U7146 (N_7146,In_2133,In_2780);
and U7147 (N_7147,In_742,In_1761);
and U7148 (N_7148,In_808,In_3688);
or U7149 (N_7149,In_4507,In_1684);
or U7150 (N_7150,In_4352,In_242);
and U7151 (N_7151,In_2718,In_4335);
or U7152 (N_7152,In_3697,In_1168);
nand U7153 (N_7153,In_3513,In_1551);
and U7154 (N_7154,In_3489,In_2751);
and U7155 (N_7155,In_1610,In_3341);
or U7156 (N_7156,In_4921,In_2701);
or U7157 (N_7157,In_2626,In_905);
and U7158 (N_7158,In_1883,In_1000);
xnor U7159 (N_7159,In_360,In_1495);
or U7160 (N_7160,In_2062,In_3541);
and U7161 (N_7161,In_4877,In_4909);
nand U7162 (N_7162,In_2013,In_2092);
or U7163 (N_7163,In_175,In_4098);
and U7164 (N_7164,In_3112,In_3395);
and U7165 (N_7165,In_1180,In_3517);
and U7166 (N_7166,In_1949,In_418);
or U7167 (N_7167,In_1112,In_4278);
and U7168 (N_7168,In_1740,In_3456);
nor U7169 (N_7169,In_4029,In_4177);
nand U7170 (N_7170,In_4904,In_3082);
or U7171 (N_7171,In_4808,In_1984);
nand U7172 (N_7172,In_3138,In_3931);
nand U7173 (N_7173,In_4293,In_3763);
nor U7174 (N_7174,In_1122,In_3247);
nand U7175 (N_7175,In_4092,In_715);
nor U7176 (N_7176,In_4816,In_2573);
and U7177 (N_7177,In_3822,In_1855);
or U7178 (N_7178,In_3639,In_355);
nand U7179 (N_7179,In_1324,In_4336);
nand U7180 (N_7180,In_3981,In_1627);
or U7181 (N_7181,In_2627,In_2346);
nor U7182 (N_7182,In_3427,In_4210);
and U7183 (N_7183,In_3433,In_1640);
nand U7184 (N_7184,In_405,In_3382);
nand U7185 (N_7185,In_1253,In_1331);
nor U7186 (N_7186,In_2346,In_1790);
nand U7187 (N_7187,In_4350,In_3504);
nor U7188 (N_7188,In_4088,In_2989);
nand U7189 (N_7189,In_3744,In_494);
nor U7190 (N_7190,In_3803,In_4942);
or U7191 (N_7191,In_2551,In_1820);
or U7192 (N_7192,In_4524,In_500);
nor U7193 (N_7193,In_179,In_4059);
and U7194 (N_7194,In_1848,In_2689);
nor U7195 (N_7195,In_2287,In_1498);
or U7196 (N_7196,In_2538,In_943);
and U7197 (N_7197,In_4771,In_3983);
or U7198 (N_7198,In_1971,In_3406);
nand U7199 (N_7199,In_495,In_2463);
and U7200 (N_7200,In_212,In_1648);
and U7201 (N_7201,In_4290,In_2130);
xnor U7202 (N_7202,In_1347,In_3814);
xnor U7203 (N_7203,In_4541,In_190);
and U7204 (N_7204,In_728,In_4424);
nor U7205 (N_7205,In_4789,In_688);
or U7206 (N_7206,In_1162,In_282);
nor U7207 (N_7207,In_1894,In_739);
or U7208 (N_7208,In_4854,In_4744);
nor U7209 (N_7209,In_521,In_3335);
or U7210 (N_7210,In_2784,In_4932);
and U7211 (N_7211,In_3,In_4711);
nor U7212 (N_7212,In_2337,In_1536);
or U7213 (N_7213,In_2909,In_1701);
nor U7214 (N_7214,In_890,In_3074);
nor U7215 (N_7215,In_3173,In_1319);
or U7216 (N_7216,In_1520,In_1062);
xor U7217 (N_7217,In_1085,In_3725);
nand U7218 (N_7218,In_4572,In_4437);
or U7219 (N_7219,In_4389,In_2826);
and U7220 (N_7220,In_1573,In_2371);
or U7221 (N_7221,In_286,In_44);
and U7222 (N_7222,In_425,In_4643);
or U7223 (N_7223,In_2595,In_972);
nor U7224 (N_7224,In_3002,In_4274);
and U7225 (N_7225,In_4103,In_2287);
nor U7226 (N_7226,In_814,In_1774);
or U7227 (N_7227,In_1005,In_2156);
and U7228 (N_7228,In_703,In_2592);
xnor U7229 (N_7229,In_1250,In_4774);
nor U7230 (N_7230,In_1014,In_1354);
and U7231 (N_7231,In_2825,In_1468);
or U7232 (N_7232,In_3139,In_1049);
and U7233 (N_7233,In_2736,In_951);
or U7234 (N_7234,In_4521,In_1597);
nand U7235 (N_7235,In_3527,In_3248);
nor U7236 (N_7236,In_4527,In_2912);
and U7237 (N_7237,In_4277,In_1449);
and U7238 (N_7238,In_885,In_751);
and U7239 (N_7239,In_1360,In_3795);
nor U7240 (N_7240,In_4546,In_1663);
nor U7241 (N_7241,In_650,In_2405);
and U7242 (N_7242,In_1415,In_555);
and U7243 (N_7243,In_4080,In_2549);
or U7244 (N_7244,In_1467,In_1069);
or U7245 (N_7245,In_927,In_1995);
nand U7246 (N_7246,In_2422,In_764);
xnor U7247 (N_7247,In_4933,In_1566);
and U7248 (N_7248,In_4422,In_4647);
nor U7249 (N_7249,In_4934,In_2559);
nand U7250 (N_7250,In_3819,In_422);
and U7251 (N_7251,In_1517,In_2187);
or U7252 (N_7252,In_1868,In_3817);
nor U7253 (N_7253,In_4095,In_3139);
and U7254 (N_7254,In_4552,In_1577);
nand U7255 (N_7255,In_4466,In_4326);
or U7256 (N_7256,In_1018,In_4838);
or U7257 (N_7257,In_464,In_3115);
or U7258 (N_7258,In_3335,In_4635);
nand U7259 (N_7259,In_4063,In_4777);
nor U7260 (N_7260,In_1023,In_2711);
or U7261 (N_7261,In_1054,In_199);
or U7262 (N_7262,In_4424,In_2941);
nand U7263 (N_7263,In_485,In_2112);
nand U7264 (N_7264,In_2002,In_1562);
or U7265 (N_7265,In_4358,In_2311);
nand U7266 (N_7266,In_3098,In_1649);
nor U7267 (N_7267,In_487,In_2242);
nand U7268 (N_7268,In_2157,In_890);
nor U7269 (N_7269,In_4072,In_4535);
and U7270 (N_7270,In_4847,In_3992);
and U7271 (N_7271,In_1694,In_2373);
and U7272 (N_7272,In_4361,In_3975);
or U7273 (N_7273,In_2956,In_2855);
nor U7274 (N_7274,In_4051,In_1125);
nand U7275 (N_7275,In_2643,In_579);
nor U7276 (N_7276,In_4997,In_3687);
and U7277 (N_7277,In_3718,In_1443);
and U7278 (N_7278,In_3151,In_1449);
and U7279 (N_7279,In_3035,In_1741);
or U7280 (N_7280,In_2798,In_3992);
and U7281 (N_7281,In_3279,In_4918);
nor U7282 (N_7282,In_471,In_564);
nor U7283 (N_7283,In_156,In_3957);
or U7284 (N_7284,In_4448,In_3315);
nand U7285 (N_7285,In_2667,In_2066);
or U7286 (N_7286,In_47,In_3103);
and U7287 (N_7287,In_4022,In_970);
nor U7288 (N_7288,In_2797,In_3045);
nand U7289 (N_7289,In_348,In_1933);
or U7290 (N_7290,In_112,In_3646);
nor U7291 (N_7291,In_3523,In_4162);
or U7292 (N_7292,In_3473,In_2925);
and U7293 (N_7293,In_2062,In_4209);
nand U7294 (N_7294,In_795,In_1430);
nand U7295 (N_7295,In_1572,In_2916);
and U7296 (N_7296,In_4378,In_962);
and U7297 (N_7297,In_530,In_2875);
and U7298 (N_7298,In_2731,In_177);
nand U7299 (N_7299,In_1041,In_2487);
nand U7300 (N_7300,In_1117,In_1371);
and U7301 (N_7301,In_559,In_1477);
nand U7302 (N_7302,In_11,In_2214);
nand U7303 (N_7303,In_4885,In_661);
and U7304 (N_7304,In_2393,In_4976);
or U7305 (N_7305,In_1482,In_1804);
nor U7306 (N_7306,In_4795,In_2529);
and U7307 (N_7307,In_615,In_61);
xnor U7308 (N_7308,In_4556,In_1134);
nand U7309 (N_7309,In_1234,In_3596);
nor U7310 (N_7310,In_3010,In_460);
and U7311 (N_7311,In_997,In_1964);
nand U7312 (N_7312,In_2091,In_1090);
nand U7313 (N_7313,In_1889,In_4270);
and U7314 (N_7314,In_850,In_3517);
or U7315 (N_7315,In_343,In_4950);
and U7316 (N_7316,In_678,In_3320);
xnor U7317 (N_7317,In_3680,In_10);
or U7318 (N_7318,In_3255,In_1354);
or U7319 (N_7319,In_1828,In_116);
nand U7320 (N_7320,In_537,In_3886);
or U7321 (N_7321,In_3770,In_4801);
nor U7322 (N_7322,In_3571,In_2817);
xnor U7323 (N_7323,In_1938,In_1111);
nand U7324 (N_7324,In_1144,In_4416);
or U7325 (N_7325,In_1432,In_2592);
nand U7326 (N_7326,In_2712,In_854);
nand U7327 (N_7327,In_1312,In_2357);
nand U7328 (N_7328,In_729,In_1307);
xor U7329 (N_7329,In_4837,In_2706);
nor U7330 (N_7330,In_1975,In_40);
and U7331 (N_7331,In_2225,In_1141);
or U7332 (N_7332,In_2700,In_4812);
nor U7333 (N_7333,In_1048,In_1816);
or U7334 (N_7334,In_940,In_1498);
nand U7335 (N_7335,In_729,In_4153);
xnor U7336 (N_7336,In_1488,In_1340);
and U7337 (N_7337,In_4585,In_3844);
xor U7338 (N_7338,In_4327,In_3700);
and U7339 (N_7339,In_326,In_4116);
nand U7340 (N_7340,In_1586,In_2790);
or U7341 (N_7341,In_2764,In_524);
and U7342 (N_7342,In_3589,In_693);
or U7343 (N_7343,In_1195,In_3308);
and U7344 (N_7344,In_2199,In_4677);
nand U7345 (N_7345,In_1684,In_565);
or U7346 (N_7346,In_1853,In_1747);
and U7347 (N_7347,In_1760,In_224);
nor U7348 (N_7348,In_2713,In_1792);
nor U7349 (N_7349,In_46,In_2477);
and U7350 (N_7350,In_1932,In_1797);
nand U7351 (N_7351,In_1302,In_2684);
nand U7352 (N_7352,In_3277,In_845);
nor U7353 (N_7353,In_456,In_1220);
nand U7354 (N_7354,In_2626,In_3034);
xor U7355 (N_7355,In_534,In_1044);
or U7356 (N_7356,In_1731,In_3468);
nand U7357 (N_7357,In_71,In_3268);
or U7358 (N_7358,In_585,In_2859);
nand U7359 (N_7359,In_227,In_2445);
and U7360 (N_7360,In_3485,In_94);
or U7361 (N_7361,In_3046,In_1083);
and U7362 (N_7362,In_22,In_3792);
nor U7363 (N_7363,In_2237,In_3612);
nand U7364 (N_7364,In_4067,In_910);
xor U7365 (N_7365,In_374,In_1020);
and U7366 (N_7366,In_1944,In_1994);
and U7367 (N_7367,In_930,In_3955);
nor U7368 (N_7368,In_4208,In_4689);
and U7369 (N_7369,In_1839,In_4964);
and U7370 (N_7370,In_2918,In_733);
or U7371 (N_7371,In_2707,In_3619);
nor U7372 (N_7372,In_1645,In_2261);
or U7373 (N_7373,In_1567,In_955);
nand U7374 (N_7374,In_4657,In_1610);
nand U7375 (N_7375,In_2795,In_3251);
xnor U7376 (N_7376,In_2617,In_802);
xor U7377 (N_7377,In_917,In_2724);
or U7378 (N_7378,In_1678,In_3318);
nand U7379 (N_7379,In_4456,In_3125);
and U7380 (N_7380,In_3365,In_4888);
nand U7381 (N_7381,In_4181,In_1492);
and U7382 (N_7382,In_891,In_21);
or U7383 (N_7383,In_1565,In_2798);
nand U7384 (N_7384,In_405,In_4045);
nor U7385 (N_7385,In_4058,In_1814);
nor U7386 (N_7386,In_3686,In_4069);
or U7387 (N_7387,In_2823,In_2142);
nor U7388 (N_7388,In_4688,In_1730);
xnor U7389 (N_7389,In_3081,In_1180);
and U7390 (N_7390,In_3853,In_54);
or U7391 (N_7391,In_2642,In_3162);
and U7392 (N_7392,In_2120,In_1313);
or U7393 (N_7393,In_3604,In_1811);
and U7394 (N_7394,In_2195,In_4354);
nand U7395 (N_7395,In_1340,In_1432);
nor U7396 (N_7396,In_920,In_1788);
xnor U7397 (N_7397,In_3836,In_3265);
and U7398 (N_7398,In_4609,In_4464);
nand U7399 (N_7399,In_4117,In_2202);
or U7400 (N_7400,In_3230,In_3917);
nand U7401 (N_7401,In_1275,In_1003);
and U7402 (N_7402,In_4607,In_3087);
nor U7403 (N_7403,In_1561,In_3167);
or U7404 (N_7404,In_828,In_1698);
nand U7405 (N_7405,In_1693,In_3751);
nand U7406 (N_7406,In_2497,In_3615);
xnor U7407 (N_7407,In_850,In_1564);
and U7408 (N_7408,In_2763,In_4476);
or U7409 (N_7409,In_68,In_4015);
or U7410 (N_7410,In_291,In_2579);
nand U7411 (N_7411,In_322,In_1965);
and U7412 (N_7412,In_1835,In_1108);
nand U7413 (N_7413,In_413,In_1088);
and U7414 (N_7414,In_4146,In_2332);
nor U7415 (N_7415,In_217,In_472);
nor U7416 (N_7416,In_2322,In_545);
nor U7417 (N_7417,In_2694,In_3909);
and U7418 (N_7418,In_1816,In_4396);
and U7419 (N_7419,In_2785,In_1657);
nor U7420 (N_7420,In_2994,In_4902);
nand U7421 (N_7421,In_81,In_4193);
xnor U7422 (N_7422,In_3968,In_2289);
nor U7423 (N_7423,In_3561,In_1962);
nor U7424 (N_7424,In_4278,In_1919);
and U7425 (N_7425,In_1140,In_3088);
nor U7426 (N_7426,In_3198,In_3090);
or U7427 (N_7427,In_2101,In_1550);
nand U7428 (N_7428,In_1350,In_3855);
nor U7429 (N_7429,In_3437,In_79);
or U7430 (N_7430,In_2757,In_4860);
nand U7431 (N_7431,In_237,In_2122);
or U7432 (N_7432,In_3321,In_1241);
nor U7433 (N_7433,In_542,In_1119);
nor U7434 (N_7434,In_2258,In_2605);
nand U7435 (N_7435,In_9,In_2502);
or U7436 (N_7436,In_904,In_4538);
nor U7437 (N_7437,In_2908,In_1972);
and U7438 (N_7438,In_2292,In_973);
nor U7439 (N_7439,In_388,In_656);
nand U7440 (N_7440,In_1260,In_4492);
and U7441 (N_7441,In_2750,In_138);
nand U7442 (N_7442,In_945,In_1976);
and U7443 (N_7443,In_2931,In_2928);
nand U7444 (N_7444,In_1218,In_4835);
nor U7445 (N_7445,In_2096,In_1325);
nand U7446 (N_7446,In_2212,In_2931);
and U7447 (N_7447,In_1821,In_1762);
or U7448 (N_7448,In_619,In_3853);
xnor U7449 (N_7449,In_535,In_1506);
nor U7450 (N_7450,In_4928,In_2358);
or U7451 (N_7451,In_4364,In_1112);
and U7452 (N_7452,In_3587,In_2746);
or U7453 (N_7453,In_3994,In_4021);
nor U7454 (N_7454,In_4298,In_3391);
and U7455 (N_7455,In_2393,In_2282);
or U7456 (N_7456,In_62,In_1035);
nor U7457 (N_7457,In_1284,In_4025);
nand U7458 (N_7458,In_4948,In_4116);
nor U7459 (N_7459,In_2661,In_4425);
nand U7460 (N_7460,In_620,In_3658);
or U7461 (N_7461,In_4575,In_3452);
and U7462 (N_7462,In_4862,In_4616);
nand U7463 (N_7463,In_1500,In_3783);
nor U7464 (N_7464,In_604,In_4233);
nor U7465 (N_7465,In_495,In_1226);
and U7466 (N_7466,In_1786,In_4626);
xor U7467 (N_7467,In_297,In_4168);
or U7468 (N_7468,In_3150,In_4581);
nand U7469 (N_7469,In_3324,In_2147);
or U7470 (N_7470,In_4886,In_1438);
nor U7471 (N_7471,In_1947,In_4698);
nor U7472 (N_7472,In_3541,In_2559);
or U7473 (N_7473,In_3243,In_2915);
and U7474 (N_7474,In_2414,In_3744);
nand U7475 (N_7475,In_4082,In_3404);
nor U7476 (N_7476,In_3081,In_1312);
xor U7477 (N_7477,In_2445,In_3865);
and U7478 (N_7478,In_4891,In_2956);
and U7479 (N_7479,In_2784,In_969);
xnor U7480 (N_7480,In_2151,In_2763);
xnor U7481 (N_7481,In_4897,In_717);
or U7482 (N_7482,In_2509,In_2884);
and U7483 (N_7483,In_3708,In_1347);
and U7484 (N_7484,In_4195,In_329);
or U7485 (N_7485,In_2132,In_1442);
and U7486 (N_7486,In_1275,In_2631);
nand U7487 (N_7487,In_4251,In_1700);
xor U7488 (N_7488,In_3305,In_324);
or U7489 (N_7489,In_231,In_3558);
and U7490 (N_7490,In_3503,In_2815);
nor U7491 (N_7491,In_2775,In_4092);
nor U7492 (N_7492,In_672,In_3596);
and U7493 (N_7493,In_1693,In_1575);
nand U7494 (N_7494,In_2325,In_437);
or U7495 (N_7495,In_143,In_1674);
nor U7496 (N_7496,In_4243,In_1268);
or U7497 (N_7497,In_1346,In_4531);
and U7498 (N_7498,In_4331,In_2893);
nor U7499 (N_7499,In_2656,In_1819);
xor U7500 (N_7500,In_237,In_2230);
or U7501 (N_7501,In_4072,In_4170);
nand U7502 (N_7502,In_1520,In_750);
or U7503 (N_7503,In_833,In_202);
nor U7504 (N_7504,In_4634,In_3550);
and U7505 (N_7505,In_3796,In_2669);
or U7506 (N_7506,In_155,In_2448);
or U7507 (N_7507,In_3676,In_571);
and U7508 (N_7508,In_2710,In_384);
nand U7509 (N_7509,In_461,In_141);
xnor U7510 (N_7510,In_1838,In_4715);
xnor U7511 (N_7511,In_2559,In_1330);
and U7512 (N_7512,In_1424,In_1809);
and U7513 (N_7513,In_4591,In_3083);
nor U7514 (N_7514,In_3891,In_1718);
nor U7515 (N_7515,In_2729,In_1735);
nor U7516 (N_7516,In_604,In_1981);
or U7517 (N_7517,In_2440,In_276);
or U7518 (N_7518,In_707,In_4653);
nor U7519 (N_7519,In_799,In_1385);
nor U7520 (N_7520,In_4809,In_3941);
and U7521 (N_7521,In_2967,In_4779);
nand U7522 (N_7522,In_5,In_267);
nor U7523 (N_7523,In_764,In_3141);
nand U7524 (N_7524,In_2108,In_585);
nand U7525 (N_7525,In_329,In_1663);
nand U7526 (N_7526,In_3976,In_3562);
or U7527 (N_7527,In_3551,In_4094);
nor U7528 (N_7528,In_3338,In_1933);
nor U7529 (N_7529,In_2038,In_1527);
nor U7530 (N_7530,In_4834,In_2634);
or U7531 (N_7531,In_242,In_1628);
xnor U7532 (N_7532,In_1849,In_2922);
nor U7533 (N_7533,In_4112,In_4684);
xor U7534 (N_7534,In_1868,In_3047);
and U7535 (N_7535,In_3107,In_3780);
or U7536 (N_7536,In_4706,In_1552);
nor U7537 (N_7537,In_4336,In_1631);
nor U7538 (N_7538,In_3507,In_2644);
and U7539 (N_7539,In_3817,In_4917);
and U7540 (N_7540,In_4742,In_4005);
nor U7541 (N_7541,In_497,In_4961);
xnor U7542 (N_7542,In_218,In_4475);
nor U7543 (N_7543,In_2962,In_3434);
nor U7544 (N_7544,In_3611,In_2851);
or U7545 (N_7545,In_4826,In_3929);
nor U7546 (N_7546,In_4248,In_2985);
and U7547 (N_7547,In_3395,In_1229);
nor U7548 (N_7548,In_3277,In_1592);
or U7549 (N_7549,In_4764,In_3003);
nor U7550 (N_7550,In_3509,In_477);
nor U7551 (N_7551,In_4709,In_477);
xnor U7552 (N_7552,In_3577,In_2059);
and U7553 (N_7553,In_2379,In_3027);
nand U7554 (N_7554,In_1260,In_1889);
and U7555 (N_7555,In_3386,In_125);
nor U7556 (N_7556,In_4350,In_2660);
or U7557 (N_7557,In_1551,In_564);
and U7558 (N_7558,In_1645,In_4713);
and U7559 (N_7559,In_1765,In_325);
nand U7560 (N_7560,In_309,In_4753);
nor U7561 (N_7561,In_918,In_4552);
or U7562 (N_7562,In_2973,In_3669);
and U7563 (N_7563,In_2407,In_2243);
nand U7564 (N_7564,In_4394,In_3621);
nand U7565 (N_7565,In_1386,In_4777);
nor U7566 (N_7566,In_475,In_1914);
or U7567 (N_7567,In_4002,In_2066);
xnor U7568 (N_7568,In_1159,In_840);
nand U7569 (N_7569,In_977,In_525);
or U7570 (N_7570,In_4143,In_2318);
and U7571 (N_7571,In_3247,In_1319);
nor U7572 (N_7572,In_4870,In_775);
nor U7573 (N_7573,In_562,In_3370);
xor U7574 (N_7574,In_194,In_3339);
or U7575 (N_7575,In_1758,In_3678);
nor U7576 (N_7576,In_3389,In_827);
nand U7577 (N_7577,In_3622,In_1788);
xnor U7578 (N_7578,In_3154,In_1307);
nand U7579 (N_7579,In_1482,In_3035);
nand U7580 (N_7580,In_3038,In_3873);
nor U7581 (N_7581,In_4052,In_1331);
and U7582 (N_7582,In_4665,In_923);
nand U7583 (N_7583,In_4292,In_3408);
xnor U7584 (N_7584,In_80,In_3823);
and U7585 (N_7585,In_3331,In_3556);
nand U7586 (N_7586,In_1314,In_872);
nand U7587 (N_7587,In_504,In_3507);
and U7588 (N_7588,In_3973,In_3698);
or U7589 (N_7589,In_4769,In_4188);
nand U7590 (N_7590,In_270,In_1068);
nand U7591 (N_7591,In_1314,In_1023);
xnor U7592 (N_7592,In_1152,In_4769);
or U7593 (N_7593,In_549,In_3004);
or U7594 (N_7594,In_3474,In_1585);
nand U7595 (N_7595,In_287,In_1417);
nand U7596 (N_7596,In_24,In_1898);
or U7597 (N_7597,In_2263,In_4772);
and U7598 (N_7598,In_1682,In_145);
or U7599 (N_7599,In_2171,In_3905);
xnor U7600 (N_7600,In_1484,In_1569);
xor U7601 (N_7601,In_2112,In_2325);
xnor U7602 (N_7602,In_917,In_1317);
or U7603 (N_7603,In_1774,In_1103);
or U7604 (N_7604,In_3966,In_559);
and U7605 (N_7605,In_3101,In_1488);
nor U7606 (N_7606,In_3194,In_1364);
nand U7607 (N_7607,In_2317,In_755);
or U7608 (N_7608,In_2430,In_277);
and U7609 (N_7609,In_1187,In_4036);
xor U7610 (N_7610,In_574,In_3359);
or U7611 (N_7611,In_4208,In_4277);
or U7612 (N_7612,In_1319,In_405);
xor U7613 (N_7613,In_1539,In_679);
or U7614 (N_7614,In_2815,In_3753);
nand U7615 (N_7615,In_1914,In_636);
and U7616 (N_7616,In_2840,In_724);
and U7617 (N_7617,In_2425,In_3663);
xnor U7618 (N_7618,In_884,In_3822);
nor U7619 (N_7619,In_4702,In_2143);
and U7620 (N_7620,In_2612,In_23);
or U7621 (N_7621,In_2540,In_4693);
nand U7622 (N_7622,In_3399,In_2393);
or U7623 (N_7623,In_550,In_2549);
nor U7624 (N_7624,In_3781,In_1298);
or U7625 (N_7625,In_3642,In_1681);
or U7626 (N_7626,In_1692,In_2866);
or U7627 (N_7627,In_2362,In_4288);
nand U7628 (N_7628,In_2664,In_4456);
nand U7629 (N_7629,In_3511,In_1305);
xnor U7630 (N_7630,In_2973,In_39);
nor U7631 (N_7631,In_632,In_4286);
xor U7632 (N_7632,In_2916,In_1008);
nor U7633 (N_7633,In_4230,In_3259);
xor U7634 (N_7634,In_3523,In_1587);
nand U7635 (N_7635,In_3347,In_2855);
and U7636 (N_7636,In_1655,In_2573);
and U7637 (N_7637,In_1151,In_436);
and U7638 (N_7638,In_3515,In_3667);
nand U7639 (N_7639,In_1410,In_4384);
and U7640 (N_7640,In_1561,In_2198);
and U7641 (N_7641,In_1930,In_1676);
nor U7642 (N_7642,In_3523,In_1400);
nor U7643 (N_7643,In_4537,In_1574);
nand U7644 (N_7644,In_2945,In_144);
or U7645 (N_7645,In_3230,In_642);
and U7646 (N_7646,In_423,In_631);
or U7647 (N_7647,In_4881,In_2520);
nand U7648 (N_7648,In_295,In_4768);
or U7649 (N_7649,In_4719,In_4248);
nand U7650 (N_7650,In_4970,In_3136);
nor U7651 (N_7651,In_1331,In_1657);
or U7652 (N_7652,In_4151,In_1178);
nand U7653 (N_7653,In_3376,In_2976);
xor U7654 (N_7654,In_2676,In_2081);
nor U7655 (N_7655,In_4425,In_1261);
nand U7656 (N_7656,In_868,In_301);
and U7657 (N_7657,In_2396,In_661);
nand U7658 (N_7658,In_2755,In_1473);
nor U7659 (N_7659,In_3463,In_650);
or U7660 (N_7660,In_2322,In_601);
nand U7661 (N_7661,In_3457,In_710);
nand U7662 (N_7662,In_1598,In_1834);
and U7663 (N_7663,In_19,In_1226);
nand U7664 (N_7664,In_2053,In_2731);
or U7665 (N_7665,In_565,In_4874);
or U7666 (N_7666,In_4021,In_3639);
nand U7667 (N_7667,In_3511,In_4717);
and U7668 (N_7668,In_3332,In_1658);
and U7669 (N_7669,In_3392,In_239);
nor U7670 (N_7670,In_606,In_4967);
nor U7671 (N_7671,In_3589,In_2867);
nand U7672 (N_7672,In_2227,In_3119);
xor U7673 (N_7673,In_1683,In_1745);
or U7674 (N_7674,In_2567,In_296);
and U7675 (N_7675,In_2318,In_3655);
nor U7676 (N_7676,In_4046,In_1893);
xnor U7677 (N_7677,In_2226,In_4566);
nand U7678 (N_7678,In_3012,In_261);
nand U7679 (N_7679,In_3214,In_2644);
and U7680 (N_7680,In_1096,In_4125);
or U7681 (N_7681,In_2633,In_1134);
nor U7682 (N_7682,In_3908,In_3133);
xnor U7683 (N_7683,In_2345,In_1354);
or U7684 (N_7684,In_215,In_3363);
and U7685 (N_7685,In_2781,In_438);
nand U7686 (N_7686,In_2491,In_394);
nor U7687 (N_7687,In_2217,In_3351);
nor U7688 (N_7688,In_2098,In_95);
and U7689 (N_7689,In_1935,In_2789);
and U7690 (N_7690,In_532,In_2873);
nor U7691 (N_7691,In_1047,In_4341);
nand U7692 (N_7692,In_2519,In_4299);
xor U7693 (N_7693,In_3059,In_3907);
and U7694 (N_7694,In_645,In_1172);
and U7695 (N_7695,In_2207,In_1738);
nor U7696 (N_7696,In_3214,In_4031);
nor U7697 (N_7697,In_4714,In_1422);
nor U7698 (N_7698,In_4701,In_4094);
nand U7699 (N_7699,In_4511,In_4403);
nor U7700 (N_7700,In_2546,In_1375);
nor U7701 (N_7701,In_2093,In_262);
and U7702 (N_7702,In_4143,In_2202);
xnor U7703 (N_7703,In_3809,In_781);
and U7704 (N_7704,In_4541,In_1803);
or U7705 (N_7705,In_776,In_1808);
nor U7706 (N_7706,In_2393,In_1489);
or U7707 (N_7707,In_2789,In_4865);
or U7708 (N_7708,In_312,In_2499);
and U7709 (N_7709,In_1021,In_2999);
nor U7710 (N_7710,In_3441,In_440);
nand U7711 (N_7711,In_2675,In_1822);
or U7712 (N_7712,In_874,In_2995);
or U7713 (N_7713,In_4431,In_4873);
nor U7714 (N_7714,In_2852,In_269);
and U7715 (N_7715,In_2464,In_2522);
or U7716 (N_7716,In_746,In_3367);
and U7717 (N_7717,In_215,In_2856);
nor U7718 (N_7718,In_4903,In_598);
xnor U7719 (N_7719,In_143,In_3663);
or U7720 (N_7720,In_584,In_4817);
nand U7721 (N_7721,In_211,In_4950);
xnor U7722 (N_7722,In_2894,In_3484);
or U7723 (N_7723,In_2541,In_171);
nor U7724 (N_7724,In_237,In_1446);
nor U7725 (N_7725,In_1449,In_3783);
nand U7726 (N_7726,In_4766,In_638);
and U7727 (N_7727,In_2915,In_2049);
nand U7728 (N_7728,In_3378,In_4070);
and U7729 (N_7729,In_470,In_2261);
nand U7730 (N_7730,In_1301,In_112);
nand U7731 (N_7731,In_419,In_763);
nor U7732 (N_7732,In_4469,In_118);
and U7733 (N_7733,In_3319,In_1214);
or U7734 (N_7734,In_1136,In_4119);
or U7735 (N_7735,In_1691,In_981);
nand U7736 (N_7736,In_1335,In_557);
nor U7737 (N_7737,In_3612,In_2444);
nand U7738 (N_7738,In_4036,In_4550);
nand U7739 (N_7739,In_478,In_1930);
and U7740 (N_7740,In_894,In_4467);
nand U7741 (N_7741,In_4181,In_1409);
and U7742 (N_7742,In_1160,In_2671);
xnor U7743 (N_7743,In_3819,In_1058);
nor U7744 (N_7744,In_3519,In_3239);
or U7745 (N_7745,In_3574,In_2838);
nor U7746 (N_7746,In_3689,In_673);
nor U7747 (N_7747,In_2308,In_3034);
nor U7748 (N_7748,In_638,In_454);
and U7749 (N_7749,In_225,In_2327);
and U7750 (N_7750,In_3204,In_2244);
or U7751 (N_7751,In_4436,In_4080);
and U7752 (N_7752,In_2875,In_3869);
xor U7753 (N_7753,In_2312,In_2933);
nand U7754 (N_7754,In_256,In_3831);
nand U7755 (N_7755,In_4809,In_2756);
and U7756 (N_7756,In_3589,In_2100);
or U7757 (N_7757,In_2039,In_3423);
nand U7758 (N_7758,In_718,In_3491);
or U7759 (N_7759,In_523,In_3248);
nor U7760 (N_7760,In_326,In_1319);
nor U7761 (N_7761,In_3939,In_1115);
nor U7762 (N_7762,In_348,In_2742);
nand U7763 (N_7763,In_4110,In_2674);
nor U7764 (N_7764,In_4159,In_4947);
nor U7765 (N_7765,In_486,In_3873);
and U7766 (N_7766,In_540,In_1377);
or U7767 (N_7767,In_3826,In_3861);
or U7768 (N_7768,In_972,In_1594);
or U7769 (N_7769,In_966,In_3523);
and U7770 (N_7770,In_1050,In_2571);
or U7771 (N_7771,In_3649,In_4043);
and U7772 (N_7772,In_3139,In_1424);
or U7773 (N_7773,In_562,In_3353);
or U7774 (N_7774,In_730,In_1890);
or U7775 (N_7775,In_3156,In_1939);
or U7776 (N_7776,In_2906,In_715);
nor U7777 (N_7777,In_4295,In_2558);
and U7778 (N_7778,In_4569,In_2315);
nor U7779 (N_7779,In_1954,In_3998);
and U7780 (N_7780,In_4841,In_2269);
and U7781 (N_7781,In_1265,In_3414);
xor U7782 (N_7782,In_975,In_71);
nor U7783 (N_7783,In_194,In_794);
and U7784 (N_7784,In_29,In_3662);
and U7785 (N_7785,In_1582,In_811);
nand U7786 (N_7786,In_2967,In_4229);
nand U7787 (N_7787,In_4492,In_584);
or U7788 (N_7788,In_4486,In_1418);
nand U7789 (N_7789,In_2138,In_4668);
nand U7790 (N_7790,In_4278,In_2076);
nor U7791 (N_7791,In_2477,In_3819);
nor U7792 (N_7792,In_4279,In_1645);
nor U7793 (N_7793,In_1026,In_4422);
or U7794 (N_7794,In_1950,In_4234);
xnor U7795 (N_7795,In_1367,In_520);
nor U7796 (N_7796,In_316,In_334);
and U7797 (N_7797,In_4317,In_501);
or U7798 (N_7798,In_1783,In_2407);
nand U7799 (N_7799,In_3583,In_1791);
xor U7800 (N_7800,In_3409,In_2642);
nand U7801 (N_7801,In_2276,In_4844);
and U7802 (N_7802,In_3,In_1171);
or U7803 (N_7803,In_983,In_968);
nand U7804 (N_7804,In_4830,In_2735);
nand U7805 (N_7805,In_413,In_2461);
nand U7806 (N_7806,In_4733,In_4351);
nand U7807 (N_7807,In_4214,In_1766);
and U7808 (N_7808,In_3950,In_885);
nor U7809 (N_7809,In_1476,In_4058);
and U7810 (N_7810,In_2081,In_482);
or U7811 (N_7811,In_4768,In_215);
nor U7812 (N_7812,In_4849,In_3235);
xor U7813 (N_7813,In_766,In_1915);
nand U7814 (N_7814,In_867,In_2063);
nand U7815 (N_7815,In_1541,In_2573);
and U7816 (N_7816,In_4366,In_3889);
nand U7817 (N_7817,In_3492,In_2493);
xor U7818 (N_7818,In_695,In_801);
or U7819 (N_7819,In_2775,In_4026);
and U7820 (N_7820,In_4468,In_864);
nand U7821 (N_7821,In_1438,In_1575);
nand U7822 (N_7822,In_3120,In_2242);
nor U7823 (N_7823,In_1093,In_278);
nand U7824 (N_7824,In_4830,In_753);
or U7825 (N_7825,In_4481,In_4699);
or U7826 (N_7826,In_442,In_1299);
xnor U7827 (N_7827,In_3163,In_2460);
and U7828 (N_7828,In_228,In_4637);
nand U7829 (N_7829,In_1804,In_4703);
and U7830 (N_7830,In_2942,In_2634);
or U7831 (N_7831,In_1634,In_4650);
and U7832 (N_7832,In_2041,In_2446);
nand U7833 (N_7833,In_3223,In_3923);
nor U7834 (N_7834,In_2817,In_1810);
nor U7835 (N_7835,In_4386,In_4405);
and U7836 (N_7836,In_2964,In_2159);
xnor U7837 (N_7837,In_1258,In_3847);
and U7838 (N_7838,In_1567,In_3945);
and U7839 (N_7839,In_4508,In_1371);
nor U7840 (N_7840,In_3904,In_2005);
or U7841 (N_7841,In_3424,In_1273);
nor U7842 (N_7842,In_2777,In_1122);
nor U7843 (N_7843,In_4003,In_2357);
xnor U7844 (N_7844,In_1703,In_3410);
xnor U7845 (N_7845,In_3997,In_3735);
nor U7846 (N_7846,In_436,In_3523);
nor U7847 (N_7847,In_4523,In_987);
nand U7848 (N_7848,In_149,In_4105);
or U7849 (N_7849,In_1348,In_4239);
nand U7850 (N_7850,In_2508,In_2689);
xnor U7851 (N_7851,In_4545,In_2270);
or U7852 (N_7852,In_419,In_4188);
or U7853 (N_7853,In_2158,In_780);
nor U7854 (N_7854,In_1656,In_2656);
nand U7855 (N_7855,In_4637,In_3887);
nor U7856 (N_7856,In_1473,In_468);
or U7857 (N_7857,In_1696,In_2408);
or U7858 (N_7858,In_1615,In_1598);
xor U7859 (N_7859,In_3058,In_2922);
or U7860 (N_7860,In_2009,In_50);
and U7861 (N_7861,In_3309,In_2337);
xor U7862 (N_7862,In_2652,In_2273);
and U7863 (N_7863,In_1113,In_1839);
nor U7864 (N_7864,In_2766,In_146);
nor U7865 (N_7865,In_572,In_1571);
and U7866 (N_7866,In_4839,In_4482);
nor U7867 (N_7867,In_2271,In_3467);
xor U7868 (N_7868,In_909,In_1048);
and U7869 (N_7869,In_710,In_4994);
and U7870 (N_7870,In_913,In_247);
or U7871 (N_7871,In_1996,In_2755);
or U7872 (N_7872,In_3494,In_4433);
nor U7873 (N_7873,In_2299,In_4876);
nand U7874 (N_7874,In_4168,In_4784);
nand U7875 (N_7875,In_273,In_251);
nand U7876 (N_7876,In_3400,In_4801);
or U7877 (N_7877,In_2720,In_2444);
nor U7878 (N_7878,In_3210,In_2749);
and U7879 (N_7879,In_4150,In_2062);
or U7880 (N_7880,In_2698,In_2555);
nor U7881 (N_7881,In_2961,In_2079);
and U7882 (N_7882,In_4024,In_3373);
nand U7883 (N_7883,In_3882,In_2258);
nand U7884 (N_7884,In_2778,In_977);
and U7885 (N_7885,In_2500,In_2976);
nand U7886 (N_7886,In_4708,In_2953);
or U7887 (N_7887,In_448,In_75);
nor U7888 (N_7888,In_446,In_1653);
or U7889 (N_7889,In_2570,In_4398);
nand U7890 (N_7890,In_718,In_910);
nor U7891 (N_7891,In_3319,In_4202);
nand U7892 (N_7892,In_4547,In_2291);
nand U7893 (N_7893,In_917,In_2657);
or U7894 (N_7894,In_2496,In_1902);
nor U7895 (N_7895,In_446,In_2736);
xnor U7896 (N_7896,In_991,In_882);
nand U7897 (N_7897,In_3591,In_1382);
and U7898 (N_7898,In_2915,In_4404);
nand U7899 (N_7899,In_2443,In_2211);
and U7900 (N_7900,In_2664,In_4130);
nor U7901 (N_7901,In_1314,In_2834);
nand U7902 (N_7902,In_4740,In_3740);
or U7903 (N_7903,In_1241,In_4722);
and U7904 (N_7904,In_1172,In_817);
and U7905 (N_7905,In_4077,In_4258);
or U7906 (N_7906,In_4198,In_652);
and U7907 (N_7907,In_4468,In_569);
or U7908 (N_7908,In_4778,In_3223);
and U7909 (N_7909,In_3533,In_3364);
xnor U7910 (N_7910,In_1653,In_2210);
nor U7911 (N_7911,In_689,In_976);
xor U7912 (N_7912,In_1808,In_364);
nand U7913 (N_7913,In_700,In_1180);
or U7914 (N_7914,In_567,In_3310);
nand U7915 (N_7915,In_3299,In_3506);
nand U7916 (N_7916,In_1865,In_835);
and U7917 (N_7917,In_3426,In_3655);
nand U7918 (N_7918,In_4890,In_2350);
and U7919 (N_7919,In_4584,In_2092);
and U7920 (N_7920,In_3876,In_586);
nor U7921 (N_7921,In_1559,In_4587);
nand U7922 (N_7922,In_3925,In_2605);
or U7923 (N_7923,In_1824,In_308);
nand U7924 (N_7924,In_4283,In_2312);
nand U7925 (N_7925,In_4272,In_4218);
nand U7926 (N_7926,In_1727,In_1636);
nor U7927 (N_7927,In_3347,In_84);
and U7928 (N_7928,In_1210,In_3010);
nand U7929 (N_7929,In_648,In_4465);
or U7930 (N_7930,In_2205,In_2131);
nor U7931 (N_7931,In_4383,In_2252);
xnor U7932 (N_7932,In_916,In_4671);
and U7933 (N_7933,In_2492,In_2723);
and U7934 (N_7934,In_563,In_4060);
nor U7935 (N_7935,In_4463,In_3313);
nor U7936 (N_7936,In_4489,In_2665);
nand U7937 (N_7937,In_4937,In_24);
nand U7938 (N_7938,In_4764,In_2076);
nor U7939 (N_7939,In_4287,In_2935);
and U7940 (N_7940,In_874,In_1784);
nand U7941 (N_7941,In_2177,In_1909);
and U7942 (N_7942,In_747,In_4251);
and U7943 (N_7943,In_2891,In_3554);
nor U7944 (N_7944,In_3059,In_1058);
and U7945 (N_7945,In_818,In_1495);
nor U7946 (N_7946,In_560,In_532);
nor U7947 (N_7947,In_4331,In_3132);
and U7948 (N_7948,In_3352,In_3559);
and U7949 (N_7949,In_2382,In_901);
nor U7950 (N_7950,In_2378,In_213);
nor U7951 (N_7951,In_4092,In_3491);
nor U7952 (N_7952,In_2588,In_4089);
or U7953 (N_7953,In_297,In_3614);
and U7954 (N_7954,In_897,In_2122);
or U7955 (N_7955,In_4806,In_4603);
xor U7956 (N_7956,In_3974,In_1964);
nor U7957 (N_7957,In_979,In_2535);
xnor U7958 (N_7958,In_3954,In_1942);
nand U7959 (N_7959,In_522,In_419);
and U7960 (N_7960,In_2946,In_4054);
nor U7961 (N_7961,In_4506,In_384);
xnor U7962 (N_7962,In_2977,In_2622);
or U7963 (N_7963,In_4279,In_3846);
and U7964 (N_7964,In_1676,In_1254);
nor U7965 (N_7965,In_4889,In_3178);
or U7966 (N_7966,In_3835,In_4297);
nor U7967 (N_7967,In_946,In_2193);
xor U7968 (N_7968,In_3359,In_1784);
or U7969 (N_7969,In_2511,In_2766);
or U7970 (N_7970,In_2834,In_10);
nand U7971 (N_7971,In_4114,In_1784);
nand U7972 (N_7972,In_1133,In_2565);
and U7973 (N_7973,In_192,In_2102);
nor U7974 (N_7974,In_3861,In_792);
and U7975 (N_7975,In_3765,In_3327);
or U7976 (N_7976,In_3073,In_4441);
nor U7977 (N_7977,In_1756,In_4069);
and U7978 (N_7978,In_2923,In_1020);
or U7979 (N_7979,In_4419,In_2555);
or U7980 (N_7980,In_2380,In_2752);
and U7981 (N_7981,In_4901,In_573);
nand U7982 (N_7982,In_3466,In_737);
nor U7983 (N_7983,In_3238,In_2646);
nand U7984 (N_7984,In_2493,In_3215);
and U7985 (N_7985,In_2172,In_1994);
and U7986 (N_7986,In_4708,In_4822);
nand U7987 (N_7987,In_1377,In_2071);
or U7988 (N_7988,In_189,In_163);
nand U7989 (N_7989,In_1937,In_1297);
nor U7990 (N_7990,In_1054,In_290);
nand U7991 (N_7991,In_3875,In_2084);
nand U7992 (N_7992,In_1094,In_3628);
or U7993 (N_7993,In_4012,In_1458);
or U7994 (N_7994,In_313,In_1914);
nand U7995 (N_7995,In_3445,In_3857);
and U7996 (N_7996,In_866,In_3946);
and U7997 (N_7997,In_4044,In_1658);
nand U7998 (N_7998,In_967,In_4486);
nand U7999 (N_7999,In_635,In_2081);
or U8000 (N_8000,In_288,In_91);
or U8001 (N_8001,In_4510,In_3197);
nor U8002 (N_8002,In_4377,In_2097);
and U8003 (N_8003,In_3202,In_2162);
nor U8004 (N_8004,In_2143,In_4922);
or U8005 (N_8005,In_373,In_4484);
nand U8006 (N_8006,In_224,In_3587);
nand U8007 (N_8007,In_442,In_63);
nand U8008 (N_8008,In_657,In_4642);
nand U8009 (N_8009,In_3325,In_323);
xnor U8010 (N_8010,In_2553,In_4099);
nor U8011 (N_8011,In_1606,In_4557);
nand U8012 (N_8012,In_1859,In_2516);
or U8013 (N_8013,In_3345,In_662);
nand U8014 (N_8014,In_309,In_3925);
nor U8015 (N_8015,In_4288,In_459);
and U8016 (N_8016,In_4636,In_3391);
or U8017 (N_8017,In_407,In_617);
or U8018 (N_8018,In_3087,In_2517);
and U8019 (N_8019,In_936,In_4053);
and U8020 (N_8020,In_128,In_3576);
and U8021 (N_8021,In_1132,In_4658);
nand U8022 (N_8022,In_3231,In_2187);
nand U8023 (N_8023,In_1395,In_1967);
xor U8024 (N_8024,In_3017,In_565);
nand U8025 (N_8025,In_4663,In_3060);
nand U8026 (N_8026,In_115,In_2937);
and U8027 (N_8027,In_1614,In_1491);
and U8028 (N_8028,In_1069,In_2005);
or U8029 (N_8029,In_2544,In_1076);
or U8030 (N_8030,In_4450,In_1976);
and U8031 (N_8031,In_1778,In_4491);
xor U8032 (N_8032,In_988,In_2888);
nor U8033 (N_8033,In_671,In_1182);
nor U8034 (N_8034,In_1554,In_1882);
nor U8035 (N_8035,In_2331,In_3023);
nor U8036 (N_8036,In_3385,In_3433);
nand U8037 (N_8037,In_4408,In_1063);
or U8038 (N_8038,In_112,In_1362);
nor U8039 (N_8039,In_1887,In_4858);
nand U8040 (N_8040,In_4855,In_600);
nor U8041 (N_8041,In_4148,In_4687);
nand U8042 (N_8042,In_1529,In_1574);
xnor U8043 (N_8043,In_1639,In_4433);
nor U8044 (N_8044,In_648,In_1448);
nand U8045 (N_8045,In_3422,In_4284);
and U8046 (N_8046,In_915,In_1929);
or U8047 (N_8047,In_1464,In_1938);
nor U8048 (N_8048,In_3507,In_4391);
nor U8049 (N_8049,In_34,In_1836);
nor U8050 (N_8050,In_4016,In_4568);
nor U8051 (N_8051,In_3018,In_4262);
or U8052 (N_8052,In_1320,In_4835);
or U8053 (N_8053,In_3555,In_2408);
or U8054 (N_8054,In_1998,In_4318);
or U8055 (N_8055,In_471,In_3859);
or U8056 (N_8056,In_3521,In_4279);
nor U8057 (N_8057,In_3097,In_4869);
or U8058 (N_8058,In_4268,In_2423);
nand U8059 (N_8059,In_909,In_4882);
or U8060 (N_8060,In_1625,In_908);
nor U8061 (N_8061,In_140,In_3676);
and U8062 (N_8062,In_3178,In_3687);
xnor U8063 (N_8063,In_4462,In_3889);
nor U8064 (N_8064,In_3588,In_3074);
or U8065 (N_8065,In_4749,In_1612);
or U8066 (N_8066,In_2547,In_3275);
nand U8067 (N_8067,In_2225,In_2345);
and U8068 (N_8068,In_2214,In_2603);
nand U8069 (N_8069,In_3275,In_2668);
nand U8070 (N_8070,In_96,In_3411);
xor U8071 (N_8071,In_802,In_4751);
nor U8072 (N_8072,In_3446,In_4336);
nor U8073 (N_8073,In_2818,In_1812);
and U8074 (N_8074,In_2677,In_4101);
nor U8075 (N_8075,In_98,In_3700);
or U8076 (N_8076,In_3098,In_2743);
and U8077 (N_8077,In_3451,In_4379);
nand U8078 (N_8078,In_4912,In_4557);
or U8079 (N_8079,In_3515,In_62);
nor U8080 (N_8080,In_1029,In_1030);
or U8081 (N_8081,In_3643,In_2310);
and U8082 (N_8082,In_4060,In_76);
xor U8083 (N_8083,In_4878,In_824);
nor U8084 (N_8084,In_120,In_784);
xor U8085 (N_8085,In_360,In_3691);
nand U8086 (N_8086,In_74,In_1016);
nor U8087 (N_8087,In_2327,In_2991);
or U8088 (N_8088,In_1219,In_1268);
nand U8089 (N_8089,In_4078,In_4597);
nor U8090 (N_8090,In_1174,In_3156);
and U8091 (N_8091,In_4847,In_1416);
nand U8092 (N_8092,In_3433,In_2070);
and U8093 (N_8093,In_2024,In_184);
or U8094 (N_8094,In_654,In_3922);
nand U8095 (N_8095,In_196,In_1533);
and U8096 (N_8096,In_2292,In_2374);
nor U8097 (N_8097,In_2188,In_500);
nand U8098 (N_8098,In_4835,In_4697);
or U8099 (N_8099,In_1765,In_1255);
and U8100 (N_8100,In_4507,In_3069);
and U8101 (N_8101,In_4096,In_3940);
nand U8102 (N_8102,In_689,In_4560);
nand U8103 (N_8103,In_248,In_2349);
nor U8104 (N_8104,In_1903,In_325);
or U8105 (N_8105,In_2679,In_4366);
nor U8106 (N_8106,In_1246,In_2260);
or U8107 (N_8107,In_3401,In_112);
or U8108 (N_8108,In_936,In_34);
or U8109 (N_8109,In_4908,In_2816);
and U8110 (N_8110,In_4680,In_2925);
nor U8111 (N_8111,In_2514,In_1519);
nor U8112 (N_8112,In_1629,In_4580);
xor U8113 (N_8113,In_1824,In_1238);
or U8114 (N_8114,In_1728,In_2056);
or U8115 (N_8115,In_1987,In_419);
and U8116 (N_8116,In_224,In_3549);
or U8117 (N_8117,In_2717,In_1313);
and U8118 (N_8118,In_714,In_3589);
nand U8119 (N_8119,In_4539,In_4933);
nor U8120 (N_8120,In_464,In_3687);
and U8121 (N_8121,In_3951,In_3694);
nand U8122 (N_8122,In_1801,In_1904);
nor U8123 (N_8123,In_1233,In_4484);
nor U8124 (N_8124,In_2024,In_2842);
nand U8125 (N_8125,In_1895,In_4639);
xnor U8126 (N_8126,In_304,In_2669);
or U8127 (N_8127,In_1212,In_1565);
nand U8128 (N_8128,In_4870,In_2159);
xor U8129 (N_8129,In_3079,In_3597);
nor U8130 (N_8130,In_3215,In_1988);
and U8131 (N_8131,In_3735,In_3495);
nand U8132 (N_8132,In_4093,In_2199);
nor U8133 (N_8133,In_2848,In_4017);
nand U8134 (N_8134,In_3111,In_2711);
xnor U8135 (N_8135,In_4302,In_2239);
xnor U8136 (N_8136,In_2965,In_2544);
or U8137 (N_8137,In_4985,In_4679);
nor U8138 (N_8138,In_989,In_69);
nor U8139 (N_8139,In_2073,In_105);
or U8140 (N_8140,In_3222,In_3112);
xnor U8141 (N_8141,In_828,In_3873);
nand U8142 (N_8142,In_910,In_4416);
nand U8143 (N_8143,In_4698,In_3570);
and U8144 (N_8144,In_1776,In_3352);
nor U8145 (N_8145,In_2114,In_4014);
and U8146 (N_8146,In_1079,In_4131);
and U8147 (N_8147,In_1237,In_1900);
nand U8148 (N_8148,In_3828,In_3870);
nor U8149 (N_8149,In_2008,In_4719);
nand U8150 (N_8150,In_634,In_3714);
nand U8151 (N_8151,In_2535,In_3202);
nand U8152 (N_8152,In_741,In_653);
xor U8153 (N_8153,In_1223,In_1272);
nor U8154 (N_8154,In_3966,In_4904);
or U8155 (N_8155,In_1061,In_2162);
or U8156 (N_8156,In_2467,In_4068);
or U8157 (N_8157,In_1352,In_2217);
or U8158 (N_8158,In_2612,In_2451);
and U8159 (N_8159,In_3350,In_4049);
nand U8160 (N_8160,In_1767,In_3749);
and U8161 (N_8161,In_1358,In_3035);
or U8162 (N_8162,In_2173,In_808);
and U8163 (N_8163,In_960,In_3000);
or U8164 (N_8164,In_1403,In_1934);
nor U8165 (N_8165,In_3013,In_1753);
or U8166 (N_8166,In_2221,In_588);
xor U8167 (N_8167,In_996,In_868);
or U8168 (N_8168,In_1136,In_3355);
nor U8169 (N_8169,In_4426,In_762);
nand U8170 (N_8170,In_3021,In_1900);
and U8171 (N_8171,In_4470,In_2681);
nor U8172 (N_8172,In_475,In_3895);
nor U8173 (N_8173,In_4866,In_2556);
nand U8174 (N_8174,In_2694,In_3797);
and U8175 (N_8175,In_902,In_658);
or U8176 (N_8176,In_1841,In_4356);
and U8177 (N_8177,In_1226,In_313);
nand U8178 (N_8178,In_637,In_3970);
and U8179 (N_8179,In_2321,In_949);
or U8180 (N_8180,In_2860,In_451);
and U8181 (N_8181,In_959,In_3793);
and U8182 (N_8182,In_3407,In_4315);
or U8183 (N_8183,In_4752,In_3803);
nand U8184 (N_8184,In_2340,In_4021);
xnor U8185 (N_8185,In_2053,In_3104);
nor U8186 (N_8186,In_4223,In_590);
and U8187 (N_8187,In_3761,In_3918);
and U8188 (N_8188,In_2741,In_1664);
nand U8189 (N_8189,In_4797,In_2091);
or U8190 (N_8190,In_1095,In_1861);
and U8191 (N_8191,In_399,In_4843);
or U8192 (N_8192,In_3653,In_1748);
or U8193 (N_8193,In_1171,In_3321);
nand U8194 (N_8194,In_3919,In_2116);
and U8195 (N_8195,In_3708,In_4715);
nand U8196 (N_8196,In_641,In_1021);
nand U8197 (N_8197,In_1537,In_1564);
nor U8198 (N_8198,In_1171,In_1417);
xnor U8199 (N_8199,In_1946,In_3322);
and U8200 (N_8200,In_2089,In_4756);
nor U8201 (N_8201,In_3334,In_3116);
and U8202 (N_8202,In_3075,In_231);
or U8203 (N_8203,In_476,In_2455);
nand U8204 (N_8204,In_2523,In_3528);
or U8205 (N_8205,In_1756,In_2686);
or U8206 (N_8206,In_3423,In_1446);
nand U8207 (N_8207,In_1616,In_3509);
and U8208 (N_8208,In_2996,In_3066);
nor U8209 (N_8209,In_3637,In_1298);
and U8210 (N_8210,In_1560,In_3829);
or U8211 (N_8211,In_3705,In_1627);
nand U8212 (N_8212,In_1893,In_3602);
nand U8213 (N_8213,In_1263,In_4443);
nor U8214 (N_8214,In_1739,In_517);
and U8215 (N_8215,In_1846,In_509);
nand U8216 (N_8216,In_2986,In_3331);
nand U8217 (N_8217,In_1618,In_3653);
or U8218 (N_8218,In_2013,In_1272);
and U8219 (N_8219,In_3028,In_1062);
and U8220 (N_8220,In_4286,In_3784);
or U8221 (N_8221,In_4626,In_3393);
xor U8222 (N_8222,In_3699,In_1552);
nor U8223 (N_8223,In_1724,In_3846);
nor U8224 (N_8224,In_4863,In_3229);
xor U8225 (N_8225,In_1076,In_910);
nor U8226 (N_8226,In_4148,In_4008);
or U8227 (N_8227,In_2900,In_2386);
nor U8228 (N_8228,In_4306,In_1551);
or U8229 (N_8229,In_379,In_220);
and U8230 (N_8230,In_4330,In_3249);
nor U8231 (N_8231,In_2779,In_4842);
nor U8232 (N_8232,In_2479,In_2669);
and U8233 (N_8233,In_478,In_4587);
nor U8234 (N_8234,In_4138,In_406);
or U8235 (N_8235,In_1748,In_4749);
nor U8236 (N_8236,In_2873,In_1669);
nor U8237 (N_8237,In_4423,In_3134);
and U8238 (N_8238,In_2849,In_3597);
or U8239 (N_8239,In_4755,In_4752);
or U8240 (N_8240,In_3926,In_3254);
and U8241 (N_8241,In_1053,In_3980);
nand U8242 (N_8242,In_4587,In_4057);
or U8243 (N_8243,In_1509,In_145);
xor U8244 (N_8244,In_2422,In_778);
or U8245 (N_8245,In_1238,In_3089);
and U8246 (N_8246,In_3748,In_4555);
and U8247 (N_8247,In_548,In_1574);
nand U8248 (N_8248,In_3331,In_2024);
nor U8249 (N_8249,In_785,In_4797);
or U8250 (N_8250,In_2335,In_4180);
and U8251 (N_8251,In_4097,In_498);
xor U8252 (N_8252,In_2067,In_3127);
or U8253 (N_8253,In_1221,In_4986);
nor U8254 (N_8254,In_1569,In_4714);
and U8255 (N_8255,In_927,In_2600);
or U8256 (N_8256,In_1991,In_1882);
and U8257 (N_8257,In_3607,In_894);
xnor U8258 (N_8258,In_2422,In_2176);
xnor U8259 (N_8259,In_1694,In_849);
or U8260 (N_8260,In_4415,In_3192);
or U8261 (N_8261,In_3563,In_4380);
nor U8262 (N_8262,In_3418,In_4973);
nand U8263 (N_8263,In_3999,In_4014);
and U8264 (N_8264,In_3337,In_1705);
or U8265 (N_8265,In_3878,In_4667);
nor U8266 (N_8266,In_3060,In_1375);
nand U8267 (N_8267,In_722,In_2293);
or U8268 (N_8268,In_2486,In_4466);
nor U8269 (N_8269,In_2459,In_1668);
nand U8270 (N_8270,In_2780,In_2098);
and U8271 (N_8271,In_2901,In_1894);
and U8272 (N_8272,In_766,In_2753);
xnor U8273 (N_8273,In_3705,In_2321);
or U8274 (N_8274,In_3007,In_4426);
nand U8275 (N_8275,In_2536,In_4213);
nor U8276 (N_8276,In_1586,In_4991);
and U8277 (N_8277,In_1987,In_1369);
nor U8278 (N_8278,In_66,In_592);
or U8279 (N_8279,In_1217,In_2792);
nand U8280 (N_8280,In_3907,In_3270);
nand U8281 (N_8281,In_2055,In_1677);
xnor U8282 (N_8282,In_78,In_165);
and U8283 (N_8283,In_2997,In_10);
nand U8284 (N_8284,In_3334,In_3427);
nor U8285 (N_8285,In_4204,In_477);
or U8286 (N_8286,In_1350,In_1523);
nor U8287 (N_8287,In_66,In_2984);
xnor U8288 (N_8288,In_4169,In_3012);
or U8289 (N_8289,In_801,In_1987);
nand U8290 (N_8290,In_1789,In_4729);
or U8291 (N_8291,In_2721,In_3707);
or U8292 (N_8292,In_751,In_1931);
and U8293 (N_8293,In_4290,In_4340);
and U8294 (N_8294,In_30,In_4371);
nor U8295 (N_8295,In_4336,In_1806);
and U8296 (N_8296,In_765,In_4653);
nor U8297 (N_8297,In_3259,In_2684);
or U8298 (N_8298,In_2287,In_3391);
and U8299 (N_8299,In_4908,In_1510);
nor U8300 (N_8300,In_1328,In_2066);
nor U8301 (N_8301,In_2191,In_3862);
nor U8302 (N_8302,In_1915,In_1996);
or U8303 (N_8303,In_124,In_4654);
or U8304 (N_8304,In_422,In_1413);
nor U8305 (N_8305,In_3819,In_2760);
nand U8306 (N_8306,In_1439,In_4697);
or U8307 (N_8307,In_3077,In_2360);
or U8308 (N_8308,In_4622,In_155);
xor U8309 (N_8309,In_2381,In_1689);
or U8310 (N_8310,In_69,In_2673);
nand U8311 (N_8311,In_2687,In_4819);
nand U8312 (N_8312,In_4673,In_2616);
nand U8313 (N_8313,In_4137,In_353);
nand U8314 (N_8314,In_2298,In_2257);
nand U8315 (N_8315,In_2376,In_2867);
and U8316 (N_8316,In_3246,In_4113);
xnor U8317 (N_8317,In_636,In_981);
or U8318 (N_8318,In_4031,In_70);
xnor U8319 (N_8319,In_931,In_3055);
nand U8320 (N_8320,In_4563,In_4847);
or U8321 (N_8321,In_1547,In_2822);
and U8322 (N_8322,In_1661,In_1576);
or U8323 (N_8323,In_1883,In_3168);
nand U8324 (N_8324,In_4791,In_1754);
or U8325 (N_8325,In_1033,In_673);
or U8326 (N_8326,In_1327,In_2622);
nand U8327 (N_8327,In_3520,In_1042);
nor U8328 (N_8328,In_3906,In_2853);
nand U8329 (N_8329,In_3807,In_4253);
and U8330 (N_8330,In_2820,In_2580);
nand U8331 (N_8331,In_639,In_1463);
and U8332 (N_8332,In_557,In_259);
nand U8333 (N_8333,In_694,In_1981);
nor U8334 (N_8334,In_4229,In_45);
or U8335 (N_8335,In_4738,In_1826);
nor U8336 (N_8336,In_843,In_493);
and U8337 (N_8337,In_520,In_1023);
nand U8338 (N_8338,In_3735,In_3719);
or U8339 (N_8339,In_4036,In_1696);
and U8340 (N_8340,In_201,In_3780);
and U8341 (N_8341,In_4082,In_4367);
xnor U8342 (N_8342,In_3264,In_3763);
xnor U8343 (N_8343,In_1985,In_1910);
nand U8344 (N_8344,In_1284,In_409);
and U8345 (N_8345,In_3493,In_1415);
nand U8346 (N_8346,In_1779,In_3332);
nor U8347 (N_8347,In_1149,In_2301);
or U8348 (N_8348,In_1447,In_718);
nor U8349 (N_8349,In_768,In_886);
nor U8350 (N_8350,In_4721,In_2903);
or U8351 (N_8351,In_3719,In_4604);
nor U8352 (N_8352,In_3520,In_2668);
nor U8353 (N_8353,In_1941,In_2821);
or U8354 (N_8354,In_1468,In_1066);
xor U8355 (N_8355,In_1379,In_1266);
nand U8356 (N_8356,In_1690,In_3400);
nor U8357 (N_8357,In_2375,In_1357);
nor U8358 (N_8358,In_708,In_153);
and U8359 (N_8359,In_2629,In_4008);
xnor U8360 (N_8360,In_1708,In_2644);
or U8361 (N_8361,In_4422,In_1503);
xnor U8362 (N_8362,In_2504,In_3922);
and U8363 (N_8363,In_1796,In_4590);
xnor U8364 (N_8364,In_3005,In_4218);
nor U8365 (N_8365,In_2136,In_4422);
nor U8366 (N_8366,In_3642,In_618);
or U8367 (N_8367,In_3758,In_4736);
or U8368 (N_8368,In_4198,In_2374);
or U8369 (N_8369,In_1334,In_2988);
nand U8370 (N_8370,In_175,In_4563);
nand U8371 (N_8371,In_540,In_1603);
nor U8372 (N_8372,In_1563,In_1639);
xor U8373 (N_8373,In_709,In_2322);
nor U8374 (N_8374,In_1171,In_1348);
nor U8375 (N_8375,In_4264,In_1687);
nor U8376 (N_8376,In_3200,In_201);
nor U8377 (N_8377,In_2308,In_3147);
and U8378 (N_8378,In_2504,In_2173);
and U8379 (N_8379,In_422,In_360);
and U8380 (N_8380,In_1040,In_93);
xnor U8381 (N_8381,In_2313,In_3810);
and U8382 (N_8382,In_537,In_3452);
and U8383 (N_8383,In_164,In_4115);
nand U8384 (N_8384,In_84,In_1473);
or U8385 (N_8385,In_4555,In_734);
nand U8386 (N_8386,In_4672,In_454);
nor U8387 (N_8387,In_330,In_3681);
nor U8388 (N_8388,In_3852,In_2842);
xor U8389 (N_8389,In_2866,In_1468);
or U8390 (N_8390,In_2023,In_136);
or U8391 (N_8391,In_2324,In_1511);
nor U8392 (N_8392,In_1666,In_3393);
nor U8393 (N_8393,In_1506,In_2353);
and U8394 (N_8394,In_572,In_3640);
nand U8395 (N_8395,In_3977,In_108);
xnor U8396 (N_8396,In_3563,In_3216);
and U8397 (N_8397,In_763,In_4859);
and U8398 (N_8398,In_2810,In_4990);
and U8399 (N_8399,In_1466,In_233);
or U8400 (N_8400,In_3866,In_4356);
or U8401 (N_8401,In_3273,In_1311);
or U8402 (N_8402,In_2614,In_2820);
or U8403 (N_8403,In_3515,In_3551);
xor U8404 (N_8404,In_1266,In_1441);
or U8405 (N_8405,In_2728,In_4964);
and U8406 (N_8406,In_236,In_3202);
nand U8407 (N_8407,In_1225,In_3681);
and U8408 (N_8408,In_3108,In_3765);
nand U8409 (N_8409,In_76,In_3137);
nor U8410 (N_8410,In_4382,In_3760);
or U8411 (N_8411,In_3967,In_637);
nand U8412 (N_8412,In_4509,In_3077);
nor U8413 (N_8413,In_3240,In_1039);
nand U8414 (N_8414,In_566,In_4575);
and U8415 (N_8415,In_779,In_3956);
and U8416 (N_8416,In_3916,In_658);
nor U8417 (N_8417,In_1347,In_1346);
nand U8418 (N_8418,In_3724,In_854);
nand U8419 (N_8419,In_460,In_1785);
nor U8420 (N_8420,In_3880,In_4364);
nor U8421 (N_8421,In_3479,In_3216);
and U8422 (N_8422,In_4200,In_3953);
and U8423 (N_8423,In_3799,In_442);
nor U8424 (N_8424,In_1333,In_2016);
nand U8425 (N_8425,In_2471,In_2364);
and U8426 (N_8426,In_541,In_2814);
xnor U8427 (N_8427,In_2619,In_2497);
nand U8428 (N_8428,In_2950,In_3035);
and U8429 (N_8429,In_1106,In_4845);
nand U8430 (N_8430,In_1534,In_2824);
or U8431 (N_8431,In_2097,In_2417);
or U8432 (N_8432,In_4117,In_4498);
nand U8433 (N_8433,In_2358,In_176);
nand U8434 (N_8434,In_555,In_4513);
or U8435 (N_8435,In_2350,In_1298);
and U8436 (N_8436,In_295,In_2066);
nor U8437 (N_8437,In_2198,In_2866);
nand U8438 (N_8438,In_390,In_2020);
nand U8439 (N_8439,In_1647,In_2224);
xor U8440 (N_8440,In_3076,In_125);
or U8441 (N_8441,In_3125,In_4957);
or U8442 (N_8442,In_606,In_1925);
nor U8443 (N_8443,In_4999,In_3818);
nand U8444 (N_8444,In_2834,In_1704);
nor U8445 (N_8445,In_4922,In_3246);
or U8446 (N_8446,In_4326,In_2213);
nor U8447 (N_8447,In_158,In_2306);
xor U8448 (N_8448,In_3740,In_1941);
nand U8449 (N_8449,In_733,In_1584);
nor U8450 (N_8450,In_1197,In_3026);
nand U8451 (N_8451,In_1890,In_434);
nand U8452 (N_8452,In_2664,In_3331);
xnor U8453 (N_8453,In_2257,In_4003);
or U8454 (N_8454,In_4350,In_31);
nand U8455 (N_8455,In_4639,In_3927);
nor U8456 (N_8456,In_2701,In_3902);
nor U8457 (N_8457,In_4231,In_753);
and U8458 (N_8458,In_2471,In_1329);
or U8459 (N_8459,In_2844,In_4720);
nand U8460 (N_8460,In_1282,In_3897);
and U8461 (N_8461,In_2916,In_2713);
or U8462 (N_8462,In_1014,In_4285);
nor U8463 (N_8463,In_3220,In_4911);
nor U8464 (N_8464,In_3448,In_1387);
and U8465 (N_8465,In_743,In_233);
xor U8466 (N_8466,In_4293,In_1843);
nor U8467 (N_8467,In_1011,In_4636);
nand U8468 (N_8468,In_1938,In_742);
nor U8469 (N_8469,In_4877,In_3264);
or U8470 (N_8470,In_2592,In_2905);
or U8471 (N_8471,In_2217,In_2757);
nand U8472 (N_8472,In_3639,In_2561);
nand U8473 (N_8473,In_3610,In_1971);
nand U8474 (N_8474,In_1843,In_2522);
xor U8475 (N_8475,In_4128,In_399);
nor U8476 (N_8476,In_3291,In_4898);
and U8477 (N_8477,In_138,In_1387);
and U8478 (N_8478,In_4218,In_2478);
nor U8479 (N_8479,In_1714,In_3653);
nand U8480 (N_8480,In_2956,In_3034);
or U8481 (N_8481,In_2094,In_3609);
and U8482 (N_8482,In_7,In_3826);
and U8483 (N_8483,In_2054,In_3166);
or U8484 (N_8484,In_1300,In_3971);
nor U8485 (N_8485,In_3451,In_1036);
nor U8486 (N_8486,In_1658,In_862);
nand U8487 (N_8487,In_4255,In_3310);
or U8488 (N_8488,In_999,In_2175);
nor U8489 (N_8489,In_2547,In_3986);
nor U8490 (N_8490,In_2975,In_628);
and U8491 (N_8491,In_1155,In_2465);
or U8492 (N_8492,In_3384,In_4544);
xnor U8493 (N_8493,In_2882,In_1715);
and U8494 (N_8494,In_4099,In_3709);
and U8495 (N_8495,In_2316,In_2910);
or U8496 (N_8496,In_4506,In_1463);
nand U8497 (N_8497,In_904,In_3028);
or U8498 (N_8498,In_543,In_2635);
xnor U8499 (N_8499,In_3891,In_2251);
nand U8500 (N_8500,In_3528,In_2750);
or U8501 (N_8501,In_31,In_3138);
nor U8502 (N_8502,In_3850,In_4075);
nand U8503 (N_8503,In_1761,In_784);
and U8504 (N_8504,In_370,In_3902);
or U8505 (N_8505,In_2170,In_518);
nor U8506 (N_8506,In_3409,In_78);
nor U8507 (N_8507,In_4817,In_1371);
and U8508 (N_8508,In_1038,In_4659);
nor U8509 (N_8509,In_2508,In_3858);
nand U8510 (N_8510,In_1547,In_2861);
nor U8511 (N_8511,In_3148,In_3272);
nand U8512 (N_8512,In_2345,In_4262);
or U8513 (N_8513,In_2449,In_4689);
or U8514 (N_8514,In_1919,In_4811);
and U8515 (N_8515,In_3151,In_305);
nor U8516 (N_8516,In_1036,In_2813);
nand U8517 (N_8517,In_1760,In_4310);
and U8518 (N_8518,In_123,In_1787);
or U8519 (N_8519,In_1224,In_4881);
nand U8520 (N_8520,In_1295,In_2538);
or U8521 (N_8521,In_2113,In_4067);
nor U8522 (N_8522,In_447,In_1902);
nor U8523 (N_8523,In_1319,In_4674);
xnor U8524 (N_8524,In_1533,In_49);
nand U8525 (N_8525,In_3162,In_4408);
nor U8526 (N_8526,In_270,In_4327);
nand U8527 (N_8527,In_685,In_164);
or U8528 (N_8528,In_411,In_4034);
nand U8529 (N_8529,In_4503,In_3684);
nand U8530 (N_8530,In_4689,In_290);
xnor U8531 (N_8531,In_3821,In_3532);
nand U8532 (N_8532,In_1082,In_2766);
xnor U8533 (N_8533,In_4306,In_526);
xor U8534 (N_8534,In_4908,In_2024);
or U8535 (N_8535,In_3191,In_4318);
nand U8536 (N_8536,In_3058,In_2203);
nor U8537 (N_8537,In_1533,In_2372);
nand U8538 (N_8538,In_3899,In_4425);
nor U8539 (N_8539,In_1510,In_1170);
xnor U8540 (N_8540,In_1413,In_4585);
or U8541 (N_8541,In_3858,In_1164);
and U8542 (N_8542,In_1633,In_2115);
or U8543 (N_8543,In_1912,In_3521);
xnor U8544 (N_8544,In_2254,In_1700);
nor U8545 (N_8545,In_2833,In_393);
or U8546 (N_8546,In_3139,In_4725);
or U8547 (N_8547,In_3652,In_2441);
nand U8548 (N_8548,In_2333,In_2311);
or U8549 (N_8549,In_8,In_4903);
nor U8550 (N_8550,In_1009,In_3348);
nor U8551 (N_8551,In_3893,In_113);
nand U8552 (N_8552,In_1565,In_1626);
and U8553 (N_8553,In_1680,In_1707);
and U8554 (N_8554,In_1275,In_3676);
or U8555 (N_8555,In_3821,In_451);
xor U8556 (N_8556,In_2276,In_4688);
nor U8557 (N_8557,In_1329,In_3072);
nand U8558 (N_8558,In_4752,In_1556);
nand U8559 (N_8559,In_2759,In_965);
and U8560 (N_8560,In_3300,In_2914);
xnor U8561 (N_8561,In_1181,In_1978);
nand U8562 (N_8562,In_3422,In_1524);
nand U8563 (N_8563,In_3802,In_270);
nand U8564 (N_8564,In_4772,In_2333);
nand U8565 (N_8565,In_3071,In_3452);
or U8566 (N_8566,In_4883,In_4084);
and U8567 (N_8567,In_268,In_2049);
nor U8568 (N_8568,In_800,In_1069);
nand U8569 (N_8569,In_1979,In_2809);
nor U8570 (N_8570,In_4934,In_3428);
nor U8571 (N_8571,In_3983,In_1672);
or U8572 (N_8572,In_2334,In_398);
xnor U8573 (N_8573,In_2400,In_1138);
and U8574 (N_8574,In_4342,In_3828);
or U8575 (N_8575,In_3723,In_4894);
and U8576 (N_8576,In_2976,In_4030);
nand U8577 (N_8577,In_2971,In_4248);
and U8578 (N_8578,In_4792,In_793);
and U8579 (N_8579,In_3997,In_715);
nor U8580 (N_8580,In_2920,In_4505);
nand U8581 (N_8581,In_292,In_4125);
or U8582 (N_8582,In_3941,In_2347);
nor U8583 (N_8583,In_2983,In_3448);
and U8584 (N_8584,In_1183,In_1290);
nor U8585 (N_8585,In_4360,In_3632);
nor U8586 (N_8586,In_2928,In_2417);
or U8587 (N_8587,In_1882,In_4176);
xor U8588 (N_8588,In_43,In_360);
nor U8589 (N_8589,In_896,In_4112);
or U8590 (N_8590,In_1357,In_3644);
nor U8591 (N_8591,In_4446,In_2966);
or U8592 (N_8592,In_721,In_3224);
xnor U8593 (N_8593,In_1736,In_3757);
nor U8594 (N_8594,In_4518,In_3526);
nor U8595 (N_8595,In_1952,In_2452);
or U8596 (N_8596,In_3299,In_4836);
nor U8597 (N_8597,In_1229,In_2879);
or U8598 (N_8598,In_2082,In_791);
nor U8599 (N_8599,In_3359,In_2083);
nand U8600 (N_8600,In_791,In_4276);
nor U8601 (N_8601,In_1960,In_3078);
and U8602 (N_8602,In_3966,In_1592);
and U8603 (N_8603,In_4844,In_704);
xor U8604 (N_8604,In_1092,In_2297);
or U8605 (N_8605,In_1195,In_3671);
or U8606 (N_8606,In_3070,In_2117);
xnor U8607 (N_8607,In_1064,In_3839);
or U8608 (N_8608,In_2842,In_3946);
or U8609 (N_8609,In_1032,In_3058);
and U8610 (N_8610,In_3303,In_2925);
nor U8611 (N_8611,In_140,In_4957);
and U8612 (N_8612,In_4377,In_4992);
or U8613 (N_8613,In_2487,In_767);
and U8614 (N_8614,In_3045,In_3621);
xor U8615 (N_8615,In_1045,In_3835);
xnor U8616 (N_8616,In_2010,In_987);
and U8617 (N_8617,In_2557,In_4009);
nor U8618 (N_8618,In_1214,In_174);
xnor U8619 (N_8619,In_1386,In_1486);
nand U8620 (N_8620,In_2315,In_476);
nand U8621 (N_8621,In_2693,In_4989);
nand U8622 (N_8622,In_4971,In_881);
xnor U8623 (N_8623,In_1666,In_4336);
nand U8624 (N_8624,In_1394,In_1487);
and U8625 (N_8625,In_1265,In_581);
nand U8626 (N_8626,In_2637,In_3157);
xnor U8627 (N_8627,In_3348,In_4556);
and U8628 (N_8628,In_3539,In_4908);
nand U8629 (N_8629,In_1937,In_184);
xnor U8630 (N_8630,In_4479,In_3826);
or U8631 (N_8631,In_214,In_3973);
nand U8632 (N_8632,In_4271,In_419);
nand U8633 (N_8633,In_1427,In_2326);
or U8634 (N_8634,In_3851,In_4910);
nand U8635 (N_8635,In_2862,In_3023);
or U8636 (N_8636,In_2757,In_3613);
and U8637 (N_8637,In_2587,In_1560);
nand U8638 (N_8638,In_3715,In_2340);
nand U8639 (N_8639,In_1541,In_4129);
nand U8640 (N_8640,In_2663,In_4243);
nand U8641 (N_8641,In_4321,In_4924);
xor U8642 (N_8642,In_3368,In_1690);
and U8643 (N_8643,In_4298,In_1093);
or U8644 (N_8644,In_3699,In_106);
or U8645 (N_8645,In_4781,In_2565);
nor U8646 (N_8646,In_4838,In_3504);
nor U8647 (N_8647,In_1450,In_913);
nor U8648 (N_8648,In_4547,In_4097);
nand U8649 (N_8649,In_4757,In_2865);
and U8650 (N_8650,In_2106,In_1345);
nor U8651 (N_8651,In_2169,In_195);
nor U8652 (N_8652,In_2395,In_4039);
and U8653 (N_8653,In_4065,In_3294);
and U8654 (N_8654,In_247,In_2268);
xnor U8655 (N_8655,In_4699,In_4817);
nor U8656 (N_8656,In_3829,In_4293);
xnor U8657 (N_8657,In_699,In_1648);
and U8658 (N_8658,In_2309,In_2240);
and U8659 (N_8659,In_4617,In_3147);
and U8660 (N_8660,In_1941,In_4046);
nor U8661 (N_8661,In_4321,In_2455);
nand U8662 (N_8662,In_3594,In_857);
or U8663 (N_8663,In_2212,In_850);
xor U8664 (N_8664,In_3655,In_1018);
nand U8665 (N_8665,In_350,In_2180);
or U8666 (N_8666,In_3040,In_673);
nor U8667 (N_8667,In_2777,In_1551);
nand U8668 (N_8668,In_3249,In_3978);
or U8669 (N_8669,In_872,In_908);
nor U8670 (N_8670,In_2109,In_3341);
nand U8671 (N_8671,In_4719,In_3704);
or U8672 (N_8672,In_361,In_2128);
nand U8673 (N_8673,In_2014,In_3080);
or U8674 (N_8674,In_1414,In_4879);
nor U8675 (N_8675,In_4959,In_790);
nor U8676 (N_8676,In_3878,In_2283);
nor U8677 (N_8677,In_4685,In_1387);
and U8678 (N_8678,In_4659,In_680);
or U8679 (N_8679,In_1298,In_1743);
nand U8680 (N_8680,In_995,In_858);
xor U8681 (N_8681,In_2682,In_2541);
nor U8682 (N_8682,In_1307,In_913);
or U8683 (N_8683,In_1023,In_2966);
nand U8684 (N_8684,In_1199,In_3856);
nand U8685 (N_8685,In_3970,In_4295);
or U8686 (N_8686,In_4562,In_622);
and U8687 (N_8687,In_4258,In_801);
and U8688 (N_8688,In_2965,In_3720);
and U8689 (N_8689,In_661,In_4895);
or U8690 (N_8690,In_555,In_249);
and U8691 (N_8691,In_2493,In_1935);
xor U8692 (N_8692,In_2142,In_1771);
and U8693 (N_8693,In_3801,In_2649);
or U8694 (N_8694,In_2121,In_4891);
or U8695 (N_8695,In_639,In_4265);
xnor U8696 (N_8696,In_4853,In_4857);
or U8697 (N_8697,In_986,In_2763);
and U8698 (N_8698,In_1145,In_1982);
nor U8699 (N_8699,In_4176,In_4309);
and U8700 (N_8700,In_4747,In_3661);
xnor U8701 (N_8701,In_946,In_1631);
nor U8702 (N_8702,In_4814,In_3811);
and U8703 (N_8703,In_2068,In_3809);
or U8704 (N_8704,In_1659,In_2509);
nand U8705 (N_8705,In_1250,In_4264);
nand U8706 (N_8706,In_344,In_4002);
or U8707 (N_8707,In_1929,In_1142);
and U8708 (N_8708,In_2843,In_3715);
nand U8709 (N_8709,In_2936,In_2245);
nor U8710 (N_8710,In_4465,In_3271);
xor U8711 (N_8711,In_3475,In_4832);
or U8712 (N_8712,In_4914,In_4334);
nor U8713 (N_8713,In_2847,In_84);
and U8714 (N_8714,In_1537,In_999);
or U8715 (N_8715,In_210,In_4765);
xor U8716 (N_8716,In_2307,In_2083);
nor U8717 (N_8717,In_3040,In_4193);
nand U8718 (N_8718,In_2300,In_891);
nor U8719 (N_8719,In_119,In_607);
nand U8720 (N_8720,In_2156,In_387);
and U8721 (N_8721,In_3090,In_1336);
nor U8722 (N_8722,In_3727,In_4802);
nor U8723 (N_8723,In_2779,In_524);
and U8724 (N_8724,In_3068,In_368);
or U8725 (N_8725,In_4661,In_2095);
or U8726 (N_8726,In_281,In_4719);
nand U8727 (N_8727,In_1109,In_2368);
nor U8728 (N_8728,In_4057,In_3973);
and U8729 (N_8729,In_846,In_1241);
or U8730 (N_8730,In_4097,In_1521);
nand U8731 (N_8731,In_1953,In_4267);
nand U8732 (N_8732,In_1513,In_2269);
or U8733 (N_8733,In_711,In_101);
or U8734 (N_8734,In_3847,In_4689);
or U8735 (N_8735,In_101,In_687);
and U8736 (N_8736,In_2880,In_1808);
and U8737 (N_8737,In_4015,In_3949);
nand U8738 (N_8738,In_1962,In_2042);
nor U8739 (N_8739,In_4863,In_3924);
nand U8740 (N_8740,In_4240,In_4357);
nand U8741 (N_8741,In_3201,In_1642);
nor U8742 (N_8742,In_1464,In_234);
xor U8743 (N_8743,In_1754,In_2422);
nor U8744 (N_8744,In_3299,In_1664);
xor U8745 (N_8745,In_4351,In_3615);
nor U8746 (N_8746,In_4957,In_407);
and U8747 (N_8747,In_4959,In_1989);
or U8748 (N_8748,In_1505,In_3260);
or U8749 (N_8749,In_1984,In_3917);
and U8750 (N_8750,In_1132,In_941);
or U8751 (N_8751,In_3395,In_2888);
and U8752 (N_8752,In_4213,In_623);
nand U8753 (N_8753,In_3469,In_4712);
nand U8754 (N_8754,In_1835,In_3791);
xnor U8755 (N_8755,In_3011,In_1539);
nand U8756 (N_8756,In_2358,In_716);
and U8757 (N_8757,In_2425,In_75);
nand U8758 (N_8758,In_1738,In_202);
nand U8759 (N_8759,In_1849,In_4357);
nand U8760 (N_8760,In_510,In_1957);
and U8761 (N_8761,In_2843,In_2078);
nor U8762 (N_8762,In_1520,In_4574);
or U8763 (N_8763,In_1405,In_3294);
and U8764 (N_8764,In_393,In_67);
nand U8765 (N_8765,In_346,In_4985);
and U8766 (N_8766,In_2254,In_4995);
and U8767 (N_8767,In_4263,In_4927);
or U8768 (N_8768,In_2203,In_3406);
and U8769 (N_8769,In_3492,In_769);
nor U8770 (N_8770,In_749,In_2904);
nor U8771 (N_8771,In_4796,In_2791);
nor U8772 (N_8772,In_257,In_2124);
xor U8773 (N_8773,In_4316,In_1024);
xor U8774 (N_8774,In_1274,In_91);
nor U8775 (N_8775,In_3827,In_4411);
nand U8776 (N_8776,In_4792,In_1298);
or U8777 (N_8777,In_3551,In_310);
nor U8778 (N_8778,In_4167,In_822);
xor U8779 (N_8779,In_4678,In_1363);
xnor U8780 (N_8780,In_2359,In_4631);
or U8781 (N_8781,In_3140,In_4985);
or U8782 (N_8782,In_4711,In_163);
or U8783 (N_8783,In_1457,In_4274);
nor U8784 (N_8784,In_4153,In_4621);
nand U8785 (N_8785,In_4404,In_2895);
and U8786 (N_8786,In_2290,In_3639);
xnor U8787 (N_8787,In_4614,In_3511);
nand U8788 (N_8788,In_2236,In_2340);
or U8789 (N_8789,In_1006,In_3124);
nand U8790 (N_8790,In_3699,In_1384);
nor U8791 (N_8791,In_4360,In_164);
and U8792 (N_8792,In_3931,In_1342);
xnor U8793 (N_8793,In_1796,In_1923);
nand U8794 (N_8794,In_3954,In_2671);
nor U8795 (N_8795,In_632,In_4396);
nand U8796 (N_8796,In_2613,In_2083);
nor U8797 (N_8797,In_3459,In_567);
nor U8798 (N_8798,In_3009,In_1490);
nand U8799 (N_8799,In_557,In_508);
or U8800 (N_8800,In_1498,In_3603);
and U8801 (N_8801,In_2366,In_30);
nand U8802 (N_8802,In_2364,In_3107);
nor U8803 (N_8803,In_2027,In_2665);
nand U8804 (N_8804,In_517,In_1335);
nand U8805 (N_8805,In_1073,In_2162);
and U8806 (N_8806,In_1906,In_2286);
and U8807 (N_8807,In_4323,In_215);
nor U8808 (N_8808,In_2499,In_1579);
and U8809 (N_8809,In_3500,In_4652);
and U8810 (N_8810,In_698,In_2563);
nor U8811 (N_8811,In_2253,In_1272);
xnor U8812 (N_8812,In_2776,In_4386);
nor U8813 (N_8813,In_4298,In_1290);
and U8814 (N_8814,In_474,In_3997);
xnor U8815 (N_8815,In_3524,In_2233);
or U8816 (N_8816,In_1074,In_3004);
xnor U8817 (N_8817,In_4754,In_4896);
and U8818 (N_8818,In_1144,In_203);
xnor U8819 (N_8819,In_2748,In_474);
and U8820 (N_8820,In_2159,In_3688);
or U8821 (N_8821,In_1422,In_830);
or U8822 (N_8822,In_368,In_4836);
or U8823 (N_8823,In_2081,In_4265);
nand U8824 (N_8824,In_2884,In_4700);
nor U8825 (N_8825,In_3820,In_543);
or U8826 (N_8826,In_1466,In_678);
xnor U8827 (N_8827,In_180,In_3236);
and U8828 (N_8828,In_2987,In_4319);
and U8829 (N_8829,In_1316,In_1105);
or U8830 (N_8830,In_2378,In_1354);
and U8831 (N_8831,In_2767,In_3858);
and U8832 (N_8832,In_1039,In_1138);
nand U8833 (N_8833,In_4458,In_4135);
nor U8834 (N_8834,In_4466,In_4202);
xor U8835 (N_8835,In_1867,In_1333);
and U8836 (N_8836,In_769,In_2639);
nor U8837 (N_8837,In_2941,In_4615);
xnor U8838 (N_8838,In_3265,In_1997);
nand U8839 (N_8839,In_463,In_2493);
and U8840 (N_8840,In_2301,In_4756);
nor U8841 (N_8841,In_3447,In_3890);
nand U8842 (N_8842,In_1272,In_3705);
or U8843 (N_8843,In_3741,In_3030);
nor U8844 (N_8844,In_2030,In_999);
xnor U8845 (N_8845,In_656,In_205);
nor U8846 (N_8846,In_3789,In_1763);
xnor U8847 (N_8847,In_2270,In_3721);
or U8848 (N_8848,In_3794,In_2210);
or U8849 (N_8849,In_2611,In_515);
and U8850 (N_8850,In_277,In_2898);
or U8851 (N_8851,In_3362,In_4044);
or U8852 (N_8852,In_3008,In_4812);
or U8853 (N_8853,In_390,In_3181);
xnor U8854 (N_8854,In_4169,In_3999);
nor U8855 (N_8855,In_3920,In_2691);
and U8856 (N_8856,In_1679,In_1125);
and U8857 (N_8857,In_3193,In_1277);
nor U8858 (N_8858,In_502,In_4208);
nor U8859 (N_8859,In_1632,In_928);
nor U8860 (N_8860,In_3422,In_43);
and U8861 (N_8861,In_2943,In_2836);
and U8862 (N_8862,In_2035,In_1855);
nand U8863 (N_8863,In_81,In_1323);
and U8864 (N_8864,In_2087,In_434);
or U8865 (N_8865,In_2660,In_45);
nand U8866 (N_8866,In_4964,In_3611);
nand U8867 (N_8867,In_2743,In_326);
nand U8868 (N_8868,In_1610,In_2949);
nand U8869 (N_8869,In_1512,In_2853);
nor U8870 (N_8870,In_4673,In_1100);
nand U8871 (N_8871,In_4802,In_474);
nor U8872 (N_8872,In_3956,In_3584);
xor U8873 (N_8873,In_3391,In_3460);
nor U8874 (N_8874,In_1652,In_1020);
nor U8875 (N_8875,In_4907,In_4494);
nand U8876 (N_8876,In_510,In_3732);
nor U8877 (N_8877,In_4936,In_4868);
and U8878 (N_8878,In_1640,In_2394);
nand U8879 (N_8879,In_524,In_4427);
nand U8880 (N_8880,In_1387,In_3974);
nor U8881 (N_8881,In_2149,In_4930);
nor U8882 (N_8882,In_3902,In_3566);
nor U8883 (N_8883,In_3368,In_601);
and U8884 (N_8884,In_2773,In_3014);
or U8885 (N_8885,In_1236,In_906);
nor U8886 (N_8886,In_1391,In_2991);
nor U8887 (N_8887,In_296,In_3790);
and U8888 (N_8888,In_2627,In_921);
and U8889 (N_8889,In_1682,In_757);
and U8890 (N_8890,In_2040,In_2122);
xor U8891 (N_8891,In_4175,In_3925);
nor U8892 (N_8892,In_1580,In_1416);
xor U8893 (N_8893,In_4527,In_2838);
and U8894 (N_8894,In_2144,In_2644);
nor U8895 (N_8895,In_403,In_4684);
and U8896 (N_8896,In_3646,In_2097);
nor U8897 (N_8897,In_2100,In_1422);
and U8898 (N_8898,In_622,In_1944);
nor U8899 (N_8899,In_2618,In_1751);
nand U8900 (N_8900,In_4562,In_3291);
nand U8901 (N_8901,In_4305,In_1187);
nand U8902 (N_8902,In_3785,In_4139);
and U8903 (N_8903,In_127,In_3171);
or U8904 (N_8904,In_1127,In_2724);
or U8905 (N_8905,In_458,In_970);
xnor U8906 (N_8906,In_4988,In_1531);
and U8907 (N_8907,In_834,In_2117);
xor U8908 (N_8908,In_3119,In_1381);
xor U8909 (N_8909,In_1142,In_1321);
nand U8910 (N_8910,In_4042,In_3584);
nor U8911 (N_8911,In_4672,In_534);
nand U8912 (N_8912,In_3697,In_510);
or U8913 (N_8913,In_2948,In_4867);
nor U8914 (N_8914,In_1331,In_3722);
and U8915 (N_8915,In_2806,In_2322);
or U8916 (N_8916,In_4079,In_4293);
nor U8917 (N_8917,In_639,In_3038);
nor U8918 (N_8918,In_457,In_4306);
and U8919 (N_8919,In_4758,In_2459);
and U8920 (N_8920,In_4322,In_3173);
or U8921 (N_8921,In_1241,In_217);
xnor U8922 (N_8922,In_3963,In_3444);
nor U8923 (N_8923,In_2878,In_2888);
and U8924 (N_8924,In_4817,In_1835);
nor U8925 (N_8925,In_1298,In_467);
nand U8926 (N_8926,In_2394,In_2678);
xnor U8927 (N_8927,In_3249,In_1906);
nor U8928 (N_8928,In_2908,In_2119);
and U8929 (N_8929,In_3199,In_1788);
xor U8930 (N_8930,In_2370,In_2278);
nand U8931 (N_8931,In_2966,In_4973);
nand U8932 (N_8932,In_1266,In_4372);
xnor U8933 (N_8933,In_2665,In_2589);
and U8934 (N_8934,In_2563,In_3001);
or U8935 (N_8935,In_2814,In_4913);
or U8936 (N_8936,In_1556,In_3417);
nor U8937 (N_8937,In_4808,In_4124);
and U8938 (N_8938,In_2306,In_4436);
nand U8939 (N_8939,In_3418,In_2793);
xor U8940 (N_8940,In_1215,In_3584);
and U8941 (N_8941,In_1293,In_4915);
xor U8942 (N_8942,In_3996,In_2952);
and U8943 (N_8943,In_2166,In_493);
nand U8944 (N_8944,In_4365,In_3084);
nor U8945 (N_8945,In_714,In_867);
or U8946 (N_8946,In_4889,In_3260);
nor U8947 (N_8947,In_1317,In_2896);
nor U8948 (N_8948,In_3958,In_883);
and U8949 (N_8949,In_811,In_1671);
xor U8950 (N_8950,In_2395,In_2735);
and U8951 (N_8951,In_2314,In_1792);
nand U8952 (N_8952,In_187,In_3862);
nor U8953 (N_8953,In_4822,In_2414);
and U8954 (N_8954,In_3191,In_1304);
xor U8955 (N_8955,In_905,In_1632);
nor U8956 (N_8956,In_3247,In_4796);
or U8957 (N_8957,In_4428,In_4192);
and U8958 (N_8958,In_2818,In_2671);
nor U8959 (N_8959,In_3884,In_1428);
nor U8960 (N_8960,In_1588,In_4060);
nor U8961 (N_8961,In_855,In_95);
nand U8962 (N_8962,In_3166,In_4622);
nor U8963 (N_8963,In_1453,In_1091);
nand U8964 (N_8964,In_3223,In_3049);
nor U8965 (N_8965,In_4618,In_2267);
nand U8966 (N_8966,In_3985,In_1500);
nand U8967 (N_8967,In_183,In_4846);
nor U8968 (N_8968,In_2714,In_1908);
xnor U8969 (N_8969,In_4256,In_3279);
nor U8970 (N_8970,In_3069,In_3080);
or U8971 (N_8971,In_3987,In_3709);
or U8972 (N_8972,In_1610,In_424);
and U8973 (N_8973,In_787,In_2463);
nand U8974 (N_8974,In_1720,In_261);
or U8975 (N_8975,In_1801,In_467);
xor U8976 (N_8976,In_4387,In_1609);
or U8977 (N_8977,In_1295,In_1918);
and U8978 (N_8978,In_1171,In_1545);
or U8979 (N_8979,In_2369,In_4358);
or U8980 (N_8980,In_2996,In_3162);
and U8981 (N_8981,In_334,In_3282);
nand U8982 (N_8982,In_3709,In_4784);
or U8983 (N_8983,In_197,In_2683);
or U8984 (N_8984,In_2816,In_589);
or U8985 (N_8985,In_4273,In_1723);
and U8986 (N_8986,In_4060,In_952);
nor U8987 (N_8987,In_2278,In_862);
nand U8988 (N_8988,In_3220,In_2773);
and U8989 (N_8989,In_3260,In_4352);
or U8990 (N_8990,In_1757,In_1977);
nor U8991 (N_8991,In_954,In_854);
or U8992 (N_8992,In_3251,In_260);
nand U8993 (N_8993,In_1056,In_534);
and U8994 (N_8994,In_4668,In_1651);
nand U8995 (N_8995,In_3348,In_2285);
xor U8996 (N_8996,In_4073,In_1210);
and U8997 (N_8997,In_2774,In_37);
or U8998 (N_8998,In_350,In_2054);
or U8999 (N_8999,In_713,In_3250);
or U9000 (N_9000,In_4487,In_3889);
nand U9001 (N_9001,In_3587,In_1897);
nand U9002 (N_9002,In_2993,In_2705);
nor U9003 (N_9003,In_4099,In_2478);
nand U9004 (N_9004,In_1642,In_4466);
nor U9005 (N_9005,In_736,In_3142);
xor U9006 (N_9006,In_1249,In_1659);
or U9007 (N_9007,In_3786,In_1468);
and U9008 (N_9008,In_3170,In_3246);
and U9009 (N_9009,In_2567,In_3047);
and U9010 (N_9010,In_3302,In_201);
and U9011 (N_9011,In_2641,In_298);
or U9012 (N_9012,In_725,In_262);
nand U9013 (N_9013,In_4352,In_4514);
or U9014 (N_9014,In_11,In_4176);
nand U9015 (N_9015,In_3576,In_398);
and U9016 (N_9016,In_3393,In_846);
nor U9017 (N_9017,In_1948,In_4409);
or U9018 (N_9018,In_2134,In_432);
nor U9019 (N_9019,In_36,In_3684);
and U9020 (N_9020,In_4633,In_4003);
xor U9021 (N_9021,In_4817,In_610);
or U9022 (N_9022,In_2449,In_792);
or U9023 (N_9023,In_3822,In_2960);
or U9024 (N_9024,In_514,In_1353);
nand U9025 (N_9025,In_3692,In_2115);
nand U9026 (N_9026,In_304,In_3619);
and U9027 (N_9027,In_3267,In_3489);
nand U9028 (N_9028,In_3791,In_654);
and U9029 (N_9029,In_2291,In_3332);
and U9030 (N_9030,In_3452,In_1167);
or U9031 (N_9031,In_982,In_2524);
xnor U9032 (N_9032,In_168,In_2846);
xnor U9033 (N_9033,In_2816,In_3144);
xnor U9034 (N_9034,In_922,In_4600);
and U9035 (N_9035,In_2584,In_2317);
nor U9036 (N_9036,In_2671,In_1944);
nor U9037 (N_9037,In_2420,In_2315);
or U9038 (N_9038,In_2896,In_1570);
nand U9039 (N_9039,In_2116,In_1450);
nand U9040 (N_9040,In_3820,In_1549);
and U9041 (N_9041,In_4933,In_54);
nor U9042 (N_9042,In_4936,In_1656);
nand U9043 (N_9043,In_2287,In_4131);
nand U9044 (N_9044,In_3039,In_1664);
nand U9045 (N_9045,In_4435,In_11);
or U9046 (N_9046,In_1172,In_2499);
nand U9047 (N_9047,In_2881,In_215);
and U9048 (N_9048,In_0,In_1751);
or U9049 (N_9049,In_1803,In_2560);
nor U9050 (N_9050,In_1543,In_4710);
xor U9051 (N_9051,In_1392,In_3972);
or U9052 (N_9052,In_948,In_2080);
and U9053 (N_9053,In_4140,In_1919);
xnor U9054 (N_9054,In_2957,In_4373);
xnor U9055 (N_9055,In_1025,In_1893);
nor U9056 (N_9056,In_4439,In_3055);
xnor U9057 (N_9057,In_2005,In_3237);
or U9058 (N_9058,In_1983,In_4626);
and U9059 (N_9059,In_3324,In_3445);
and U9060 (N_9060,In_3871,In_1092);
nor U9061 (N_9061,In_454,In_85);
nand U9062 (N_9062,In_2459,In_3831);
or U9063 (N_9063,In_2855,In_3657);
or U9064 (N_9064,In_274,In_4980);
and U9065 (N_9065,In_860,In_2268);
nor U9066 (N_9066,In_4913,In_3092);
nor U9067 (N_9067,In_861,In_2961);
or U9068 (N_9068,In_3945,In_3280);
nand U9069 (N_9069,In_2490,In_1875);
xor U9070 (N_9070,In_2149,In_2440);
and U9071 (N_9071,In_2305,In_1122);
and U9072 (N_9072,In_2697,In_2116);
nor U9073 (N_9073,In_841,In_3827);
and U9074 (N_9074,In_3666,In_3210);
nand U9075 (N_9075,In_4630,In_3889);
nor U9076 (N_9076,In_3507,In_1519);
and U9077 (N_9077,In_901,In_1226);
xnor U9078 (N_9078,In_315,In_3851);
or U9079 (N_9079,In_4744,In_1527);
or U9080 (N_9080,In_1088,In_4082);
nand U9081 (N_9081,In_85,In_1006);
nor U9082 (N_9082,In_1735,In_538);
and U9083 (N_9083,In_4369,In_1440);
or U9084 (N_9084,In_3122,In_2606);
or U9085 (N_9085,In_2944,In_874);
or U9086 (N_9086,In_1872,In_4547);
and U9087 (N_9087,In_1813,In_820);
nor U9088 (N_9088,In_3616,In_1053);
nor U9089 (N_9089,In_1836,In_3799);
xnor U9090 (N_9090,In_2422,In_494);
nand U9091 (N_9091,In_2134,In_4138);
nor U9092 (N_9092,In_810,In_2505);
and U9093 (N_9093,In_1471,In_1830);
or U9094 (N_9094,In_2216,In_3420);
xnor U9095 (N_9095,In_3137,In_2996);
xnor U9096 (N_9096,In_2868,In_2683);
xnor U9097 (N_9097,In_3013,In_1205);
nand U9098 (N_9098,In_1047,In_373);
nor U9099 (N_9099,In_4083,In_2009);
nand U9100 (N_9100,In_946,In_1088);
or U9101 (N_9101,In_2917,In_828);
nor U9102 (N_9102,In_1142,In_2294);
and U9103 (N_9103,In_4145,In_4067);
nor U9104 (N_9104,In_781,In_2709);
and U9105 (N_9105,In_4459,In_249);
nor U9106 (N_9106,In_4286,In_4899);
nand U9107 (N_9107,In_3820,In_3946);
and U9108 (N_9108,In_4450,In_976);
nand U9109 (N_9109,In_3871,In_449);
and U9110 (N_9110,In_3514,In_3229);
or U9111 (N_9111,In_2852,In_927);
nor U9112 (N_9112,In_4626,In_726);
and U9113 (N_9113,In_3948,In_4728);
nor U9114 (N_9114,In_4493,In_4329);
or U9115 (N_9115,In_3518,In_2452);
nor U9116 (N_9116,In_540,In_1937);
or U9117 (N_9117,In_1907,In_1680);
nor U9118 (N_9118,In_3984,In_2342);
xor U9119 (N_9119,In_4405,In_4226);
xor U9120 (N_9120,In_4449,In_2677);
nand U9121 (N_9121,In_671,In_3567);
xnor U9122 (N_9122,In_3244,In_1099);
and U9123 (N_9123,In_3546,In_1602);
and U9124 (N_9124,In_4170,In_936);
and U9125 (N_9125,In_2105,In_1995);
nand U9126 (N_9126,In_4455,In_4384);
or U9127 (N_9127,In_2510,In_4798);
and U9128 (N_9128,In_1613,In_2497);
or U9129 (N_9129,In_622,In_4276);
nor U9130 (N_9130,In_3558,In_68);
xnor U9131 (N_9131,In_4548,In_2930);
or U9132 (N_9132,In_3731,In_1019);
nand U9133 (N_9133,In_2079,In_3166);
and U9134 (N_9134,In_3238,In_458);
nor U9135 (N_9135,In_3741,In_377);
xor U9136 (N_9136,In_1762,In_1935);
nor U9137 (N_9137,In_2354,In_2098);
nand U9138 (N_9138,In_4157,In_4634);
or U9139 (N_9139,In_2457,In_2332);
or U9140 (N_9140,In_3441,In_3175);
and U9141 (N_9141,In_968,In_2142);
and U9142 (N_9142,In_1225,In_4645);
and U9143 (N_9143,In_4650,In_1969);
nor U9144 (N_9144,In_3496,In_1886);
and U9145 (N_9145,In_1411,In_3433);
nor U9146 (N_9146,In_1835,In_1209);
or U9147 (N_9147,In_242,In_2116);
nand U9148 (N_9148,In_3742,In_240);
nor U9149 (N_9149,In_3886,In_2552);
and U9150 (N_9150,In_4929,In_3208);
nand U9151 (N_9151,In_780,In_4555);
nand U9152 (N_9152,In_2344,In_4740);
and U9153 (N_9153,In_4886,In_4144);
nor U9154 (N_9154,In_3933,In_3150);
nor U9155 (N_9155,In_4143,In_1326);
nand U9156 (N_9156,In_1194,In_2375);
nand U9157 (N_9157,In_943,In_3854);
nor U9158 (N_9158,In_3752,In_2079);
nand U9159 (N_9159,In_817,In_1373);
nand U9160 (N_9160,In_2685,In_2062);
and U9161 (N_9161,In_804,In_1920);
or U9162 (N_9162,In_870,In_4951);
xor U9163 (N_9163,In_3758,In_4043);
or U9164 (N_9164,In_949,In_4037);
nor U9165 (N_9165,In_3894,In_1060);
nor U9166 (N_9166,In_935,In_3888);
or U9167 (N_9167,In_4950,In_4561);
xnor U9168 (N_9168,In_2632,In_4789);
and U9169 (N_9169,In_710,In_2952);
or U9170 (N_9170,In_1260,In_2835);
or U9171 (N_9171,In_3275,In_4077);
and U9172 (N_9172,In_4497,In_3727);
and U9173 (N_9173,In_3002,In_3543);
xor U9174 (N_9174,In_802,In_897);
xor U9175 (N_9175,In_4460,In_4616);
xor U9176 (N_9176,In_3873,In_966);
nor U9177 (N_9177,In_3638,In_3092);
and U9178 (N_9178,In_1820,In_2524);
or U9179 (N_9179,In_2564,In_1204);
nand U9180 (N_9180,In_1818,In_1702);
or U9181 (N_9181,In_2006,In_1274);
or U9182 (N_9182,In_2552,In_3930);
nand U9183 (N_9183,In_609,In_2727);
or U9184 (N_9184,In_1524,In_4457);
and U9185 (N_9185,In_4683,In_2947);
and U9186 (N_9186,In_4497,In_4482);
nor U9187 (N_9187,In_81,In_3872);
nor U9188 (N_9188,In_816,In_2151);
nand U9189 (N_9189,In_827,In_2685);
or U9190 (N_9190,In_830,In_2681);
or U9191 (N_9191,In_1064,In_957);
or U9192 (N_9192,In_4439,In_388);
or U9193 (N_9193,In_3907,In_96);
nand U9194 (N_9194,In_2643,In_923);
nor U9195 (N_9195,In_618,In_2892);
nand U9196 (N_9196,In_3612,In_4253);
and U9197 (N_9197,In_4814,In_993);
nor U9198 (N_9198,In_1411,In_4305);
nand U9199 (N_9199,In_2525,In_2112);
nor U9200 (N_9200,In_235,In_2401);
nor U9201 (N_9201,In_3758,In_691);
xor U9202 (N_9202,In_2660,In_4691);
or U9203 (N_9203,In_1158,In_407);
nor U9204 (N_9204,In_1663,In_1353);
nand U9205 (N_9205,In_4283,In_3014);
nor U9206 (N_9206,In_449,In_98);
or U9207 (N_9207,In_2333,In_4695);
and U9208 (N_9208,In_4897,In_3287);
nand U9209 (N_9209,In_3503,In_4695);
xor U9210 (N_9210,In_1314,In_2730);
or U9211 (N_9211,In_4102,In_923);
and U9212 (N_9212,In_4910,In_695);
nor U9213 (N_9213,In_135,In_3165);
and U9214 (N_9214,In_1366,In_4556);
and U9215 (N_9215,In_1500,In_4038);
xnor U9216 (N_9216,In_3460,In_2042);
and U9217 (N_9217,In_2710,In_3329);
and U9218 (N_9218,In_2126,In_3169);
xnor U9219 (N_9219,In_3285,In_4776);
nor U9220 (N_9220,In_90,In_1110);
nand U9221 (N_9221,In_2226,In_3729);
or U9222 (N_9222,In_3416,In_2536);
nor U9223 (N_9223,In_2209,In_2860);
nor U9224 (N_9224,In_4598,In_4596);
xnor U9225 (N_9225,In_2640,In_4358);
or U9226 (N_9226,In_1859,In_3747);
xnor U9227 (N_9227,In_3775,In_3197);
nor U9228 (N_9228,In_1219,In_4018);
nand U9229 (N_9229,In_3723,In_1844);
or U9230 (N_9230,In_364,In_1608);
or U9231 (N_9231,In_1733,In_2018);
nor U9232 (N_9232,In_370,In_4266);
nor U9233 (N_9233,In_476,In_3635);
and U9234 (N_9234,In_4464,In_184);
or U9235 (N_9235,In_4383,In_3814);
nor U9236 (N_9236,In_3863,In_1097);
and U9237 (N_9237,In_4692,In_4814);
nand U9238 (N_9238,In_174,In_626);
nand U9239 (N_9239,In_1696,In_3007);
nor U9240 (N_9240,In_277,In_3299);
nor U9241 (N_9241,In_1075,In_1451);
or U9242 (N_9242,In_1920,In_286);
and U9243 (N_9243,In_2431,In_2184);
and U9244 (N_9244,In_4182,In_2745);
nand U9245 (N_9245,In_4352,In_230);
nor U9246 (N_9246,In_2698,In_1852);
nand U9247 (N_9247,In_4674,In_523);
nand U9248 (N_9248,In_4468,In_3681);
nor U9249 (N_9249,In_3192,In_1166);
or U9250 (N_9250,In_1503,In_2881);
or U9251 (N_9251,In_3186,In_4938);
xnor U9252 (N_9252,In_875,In_301);
nand U9253 (N_9253,In_4842,In_1030);
nor U9254 (N_9254,In_657,In_2504);
nand U9255 (N_9255,In_4206,In_1039);
and U9256 (N_9256,In_4212,In_601);
nand U9257 (N_9257,In_100,In_3842);
nor U9258 (N_9258,In_3697,In_4566);
and U9259 (N_9259,In_3263,In_2091);
nor U9260 (N_9260,In_4902,In_2544);
or U9261 (N_9261,In_4251,In_637);
and U9262 (N_9262,In_3856,In_4352);
or U9263 (N_9263,In_910,In_1125);
nand U9264 (N_9264,In_2174,In_2052);
and U9265 (N_9265,In_3840,In_820);
and U9266 (N_9266,In_661,In_944);
nand U9267 (N_9267,In_4353,In_2772);
or U9268 (N_9268,In_1337,In_1589);
or U9269 (N_9269,In_2886,In_1814);
or U9270 (N_9270,In_853,In_4908);
nor U9271 (N_9271,In_2412,In_4551);
xnor U9272 (N_9272,In_3105,In_4749);
and U9273 (N_9273,In_3754,In_531);
nand U9274 (N_9274,In_4648,In_3049);
nor U9275 (N_9275,In_409,In_1257);
or U9276 (N_9276,In_4694,In_1728);
and U9277 (N_9277,In_3673,In_1014);
and U9278 (N_9278,In_4175,In_422);
xor U9279 (N_9279,In_1984,In_4753);
nand U9280 (N_9280,In_2653,In_2095);
nor U9281 (N_9281,In_433,In_2525);
nand U9282 (N_9282,In_1298,In_3732);
or U9283 (N_9283,In_542,In_2118);
nand U9284 (N_9284,In_3852,In_4102);
or U9285 (N_9285,In_2177,In_30);
nor U9286 (N_9286,In_4419,In_2499);
or U9287 (N_9287,In_3961,In_3229);
nand U9288 (N_9288,In_4265,In_2879);
or U9289 (N_9289,In_4046,In_3833);
or U9290 (N_9290,In_997,In_2568);
nand U9291 (N_9291,In_2369,In_2800);
or U9292 (N_9292,In_3381,In_4589);
nor U9293 (N_9293,In_1817,In_2313);
and U9294 (N_9294,In_1797,In_3723);
or U9295 (N_9295,In_3690,In_1561);
or U9296 (N_9296,In_3114,In_3457);
nor U9297 (N_9297,In_2769,In_4865);
nand U9298 (N_9298,In_3078,In_607);
xor U9299 (N_9299,In_1853,In_4906);
nor U9300 (N_9300,In_370,In_103);
or U9301 (N_9301,In_3174,In_2954);
nor U9302 (N_9302,In_4252,In_970);
or U9303 (N_9303,In_4012,In_3746);
xor U9304 (N_9304,In_1468,In_704);
nor U9305 (N_9305,In_3513,In_4639);
nand U9306 (N_9306,In_4418,In_2746);
xnor U9307 (N_9307,In_2728,In_598);
and U9308 (N_9308,In_3304,In_2850);
and U9309 (N_9309,In_2286,In_202);
and U9310 (N_9310,In_2212,In_356);
nor U9311 (N_9311,In_3128,In_3230);
nor U9312 (N_9312,In_1360,In_2485);
or U9313 (N_9313,In_1837,In_2194);
nand U9314 (N_9314,In_311,In_1378);
or U9315 (N_9315,In_4213,In_3282);
nand U9316 (N_9316,In_1539,In_322);
nor U9317 (N_9317,In_4438,In_3640);
xor U9318 (N_9318,In_4395,In_2113);
and U9319 (N_9319,In_1011,In_638);
nand U9320 (N_9320,In_431,In_4725);
nand U9321 (N_9321,In_1656,In_4274);
nand U9322 (N_9322,In_539,In_2213);
nor U9323 (N_9323,In_2777,In_4014);
nand U9324 (N_9324,In_2380,In_3813);
nor U9325 (N_9325,In_2620,In_1405);
nor U9326 (N_9326,In_2958,In_1518);
nor U9327 (N_9327,In_6,In_3666);
or U9328 (N_9328,In_2157,In_2673);
xnor U9329 (N_9329,In_1670,In_2551);
and U9330 (N_9330,In_1335,In_4336);
or U9331 (N_9331,In_3757,In_1878);
nand U9332 (N_9332,In_3912,In_2843);
and U9333 (N_9333,In_2738,In_884);
nand U9334 (N_9334,In_486,In_2380);
nand U9335 (N_9335,In_346,In_1688);
nand U9336 (N_9336,In_1127,In_2954);
and U9337 (N_9337,In_2322,In_2191);
or U9338 (N_9338,In_43,In_2357);
and U9339 (N_9339,In_2758,In_413);
and U9340 (N_9340,In_4126,In_2831);
nor U9341 (N_9341,In_2507,In_3132);
nor U9342 (N_9342,In_3479,In_3016);
and U9343 (N_9343,In_3539,In_2561);
and U9344 (N_9344,In_2526,In_933);
nor U9345 (N_9345,In_2159,In_858);
xnor U9346 (N_9346,In_1815,In_2501);
nand U9347 (N_9347,In_233,In_3745);
nor U9348 (N_9348,In_3888,In_4185);
or U9349 (N_9349,In_1836,In_3774);
or U9350 (N_9350,In_380,In_2291);
xor U9351 (N_9351,In_3352,In_3315);
nand U9352 (N_9352,In_3007,In_3312);
xnor U9353 (N_9353,In_3351,In_2170);
nor U9354 (N_9354,In_1829,In_1662);
xnor U9355 (N_9355,In_3908,In_4691);
and U9356 (N_9356,In_2722,In_4929);
or U9357 (N_9357,In_2753,In_3571);
and U9358 (N_9358,In_4588,In_212);
and U9359 (N_9359,In_1160,In_540);
nor U9360 (N_9360,In_1066,In_2960);
and U9361 (N_9361,In_842,In_4560);
nor U9362 (N_9362,In_951,In_1731);
nor U9363 (N_9363,In_2728,In_1300);
nand U9364 (N_9364,In_2412,In_115);
nand U9365 (N_9365,In_4793,In_1148);
nand U9366 (N_9366,In_2598,In_4330);
nand U9367 (N_9367,In_4049,In_1529);
nand U9368 (N_9368,In_149,In_2164);
nor U9369 (N_9369,In_2809,In_1708);
nor U9370 (N_9370,In_4456,In_2928);
and U9371 (N_9371,In_3673,In_900);
and U9372 (N_9372,In_144,In_1879);
nor U9373 (N_9373,In_776,In_1654);
nand U9374 (N_9374,In_361,In_218);
xor U9375 (N_9375,In_235,In_678);
and U9376 (N_9376,In_1436,In_2410);
and U9377 (N_9377,In_3122,In_2919);
or U9378 (N_9378,In_4005,In_452);
or U9379 (N_9379,In_3240,In_2090);
nor U9380 (N_9380,In_2337,In_1486);
or U9381 (N_9381,In_244,In_3323);
or U9382 (N_9382,In_1422,In_3522);
and U9383 (N_9383,In_3272,In_2825);
nand U9384 (N_9384,In_3241,In_4296);
and U9385 (N_9385,In_2178,In_2338);
and U9386 (N_9386,In_4360,In_2452);
xor U9387 (N_9387,In_1469,In_984);
nand U9388 (N_9388,In_1647,In_4144);
nand U9389 (N_9389,In_159,In_600);
or U9390 (N_9390,In_4084,In_4580);
nor U9391 (N_9391,In_1348,In_726);
nand U9392 (N_9392,In_3737,In_2475);
nand U9393 (N_9393,In_77,In_1148);
nor U9394 (N_9394,In_1217,In_866);
and U9395 (N_9395,In_4763,In_1302);
nor U9396 (N_9396,In_4012,In_3797);
and U9397 (N_9397,In_1015,In_1636);
nor U9398 (N_9398,In_1819,In_1284);
and U9399 (N_9399,In_1145,In_1576);
and U9400 (N_9400,In_2257,In_2256);
nor U9401 (N_9401,In_2422,In_3020);
nor U9402 (N_9402,In_3589,In_2155);
nor U9403 (N_9403,In_2663,In_1931);
or U9404 (N_9404,In_3560,In_2595);
nand U9405 (N_9405,In_3718,In_1572);
and U9406 (N_9406,In_886,In_55);
xor U9407 (N_9407,In_2745,In_1238);
or U9408 (N_9408,In_4725,In_1920);
xnor U9409 (N_9409,In_2156,In_2354);
and U9410 (N_9410,In_4559,In_2725);
and U9411 (N_9411,In_2700,In_685);
or U9412 (N_9412,In_2431,In_2745);
or U9413 (N_9413,In_3020,In_898);
xnor U9414 (N_9414,In_1091,In_1115);
or U9415 (N_9415,In_3409,In_2948);
nand U9416 (N_9416,In_1510,In_355);
nor U9417 (N_9417,In_536,In_2656);
nand U9418 (N_9418,In_3577,In_1239);
nor U9419 (N_9419,In_4435,In_4080);
and U9420 (N_9420,In_3992,In_1990);
and U9421 (N_9421,In_4646,In_2437);
or U9422 (N_9422,In_2114,In_3564);
and U9423 (N_9423,In_626,In_3546);
nor U9424 (N_9424,In_1897,In_2096);
or U9425 (N_9425,In_451,In_69);
or U9426 (N_9426,In_782,In_1618);
xor U9427 (N_9427,In_630,In_1306);
and U9428 (N_9428,In_157,In_656);
nand U9429 (N_9429,In_2726,In_1415);
nand U9430 (N_9430,In_1024,In_2585);
nor U9431 (N_9431,In_3999,In_3022);
or U9432 (N_9432,In_3007,In_2276);
or U9433 (N_9433,In_4109,In_4276);
nand U9434 (N_9434,In_1134,In_4665);
and U9435 (N_9435,In_1876,In_1191);
nor U9436 (N_9436,In_1246,In_3284);
and U9437 (N_9437,In_4158,In_4524);
and U9438 (N_9438,In_4563,In_3424);
nor U9439 (N_9439,In_3085,In_2014);
or U9440 (N_9440,In_33,In_3454);
or U9441 (N_9441,In_4804,In_2668);
and U9442 (N_9442,In_4844,In_1073);
nor U9443 (N_9443,In_1774,In_1729);
or U9444 (N_9444,In_2106,In_2000);
and U9445 (N_9445,In_2676,In_3239);
nand U9446 (N_9446,In_3403,In_256);
and U9447 (N_9447,In_866,In_498);
nand U9448 (N_9448,In_3949,In_4735);
or U9449 (N_9449,In_1633,In_3602);
nor U9450 (N_9450,In_1216,In_4072);
and U9451 (N_9451,In_108,In_3080);
and U9452 (N_9452,In_448,In_3185);
xor U9453 (N_9453,In_3313,In_1237);
or U9454 (N_9454,In_1488,In_1794);
or U9455 (N_9455,In_1068,In_2439);
nand U9456 (N_9456,In_4857,In_596);
nor U9457 (N_9457,In_4713,In_2021);
nand U9458 (N_9458,In_2273,In_3070);
nand U9459 (N_9459,In_2945,In_3969);
and U9460 (N_9460,In_3286,In_2026);
or U9461 (N_9461,In_2231,In_1368);
nor U9462 (N_9462,In_3229,In_4230);
nand U9463 (N_9463,In_3954,In_4815);
nand U9464 (N_9464,In_3774,In_1956);
nand U9465 (N_9465,In_407,In_47);
xor U9466 (N_9466,In_4295,In_272);
nor U9467 (N_9467,In_1758,In_4960);
nor U9468 (N_9468,In_2205,In_1690);
and U9469 (N_9469,In_1421,In_126);
or U9470 (N_9470,In_2853,In_1049);
xnor U9471 (N_9471,In_79,In_3202);
nand U9472 (N_9472,In_3997,In_1510);
or U9473 (N_9473,In_1717,In_2001);
nand U9474 (N_9474,In_384,In_997);
xor U9475 (N_9475,In_2494,In_4274);
nand U9476 (N_9476,In_2211,In_4303);
nand U9477 (N_9477,In_2120,In_2840);
or U9478 (N_9478,In_2320,In_1117);
nand U9479 (N_9479,In_4581,In_1357);
nand U9480 (N_9480,In_2988,In_2058);
nand U9481 (N_9481,In_4003,In_4911);
nand U9482 (N_9482,In_4168,In_3970);
xnor U9483 (N_9483,In_4973,In_2255);
nor U9484 (N_9484,In_4535,In_981);
nor U9485 (N_9485,In_646,In_4969);
nand U9486 (N_9486,In_1692,In_4581);
or U9487 (N_9487,In_841,In_580);
nor U9488 (N_9488,In_1906,In_1417);
nor U9489 (N_9489,In_3896,In_345);
nand U9490 (N_9490,In_2814,In_509);
or U9491 (N_9491,In_3479,In_1021);
and U9492 (N_9492,In_2221,In_3982);
nand U9493 (N_9493,In_4693,In_2723);
and U9494 (N_9494,In_1867,In_918);
xnor U9495 (N_9495,In_845,In_582);
nand U9496 (N_9496,In_2131,In_3463);
nand U9497 (N_9497,In_2709,In_4143);
nand U9498 (N_9498,In_1649,In_4520);
nor U9499 (N_9499,In_2396,In_2354);
nand U9500 (N_9500,In_4637,In_3108);
and U9501 (N_9501,In_776,In_1623);
or U9502 (N_9502,In_3638,In_4596);
or U9503 (N_9503,In_4390,In_2327);
and U9504 (N_9504,In_4401,In_1632);
and U9505 (N_9505,In_2263,In_2261);
or U9506 (N_9506,In_4351,In_806);
or U9507 (N_9507,In_1156,In_286);
nand U9508 (N_9508,In_4651,In_1440);
or U9509 (N_9509,In_1134,In_1764);
nand U9510 (N_9510,In_1457,In_3965);
nand U9511 (N_9511,In_4788,In_1136);
nor U9512 (N_9512,In_2390,In_2078);
or U9513 (N_9513,In_144,In_2405);
nand U9514 (N_9514,In_4770,In_1476);
or U9515 (N_9515,In_1312,In_2029);
nor U9516 (N_9516,In_3974,In_925);
and U9517 (N_9517,In_4595,In_1100);
nor U9518 (N_9518,In_8,In_2725);
nor U9519 (N_9519,In_2919,In_2429);
xor U9520 (N_9520,In_4465,In_3409);
or U9521 (N_9521,In_2047,In_4675);
nor U9522 (N_9522,In_2640,In_1413);
xor U9523 (N_9523,In_4233,In_1332);
or U9524 (N_9524,In_4237,In_4956);
xnor U9525 (N_9525,In_1437,In_3973);
nor U9526 (N_9526,In_1692,In_4990);
nand U9527 (N_9527,In_1646,In_882);
or U9528 (N_9528,In_4218,In_3575);
or U9529 (N_9529,In_2507,In_557);
or U9530 (N_9530,In_3963,In_247);
xor U9531 (N_9531,In_602,In_3204);
nand U9532 (N_9532,In_1283,In_2928);
nand U9533 (N_9533,In_1053,In_4933);
nand U9534 (N_9534,In_2973,In_4720);
or U9535 (N_9535,In_385,In_3983);
xor U9536 (N_9536,In_4281,In_143);
or U9537 (N_9537,In_2292,In_2975);
nor U9538 (N_9538,In_3764,In_3956);
or U9539 (N_9539,In_4082,In_891);
nor U9540 (N_9540,In_2853,In_4093);
and U9541 (N_9541,In_1813,In_3743);
nand U9542 (N_9542,In_3164,In_464);
nand U9543 (N_9543,In_2422,In_514);
nor U9544 (N_9544,In_3694,In_4870);
xnor U9545 (N_9545,In_1139,In_1822);
and U9546 (N_9546,In_3104,In_4100);
or U9547 (N_9547,In_4453,In_1131);
and U9548 (N_9548,In_3041,In_1073);
nand U9549 (N_9549,In_229,In_204);
nand U9550 (N_9550,In_64,In_3889);
nand U9551 (N_9551,In_302,In_4321);
nor U9552 (N_9552,In_1607,In_2625);
nand U9553 (N_9553,In_1954,In_3484);
xor U9554 (N_9554,In_3327,In_4186);
nor U9555 (N_9555,In_639,In_4846);
or U9556 (N_9556,In_434,In_3460);
nand U9557 (N_9557,In_2080,In_2609);
nand U9558 (N_9558,In_1867,In_531);
nor U9559 (N_9559,In_3682,In_1399);
or U9560 (N_9560,In_3727,In_2787);
nor U9561 (N_9561,In_1929,In_3945);
and U9562 (N_9562,In_1826,In_4329);
nor U9563 (N_9563,In_4757,In_1307);
and U9564 (N_9564,In_1414,In_2446);
and U9565 (N_9565,In_3916,In_2712);
nand U9566 (N_9566,In_1916,In_2083);
nand U9567 (N_9567,In_2457,In_2126);
nand U9568 (N_9568,In_2978,In_3621);
nor U9569 (N_9569,In_4464,In_2394);
and U9570 (N_9570,In_3097,In_732);
nor U9571 (N_9571,In_4063,In_4132);
or U9572 (N_9572,In_4987,In_1595);
or U9573 (N_9573,In_4287,In_4493);
nor U9574 (N_9574,In_91,In_435);
or U9575 (N_9575,In_3655,In_881);
nor U9576 (N_9576,In_4558,In_3600);
xnor U9577 (N_9577,In_3449,In_3758);
nand U9578 (N_9578,In_75,In_3755);
nor U9579 (N_9579,In_2559,In_2028);
nand U9580 (N_9580,In_3644,In_2149);
and U9581 (N_9581,In_2370,In_2880);
nand U9582 (N_9582,In_2207,In_2411);
nor U9583 (N_9583,In_65,In_794);
nand U9584 (N_9584,In_623,In_1590);
nor U9585 (N_9585,In_1974,In_2246);
nand U9586 (N_9586,In_1208,In_144);
or U9587 (N_9587,In_3891,In_1329);
nor U9588 (N_9588,In_467,In_3026);
nor U9589 (N_9589,In_4111,In_1496);
or U9590 (N_9590,In_4092,In_574);
nand U9591 (N_9591,In_2031,In_924);
nor U9592 (N_9592,In_2850,In_643);
nor U9593 (N_9593,In_1355,In_4074);
or U9594 (N_9594,In_4143,In_3976);
or U9595 (N_9595,In_2764,In_1528);
and U9596 (N_9596,In_4565,In_4502);
nor U9597 (N_9597,In_2543,In_2437);
or U9598 (N_9598,In_2650,In_2301);
or U9599 (N_9599,In_3077,In_4746);
nand U9600 (N_9600,In_4711,In_1265);
and U9601 (N_9601,In_322,In_2397);
nor U9602 (N_9602,In_3756,In_277);
or U9603 (N_9603,In_1313,In_1375);
nand U9604 (N_9604,In_3789,In_1867);
nor U9605 (N_9605,In_1306,In_3222);
nor U9606 (N_9606,In_4981,In_2441);
nand U9607 (N_9607,In_1648,In_13);
xnor U9608 (N_9608,In_1070,In_999);
or U9609 (N_9609,In_4866,In_3419);
and U9610 (N_9610,In_35,In_2064);
or U9611 (N_9611,In_631,In_1262);
or U9612 (N_9612,In_1248,In_4839);
nor U9613 (N_9613,In_3050,In_4019);
nor U9614 (N_9614,In_1019,In_1276);
or U9615 (N_9615,In_3451,In_4670);
and U9616 (N_9616,In_4803,In_836);
xor U9617 (N_9617,In_3713,In_190);
nor U9618 (N_9618,In_2955,In_3808);
or U9619 (N_9619,In_4185,In_2828);
xor U9620 (N_9620,In_3647,In_2877);
xor U9621 (N_9621,In_1332,In_4409);
and U9622 (N_9622,In_1283,In_1448);
nand U9623 (N_9623,In_2439,In_990);
and U9624 (N_9624,In_2652,In_1579);
nand U9625 (N_9625,In_4967,In_1509);
nand U9626 (N_9626,In_2880,In_3109);
nand U9627 (N_9627,In_3584,In_2978);
or U9628 (N_9628,In_1590,In_703);
nor U9629 (N_9629,In_4823,In_1935);
xor U9630 (N_9630,In_535,In_1293);
or U9631 (N_9631,In_2303,In_4146);
xor U9632 (N_9632,In_1246,In_1622);
nand U9633 (N_9633,In_4260,In_1629);
xor U9634 (N_9634,In_930,In_523);
or U9635 (N_9635,In_353,In_1576);
nor U9636 (N_9636,In_2481,In_3625);
or U9637 (N_9637,In_4777,In_4731);
and U9638 (N_9638,In_2476,In_381);
and U9639 (N_9639,In_3331,In_847);
nand U9640 (N_9640,In_2734,In_3060);
or U9641 (N_9641,In_2666,In_854);
xnor U9642 (N_9642,In_449,In_499);
nand U9643 (N_9643,In_1328,In_4505);
or U9644 (N_9644,In_4077,In_3438);
or U9645 (N_9645,In_503,In_946);
nand U9646 (N_9646,In_4668,In_2458);
nand U9647 (N_9647,In_1762,In_886);
or U9648 (N_9648,In_3567,In_4797);
or U9649 (N_9649,In_3965,In_4547);
and U9650 (N_9650,In_439,In_1949);
nand U9651 (N_9651,In_342,In_3561);
xor U9652 (N_9652,In_2161,In_3995);
and U9653 (N_9653,In_3615,In_4608);
nor U9654 (N_9654,In_1334,In_2139);
xnor U9655 (N_9655,In_4484,In_4037);
or U9656 (N_9656,In_3544,In_3455);
nand U9657 (N_9657,In_3141,In_1482);
or U9658 (N_9658,In_3640,In_3288);
nand U9659 (N_9659,In_521,In_3480);
and U9660 (N_9660,In_3101,In_487);
or U9661 (N_9661,In_2292,In_4267);
nand U9662 (N_9662,In_4240,In_1364);
or U9663 (N_9663,In_4353,In_4703);
and U9664 (N_9664,In_382,In_2700);
or U9665 (N_9665,In_4787,In_2978);
xor U9666 (N_9666,In_193,In_1443);
and U9667 (N_9667,In_508,In_1379);
or U9668 (N_9668,In_4455,In_4906);
or U9669 (N_9669,In_4225,In_1960);
xnor U9670 (N_9670,In_1422,In_492);
nor U9671 (N_9671,In_2038,In_4665);
and U9672 (N_9672,In_2806,In_2844);
or U9673 (N_9673,In_426,In_3962);
xor U9674 (N_9674,In_4822,In_1250);
nor U9675 (N_9675,In_2687,In_352);
or U9676 (N_9676,In_4193,In_3395);
or U9677 (N_9677,In_4210,In_4870);
and U9678 (N_9678,In_3701,In_781);
and U9679 (N_9679,In_1685,In_4307);
xnor U9680 (N_9680,In_4754,In_3755);
and U9681 (N_9681,In_2787,In_2076);
and U9682 (N_9682,In_2294,In_2752);
nor U9683 (N_9683,In_872,In_1442);
or U9684 (N_9684,In_4582,In_28);
and U9685 (N_9685,In_3588,In_1747);
and U9686 (N_9686,In_4447,In_2278);
nand U9687 (N_9687,In_4899,In_4973);
or U9688 (N_9688,In_30,In_1133);
or U9689 (N_9689,In_90,In_1465);
and U9690 (N_9690,In_4879,In_3227);
or U9691 (N_9691,In_4223,In_3747);
or U9692 (N_9692,In_4480,In_570);
nor U9693 (N_9693,In_1291,In_3237);
and U9694 (N_9694,In_4182,In_4266);
nand U9695 (N_9695,In_2041,In_992);
nor U9696 (N_9696,In_2944,In_1531);
nor U9697 (N_9697,In_1527,In_1733);
or U9698 (N_9698,In_2539,In_1509);
and U9699 (N_9699,In_2567,In_2162);
xor U9700 (N_9700,In_386,In_1695);
nand U9701 (N_9701,In_300,In_298);
nand U9702 (N_9702,In_1402,In_1760);
nand U9703 (N_9703,In_4037,In_4215);
and U9704 (N_9704,In_1234,In_4288);
nor U9705 (N_9705,In_89,In_3109);
nor U9706 (N_9706,In_4925,In_4396);
nor U9707 (N_9707,In_3766,In_4868);
nor U9708 (N_9708,In_4885,In_3537);
nand U9709 (N_9709,In_1029,In_3486);
nand U9710 (N_9710,In_4753,In_3533);
nor U9711 (N_9711,In_3746,In_384);
and U9712 (N_9712,In_1916,In_3094);
and U9713 (N_9713,In_309,In_3048);
and U9714 (N_9714,In_1086,In_1534);
and U9715 (N_9715,In_4267,In_4941);
and U9716 (N_9716,In_4308,In_4863);
or U9717 (N_9717,In_4627,In_1117);
nor U9718 (N_9718,In_2990,In_2948);
or U9719 (N_9719,In_1912,In_714);
nand U9720 (N_9720,In_2071,In_2364);
nor U9721 (N_9721,In_542,In_2636);
and U9722 (N_9722,In_1391,In_1914);
nor U9723 (N_9723,In_2066,In_2062);
and U9724 (N_9724,In_4097,In_2346);
or U9725 (N_9725,In_2285,In_2014);
xnor U9726 (N_9726,In_4898,In_3910);
and U9727 (N_9727,In_3370,In_2421);
nor U9728 (N_9728,In_2286,In_3069);
nor U9729 (N_9729,In_1633,In_2700);
xor U9730 (N_9730,In_2418,In_4484);
nand U9731 (N_9731,In_4736,In_1691);
nand U9732 (N_9732,In_4643,In_2034);
and U9733 (N_9733,In_2101,In_1646);
nor U9734 (N_9734,In_4156,In_1047);
nand U9735 (N_9735,In_3030,In_2620);
and U9736 (N_9736,In_1249,In_4516);
nand U9737 (N_9737,In_3852,In_4853);
or U9738 (N_9738,In_284,In_951);
and U9739 (N_9739,In_2456,In_1332);
and U9740 (N_9740,In_830,In_1250);
or U9741 (N_9741,In_808,In_3428);
and U9742 (N_9742,In_804,In_2872);
nor U9743 (N_9743,In_3099,In_2577);
xor U9744 (N_9744,In_3717,In_1650);
or U9745 (N_9745,In_3964,In_4122);
nor U9746 (N_9746,In_519,In_576);
nand U9747 (N_9747,In_2277,In_1365);
and U9748 (N_9748,In_3974,In_375);
and U9749 (N_9749,In_977,In_1171);
and U9750 (N_9750,In_2036,In_1140);
nor U9751 (N_9751,In_2183,In_1996);
nor U9752 (N_9752,In_2189,In_3977);
nor U9753 (N_9753,In_4740,In_2942);
nor U9754 (N_9754,In_2408,In_1536);
nand U9755 (N_9755,In_3076,In_3684);
or U9756 (N_9756,In_241,In_1444);
nor U9757 (N_9757,In_1608,In_2362);
xnor U9758 (N_9758,In_948,In_4626);
nor U9759 (N_9759,In_2034,In_1374);
nor U9760 (N_9760,In_1852,In_4414);
nor U9761 (N_9761,In_4265,In_4572);
nor U9762 (N_9762,In_2662,In_506);
nor U9763 (N_9763,In_4832,In_3007);
xor U9764 (N_9764,In_1347,In_2979);
or U9765 (N_9765,In_4209,In_688);
or U9766 (N_9766,In_3205,In_4913);
nand U9767 (N_9767,In_469,In_1299);
nor U9768 (N_9768,In_1556,In_1422);
nor U9769 (N_9769,In_3731,In_656);
or U9770 (N_9770,In_2149,In_3918);
nand U9771 (N_9771,In_3396,In_4768);
and U9772 (N_9772,In_2606,In_3372);
nor U9773 (N_9773,In_4217,In_3387);
nor U9774 (N_9774,In_3331,In_1252);
and U9775 (N_9775,In_2146,In_342);
nor U9776 (N_9776,In_5,In_1386);
or U9777 (N_9777,In_4717,In_1700);
and U9778 (N_9778,In_1480,In_2825);
nand U9779 (N_9779,In_275,In_2244);
or U9780 (N_9780,In_2095,In_3160);
nand U9781 (N_9781,In_3140,In_2956);
and U9782 (N_9782,In_4258,In_4187);
or U9783 (N_9783,In_3136,In_2627);
nor U9784 (N_9784,In_4845,In_1950);
or U9785 (N_9785,In_3762,In_1218);
nand U9786 (N_9786,In_2725,In_1532);
xor U9787 (N_9787,In_4314,In_1664);
and U9788 (N_9788,In_4911,In_2211);
nand U9789 (N_9789,In_298,In_4399);
nor U9790 (N_9790,In_152,In_282);
xor U9791 (N_9791,In_1148,In_1548);
or U9792 (N_9792,In_221,In_1185);
nand U9793 (N_9793,In_1497,In_4005);
xnor U9794 (N_9794,In_1137,In_2196);
xnor U9795 (N_9795,In_3802,In_1990);
xnor U9796 (N_9796,In_2914,In_4225);
xnor U9797 (N_9797,In_4632,In_927);
nor U9798 (N_9798,In_3191,In_473);
xor U9799 (N_9799,In_2399,In_4675);
nor U9800 (N_9800,In_4444,In_454);
and U9801 (N_9801,In_2033,In_4929);
nor U9802 (N_9802,In_4336,In_4380);
and U9803 (N_9803,In_1055,In_2612);
nor U9804 (N_9804,In_1512,In_3999);
and U9805 (N_9805,In_3210,In_2494);
xor U9806 (N_9806,In_3008,In_3854);
and U9807 (N_9807,In_4848,In_3660);
or U9808 (N_9808,In_1161,In_4758);
and U9809 (N_9809,In_1259,In_4677);
and U9810 (N_9810,In_4461,In_1258);
and U9811 (N_9811,In_3742,In_4403);
or U9812 (N_9812,In_2914,In_142);
nor U9813 (N_9813,In_4035,In_1043);
nand U9814 (N_9814,In_4092,In_1995);
nand U9815 (N_9815,In_4557,In_3975);
nor U9816 (N_9816,In_4551,In_271);
and U9817 (N_9817,In_2012,In_3543);
and U9818 (N_9818,In_2977,In_2952);
nor U9819 (N_9819,In_4809,In_2998);
or U9820 (N_9820,In_2993,In_895);
nor U9821 (N_9821,In_3398,In_2610);
or U9822 (N_9822,In_1617,In_1993);
nor U9823 (N_9823,In_1628,In_1077);
xnor U9824 (N_9824,In_3546,In_1991);
or U9825 (N_9825,In_1826,In_3803);
nor U9826 (N_9826,In_1386,In_659);
nand U9827 (N_9827,In_4612,In_2938);
nand U9828 (N_9828,In_949,In_3345);
and U9829 (N_9829,In_3237,In_1089);
nand U9830 (N_9830,In_1146,In_3014);
nand U9831 (N_9831,In_4908,In_4937);
nand U9832 (N_9832,In_3498,In_3757);
nand U9833 (N_9833,In_510,In_1500);
nand U9834 (N_9834,In_2461,In_220);
nor U9835 (N_9835,In_4913,In_2991);
nor U9836 (N_9836,In_750,In_3834);
nand U9837 (N_9837,In_1890,In_2711);
nor U9838 (N_9838,In_4960,In_3117);
nor U9839 (N_9839,In_2178,In_4544);
xnor U9840 (N_9840,In_835,In_1632);
nor U9841 (N_9841,In_165,In_3913);
nor U9842 (N_9842,In_33,In_3538);
nor U9843 (N_9843,In_2082,In_2055);
xnor U9844 (N_9844,In_1886,In_90);
or U9845 (N_9845,In_2011,In_1290);
or U9846 (N_9846,In_3327,In_41);
nand U9847 (N_9847,In_4872,In_1495);
and U9848 (N_9848,In_4075,In_3004);
nand U9849 (N_9849,In_703,In_1643);
xnor U9850 (N_9850,In_4455,In_737);
nor U9851 (N_9851,In_3762,In_1509);
nand U9852 (N_9852,In_3384,In_2865);
nor U9853 (N_9853,In_3865,In_686);
nor U9854 (N_9854,In_340,In_504);
and U9855 (N_9855,In_3202,In_3295);
or U9856 (N_9856,In_1916,In_4414);
and U9857 (N_9857,In_3762,In_2921);
nor U9858 (N_9858,In_1039,In_2422);
nand U9859 (N_9859,In_4911,In_1788);
nor U9860 (N_9860,In_2367,In_431);
and U9861 (N_9861,In_2851,In_2039);
or U9862 (N_9862,In_2180,In_2809);
or U9863 (N_9863,In_185,In_2430);
or U9864 (N_9864,In_3296,In_1035);
nor U9865 (N_9865,In_512,In_1137);
nor U9866 (N_9866,In_3115,In_3627);
xnor U9867 (N_9867,In_1279,In_1165);
nor U9868 (N_9868,In_4061,In_3562);
or U9869 (N_9869,In_4876,In_610);
nand U9870 (N_9870,In_3528,In_393);
nand U9871 (N_9871,In_4347,In_1736);
xor U9872 (N_9872,In_1832,In_2686);
nor U9873 (N_9873,In_3236,In_652);
and U9874 (N_9874,In_4037,In_1507);
nor U9875 (N_9875,In_375,In_2275);
nand U9876 (N_9876,In_2019,In_1374);
nand U9877 (N_9877,In_2094,In_1184);
and U9878 (N_9878,In_774,In_3576);
xor U9879 (N_9879,In_182,In_3684);
or U9880 (N_9880,In_3848,In_470);
nor U9881 (N_9881,In_3158,In_2727);
xnor U9882 (N_9882,In_4098,In_4725);
nor U9883 (N_9883,In_2137,In_707);
nor U9884 (N_9884,In_389,In_4154);
and U9885 (N_9885,In_124,In_964);
nor U9886 (N_9886,In_3630,In_4161);
and U9887 (N_9887,In_2116,In_4794);
nand U9888 (N_9888,In_257,In_1115);
nand U9889 (N_9889,In_1864,In_2242);
or U9890 (N_9890,In_2318,In_3947);
or U9891 (N_9891,In_1936,In_2767);
nor U9892 (N_9892,In_2989,In_4309);
and U9893 (N_9893,In_2900,In_1614);
nand U9894 (N_9894,In_2167,In_4328);
nand U9895 (N_9895,In_2095,In_1223);
or U9896 (N_9896,In_2327,In_2873);
and U9897 (N_9897,In_2858,In_1617);
and U9898 (N_9898,In_2854,In_4286);
and U9899 (N_9899,In_358,In_2016);
nand U9900 (N_9900,In_3481,In_2742);
nor U9901 (N_9901,In_1322,In_2409);
and U9902 (N_9902,In_1423,In_4217);
or U9903 (N_9903,In_3539,In_2387);
nand U9904 (N_9904,In_2191,In_1462);
and U9905 (N_9905,In_946,In_357);
nor U9906 (N_9906,In_2738,In_2804);
and U9907 (N_9907,In_2040,In_451);
and U9908 (N_9908,In_1270,In_1231);
and U9909 (N_9909,In_4605,In_183);
xor U9910 (N_9910,In_4050,In_3355);
nand U9911 (N_9911,In_2789,In_400);
xnor U9912 (N_9912,In_664,In_4378);
or U9913 (N_9913,In_4566,In_398);
nor U9914 (N_9914,In_3577,In_4057);
or U9915 (N_9915,In_4128,In_648);
or U9916 (N_9916,In_465,In_2694);
and U9917 (N_9917,In_4705,In_3349);
nor U9918 (N_9918,In_3469,In_1464);
nand U9919 (N_9919,In_4463,In_1079);
nor U9920 (N_9920,In_2357,In_3652);
and U9921 (N_9921,In_4507,In_4943);
and U9922 (N_9922,In_2541,In_4950);
and U9923 (N_9923,In_4434,In_1470);
and U9924 (N_9924,In_1401,In_993);
and U9925 (N_9925,In_4007,In_3956);
and U9926 (N_9926,In_4283,In_1569);
nand U9927 (N_9927,In_3922,In_346);
nand U9928 (N_9928,In_4523,In_1066);
nand U9929 (N_9929,In_329,In_2545);
nand U9930 (N_9930,In_3451,In_4572);
nor U9931 (N_9931,In_3065,In_2132);
nor U9932 (N_9932,In_4451,In_937);
or U9933 (N_9933,In_1970,In_3931);
xor U9934 (N_9934,In_1764,In_2108);
nor U9935 (N_9935,In_121,In_4712);
or U9936 (N_9936,In_705,In_643);
and U9937 (N_9937,In_3544,In_2022);
nand U9938 (N_9938,In_4823,In_3368);
nand U9939 (N_9939,In_362,In_3733);
or U9940 (N_9940,In_488,In_2571);
nor U9941 (N_9941,In_4776,In_2391);
and U9942 (N_9942,In_1065,In_2951);
nand U9943 (N_9943,In_4567,In_2065);
or U9944 (N_9944,In_2987,In_131);
xor U9945 (N_9945,In_3367,In_348);
nand U9946 (N_9946,In_233,In_4986);
or U9947 (N_9947,In_353,In_2711);
nand U9948 (N_9948,In_4422,In_4170);
and U9949 (N_9949,In_4271,In_2718);
xnor U9950 (N_9950,In_3650,In_1686);
nor U9951 (N_9951,In_2730,In_3990);
and U9952 (N_9952,In_652,In_1157);
nor U9953 (N_9953,In_4705,In_4993);
nor U9954 (N_9954,In_3469,In_5);
nand U9955 (N_9955,In_2863,In_2846);
and U9956 (N_9956,In_4007,In_1416);
or U9957 (N_9957,In_3701,In_4556);
nand U9958 (N_9958,In_4884,In_1260);
nand U9959 (N_9959,In_3306,In_1109);
nor U9960 (N_9960,In_2633,In_2792);
nand U9961 (N_9961,In_1421,In_2972);
nand U9962 (N_9962,In_2796,In_3498);
nor U9963 (N_9963,In_274,In_914);
and U9964 (N_9964,In_1480,In_2974);
and U9965 (N_9965,In_4357,In_3832);
or U9966 (N_9966,In_669,In_1738);
or U9967 (N_9967,In_4429,In_2666);
nor U9968 (N_9968,In_3456,In_1180);
and U9969 (N_9969,In_4243,In_4831);
nor U9970 (N_9970,In_1036,In_1509);
nand U9971 (N_9971,In_4978,In_4772);
nand U9972 (N_9972,In_70,In_2582);
and U9973 (N_9973,In_4122,In_3131);
or U9974 (N_9974,In_3182,In_595);
xor U9975 (N_9975,In_3060,In_2526);
or U9976 (N_9976,In_1682,In_4858);
nor U9977 (N_9977,In_1523,In_3294);
nand U9978 (N_9978,In_742,In_1427);
nand U9979 (N_9979,In_3846,In_3012);
or U9980 (N_9980,In_2425,In_4890);
nor U9981 (N_9981,In_3206,In_2721);
and U9982 (N_9982,In_223,In_469);
and U9983 (N_9983,In_3390,In_4359);
nor U9984 (N_9984,In_3503,In_859);
nor U9985 (N_9985,In_1182,In_2693);
xnor U9986 (N_9986,In_2202,In_2310);
nor U9987 (N_9987,In_4820,In_420);
and U9988 (N_9988,In_934,In_2356);
nor U9989 (N_9989,In_4861,In_3677);
or U9990 (N_9990,In_629,In_1505);
or U9991 (N_9991,In_1194,In_1189);
or U9992 (N_9992,In_4137,In_3216);
xor U9993 (N_9993,In_1684,In_1375);
xor U9994 (N_9994,In_1018,In_2152);
and U9995 (N_9995,In_1819,In_3053);
xnor U9996 (N_9996,In_3384,In_510);
xnor U9997 (N_9997,In_1994,In_3142);
or U9998 (N_9998,In_4034,In_389);
nand U9999 (N_9999,In_2918,In_4238);
nand U10000 (N_10000,N_4906,N_1629);
and U10001 (N_10001,N_7292,N_7863);
or U10002 (N_10002,N_7991,N_4054);
nor U10003 (N_10003,N_6384,N_4646);
or U10004 (N_10004,N_9936,N_6105);
and U10005 (N_10005,N_2340,N_4868);
or U10006 (N_10006,N_2979,N_3968);
nor U10007 (N_10007,N_1813,N_5559);
or U10008 (N_10008,N_9189,N_4071);
and U10009 (N_10009,N_2885,N_2085);
or U10010 (N_10010,N_6466,N_4376);
xnor U10011 (N_10011,N_9232,N_3119);
and U10012 (N_10012,N_2114,N_9386);
nor U10013 (N_10013,N_3614,N_8010);
and U10014 (N_10014,N_8555,N_8215);
nand U10015 (N_10015,N_9140,N_7431);
nand U10016 (N_10016,N_413,N_4973);
nor U10017 (N_10017,N_3438,N_4673);
nand U10018 (N_10018,N_823,N_2778);
and U10019 (N_10019,N_6281,N_5101);
nor U10020 (N_10020,N_3168,N_1619);
nand U10021 (N_10021,N_9336,N_451);
xnor U10022 (N_10022,N_9396,N_4445);
and U10023 (N_10023,N_3350,N_1458);
and U10024 (N_10024,N_5661,N_6920);
and U10025 (N_10025,N_9297,N_7813);
nand U10026 (N_10026,N_38,N_2545);
xnor U10027 (N_10027,N_3772,N_9553);
nand U10028 (N_10028,N_3348,N_8819);
and U10029 (N_10029,N_394,N_7047);
and U10030 (N_10030,N_5137,N_6069);
or U10031 (N_10031,N_992,N_4099);
or U10032 (N_10032,N_4755,N_1292);
xnor U10033 (N_10033,N_2763,N_4965);
and U10034 (N_10034,N_9779,N_6206);
nor U10035 (N_10035,N_9905,N_3484);
nand U10036 (N_10036,N_2380,N_9495);
and U10037 (N_10037,N_9686,N_5955);
or U10038 (N_10038,N_3396,N_1244);
nor U10039 (N_10039,N_778,N_9259);
and U10040 (N_10040,N_8489,N_4902);
nand U10041 (N_10041,N_1698,N_6500);
nand U10042 (N_10042,N_3130,N_1607);
nand U10043 (N_10043,N_8086,N_6497);
nor U10044 (N_10044,N_2384,N_3283);
nand U10045 (N_10045,N_9369,N_6633);
or U10046 (N_10046,N_8309,N_1857);
nor U10047 (N_10047,N_6072,N_1325);
or U10048 (N_10048,N_5174,N_5766);
nor U10049 (N_10049,N_5803,N_2468);
or U10050 (N_10050,N_7100,N_7909);
nand U10051 (N_10051,N_4245,N_1579);
and U10052 (N_10052,N_5587,N_2890);
or U10053 (N_10053,N_5141,N_102);
or U10054 (N_10054,N_2787,N_4760);
nor U10055 (N_10055,N_3790,N_9804);
nand U10056 (N_10056,N_4050,N_5236);
nand U10057 (N_10057,N_5456,N_5140);
and U10058 (N_10058,N_3363,N_8992);
and U10059 (N_10059,N_8035,N_2668);
and U10060 (N_10060,N_6197,N_1384);
or U10061 (N_10061,N_3224,N_8713);
or U10062 (N_10062,N_2312,N_2104);
and U10063 (N_10063,N_1433,N_4096);
or U10064 (N_10064,N_4222,N_5606);
xnor U10065 (N_10065,N_7068,N_3056);
xor U10066 (N_10066,N_5392,N_5576);
nor U10067 (N_10067,N_8330,N_1648);
or U10068 (N_10068,N_7610,N_1213);
and U10069 (N_10069,N_506,N_968);
nor U10070 (N_10070,N_5054,N_8442);
nor U10071 (N_10071,N_5956,N_4644);
nor U10072 (N_10072,N_9050,N_494);
nor U10073 (N_10073,N_7103,N_6980);
or U10074 (N_10074,N_7446,N_2212);
and U10075 (N_10075,N_81,N_7623);
or U10076 (N_10076,N_5337,N_1123);
nor U10077 (N_10077,N_2571,N_7311);
nor U10078 (N_10078,N_1917,N_3125);
xnor U10079 (N_10079,N_8244,N_1738);
or U10080 (N_10080,N_9848,N_9886);
xnor U10081 (N_10081,N_8462,N_7183);
and U10082 (N_10082,N_3910,N_9935);
or U10083 (N_10083,N_4890,N_4275);
nand U10084 (N_10084,N_6225,N_3459);
or U10085 (N_10085,N_2024,N_9696);
nor U10086 (N_10086,N_1238,N_8433);
or U10087 (N_10087,N_9481,N_9127);
nand U10088 (N_10088,N_7873,N_7439);
or U10089 (N_10089,N_8515,N_7656);
nor U10090 (N_10090,N_8943,N_8570);
nand U10091 (N_10091,N_8997,N_1312);
and U10092 (N_10092,N_207,N_7915);
xnor U10093 (N_10093,N_1686,N_1470);
and U10094 (N_10094,N_7766,N_6806);
nor U10095 (N_10095,N_1744,N_9761);
nand U10096 (N_10096,N_4009,N_9643);
nor U10097 (N_10097,N_8267,N_2796);
and U10098 (N_10098,N_7033,N_3828);
and U10099 (N_10099,N_6196,N_1199);
xor U10100 (N_10100,N_8187,N_7443);
and U10101 (N_10101,N_8340,N_678);
xnor U10102 (N_10102,N_6964,N_2965);
or U10103 (N_10103,N_6342,N_9407);
xor U10104 (N_10104,N_6698,N_9918);
nor U10105 (N_10105,N_4216,N_1309);
and U10106 (N_10106,N_1429,N_4258);
nand U10107 (N_10107,N_6351,N_8873);
or U10108 (N_10108,N_8299,N_1295);
and U10109 (N_10109,N_4190,N_5465);
nand U10110 (N_10110,N_9271,N_1832);
and U10111 (N_10111,N_5557,N_3221);
nor U10112 (N_10112,N_6236,N_5133);
nand U10113 (N_10113,N_5099,N_5274);
and U10114 (N_10114,N_2444,N_4775);
and U10115 (N_10115,N_6513,N_3845);
xor U10116 (N_10116,N_8711,N_7228);
nor U10117 (N_10117,N_3602,N_2100);
or U10118 (N_10118,N_3218,N_1631);
nor U10119 (N_10119,N_565,N_6214);
and U10120 (N_10120,N_929,N_4093);
nand U10121 (N_10121,N_1937,N_21);
or U10122 (N_10122,N_1020,N_4670);
nand U10123 (N_10123,N_3665,N_9413);
nand U10124 (N_10124,N_132,N_1904);
nand U10125 (N_10125,N_1523,N_8883);
xor U10126 (N_10126,N_4750,N_1144);
nor U10127 (N_10127,N_7801,N_3676);
nand U10128 (N_10128,N_9956,N_5713);
nand U10129 (N_10129,N_8946,N_9719);
nor U10130 (N_10130,N_9667,N_9156);
nand U10131 (N_10131,N_3329,N_526);
and U10132 (N_10132,N_6784,N_3544);
nor U10133 (N_10133,N_1259,N_234);
nor U10134 (N_10134,N_3050,N_9066);
nor U10135 (N_10135,N_2915,N_9680);
nor U10136 (N_10136,N_5076,N_7442);
and U10137 (N_10137,N_5057,N_9699);
nor U10138 (N_10138,N_753,N_6685);
and U10139 (N_10139,N_9610,N_2002);
and U10140 (N_10140,N_2168,N_4911);
xor U10141 (N_10141,N_2889,N_2487);
nor U10142 (N_10142,N_3080,N_2540);
nor U10143 (N_10143,N_6171,N_947);
and U10144 (N_10144,N_1654,N_8408);
xor U10145 (N_10145,N_673,N_9593);
nand U10146 (N_10146,N_5499,N_9952);
xor U10147 (N_10147,N_9483,N_8247);
or U10148 (N_10148,N_7283,N_5083);
and U10149 (N_10149,N_511,N_9323);
nor U10150 (N_10150,N_855,N_1159);
and U10151 (N_10151,N_1438,N_8169);
and U10152 (N_10152,N_223,N_251);
or U10153 (N_10153,N_8673,N_760);
and U10154 (N_10154,N_9475,N_7851);
nand U10155 (N_10155,N_3069,N_6865);
nand U10156 (N_10156,N_9177,N_161);
nand U10157 (N_10157,N_5998,N_8767);
or U10158 (N_10158,N_8798,N_6158);
and U10159 (N_10159,N_670,N_2190);
nand U10160 (N_10160,N_1139,N_3390);
xnor U10161 (N_10161,N_6712,N_3464);
nand U10162 (N_10162,N_4709,N_7119);
or U10163 (N_10163,N_18,N_6084);
nand U10164 (N_10164,N_2880,N_2617);
nand U10165 (N_10165,N_3193,N_7671);
or U10166 (N_10166,N_6913,N_1568);
and U10167 (N_10167,N_7265,N_2441);
and U10168 (N_10168,N_937,N_9972);
and U10169 (N_10169,N_779,N_4176);
and U10170 (N_10170,N_2434,N_9153);
and U10171 (N_10171,N_5321,N_3081);
nor U10172 (N_10172,N_6210,N_1906);
or U10173 (N_10173,N_534,N_317);
or U10174 (N_10174,N_3905,N_9912);
nand U10175 (N_10175,N_4262,N_3148);
nor U10176 (N_10176,N_2073,N_3660);
and U10177 (N_10177,N_9801,N_7073);
nand U10178 (N_10178,N_2246,N_2461);
nand U10179 (N_10179,N_7036,N_3781);
nand U10180 (N_10180,N_2450,N_6890);
or U10181 (N_10181,N_585,N_9301);
or U10182 (N_10182,N_564,N_5435);
nor U10183 (N_10183,N_2777,N_8722);
or U10184 (N_10184,N_1844,N_3755);
xor U10185 (N_10185,N_73,N_2029);
and U10186 (N_10186,N_4936,N_4719);
nor U10187 (N_10187,N_492,N_5025);
or U10188 (N_10188,N_8354,N_9178);
and U10189 (N_10189,N_6755,N_3075);
nor U10190 (N_10190,N_9046,N_5015);
and U10191 (N_10191,N_1501,N_8690);
nor U10192 (N_10192,N_3220,N_5287);
or U10193 (N_10193,N_4298,N_5039);
and U10194 (N_10194,N_2062,N_96);
and U10195 (N_10195,N_8223,N_2377);
nor U10196 (N_10196,N_133,N_1495);
and U10197 (N_10197,N_6400,N_849);
or U10198 (N_10198,N_6051,N_3733);
nand U10199 (N_10199,N_3216,N_5769);
and U10200 (N_10200,N_1282,N_6777);
xnor U10201 (N_10201,N_8119,N_7079);
and U10202 (N_10202,N_3278,N_9586);
nand U10203 (N_10203,N_1118,N_4501);
xor U10204 (N_10204,N_6602,N_2070);
or U10205 (N_10205,N_4457,N_2926);
nor U10206 (N_10206,N_894,N_3444);
and U10207 (N_10207,N_370,N_5029);
or U10208 (N_10208,N_6559,N_6771);
or U10209 (N_10209,N_7760,N_5534);
nor U10210 (N_10210,N_8033,N_3248);
nand U10211 (N_10211,N_226,N_785);
or U10212 (N_10212,N_822,N_2848);
or U10213 (N_10213,N_6732,N_6808);
nor U10214 (N_10214,N_9161,N_4167);
or U10215 (N_10215,N_13,N_3939);
and U10216 (N_10216,N_5297,N_5421);
nor U10217 (N_10217,N_8554,N_3914);
and U10218 (N_10218,N_8252,N_6015);
or U10219 (N_10219,N_7296,N_1383);
xor U10220 (N_10220,N_2589,N_5152);
nand U10221 (N_10221,N_6624,N_7763);
nand U10222 (N_10222,N_9520,N_2021);
nor U10223 (N_10223,N_3921,N_2966);
nor U10224 (N_10224,N_9174,N_1925);
nor U10225 (N_10225,N_4492,N_8763);
nand U10226 (N_10226,N_9748,N_5648);
and U10227 (N_10227,N_8709,N_1432);
nand U10228 (N_10228,N_2895,N_2249);
nand U10229 (N_10229,N_4932,N_428);
xor U10230 (N_10230,N_4074,N_5750);
and U10231 (N_10231,N_5282,N_5361);
and U10232 (N_10232,N_7665,N_9242);
and U10233 (N_10233,N_208,N_9826);
nand U10234 (N_10234,N_5393,N_5643);
and U10235 (N_10235,N_1022,N_7488);
or U10236 (N_10236,N_5284,N_7558);
or U10237 (N_10237,N_4615,N_4789);
xnor U10238 (N_10238,N_3238,N_1414);
nand U10239 (N_10239,N_6793,N_6437);
or U10240 (N_10240,N_9879,N_5857);
nor U10241 (N_10241,N_6915,N_7020);
nand U10242 (N_10242,N_5812,N_5169);
or U10243 (N_10243,N_3540,N_8027);
nor U10244 (N_10244,N_5102,N_332);
nand U10245 (N_10245,N_5860,N_3301);
and U10246 (N_10246,N_653,N_6975);
xor U10247 (N_10247,N_6818,N_1833);
or U10248 (N_10248,N_2033,N_2695);
or U10249 (N_10249,N_5125,N_6141);
or U10250 (N_10250,N_1190,N_6162);
xor U10251 (N_10251,N_5084,N_8893);
or U10252 (N_10252,N_2967,N_3748);
and U10253 (N_10253,N_3341,N_6613);
or U10254 (N_10254,N_8937,N_1721);
xnor U10255 (N_10255,N_6838,N_3129);
or U10256 (N_10256,N_9109,N_2681);
or U10257 (N_10257,N_3333,N_1952);
or U10258 (N_10258,N_3436,N_6037);
or U10259 (N_10259,N_4523,N_4388);
nand U10260 (N_10260,N_2875,N_1538);
nor U10261 (N_10261,N_953,N_1423);
nand U10262 (N_10262,N_6232,N_8944);
or U10263 (N_10263,N_4738,N_4564);
xor U10264 (N_10264,N_9221,N_3381);
nor U10265 (N_10265,N_8840,N_9438);
or U10266 (N_10266,N_2888,N_5199);
or U10267 (N_10267,N_3187,N_1046);
and U10268 (N_10268,N_4256,N_9981);
xnor U10269 (N_10269,N_5175,N_5437);
nor U10270 (N_10270,N_2288,N_4696);
nand U10271 (N_10271,N_600,N_5675);
or U10272 (N_10272,N_3761,N_5241);
or U10273 (N_10273,N_7683,N_9290);
nor U10274 (N_10274,N_7098,N_911);
or U10275 (N_10275,N_5927,N_5309);
nor U10276 (N_10276,N_7568,N_4408);
and U10277 (N_10277,N_4896,N_7510);
or U10278 (N_10278,N_384,N_3880);
xnor U10279 (N_10279,N_2413,N_9865);
or U10280 (N_10280,N_2546,N_3491);
nand U10281 (N_10281,N_3503,N_7792);
and U10282 (N_10282,N_6877,N_3683);
nor U10283 (N_10283,N_276,N_7950);
or U10284 (N_10284,N_6134,N_7942);
nor U10285 (N_10285,N_7908,N_3513);
and U10286 (N_10286,N_2274,N_9035);
or U10287 (N_10287,N_9285,N_3280);
nor U10288 (N_10288,N_9113,N_7895);
nand U10289 (N_10289,N_4379,N_4352);
nor U10290 (N_10290,N_4422,N_4373);
xnor U10291 (N_10291,N_9778,N_3999);
xnor U10292 (N_10292,N_2866,N_4165);
or U10293 (N_10293,N_3034,N_1935);
and U10294 (N_10294,N_6024,N_1499);
or U10295 (N_10295,N_7465,N_1437);
or U10296 (N_10296,N_210,N_9305);
xor U10297 (N_10297,N_3490,N_7133);
xnor U10298 (N_10298,N_3255,N_5249);
nand U10299 (N_10299,N_9404,N_4117);
nand U10300 (N_10300,N_1285,N_931);
nor U10301 (N_10301,N_1214,N_7974);
or U10302 (N_10302,N_7635,N_1574);
nand U10303 (N_10303,N_415,N_4534);
and U10304 (N_10304,N_3850,N_8001);
xor U10305 (N_10305,N_3521,N_6324);
and U10306 (N_10306,N_4987,N_7479);
and U10307 (N_10307,N_5707,N_7019);
nor U10308 (N_10308,N_4213,N_5798);
or U10309 (N_10309,N_2362,N_2193);
nor U10310 (N_10310,N_2140,N_4585);
or U10311 (N_10311,N_1203,N_5184);
and U10312 (N_10312,N_9185,N_168);
nor U10313 (N_10313,N_7236,N_7454);
or U10314 (N_10314,N_8162,N_2330);
nor U10315 (N_10315,N_48,N_9873);
nand U10316 (N_10316,N_4199,N_357);
or U10317 (N_10317,N_8525,N_6349);
nand U10318 (N_10318,N_5991,N_5397);
and U10319 (N_10319,N_6703,N_1072);
and U10320 (N_10320,N_8216,N_8350);
nand U10321 (N_10321,N_2323,N_2971);
or U10322 (N_10322,N_7747,N_1459);
or U10323 (N_10323,N_1821,N_7444);
nor U10324 (N_10324,N_5744,N_7532);
xnor U10325 (N_10325,N_4486,N_7627);
and U10326 (N_10326,N_6606,N_8300);
nor U10327 (N_10327,N_9751,N_28);
nor U10328 (N_10328,N_1504,N_867);
nor U10329 (N_10329,N_443,N_3178);
and U10330 (N_10330,N_4819,N_1419);
or U10331 (N_10331,N_3394,N_7260);
nand U10332 (N_10332,N_7231,N_6622);
nand U10333 (N_10333,N_3720,N_7484);
xor U10334 (N_10334,N_5858,N_3180);
nand U10335 (N_10335,N_2198,N_3487);
or U10336 (N_10336,N_5718,N_4101);
and U10337 (N_10337,N_824,N_6817);
nor U10338 (N_10338,N_6549,N_8407);
xor U10339 (N_10339,N_4810,N_1612);
nand U10340 (N_10340,N_369,N_3144);
or U10341 (N_10341,N_536,N_4857);
or U10342 (N_10342,N_4240,N_551);
or U10343 (N_10343,N_7298,N_8772);
or U10344 (N_10344,N_2354,N_8156);
or U10345 (N_10345,N_5034,N_1492);
nand U10346 (N_10346,N_8082,N_6426);
nor U10347 (N_10347,N_7469,N_8677);
or U10348 (N_10348,N_4925,N_9227);
nor U10349 (N_10349,N_9402,N_2069);
nand U10350 (N_10350,N_1026,N_1831);
nor U10351 (N_10351,N_7057,N_6748);
or U10352 (N_10352,N_3684,N_6246);
nand U10353 (N_10353,N_3167,N_746);
nand U10354 (N_10354,N_1092,N_2508);
nor U10355 (N_10355,N_1630,N_1897);
or U10356 (N_10356,N_5878,N_505);
nor U10357 (N_10357,N_3582,N_6753);
and U10358 (N_10358,N_2042,N_3844);
xnor U10359 (N_10359,N_5281,N_5629);
or U10360 (N_10360,N_3294,N_951);
and U10361 (N_10361,N_2884,N_5124);
nand U10362 (N_10362,N_5402,N_5271);
nor U10363 (N_10363,N_2418,N_3312);
nor U10364 (N_10364,N_8057,N_1289);
and U10365 (N_10365,N_3648,N_5463);
and U10366 (N_10366,N_283,N_1647);
nor U10367 (N_10367,N_8945,N_9637);
nand U10368 (N_10368,N_2108,N_4020);
nor U10369 (N_10369,N_1345,N_7842);
or U10370 (N_10370,N_6229,N_2802);
and U10371 (N_10371,N_8159,N_7693);
nor U10372 (N_10372,N_9432,N_4667);
nor U10373 (N_10373,N_7356,N_3332);
nand U10374 (N_10374,N_1816,N_3858);
or U10375 (N_10375,N_853,N_4358);
nand U10376 (N_10376,N_2519,N_2736);
and U10377 (N_10377,N_7989,N_8672);
nand U10378 (N_10378,N_9057,N_8541);
or U10379 (N_10379,N_8910,N_4128);
and U10380 (N_10380,N_9660,N_763);
or U10381 (N_10381,N_197,N_5637);
nor U10382 (N_10382,N_7229,N_2701);
or U10383 (N_10383,N_8984,N_142);
and U10384 (N_10384,N_9039,N_4960);
nand U10385 (N_10385,N_6003,N_1341);
and U10386 (N_10386,N_5443,N_6931);
nor U10387 (N_10387,N_697,N_1699);
nor U10388 (N_10388,N_336,N_1024);
or U10389 (N_10389,N_9280,N_5736);
and U10390 (N_10390,N_3589,N_1954);
nor U10391 (N_10391,N_6223,N_1003);
xnor U10392 (N_10392,N_2076,N_3682);
nor U10393 (N_10393,N_2946,N_3603);
and U10394 (N_10394,N_7704,N_8995);
nor U10395 (N_10395,N_7961,N_424);
xnor U10396 (N_10396,N_2740,N_8734);
nand U10397 (N_10397,N_9550,N_8304);
and U10398 (N_10398,N_1035,N_6133);
nand U10399 (N_10399,N_2120,N_1839);
nand U10400 (N_10400,N_991,N_5936);
or U10401 (N_10401,N_2244,N_3578);
or U10402 (N_10402,N_5996,N_1996);
and U10403 (N_10403,N_1921,N_8361);
or U10404 (N_10404,N_2311,N_9741);
and U10405 (N_10405,N_7549,N_4205);
xnor U10406 (N_10406,N_2432,N_2959);
nor U10407 (N_10407,N_3716,N_2426);
nor U10408 (N_10408,N_9282,N_1427);
or U10409 (N_10409,N_7826,N_8316);
and U10410 (N_10410,N_1006,N_275);
nor U10411 (N_10411,N_9331,N_6684);
nand U10412 (N_10412,N_805,N_8085);
nand U10413 (N_10413,N_4160,N_9451);
and U10414 (N_10414,N_9462,N_4414);
nor U10415 (N_10415,N_117,N_3820);
nand U10416 (N_10416,N_3202,N_8916);
nand U10417 (N_10417,N_3778,N_758);
nor U10418 (N_10418,N_157,N_574);
xor U10419 (N_10419,N_5493,N_7725);
nor U10420 (N_10420,N_1318,N_9502);
nor U10421 (N_10421,N_4758,N_7680);
or U10422 (N_10422,N_2010,N_4140);
and U10423 (N_10423,N_1263,N_3530);
xnor U10424 (N_10424,N_9670,N_1516);
or U10425 (N_10425,N_3300,N_4484);
or U10426 (N_10426,N_5919,N_99);
or U10427 (N_10427,N_6142,N_4456);
or U10428 (N_10428,N_4271,N_2313);
xor U10429 (N_10429,N_315,N_2226);
or U10430 (N_10430,N_1924,N_3630);
nor U10431 (N_10431,N_3445,N_4595);
xnor U10432 (N_10432,N_8575,N_8865);
nand U10433 (N_10433,N_6619,N_7354);
or U10434 (N_10434,N_2241,N_5968);
nor U10435 (N_10435,N_5489,N_5959);
nand U10436 (N_10436,N_8197,N_2083);
nor U10437 (N_10437,N_6848,N_8707);
nand U10438 (N_10438,N_6031,N_9914);
nor U10439 (N_10439,N_8439,N_5316);
nor U10440 (N_10440,N_5627,N_2383);
xnor U10441 (N_10441,N_7242,N_7844);
or U10442 (N_10442,N_7886,N_3404);
or U10443 (N_10443,N_3302,N_6720);
nand U10444 (N_10444,N_8807,N_979);
or U10445 (N_10445,N_4773,N_9154);
xnor U10446 (N_10446,N_4088,N_6832);
nand U10447 (N_10447,N_4179,N_1271);
nor U10448 (N_10448,N_4617,N_5980);
nand U10449 (N_10449,N_7339,N_9773);
and U10450 (N_10450,N_7687,N_9692);
nor U10451 (N_10451,N_8470,N_6679);
nor U10452 (N_10452,N_8096,N_3065);
nand U10453 (N_10453,N_6979,N_2670);
xor U10454 (N_10454,N_7486,N_2186);
nor U10455 (N_10455,N_8282,N_3678);
nand U10456 (N_10456,N_477,N_4212);
nand U10457 (N_10457,N_8728,N_9509);
or U10458 (N_10458,N_6233,N_8114);
nor U10459 (N_10459,N_713,N_2113);
xor U10460 (N_10460,N_741,N_6452);
and U10461 (N_10461,N_6539,N_3819);
nand U10462 (N_10462,N_3974,N_7823);
nor U10463 (N_10463,N_1727,N_4479);
or U10464 (N_10464,N_9160,N_7464);
nor U10465 (N_10465,N_1435,N_9745);
or U10466 (N_10466,N_3272,N_9711);
and U10467 (N_10467,N_3864,N_4531);
or U10468 (N_10468,N_6346,N_1062);
or U10469 (N_10469,N_6023,N_4046);
or U10470 (N_10470,N_5699,N_9962);
nor U10471 (N_10471,N_6179,N_5723);
nand U10472 (N_10472,N_2103,N_6541);
xor U10473 (N_10473,N_93,N_2598);
nor U10474 (N_10474,N_671,N_7528);
or U10475 (N_10475,N_1894,N_8089);
or U10476 (N_10476,N_4030,N_5677);
nor U10477 (N_10477,N_4412,N_6797);
nand U10478 (N_10478,N_2294,N_1418);
nor U10479 (N_10479,N_5378,N_4468);
nor U10480 (N_10480,N_5280,N_1790);
and U10481 (N_10481,N_6159,N_4683);
nand U10482 (N_10482,N_4286,N_8356);
and U10483 (N_10483,N_647,N_9423);
nand U10484 (N_10484,N_2337,N_1567);
or U10485 (N_10485,N_6837,N_6062);
xnor U10486 (N_10486,N_1565,N_7388);
and U10487 (N_10487,N_200,N_4183);
and U10488 (N_10488,N_1765,N_5743);
nand U10489 (N_10489,N_3696,N_8297);
nand U10490 (N_10490,N_4380,N_6563);
nor U10491 (N_10491,N_7567,N_4999);
nand U10492 (N_10492,N_4084,N_2375);
and U10493 (N_10493,N_1736,N_8671);
nand U10494 (N_10494,N_7306,N_7734);
nor U10495 (N_10495,N_87,N_3585);
nand U10496 (N_10496,N_6667,N_2822);
or U10497 (N_10497,N_5445,N_3236);
nor U10498 (N_10498,N_3738,N_7258);
or U10499 (N_10499,N_7130,N_6202);
and U10500 (N_10500,N_8724,N_2551);
and U10501 (N_10501,N_5159,N_3944);
and U10502 (N_10502,N_6180,N_1893);
nand U10503 (N_10503,N_8974,N_6375);
nor U10504 (N_10504,N_5171,N_3289);
nor U10505 (N_10505,N_7290,N_6993);
xnor U10506 (N_10506,N_8646,N_9846);
nor U10507 (N_10507,N_9187,N_293);
nand U10508 (N_10508,N_4487,N_2652);
xnor U10509 (N_10509,N_9497,N_8640);
and U10510 (N_10510,N_8168,N_5452);
xor U10511 (N_10511,N_1475,N_421);
nand U10512 (N_10512,N_5665,N_1207);
nor U10513 (N_10513,N_2352,N_6235);
nand U10514 (N_10514,N_5376,N_1351);
or U10515 (N_10515,N_9591,N_7561);
or U10516 (N_10516,N_6198,N_3298);
and U10517 (N_10517,N_7404,N_5690);
or U10518 (N_10518,N_3033,N_7770);
or U10519 (N_10519,N_3580,N_8444);
nor U10520 (N_10520,N_2960,N_1483);
nor U10521 (N_10521,N_5514,N_1267);
nand U10522 (N_10522,N_2938,N_938);
nand U10523 (N_10523,N_1836,N_6301);
nor U10524 (N_10524,N_6895,N_9312);
nor U10525 (N_10525,N_8776,N_2628);
nand U10526 (N_10526,N_2748,N_662);
nor U10527 (N_10527,N_7414,N_8314);
xor U10528 (N_10528,N_2339,N_5791);
nor U10529 (N_10529,N_7393,N_4163);
or U10530 (N_10530,N_8287,N_2094);
xnor U10531 (N_10531,N_5188,N_1624);
nor U10532 (N_10532,N_817,N_5170);
or U10533 (N_10533,N_598,N_7470);
nand U10534 (N_10534,N_5817,N_8368);
and U10535 (N_10535,N_5467,N_9490);
and U10536 (N_10536,N_1825,N_2698);
nand U10537 (N_10537,N_734,N_3826);
xor U10538 (N_10538,N_4892,N_2370);
or U10539 (N_10539,N_8383,N_8935);
and U10540 (N_10540,N_8549,N_6418);
or U10541 (N_10541,N_1059,N_9946);
xor U10542 (N_10542,N_2485,N_6227);
nor U10543 (N_10543,N_3383,N_3309);
or U10544 (N_10544,N_9925,N_4253);
or U10545 (N_10545,N_9951,N_5997);
nor U10546 (N_10546,N_8812,N_7728);
and U10547 (N_10547,N_6977,N_462);
or U10548 (N_10548,N_2779,N_6020);
or U10549 (N_10549,N_1496,N_7081);
or U10550 (N_10550,N_1422,N_8643);
and U10551 (N_10551,N_1769,N_6701);
nand U10552 (N_10552,N_3710,N_4431);
or U10553 (N_10553,N_2912,N_5420);
or U10554 (N_10554,N_2124,N_6428);
and U10555 (N_10555,N_726,N_2803);
nand U10556 (N_10556,N_4589,N_4325);
nand U10557 (N_10557,N_4904,N_801);
or U10558 (N_10558,N_9343,N_7008);
nor U10559 (N_10559,N_6804,N_8917);
and U10560 (N_10560,N_2181,N_9669);
or U10561 (N_10561,N_6243,N_148);
and U10562 (N_10562,N_9754,N_6358);
and U10563 (N_10563,N_3770,N_5447);
nor U10564 (N_10564,N_6068,N_356);
or U10565 (N_10565,N_3429,N_4504);
nor U10566 (N_10566,N_4441,N_2117);
and U10567 (N_10567,N_959,N_2836);
and U10568 (N_10568,N_1692,N_449);
nor U10569 (N_10569,N_5218,N_8817);
nor U10570 (N_10570,N_1643,N_9131);
xnor U10571 (N_10571,N_2146,N_2764);
nand U10572 (N_10572,N_4661,N_5217);
nor U10573 (N_10573,N_2009,N_4844);
or U10574 (N_10574,N_5277,N_3946);
nand U10575 (N_10575,N_6850,N_5712);
nand U10576 (N_10576,N_7887,N_6847);
or U10577 (N_10577,N_8478,N_4200);
or U10578 (N_10578,N_115,N_5873);
or U10579 (N_10579,N_8406,N_3987);
and U10580 (N_10580,N_8275,N_8546);
and U10581 (N_10581,N_3549,N_7097);
or U10582 (N_10582,N_5454,N_8034);
and U10583 (N_10583,N_8687,N_9630);
nand U10584 (N_10584,N_9965,N_2827);
xnor U10585 (N_10585,N_9102,N_3271);
nor U10586 (N_10586,N_9148,N_1007);
nand U10587 (N_10587,N_7223,N_6436);
and U10588 (N_10588,N_8502,N_3531);
or U10589 (N_10589,N_2415,N_9840);
nor U10590 (N_10590,N_2099,N_141);
or U10591 (N_10591,N_8324,N_6356);
nor U10592 (N_10592,N_5735,N_2044);
and U10593 (N_10593,N_5388,N_298);
xnor U10594 (N_10594,N_6885,N_9078);
or U10595 (N_10595,N_1378,N_8532);
nand U10596 (N_10596,N_7440,N_5702);
and U10597 (N_10597,N_8564,N_8080);
nand U10598 (N_10598,N_6207,N_9231);
or U10599 (N_10599,N_3932,N_2224);
xnor U10600 (N_10600,N_9706,N_1170);
xnor U10601 (N_10601,N_5592,N_8373);
nand U10602 (N_10602,N_3897,N_4290);
nand U10603 (N_10603,N_2091,N_1875);
nand U10604 (N_10604,N_3824,N_199);
and U10605 (N_10605,N_6846,N_1028);
xor U10606 (N_10606,N_4203,N_7550);
or U10607 (N_10607,N_4915,N_8832);
nor U10608 (N_10608,N_5145,N_2066);
or U10609 (N_10609,N_837,N_5185);
nor U10610 (N_10610,N_5505,N_3343);
and U10611 (N_10611,N_2000,N_8017);
and U10612 (N_10612,N_4138,N_2065);
or U10613 (N_10613,N_2030,N_8499);
or U10614 (N_10614,N_5588,N_6822);
or U10615 (N_10615,N_8885,N_9136);
and U10616 (N_10616,N_2972,N_8186);
nand U10617 (N_10617,N_9002,N_7261);
nand U10618 (N_10618,N_4292,N_5526);
or U10619 (N_10619,N_3904,N_7914);
nand U10620 (N_10620,N_9771,N_9656);
nor U10621 (N_10621,N_490,N_765);
and U10622 (N_10622,N_9635,N_525);
nand U10623 (N_10623,N_1918,N_5033);
xor U10624 (N_10624,N_2861,N_7938);
nand U10625 (N_10625,N_1146,N_4033);
and U10626 (N_10626,N_3622,N_5710);
and U10627 (N_10627,N_577,N_1107);
and U10628 (N_10628,N_1204,N_3299);
or U10629 (N_10629,N_4681,N_4461);
or U10630 (N_10630,N_2043,N_7672);
nor U10631 (N_10631,N_641,N_1337);
nand U10632 (N_10632,N_74,N_6723);
nand U10633 (N_10633,N_4626,N_2986);
or U10634 (N_10634,N_2162,N_3074);
and U10635 (N_10635,N_3400,N_6248);
and U10636 (N_10636,N_1817,N_5444);
and U10637 (N_10637,N_9422,N_9955);
and U10638 (N_10638,N_8569,N_130);
nand U10639 (N_10639,N_6738,N_1201);
nor U10640 (N_10640,N_194,N_4018);
or U10641 (N_10641,N_3588,N_7471);
nand U10642 (N_10642,N_6132,N_2172);
nand U10643 (N_10643,N_5839,N_3387);
nor U10644 (N_10644,N_2205,N_7104);
or U10645 (N_10645,N_7483,N_8524);
or U10646 (N_10646,N_5647,N_2481);
nor U10647 (N_10647,N_7780,N_6757);
nor U10648 (N_10648,N_9347,N_691);
or U10649 (N_10649,N_7196,N_8194);
and U10650 (N_10650,N_5313,N_6864);
and U10651 (N_10651,N_7736,N_3654);
nand U10652 (N_10652,N_3365,N_7843);
xor U10653 (N_10653,N_6728,N_9496);
or U10654 (N_10654,N_4891,N_2458);
or U10655 (N_10655,N_5985,N_2576);
nand U10656 (N_10656,N_5950,N_3038);
and U10657 (N_10657,N_5108,N_6552);
and U10658 (N_10658,N_3849,N_4736);
or U10659 (N_10659,N_6534,N_4123);
nor U10660 (N_10660,N_9749,N_3093);
or U10661 (N_10661,N_5343,N_9294);
or U10662 (N_10662,N_3500,N_5783);
or U10663 (N_10663,N_6241,N_1392);
nand U10664 (N_10664,N_295,N_4436);
xor U10665 (N_10665,N_7804,N_548);
nand U10666 (N_10666,N_4499,N_733);
nand U10667 (N_10667,N_862,N_9466);
nor U10668 (N_10668,N_1031,N_4533);
or U10669 (N_10669,N_5223,N_5085);
and U10670 (N_10670,N_2548,N_6455);
nor U10671 (N_10671,N_9619,N_8585);
nor U10672 (N_10672,N_7011,N_224);
nand U10673 (N_10673,N_4097,N_8849);
nor U10674 (N_10674,N_9213,N_9142);
nand U10675 (N_10675,N_2098,N_2879);
or U10676 (N_10676,N_8881,N_8695);
xnor U10677 (N_10677,N_2179,N_4323);
and U10678 (N_10678,N_9470,N_5845);
or U10679 (N_10679,N_4552,N_5259);
or U10680 (N_10680,N_1012,N_2215);
or U10681 (N_10681,N_4856,N_3201);
or U10682 (N_10682,N_9360,N_2250);
nand U10683 (N_10683,N_6855,N_8976);
or U10684 (N_10684,N_7058,N_2406);
or U10685 (N_10685,N_9789,N_6588);
nor U10686 (N_10686,N_6746,N_3866);
nor U10687 (N_10687,N_9084,N_3164);
or U10688 (N_10688,N_5005,N_6064);
or U10689 (N_10689,N_3360,N_7628);
nor U10690 (N_10690,N_7217,N_6640);
xnor U10691 (N_10691,N_9720,N_4503);
and U10692 (N_10692,N_4893,N_9245);
or U10693 (N_10693,N_3025,N_4080);
nand U10694 (N_10694,N_701,N_8014);
and U10695 (N_10695,N_6851,N_3273);
and U10696 (N_10696,N_4870,N_8313);
and U10697 (N_10697,N_1912,N_7048);
and U10698 (N_10698,N_6820,N_9676);
nand U10699 (N_10699,N_9612,N_3834);
nor U10700 (N_10700,N_4178,N_5181);
and U10701 (N_10701,N_7381,N_7424);
xnor U10702 (N_10702,N_680,N_4174);
nor U10703 (N_10703,N_946,N_2171);
and U10704 (N_10704,N_3803,N_901);
nor U10705 (N_10705,N_1396,N_8116);
nor U10706 (N_10706,N_113,N_299);
nor U10707 (N_10707,N_9182,N_9269);
nor U10708 (N_10708,N_2553,N_7074);
or U10709 (N_10709,N_6311,N_193);
nor U10710 (N_10710,N_5384,N_5886);
and U10711 (N_10711,N_1592,N_629);
and U10712 (N_10712,N_7504,N_3336);
nand U10713 (N_10713,N_7786,N_397);
nand U10714 (N_10714,N_5540,N_3410);
and U10715 (N_10715,N_2470,N_4356);
nor U10716 (N_10716,N_4685,N_8592);
or U10717 (N_10717,N_5494,N_403);
nor U10718 (N_10718,N_1430,N_7772);
and U10719 (N_10719,N_6186,N_9717);
or U10720 (N_10720,N_8847,N_8900);
nor U10721 (N_10721,N_2015,N_1992);
and U10722 (N_10722,N_7025,N_710);
nand U10723 (N_10723,N_3786,N_1416);
nand U10724 (N_10724,N_3257,N_7764);
nand U10725 (N_10725,N_4026,N_7936);
nand U10726 (N_10726,N_3543,N_4348);
or U10727 (N_10727,N_9150,N_4677);
or U10728 (N_10728,N_8289,N_4783);
and U10729 (N_10729,N_1645,N_6689);
or U10730 (N_10730,N_1581,N_4757);
or U10731 (N_10731,N_1970,N_8797);
or U10732 (N_10732,N_1822,N_784);
or U10733 (N_10733,N_339,N_9080);
and U10734 (N_10734,N_6770,N_9727);
nor U10735 (N_10735,N_4334,N_5365);
nor U10736 (N_10736,N_7878,N_4647);
or U10737 (N_10737,N_5450,N_7280);
xnor U10738 (N_10738,N_8820,N_3447);
nor U10739 (N_10739,N_3599,N_9537);
nor U10740 (N_10740,N_6044,N_7351);
nor U10741 (N_10741,N_8107,N_2925);
or U10742 (N_10742,N_8921,N_936);
nand U10743 (N_10743,N_3713,N_4634);
xnor U10744 (N_10744,N_8212,N_5387);
nor U10745 (N_10745,N_1962,N_8193);
xnor U10746 (N_10746,N_5572,N_1079);
nand U10747 (N_10747,N_138,N_9938);
or U10748 (N_10748,N_1999,N_2616);
and U10749 (N_10749,N_6022,N_6638);
or U10750 (N_10750,N_9644,N_6543);
or U10751 (N_10751,N_8178,N_2620);
and U10752 (N_10752,N_1168,N_8430);
nor U10753 (N_10753,N_2367,N_2017);
xor U10754 (N_10754,N_9767,N_6484);
nand U10755 (N_10755,N_8894,N_1165);
and U10756 (N_10756,N_5797,N_5273);
nor U10757 (N_10757,N_6932,N_7053);
and U10758 (N_10758,N_2556,N_9551);
or U10759 (N_10759,N_5714,N_3213);
nor U10760 (N_10760,N_3619,N_8228);
nor U10761 (N_10761,N_3210,N_7758);
nand U10762 (N_10762,N_6634,N_8500);
or U10763 (N_10763,N_1880,N_9577);
nor U10764 (N_10764,N_880,N_4888);
xnor U10765 (N_10765,N_5500,N_152);
or U10766 (N_10766,N_4027,N_2410);
and U10767 (N_10767,N_309,N_7857);
nand U10768 (N_10768,N_1615,N_7591);
and U10769 (N_10769,N_4933,N_5584);
and U10770 (N_10770,N_50,N_8731);
nand U10771 (N_10771,N_1355,N_2419);
nor U10772 (N_10772,N_3008,N_7310);
nand U10773 (N_10773,N_2258,N_1172);
nand U10774 (N_10774,N_892,N_3659);
xnor U10775 (N_10775,N_4785,N_3808);
nand U10776 (N_10776,N_504,N_7482);
or U10777 (N_10777,N_8227,N_736);
or U10778 (N_10778,N_2798,N_527);
nand U10779 (N_10779,N_8049,N_104);
and U10780 (N_10780,N_3402,N_7273);
nand U10781 (N_10781,N_1515,N_6380);
or U10782 (N_10782,N_3523,N_1584);
or U10783 (N_10783,N_8708,N_4948);
nor U10784 (N_10784,N_4975,N_6786);
nand U10785 (N_10785,N_5367,N_1734);
nand U10786 (N_10786,N_5087,N_3926);
and U10787 (N_10787,N_4588,N_8539);
or U10788 (N_10788,N_2227,N_6708);
nor U10789 (N_10789,N_6071,N_7032);
and U10790 (N_10790,N_1746,N_122);
nor U10791 (N_10791,N_2829,N_4741);
nor U10792 (N_10792,N_8618,N_2035);
nand U10793 (N_10793,N_8639,N_8198);
nor U10794 (N_10794,N_8704,N_3244);
and U10795 (N_10795,N_8522,N_869);
nand U10796 (N_10796,N_9782,N_7101);
xor U10797 (N_10797,N_4395,N_4847);
or U10798 (N_10798,N_6644,N_9292);
nand U10799 (N_10799,N_1444,N_6765);
nor U10800 (N_10800,N_6899,N_3412);
or U10801 (N_10801,N_1681,N_789);
xnor U10802 (N_10802,N_5094,N_9507);
and U10803 (N_10803,N_3789,N_7320);
nor U10804 (N_10804,N_9758,N_6992);
xor U10805 (N_10805,N_8397,N_3085);
nor U10806 (N_10806,N_8366,N_8298);
nor U10807 (N_10807,N_4404,N_3114);
and U10808 (N_10808,N_6085,N_2864);
nor U10809 (N_10809,N_9780,N_458);
or U10810 (N_10810,N_995,N_249);
nor U10811 (N_10811,N_1915,N_487);
nand U10812 (N_10812,N_8530,N_9649);
and U10813 (N_10813,N_2651,N_1130);
and U10814 (N_10814,N_6220,N_7784);
nand U10815 (N_10815,N_1556,N_177);
or U10816 (N_10816,N_8185,N_5719);
or U10817 (N_10817,N_9793,N_2304);
or U10818 (N_10818,N_3243,N_8669);
xor U10819 (N_10819,N_4707,N_9257);
and U10820 (N_10820,N_6407,N_4934);
and U10821 (N_10821,N_6309,N_3391);
or U10822 (N_10822,N_8769,N_4611);
or U10823 (N_10823,N_3749,N_6321);
and U10824 (N_10824,N_3532,N_9001);
nor U10825 (N_10825,N_1236,N_2316);
and U10826 (N_10826,N_5826,N_5424);
nand U10827 (N_10827,N_6956,N_6514);
or U10828 (N_10828,N_8956,N_3086);
and U10829 (N_10829,N_2907,N_4350);
and U10830 (N_10830,N_7411,N_2745);
or U10831 (N_10831,N_8388,N_222);
xnor U10832 (N_10832,N_3744,N_2530);
or U10833 (N_10833,N_1689,N_928);
or U10834 (N_10834,N_3823,N_88);
xnor U10835 (N_10835,N_6333,N_5767);
or U10836 (N_10836,N_9531,N_5119);
nand U10837 (N_10837,N_7340,N_1702);
nand U10838 (N_10838,N_5417,N_3908);
and U10839 (N_10839,N_3935,N_5618);
nand U10840 (N_10840,N_6562,N_1633);
nor U10841 (N_10841,N_9731,N_8496);
nor U10842 (N_10842,N_9683,N_594);
nand U10843 (N_10843,N_4947,N_2428);
nand U10844 (N_10844,N_7658,N_9264);
nand U10845 (N_10845,N_5329,N_9014);
xnor U10846 (N_10846,N_7322,N_7018);
and U10847 (N_10847,N_9940,N_9115);
nand U10848 (N_10848,N_1447,N_5131);
nor U10849 (N_10849,N_353,N_7177);
or U10850 (N_10850,N_8882,N_9121);
nand U10851 (N_10851,N_9226,N_2547);
xnor U10852 (N_10852,N_3782,N_1611);
nand U10853 (N_10853,N_9068,N_287);
nand U10854 (N_10854,N_6949,N_1766);
or U10855 (N_10855,N_9274,N_8854);
or U10856 (N_10856,N_2204,N_9358);
or U10857 (N_10857,N_2758,N_9076);
or U10858 (N_10858,N_8577,N_958);
nand U10859 (N_10859,N_820,N_2401);
nand U10860 (N_10860,N_7699,N_1533);
xnor U10861 (N_10861,N_2116,N_2040);
or U10862 (N_10862,N_3515,N_8273);
xor U10863 (N_10863,N_4914,N_6652);
nand U10864 (N_10864,N_355,N_4415);
nor U10865 (N_10865,N_1424,N_2891);
or U10866 (N_10866,N_1572,N_2795);
nand U10867 (N_10867,N_7426,N_5130);
and U10868 (N_10868,N_5717,N_6256);
or U10869 (N_10869,N_8988,N_6118);
nand U10870 (N_10870,N_7932,N_2928);
or U10871 (N_10871,N_9818,N_2189);
xor U10872 (N_10872,N_503,N_6841);
or U10873 (N_10873,N_1571,N_2921);
nand U10874 (N_10874,N_9587,N_2949);
xnor U10875 (N_10875,N_2136,N_2292);
nor U10876 (N_10876,N_6035,N_7124);
nand U10877 (N_10877,N_9828,N_5195);
nor U10878 (N_10878,N_9036,N_2794);
nor U10879 (N_10879,N_8623,N_9746);
nand U10880 (N_10880,N_8138,N_9356);
nor U10881 (N_10881,N_7476,N_1044);
or U10882 (N_10882,N_828,N_6352);
and U10883 (N_10883,N_8764,N_8688);
or U10884 (N_10884,N_2453,N_6286);
nor U10885 (N_10885,N_8042,N_7230);
or U10886 (N_10886,N_2218,N_6580);
nor U10887 (N_10887,N_6396,N_4706);
nand U10888 (N_10888,N_1352,N_2529);
xor U10889 (N_10889,N_7315,N_7694);
nand U10890 (N_10890,N_7799,N_9122);
xnor U10891 (N_10891,N_7654,N_5834);
nor U10892 (N_10892,N_1990,N_3067);
and U10893 (N_10893,N_5306,N_1364);
or U10894 (N_10894,N_4217,N_6739);
and U10895 (N_10895,N_4624,N_4187);
nand U10896 (N_10896,N_36,N_5662);
nor U10897 (N_10897,N_1745,N_4532);
or U10898 (N_10898,N_4400,N_8825);
xor U10899 (N_10899,N_1208,N_1126);
or U10900 (N_10900,N_6879,N_7811);
and U10901 (N_10901,N_4813,N_3854);
nor U10902 (N_10902,N_4430,N_2338);
xnor U10903 (N_10903,N_7512,N_2253);
nand U10904 (N_10904,N_3142,N_2573);
or U10905 (N_10905,N_8118,N_6322);
or U10906 (N_10906,N_8429,N_7580);
or U10907 (N_10907,N_1514,N_9948);
and U10908 (N_10908,N_2433,N_7744);
nor U10909 (N_10909,N_7491,N_1719);
and U10910 (N_10910,N_7358,N_440);
or U10911 (N_10911,N_363,N_6705);
or U10912 (N_10912,N_3745,N_3950);
nor U10913 (N_10913,N_8998,N_6809);
nand U10914 (N_10914,N_387,N_4853);
or U10915 (N_10915,N_7987,N_9760);
nand U10916 (N_10916,N_6374,N_3972);
nand U10917 (N_10917,N_5547,N_7797);
or U10918 (N_10918,N_836,N_151);
nand U10919 (N_10919,N_4344,N_2471);
xor U10920 (N_10920,N_8386,N_4491);
nand U10921 (N_10921,N_2232,N_9735);
nand U10922 (N_10922,N_6656,N_6470);
or U10923 (N_10923,N_2225,N_246);
nand U10924 (N_10924,N_453,N_3319);
or U10925 (N_10925,N_2878,N_761);
or U10926 (N_10926,N_1167,N_3934);
and U10927 (N_10927,N_5896,N_8143);
nor U10928 (N_10928,N_3452,N_7099);
and U10929 (N_10929,N_4972,N_7494);
nor U10930 (N_10930,N_8528,N_8631);
or U10931 (N_10931,N_9691,N_7203);
nand U10932 (N_10932,N_9236,N_6056);
nor U10933 (N_10933,N_5890,N_8077);
and U10934 (N_10934,N_831,N_8110);
xor U10935 (N_10935,N_8018,N_1397);
xnor U10936 (N_10936,N_1102,N_9890);
and U10937 (N_10937,N_8123,N_7040);
nor U10938 (N_10938,N_8437,N_8696);
nor U10939 (N_10939,N_2760,N_645);
or U10940 (N_10940,N_7869,N_2704);
and U10941 (N_10941,N_7050,N_2348);
and U10942 (N_10942,N_6668,N_4069);
and U10943 (N_10943,N_1976,N_2604);
or U10944 (N_10944,N_2469,N_5881);
nand U10945 (N_10945,N_1240,N_971);
nor U10946 (N_10946,N_9230,N_6104);
nand U10947 (N_10947,N_2504,N_3825);
or U10948 (N_10948,N_4421,N_8278);
nor U10949 (N_10949,N_2308,N_1133);
and U10950 (N_10950,N_4351,N_9469);
nor U10951 (N_10951,N_5568,N_5687);
or U10952 (N_10952,N_5453,N_1519);
xnor U10953 (N_10953,N_1729,N_7466);
and U10954 (N_10954,N_8774,N_1148);
nor U10955 (N_10955,N_9040,N_5868);
and U10956 (N_10956,N_9588,N_1907);
nand U10957 (N_10957,N_2637,N_3600);
nor U10958 (N_10958,N_8326,N_8593);
and U10959 (N_10959,N_684,N_3290);
or U10960 (N_10960,N_8970,N_9368);
and U10961 (N_10961,N_875,N_2138);
nand U10962 (N_10962,N_4307,N_1908);
xnor U10963 (N_10963,N_1718,N_8877);
nor U10964 (N_10964,N_4668,N_870);
nand U10965 (N_10965,N_532,N_637);
nand U10966 (N_10966,N_9179,N_6546);
nor U10967 (N_10967,N_4956,N_8658);
xnor U10968 (N_10968,N_3562,N_6166);
nand U10969 (N_10969,N_6683,N_4478);
or U10970 (N_10970,N_8757,N_1544);
and U10971 (N_10971,N_1591,N_7629);
and U10972 (N_10972,N_6001,N_3766);
and U10973 (N_10973,N_5075,N_858);
nand U10974 (N_10974,N_9984,N_3912);
or U10975 (N_10975,N_6524,N_615);
nand U10976 (N_10976,N_9504,N_3419);
nand U10977 (N_10977,N_1071,N_2456);
or U10978 (N_10978,N_3995,N_6659);
nor U10979 (N_10979,N_3572,N_1410);
nor U10980 (N_10980,N_7389,N_9963);
or U10981 (N_10981,N_8358,N_2489);
and U10982 (N_10982,N_2081,N_1778);
or U10983 (N_10983,N_9896,N_9364);
nand U10984 (N_10984,N_4767,N_4462);
nand U10985 (N_10985,N_8327,N_6515);
nand U10986 (N_10986,N_8989,N_6288);
nor U10987 (N_10987,N_8710,N_8235);
nand U10988 (N_10988,N_620,N_2112);
and U10989 (N_10989,N_9909,N_7248);
nor U10990 (N_10990,N_27,N_328);
nand U10991 (N_10991,N_2022,N_7502);
nor U10992 (N_10992,N_9539,N_7828);
nand U10993 (N_10993,N_4144,N_3450);
nand U10994 (N_10994,N_5364,N_7773);
xnor U10995 (N_10995,N_4113,N_9920);
xor U10996 (N_10996,N_2289,N_1441);
and U10997 (N_10997,N_2773,N_5729);
xnor U10998 (N_10998,N_1792,N_6350);
or U10999 (N_10999,N_1695,N_1638);
nand U11000 (N_11000,N_4311,N_7420);
xnor U11001 (N_11001,N_1331,N_6773);
xnor U11002 (N_11002,N_5657,N_7709);
or U11003 (N_11003,N_9067,N_70);
and U11004 (N_11004,N_5243,N_263);
nor U11005 (N_11005,N_7028,N_4765);
nand U11006 (N_11006,N_788,N_5225);
and U11007 (N_11007,N_4343,N_4815);
xnor U11008 (N_11008,N_4642,N_1750);
nand U11009 (N_11009,N_6266,N_8810);
or U11010 (N_11010,N_8219,N_3181);
and U11011 (N_11011,N_3373,N_8149);
xor U11012 (N_11012,N_7880,N_1798);
and U11013 (N_11013,N_3756,N_9659);
nor U11014 (N_11014,N_2283,N_327);
nand U11015 (N_11015,N_6095,N_183);
or U11016 (N_11016,N_7971,N_9987);
or U11017 (N_11017,N_389,N_2160);
or U11018 (N_11018,N_1524,N_8733);
nor U11019 (N_11019,N_3717,N_8691);
xor U11020 (N_11020,N_3881,N_8869);
xor U11021 (N_11021,N_6950,N_9755);
or U11022 (N_11022,N_3528,N_9239);
and U11023 (N_11023,N_6625,N_5806);
nor U11024 (N_11024,N_7152,N_8846);
and U11025 (N_11025,N_1559,N_4929);
nand U11026 (N_11026,N_2045,N_1707);
nor U11027 (N_11027,N_3918,N_2440);
nor U11028 (N_11028,N_3143,N_3431);
and U11029 (N_11029,N_9709,N_8220);
or U11030 (N_11030,N_4076,N_6589);
or U11031 (N_11031,N_3982,N_8517);
and U11032 (N_11032,N_1564,N_5382);
nand U11033 (N_11033,N_4753,N_4665);
xnor U11034 (N_11034,N_7405,N_1405);
xor U11035 (N_11035,N_1614,N_4764);
nand U11036 (N_11036,N_6042,N_4406);
or U11037 (N_11037,N_5755,N_9583);
or U11038 (N_11038,N_2585,N_4782);
and U11039 (N_11039,N_211,N_2992);
and U11040 (N_11040,N_843,N_2801);
nor U11041 (N_11041,N_3335,N_2275);
nand U11042 (N_11042,N_3492,N_7860);
or U11043 (N_11043,N_9993,N_9851);
xor U11044 (N_11044,N_5571,N_1375);
nand U11045 (N_11045,N_7912,N_9579);
nand U11046 (N_11046,N_5256,N_9541);
or U11047 (N_11047,N_6365,N_3613);
or U11048 (N_11048,N_6433,N_5155);
nand U11049 (N_11049,N_1270,N_3645);
nand U11050 (N_11050,N_9600,N_8181);
xor U11051 (N_11051,N_8783,N_9424);
xor U11052 (N_11052,N_3405,N_7788);
xor U11053 (N_11053,N_7370,N_9888);
or U11054 (N_11054,N_8755,N_1301);
nor U11055 (N_11055,N_2206,N_9206);
nand U11056 (N_11056,N_6884,N_5846);
and U11057 (N_11057,N_7123,N_9129);
nor U11058 (N_11058,N_2115,N_2727);
nor U11059 (N_11059,N_9944,N_2272);
or U11060 (N_11060,N_8887,N_5625);
xnor U11061 (N_11061,N_7332,N_1342);
and U11062 (N_11062,N_8804,N_6121);
and U11063 (N_11063,N_7149,N_9283);
and U11064 (N_11064,N_6125,N_5507);
or U11065 (N_11065,N_6896,N_2667);
and U11066 (N_11066,N_8971,N_6681);
nand U11067 (N_11067,N_2990,N_983);
nor U11068 (N_11068,N_9505,N_7451);
nand U11069 (N_11069,N_4439,N_388);
or U11070 (N_11070,N_1926,N_9163);
nor U11071 (N_11071,N_3191,N_7461);
nor U11072 (N_11072,N_7102,N_2845);
or U11073 (N_11073,N_5778,N_1478);
or U11074 (N_11074,N_6483,N_6988);
nor U11075 (N_11075,N_4993,N_4978);
nand U11076 (N_11076,N_8019,N_8369);
or U11077 (N_11077,N_3548,N_2143);
or U11078 (N_11078,N_5558,N_3608);
nor U11079 (N_11079,N_1081,N_6617);
and U11080 (N_11080,N_4918,N_9087);
xor U11081 (N_11081,N_8061,N_5016);
and U11082 (N_11082,N_6255,N_3911);
nor U11083 (N_11083,N_6259,N_5449);
nand U11084 (N_11084,N_6941,N_306);
or U11085 (N_11085,N_2079,N_7199);
and U11086 (N_11086,N_9366,N_4966);
and U11087 (N_11087,N_2239,N_945);
xnor U11088 (N_11088,N_618,N_9196);
and U11089 (N_11089,N_4717,N_1481);
and U11090 (N_11090,N_2805,N_5436);
nor U11091 (N_11091,N_4593,N_9425);
or U11092 (N_11092,N_6099,N_8036);
and U11093 (N_11093,N_2006,N_786);
or U11094 (N_11094,N_2077,N_5276);
and U11095 (N_11095,N_2742,N_5844);
and U11096 (N_11096,N_8638,N_1517);
nand U11097 (N_11097,N_1315,N_290);
nor U11098 (N_11098,N_3890,N_4024);
xnor U11099 (N_11099,N_2854,N_7982);
nand U11100 (N_11100,N_278,N_7159);
nand U11101 (N_11101,N_5954,N_185);
and U11102 (N_11102,N_1398,N_6298);
nand U11103 (N_11103,N_2973,N_1530);
and U11104 (N_11104,N_1055,N_9429);
or U11105 (N_11105,N_4616,N_9164);
and U11106 (N_11106,N_8725,N_3096);
nor U11107 (N_11107,N_7651,N_5543);
or U11108 (N_11108,N_1669,N_4433);
and U11109 (N_11109,N_2335,N_6943);
and U11110 (N_11110,N_4316,N_5963);
nand U11111 (N_11111,N_6087,N_4377);
or U11112 (N_11112,N_6192,N_1494);
xnor U11113 (N_11113,N_2770,N_438);
nand U11114 (N_11114,N_9419,N_4269);
or U11115 (N_11115,N_3865,N_2391);
and U11116 (N_11116,N_611,N_1222);
or U11117 (N_11117,N_4025,N_4038);
nand U11118 (N_11118,N_2371,N_8113);
and U11119 (N_11119,N_8088,N_8966);
xnor U11120 (N_11120,N_8321,N_4429);
and U11121 (N_11121,N_7109,N_45);
xnor U11122 (N_11122,N_4185,N_2243);
nor U11123 (N_11123,N_398,N_3165);
nor U11124 (N_11124,N_9870,N_3706);
nor U11125 (N_11125,N_9874,N_5439);
xnor U11126 (N_11126,N_1327,N_2759);
and U11127 (N_11127,N_4730,N_1969);
or U11128 (N_11128,N_8204,N_5866);
or U11129 (N_11129,N_8285,N_6387);
nand U11130 (N_11130,N_4823,N_6978);
nor U11131 (N_11131,N_7276,N_3166);
and U11132 (N_11132,N_9617,N_7746);
nor U11133 (N_11133,N_5616,N_1365);
nand U11134 (N_11134,N_9511,N_7809);
nand U11135 (N_11135,N_9756,N_1730);
or U11136 (N_11136,N_5961,N_2813);
or U11137 (N_11137,N_5820,N_2734);
nand U11138 (N_11138,N_1877,N_7368);
and U11139 (N_11139,N_8850,N_9766);
or U11140 (N_11140,N_2832,N_9460);
nor U11141 (N_11141,N_6926,N_4342);
and U11142 (N_11142,N_8360,N_5293);
nor U11143 (N_11143,N_9633,N_561);
or U11144 (N_11144,N_9073,N_9342);
nand U11145 (N_11145,N_7051,N_1382);
xnor U11146 (N_11146,N_4107,N_5044);
and U11147 (N_11147,N_2639,N_787);
nand U11148 (N_11148,N_5208,N_9013);
nor U11149 (N_11149,N_7106,N_3718);
nand U11150 (N_11150,N_1847,N_5333);
or U11151 (N_11151,N_792,N_4988);
nor U11152 (N_11152,N_6226,N_3757);
or U11153 (N_11153,N_9235,N_4545);
and U11154 (N_11154,N_7387,N_8413);
xor U11155 (N_11155,N_9000,N_2642);
and U11156 (N_11156,N_7076,N_9822);
or U11157 (N_11157,N_84,N_2953);
or U11158 (N_11158,N_53,N_6473);
nor U11159 (N_11159,N_7837,N_669);
nand U11160 (N_11160,N_4747,N_4565);
and U11161 (N_11161,N_6711,N_9434);
or U11162 (N_11162,N_98,N_9729);
or U11163 (N_11163,N_8367,N_1249);
and U11164 (N_11164,N_7093,N_6666);
nor U11165 (N_11165,N_1401,N_8261);
nor U11166 (N_11166,N_2728,N_2843);
or U11167 (N_11167,N_3859,N_9734);
or U11168 (N_11168,N_969,N_5560);
nor U11169 (N_11169,N_1578,N_4451);
and U11170 (N_11170,N_334,N_6247);
and U11171 (N_11171,N_9811,N_1552);
nand U11172 (N_11172,N_1333,N_8064);
or U11173 (N_11173,N_2424,N_2983);
and U11174 (N_11174,N_7631,N_4872);
nor U11175 (N_11175,N_1251,N_8553);
and U11176 (N_11176,N_4164,N_7004);
xnor U11177 (N_11177,N_252,N_6427);
nor U11178 (N_11178,N_8150,N_7377);
and U11179 (N_11179,N_3194,N_5357);
nor U11180 (N_11180,N_9212,N_2611);
xnor U11181 (N_11181,N_8486,N_6193);
or U11182 (N_11182,N_9704,N_9863);
or U11183 (N_11183,N_998,N_6028);
xnor U11184 (N_11184,N_5508,N_8170);
and U11185 (N_11185,N_3015,N_716);
nand U11186 (N_11186,N_3367,N_4761);
nor U11187 (N_11187,N_8828,N_9813);
xor U11188 (N_11188,N_5533,N_7118);
or U11189 (N_11189,N_447,N_2991);
or U11190 (N_11190,N_5115,N_2317);
nand U11191 (N_11191,N_1770,N_4255);
or U11192 (N_11192,N_1005,N_7622);
nand U11193 (N_11193,N_1136,N_9688);
nor U11194 (N_11194,N_1603,N_1143);
nor U11195 (N_11195,N_7520,N_9162);
xor U11196 (N_11196,N_1099,N_1672);
or U11197 (N_11197,N_7190,N_158);
nor U11198 (N_11198,N_935,N_9677);
xnor U11199 (N_11199,N_9513,N_3902);
nor U11200 (N_11200,N_5123,N_6053);
nand U11201 (N_11201,N_7609,N_9359);
nor U11202 (N_11202,N_2028,N_4296);
and U11203 (N_11203,N_9442,N_3949);
nand U11204 (N_11204,N_9092,N_8281);
xnor U11205 (N_11205,N_8650,N_4692);
and U11206 (N_11206,N_6586,N_8689);
xnor U11207 (N_11207,N_2689,N_111);
nor U11208 (N_11208,N_1025,N_4749);
nand U11209 (N_11209,N_5448,N_563);
nor U11210 (N_11210,N_702,N_3687);
nor U11211 (N_11211,N_7992,N_7090);
or U11212 (N_11212,N_9506,N_592);
and U11213 (N_11213,N_5837,N_5940);
nand U11214 (N_11214,N_3435,N_4889);
nand U11215 (N_11215,N_9723,N_9330);
xnor U11216 (N_11216,N_4672,N_1881);
xnor U11217 (N_11217,N_1359,N_8565);
or U11218 (N_11218,N_4864,N_1290);
and U11219 (N_11219,N_520,N_754);
xnor U11220 (N_11220,N_638,N_4181);
nand U11221 (N_11221,N_1995,N_3936);
nand U11222 (N_11222,N_8381,N_1879);
nand U11223 (N_11223,N_7556,N_5504);
or U11224 (N_11224,N_6768,N_7128);
nand U11225 (N_11225,N_1388,N_6636);
or U11226 (N_11226,N_5180,N_2325);
or U11227 (N_11227,N_1628,N_1363);
and U11228 (N_11228,N_8656,N_1294);
or U11229 (N_11229,N_854,N_4784);
and U11230 (N_11230,N_9114,N_2196);
nand U11231 (N_11231,N_7114,N_4597);
nand U11232 (N_11232,N_4120,N_2188);
nand U11233 (N_11233,N_9885,N_9638);
nand U11234 (N_11234,N_5926,N_4557);
and U11235 (N_11235,N_5414,N_8589);
nand U11236 (N_11236,N_8742,N_3605);
nor U11237 (N_11237,N_5022,N_7696);
and U11238 (N_11238,N_4898,N_5966);
or U11239 (N_11239,N_5482,N_8122);
nor U11240 (N_11240,N_9571,N_7252);
and U11241 (N_11241,N_6567,N_3561);
nand U11242 (N_11242,N_5006,N_3073);
or U11243 (N_11243,N_8477,N_1067);
and U11244 (N_11244,N_2564,N_9884);
or U11245 (N_11245,N_2899,N_9326);
nand U11246 (N_11246,N_6614,N_7157);
nor U11247 (N_11247,N_9027,N_9086);
or U11248 (N_11248,N_2178,N_9384);
nor U11249 (N_11249,N_4607,N_5785);
nor U11250 (N_11250,N_7897,N_9233);
or U11251 (N_11251,N_406,N_7397);
and U11252 (N_11252,N_5024,N_4034);
and U11253 (N_11253,N_8737,N_4322);
nor U11254 (N_11254,N_6282,N_8826);
nor U11255 (N_11255,N_1393,N_725);
and U11256 (N_11256,N_15,N_9082);
nand U11257 (N_11257,N_6590,N_1472);
nand U11258 (N_11258,N_6948,N_5863);
xnor U11259 (N_11259,N_1916,N_4786);
nor U11260 (N_11260,N_3649,N_9549);
or U11261 (N_11261,N_2161,N_3023);
nand U11262 (N_11262,N_3261,N_9250);
nand U11263 (N_11263,N_1555,N_3837);
and U11264 (N_11264,N_4727,N_8622);
nor U11265 (N_11265,N_7733,N_4568);
nand U11266 (N_11266,N_6898,N_9899);
nor U11267 (N_11267,N_8491,N_2297);
and U11268 (N_11268,N_2882,N_4386);
and U11269 (N_11269,N_3242,N_6582);
and U11270 (N_11270,N_6649,N_5633);
or U11271 (N_11271,N_6167,N_9263);
or U11272 (N_11272,N_7137,N_3331);
nand U11273 (N_11273,N_3636,N_9942);
and U11274 (N_11274,N_1726,N_606);
and U11275 (N_11275,N_8000,N_245);
or U11276 (N_11276,N_4754,N_7990);
or U11277 (N_11277,N_519,N_1015);
or U11278 (N_11278,N_5203,N_6876);
xnor U11279 (N_11279,N_6102,N_8874);
nor U11280 (N_11280,N_8448,N_7977);
nor U11281 (N_11281,N_7139,N_6510);
and U11282 (N_11282,N_4551,N_6734);
or U11283 (N_11283,N_237,N_8653);
xor U11284 (N_11284,N_6740,N_4950);
nor U11285 (N_11285,N_6399,N_5958);
and U11286 (N_11286,N_6878,N_5312);
xor U11287 (N_11287,N_9831,N_3624);
nand U11288 (N_11288,N_3461,N_3641);
nor U11289 (N_11289,N_3806,N_7572);
nand U11290 (N_11290,N_6682,N_176);
nand U11291 (N_11291,N_1900,N_8584);
xor U11292 (N_11292,N_9860,N_7287);
and U11293 (N_11293,N_3787,N_7408);
nand U11294 (N_11294,N_7934,N_9246);
or U11295 (N_11295,N_126,N_8471);
nand U11296 (N_11296,N_5073,N_6423);
or U11297 (N_11297,N_6531,N_1725);
and U11298 (N_11298,N_8093,N_5430);
and U11299 (N_11299,N_3132,N_8102);
nor U11300 (N_11300,N_2125,N_2119);
or U11301 (N_11301,N_4236,N_3567);
nand U11302 (N_11302,N_1561,N_6511);
nand U11303 (N_11303,N_2144,N_5098);
and U11304 (N_11304,N_9629,N_6194);
nand U11305 (N_11305,N_6412,N_3571);
xor U11306 (N_11306,N_4846,N_2939);
xor U11307 (N_11307,N_7436,N_8331);
nand U11308 (N_11308,N_595,N_5077);
or U11309 (N_11309,N_3108,N_7867);
nor U11310 (N_11310,N_9975,N_267);
or U11311 (N_11311,N_6435,N_225);
and U11312 (N_11312,N_7985,N_5553);
and U11313 (N_11313,N_688,N_1656);
or U11314 (N_11314,N_4110,N_9391);
nor U11315 (N_11315,N_1187,N_3475);
nand U11316 (N_11316,N_4639,N_3868);
nand U11317 (N_11317,N_7832,N_5192);
nand U11318 (N_11318,N_6482,N_3754);
and U11319 (N_11319,N_1932,N_1178);
nand U11320 (N_11320,N_6345,N_5917);
and U11321 (N_11321,N_9957,N_3357);
xnor U11322 (N_11322,N_2789,N_6475);
nor U11323 (N_11323,N_9088,N_5945);
nand U11324 (N_11324,N_769,N_5091);
nor U11325 (N_11325,N_4569,N_5781);
or U11326 (N_11326,N_4994,N_1938);
xor U11327 (N_11327,N_4454,N_9492);
xnor U11328 (N_11328,N_1550,N_1370);
and U11329 (N_11329,N_9133,N_597);
or U11330 (N_11330,N_1723,N_6871);
xnor U11331 (N_11331,N_66,N_1182);
nor U11332 (N_11332,N_6616,N_4664);
nand U11333 (N_11333,N_3482,N_2539);
or U11334 (N_11334,N_9722,N_9265);
or U11335 (N_11335,N_7951,N_3296);
xnor U11336 (N_11336,N_3117,N_5757);
nand U11337 (N_11337,N_4952,N_5209);
xor U11338 (N_11338,N_8751,N_7589);
nand U11339 (N_11339,N_5532,N_179);
nand U11340 (N_11340,N_1901,N_6378);
or U11341 (N_11341,N_9561,N_8207);
nand U11342 (N_11342,N_481,N_3480);
or U11343 (N_11343,N_4211,N_7910);
and U11344 (N_11344,N_2565,N_5051);
and U11345 (N_11345,N_7256,N_3853);
and U11346 (N_11346,N_2978,N_6647);
nor U11347 (N_11347,N_9060,N_719);
and U11348 (N_11348,N_9663,N_5308);
nor U11349 (N_11349,N_2408,N_7163);
nand U11350 (N_11350,N_1553,N_9883);
or U11351 (N_11351,N_8533,N_1602);
and U11352 (N_11352,N_137,N_8858);
or U11353 (N_11353,N_8464,N_8578);
or U11354 (N_11354,N_6886,N_4282);
and U11355 (N_11355,N_3746,N_9954);
xor U11356 (N_11356,N_7523,N_3235);
nor U11357 (N_11357,N_9090,N_7447);
or U11358 (N_11358,N_7056,N_9120);
xnor U11359 (N_11359,N_878,N_5813);
and U11360 (N_11360,N_2976,N_5268);
nor U11361 (N_11361,N_4332,N_661);
nand U11362 (N_11362,N_4315,N_5315);
and U11363 (N_11363,N_7318,N_1761);
or U11364 (N_11364,N_711,N_814);
nand U11365 (N_11365,N_5129,N_9083);
nand U11366 (N_11366,N_9421,N_6627);
and U11367 (N_11367,N_8754,N_4635);
nor U11368 (N_11368,N_8459,N_9444);
and U11369 (N_11369,N_9482,N_3976);
nand U11370 (N_11370,N_1768,N_5758);
and U11371 (N_11371,N_1722,N_6147);
xor U11372 (N_11372,N_4090,N_8112);
nand U11373 (N_11373,N_6965,N_2531);
nor U11374 (N_11374,N_6276,N_5366);
or U11375 (N_11375,N_4509,N_4900);
and U11376 (N_11376,N_1810,N_3059);
or U11377 (N_11377,N_8678,N_1985);
nor U11378 (N_11378,N_2201,N_9172);
nand U11379 (N_11379,N_7308,N_4957);
and U11380 (N_11380,N_748,N_4149);
or U11381 (N_11381,N_6942,N_8264);
xnor U11382 (N_11382,N_2321,N_5415);
nand U11383 (N_11383,N_2815,N_4204);
or U11384 (N_11384,N_8803,N_5546);
nand U11385 (N_11385,N_1560,N_1248);
or U11386 (N_11386,N_8662,N_2234);
or U11387 (N_11387,N_1788,N_1889);
nor U11388 (N_11388,N_8211,N_6906);
and U11389 (N_11389,N_6369,N_3674);
nor U11390 (N_11390,N_7854,N_9730);
and U11391 (N_11391,N_3734,N_7866);
or U11392 (N_11392,N_7782,N_3252);
and U11393 (N_11393,N_8510,N_8343);
nor U11394 (N_11394,N_6490,N_5303);
or U11395 (N_11395,N_940,N_5304);
and U11396 (N_11396,N_382,N_460);
nor U11397 (N_11397,N_9522,N_7037);
and U11398 (N_11398,N_2755,N_3574);
nand U11399 (N_11399,N_833,N_3268);
nor U11400 (N_11400,N_3871,N_4520);
and U11401 (N_11401,N_8266,N_7012);
xor U11402 (N_11402,N_2448,N_4513);
nor U11403 (N_11403,N_6296,N_8404);
and U11404 (N_11404,N_5808,N_5143);
xor U11405 (N_11405,N_4037,N_819);
or U11406 (N_11406,N_7127,N_1886);
or U11407 (N_11407,N_7013,N_8104);
or U11408 (N_11408,N_1174,N_5215);
or U11409 (N_11409,N_5318,N_7335);
nor U11410 (N_11410,N_2235,N_4547);
nand U11411 (N_11411,N_9193,N_9074);
nand U11412 (N_11412,N_4559,N_1387);
or U11413 (N_11413,N_282,N_3763);
nor U11414 (N_11414,N_9597,N_9671);
or U11415 (N_11415,N_8959,N_923);
nor U11416 (N_11416,N_7425,N_5464);
nand U11417 (N_11417,N_1659,N_2102);
nand U11418 (N_11418,N_9573,N_5974);
or U11419 (N_11419,N_720,N_291);
xnor U11420 (N_11420,N_5375,N_7193);
and U11421 (N_11421,N_485,N_8179);
or U11422 (N_11422,N_1097,N_6213);
nand U11423 (N_11423,N_5965,N_7376);
nand U11424 (N_11424,N_3771,N_964);
or U11425 (N_11425,N_4744,N_9491);
nor U11426 (N_11426,N_6641,N_6153);
nand U11427 (N_11427,N_7621,N_1696);
or U11428 (N_11428,N_2977,N_1353);
and U11429 (N_11429,N_8514,N_4924);
nand U11430 (N_11430,N_5970,N_5549);
and U11431 (N_11431,N_6660,N_9907);
and U11432 (N_11432,N_7077,N_8778);
and U11433 (N_11433,N_1580,N_181);
and U11434 (N_11434,N_7002,N_62);
and U11435 (N_11435,N_2057,N_2221);
nand U11436 (N_11436,N_3123,N_3952);
xnor U11437 (N_11437,N_3535,N_7850);
or U11438 (N_11438,N_7403,N_1666);
xnor U11439 (N_11439,N_3885,N_1260);
nor U11440 (N_11440,N_981,N_7391);
and U11441 (N_11441,N_7201,N_5742);
nand U11442 (N_11442,N_3392,N_65);
nor U11443 (N_11443,N_9893,N_4420);
or U11444 (N_11444,N_9190,N_5193);
nand U11445 (N_11445,N_8902,N_9401);
or U11446 (N_11446,N_3207,N_7355);
nand U11447 (N_11447,N_6713,N_6924);
xnor U11448 (N_11448,N_2684,N_1038);
and U11449 (N_11449,N_642,N_3595);
nor U11450 (N_11450,N_7755,N_4130);
or U11451 (N_11451,N_8005,N_7092);
and U11452 (N_11452,N_9440,N_700);
and U11453 (N_11453,N_9015,N_8505);
nand U11454 (N_11454,N_4294,N_2127);
or U11455 (N_11455,N_3230,N_4912);
or U11456 (N_11456,N_8292,N_2599);
nand U11457 (N_11457,N_9319,N_6355);
nand U11458 (N_11458,N_7607,N_340);
nor U11459 (N_11459,N_5058,N_472);
nor U11460 (N_11460,N_5876,N_3581);
nor U11461 (N_11461,N_7978,N_1335);
and U11462 (N_11462,N_9103,N_5269);
and U11463 (N_11463,N_5065,N_3106);
or U11464 (N_11464,N_3121,N_376);
and U11465 (N_11465,N_459,N_7946);
nand U11466 (N_11466,N_3043,N_2644);
nand U11467 (N_11467,N_771,N_2806);
and U11468 (N_11468,N_9224,N_6772);
and U11469 (N_11469,N_9867,N_6203);
and U11470 (N_11470,N_3195,N_8621);
nor U11471 (N_11471,N_4710,N_8859);
nand U11472 (N_11472,N_9641,N_3538);
nand U11473 (N_11473,N_4227,N_1491);
nand U11474 (N_11474,N_9528,N_497);
nor U11475 (N_11475,N_8777,N_2807);
nand U11476 (N_11476,N_8260,N_4735);
or U11477 (N_11477,N_496,N_7278);
and U11478 (N_11478,N_4650,N_4198);
or U11479 (N_11479,N_6219,N_5994);
xor U11480 (N_11480,N_889,N_4608);
or U11481 (N_11481,N_9762,N_3157);
and U11482 (N_11482,N_4939,N_106);
xnor U11483 (N_11483,N_5407,N_7372);
and U11484 (N_11484,N_5166,N_6444);
nand U11485 (N_11485,N_8315,N_8081);
nor U11486 (N_11486,N_6535,N_4732);
nand U11487 (N_11487,N_8069,N_6856);
nand U11488 (N_11488,N_2166,N_3518);
or U11489 (N_11489,N_8685,N_1776);
or U11490 (N_11490,N_6330,N_8619);
nand U11491 (N_11491,N_94,N_1775);
and U11492 (N_11492,N_8425,N_8079);
and U11493 (N_11493,N_9123,N_5814);
nor U11494 (N_11494,N_7055,N_7416);
nand U11495 (N_11495,N_9273,N_9218);
nor U11496 (N_11496,N_9821,N_6457);
or U11497 (N_11497,N_1468,N_950);
or U11498 (N_11498,N_2554,N_7481);
nor U11499 (N_11499,N_7080,N_1763);
nor U11500 (N_11500,N_6929,N_1466);
nor U11501 (N_11501,N_7957,N_1967);
nor U11502 (N_11502,N_3898,N_3758);
nor U11503 (N_11503,N_665,N_2968);
nor U11504 (N_11504,N_5957,N_3502);
or U11505 (N_11505,N_723,N_3558);
xor U11506 (N_11506,N_3277,N_3489);
nor U11507 (N_11507,N_3267,N_3839);
or U11508 (N_11508,N_9267,N_1068);
xnor U11509 (N_11509,N_5358,N_7806);
nor U11510 (N_11510,N_2525,N_4193);
nand U11511 (N_11511,N_9486,N_261);
nand U11512 (N_11512,N_7326,N_4460);
or U11513 (N_11513,N_4364,N_9718);
or U11514 (N_11514,N_495,N_9472);
nor U11515 (N_11515,N_8111,N_1934);
or U11516 (N_11516,N_5678,N_5653);
xnor U11517 (N_11517,N_4700,N_9803);
or U11518 (N_11518,N_1286,N_7762);
nand U11519 (N_11519,N_1054,N_1039);
or U11520 (N_11520,N_9753,N_5355);
and U11521 (N_11521,N_7838,N_7168);
nor U11522 (N_11522,N_3917,N_9296);
or U11523 (N_11523,N_8334,N_2581);
xor U11524 (N_11524,N_5079,N_5344);
and U11525 (N_11525,N_7233,N_3983);
nor U11526 (N_11526,N_2631,N_5700);
nand U11527 (N_11527,N_5721,N_6097);
nor U11528 (N_11528,N_8727,N_6626);
xor U11529 (N_11529,N_7954,N_6010);
xor U11530 (N_11530,N_2994,N_8787);
or U11531 (N_11531,N_3623,N_8604);
and U11532 (N_11532,N_4498,N_1406);
and U11533 (N_11533,N_5234,N_8855);
nor U11534 (N_11534,N_5250,N_3529);
or U11535 (N_11535,N_3657,N_205);
and U11536 (N_11536,N_9645,N_9854);
and U11537 (N_11537,N_6716,N_2501);
xor U11538 (N_11538,N_9961,N_7530);
nor U11539 (N_11539,N_848,N_1613);
and U11540 (N_11540,N_9841,N_4303);
nand U11541 (N_11541,N_916,N_4690);
or U11542 (N_11542,N_5096,N_5673);
and U11543 (N_11543,N_9106,N_6008);
xnor U11544 (N_11544,N_7587,N_4151);
nand U11545 (N_11545,N_6853,N_549);
and U11546 (N_11546,N_6326,N_8272);
and U11547 (N_11547,N_9100,N_3177);
or U11548 (N_11548,N_1838,N_435);
nor U11549 (N_11549,N_8004,N_6080);
or U11550 (N_11550,N_9478,N_6);
nand U11551 (N_11551,N_368,N_4359);
nand U11552 (N_11552,N_3740,N_9968);
and U11553 (N_11553,N_4991,N_1690);
and U11554 (N_11554,N_6671,N_5591);
or U11555 (N_11555,N_8142,N_3777);
or U11556 (N_11556,N_9566,N_6579);
nand U11557 (N_11557,N_9983,N_350);
and U11558 (N_11558,N_1651,N_9322);
nand U11559 (N_11559,N_3024,N_2213);
or U11560 (N_11560,N_6527,N_3925);
nand U11561 (N_11561,N_7918,N_7497);
xnor U11562 (N_11562,N_1100,N_8108);
nand U11563 (N_11563,N_1132,N_5154);
and U11564 (N_11564,N_1989,N_7858);
nand U11565 (N_11565,N_5564,N_751);
and U11566 (N_11566,N_5109,N_3753);
or U11567 (N_11567,N_9105,N_7927);
or U11568 (N_11568,N_1367,N_2909);
nor U11569 (N_11569,N_9991,N_5389);
and U11570 (N_11570,N_139,N_6507);
nand U11571 (N_11571,N_9824,N_4792);
nor U11572 (N_11572,N_8838,N_2624);
and U11573 (N_11573,N_6182,N_2679);
and U11574 (N_11574,N_3822,N_3801);
or U11575 (N_11575,N_2840,N_8475);
nand U11576 (N_11576,N_1053,N_1677);
xor U11577 (N_11577,N_5451,N_4136);
and U11578 (N_11578,N_5299,N_777);
or U11579 (N_11579,N_8830,N_587);
nand U11580 (N_11580,N_9341,N_9568);
nand U11581 (N_11581,N_8405,N_9169);
or U11582 (N_11582,N_5913,N_3094);
or U11583 (N_11583,N_2095,N_1771);
or U11584 (N_11584,N_7944,N_4500);
nand U11585 (N_11585,N_6849,N_7122);
xor U11586 (N_11586,N_3222,N_1851);
nand U11587 (N_11587,N_474,N_1488);
and U11588 (N_11588,N_7698,N_68);
nand U11589 (N_11589,N_502,N_6393);
or U11590 (N_11590,N_4837,N_6553);
or U11591 (N_11591,N_8351,N_3879);
and U11592 (N_11592,N_2724,N_6526);
xor U11593 (N_11593,N_9834,N_6766);
nor U11594 (N_11594,N_3552,N_2402);
nor U11595 (N_11595,N_7597,N_5226);
and U11596 (N_11596,N_5779,N_76);
nor U11597 (N_11597,N_4514,N_9737);
or U11598 (N_11598,N_5390,N_7066);
nor U11599 (N_11599,N_8611,N_3644);
nand U11600 (N_11600,N_6388,N_19);
nor U11601 (N_11601,N_5658,N_7460);
xnor U11602 (N_11602,N_2411,N_2327);
and U11603 (N_11603,N_7732,N_5114);
or U11604 (N_11604,N_8146,N_3001);
xnor U11605 (N_11605,N_6724,N_8603);
or U11606 (N_11606,N_8635,N_6200);
xor U11607 (N_11607,N_4094,N_5294);
nand U11608 (N_11608,N_8436,N_9307);
or U11609 (N_11609,N_3112,N_635);
nor U11610 (N_11610,N_8344,N_924);
nand U11611 (N_11611,N_316,N_659);
and U11612 (N_11612,N_9856,N_7619);
xnor U11613 (N_11613,N_8421,N_3397);
nor U11614 (N_11614,N_9614,N_3975);
and U11615 (N_11615,N_3199,N_3485);
nor U11616 (N_11616,N_3616,N_7324);
xor U11617 (N_11617,N_899,N_7682);
nand U11618 (N_11618,N_6866,N_8379);
or U11619 (N_11619,N_8799,N_9201);
nor U11620 (N_11620,N_7274,N_3274);
and U11621 (N_11621,N_8529,N_7999);
nor U11622 (N_11622,N_7398,N_3907);
xnor U11623 (N_11623,N_1453,N_6363);
nand U11624 (N_11624,N_8750,N_7455);
or U11625 (N_11625,N_918,N_7218);
or U11626 (N_11626,N_957,N_3842);
nand U11627 (N_11627,N_835,N_893);
nand U11628 (N_11628,N_6111,N_2185);
nor U11629 (N_11629,N_5331,N_8472);
nor U11630 (N_11630,N_4539,N_9682);
nor U11631 (N_11631,N_6672,N_6972);
nor U11632 (N_11632,N_1827,N_8608);
and U11633 (N_11633,N_5204,N_103);
nor U11634 (N_11634,N_6290,N_4243);
xor U11635 (N_11635,N_288,N_5596);
nor U11636 (N_11636,N_8612,N_9777);
nand U11637 (N_11637,N_2005,N_6927);
and U11638 (N_11638,N_2462,N_1826);
nand U11639 (N_11639,N_8536,N_7402);
and U11640 (N_11640,N_6480,N_7655);
nor U11641 (N_11641,N_5683,N_8675);
nor U11642 (N_11642,N_3152,N_9306);
nand U11643 (N_11643,N_3751,N_7615);
nand U11644 (N_11644,N_9810,N_8686);
nand U11645 (N_11645,N_7891,N_1293);
and U11646 (N_11646,N_8474,N_3305);
and U11647 (N_11647,N_5394,N_6584);
xor U11648 (N_11648,N_5947,N_3028);
nand U11649 (N_11649,N_6532,N_6163);
or U11650 (N_11650,N_2082,N_8955);
and U11651 (N_11651,N_2013,N_9276);
or U11652 (N_11652,N_9622,N_29);
nand U11653 (N_11653,N_8258,N_6175);
xor U11654 (N_11654,N_3799,N_7108);
and U11655 (N_11655,N_358,N_9433);
nor U11656 (N_11656,N_6395,N_3258);
and U11657 (N_11657,N_8829,N_3632);
and U11658 (N_11658,N_5692,N_6273);
and U11659 (N_11659,N_3279,N_6344);
nand U11660 (N_11660,N_4969,N_3690);
nor U11661 (N_11661,N_8029,N_7382);
and U11662 (N_11662,N_5551,N_7275);
nor U11663 (N_11663,N_349,N_3794);
nor U11664 (N_11664,N_6651,N_3102);
nand U11665 (N_11665,N_3504,N_5731);
nand U11666 (N_11666,N_8493,N_7524);
xnor U11667 (N_11667,N_8229,N_3371);
or U11668 (N_11668,N_1287,N_7756);
nand U11669 (N_11669,N_7846,N_7462);
xnor U11670 (N_11670,N_9058,N_8994);
nor U11671 (N_11671,N_6474,N_8099);
nor U11672 (N_11672,N_8060,N_8633);
nand U11673 (N_11673,N_9759,N_6987);
or U11674 (N_11674,N_4330,N_9362);
or U11675 (N_11675,N_4339,N_5157);
nand U11676 (N_11676,N_3573,N_5386);
nand U11677 (N_11677,N_2363,N_2709);
xnor U11678 (N_11678,N_5350,N_689);
or U11679 (N_11679,N_9146,N_5539);
and U11680 (N_11680,N_9006,N_2097);
and U11681 (N_11681,N_2584,N_559);
nand U11682 (N_11682,N_9562,N_6603);
and U11683 (N_11683,N_9950,N_7543);
nand U11684 (N_11684,N_9695,N_9784);
xor U11685 (N_11685,N_3980,N_9798);
and U11686 (N_11686,N_5664,N_7039);
or U11687 (N_11687,N_8463,N_6759);
xnor U11688 (N_11688,N_6551,N_8726);
and U11689 (N_11689,N_6021,N_6565);
nor U11690 (N_11690,N_5149,N_2675);
nor U11691 (N_11691,N_1993,N_1052);
or U11692 (N_11692,N_9051,N_5074);
or U11693 (N_11693,N_9623,N_5197);
and U11694 (N_11694,N_8588,N_980);
and U11695 (N_11695,N_2382,N_2656);
nor U11696 (N_11696,N_7468,N_9535);
and U11697 (N_11697,N_8286,N_6891);
nor U11698 (N_11698,N_8234,N_7329);
and U11699 (N_11699,N_273,N_9738);
xnor U11700 (N_11700,N_2499,N_1922);
or U11701 (N_11701,N_544,N_286);
nand U11702 (N_11702,N_3111,N_2601);
nor U11703 (N_11703,N_4139,N_7904);
xnor U11704 (N_11704,N_7166,N_9456);
or U11705 (N_11705,N_8002,N_4746);
nor U11706 (N_11706,N_5595,N_5815);
or U11707 (N_11707,N_652,N_571);
and U11708 (N_11708,N_1344,N_174);
nor U11709 (N_11709,N_6919,N_2262);
and U11710 (N_11710,N_9295,N_7664);
nand U11711 (N_11711,N_2873,N_2720);
or U11712 (N_11712,N_4023,N_9689);
nor U11713 (N_11713,N_5495,N_1034);
or U11714 (N_11714,N_895,N_1246);
nor U11715 (N_11715,N_2286,N_7);
or U11716 (N_11716,N_8007,N_4206);
and U11717 (N_11717,N_6402,N_9383);
nand U11718 (N_11718,N_4066,N_2086);
nor U11719 (N_11719,N_9225,N_3615);
or U11720 (N_11720,N_5003,N_5544);
nand U11721 (N_11721,N_4526,N_7165);
nor U11722 (N_11722,N_1980,N_9519);
nand U11723 (N_11723,N_2683,N_395);
or U11724 (N_11724,N_696,N_1549);
nand U11725 (N_11725,N_515,N_2528);
and U11726 (N_11726,N_1064,N_9145);
nor U11727 (N_11727,N_2149,N_2857);
nor U11728 (N_11728,N_8452,N_9072);
nand U11729 (N_11729,N_5951,N_1506);
nor U11730 (N_11730,N_5088,N_5403);
or U11731 (N_11731,N_5270,N_3724);
or U11732 (N_11732,N_690,N_3609);
and U11733 (N_11733,N_8904,N_2646);
or U11734 (N_11734,N_8137,N_2170);
or U11735 (N_11735,N_4127,N_2694);
nand U11736 (N_11736,N_4337,N_361);
nand U11737 (N_11737,N_8371,N_3463);
nand U11738 (N_11738,N_7881,N_8503);
nand U11739 (N_11739,N_9805,N_9395);
or U11740 (N_11740,N_8011,N_7527);
xor U11741 (N_11741,N_5369,N_1551);
nor U11742 (N_11742,N_5265,N_3403);
or U11743 (N_11743,N_8058,N_9902);
and U11744 (N_11744,N_1979,N_2298);
nor U11745 (N_11745,N_9512,N_379);
and U11746 (N_11746,N_6190,N_7169);
nor U11747 (N_11747,N_4791,N_4899);
nand U11748 (N_11748,N_9642,N_2666);
or U11749 (N_11749,N_4317,N_2700);
and U11750 (N_11750,N_5246,N_4142);
nand U11751 (N_11751,N_8599,N_6680);
and U11752 (N_11752,N_9757,N_6836);
nand U11753 (N_11753,N_8306,N_196);
nand U11754 (N_11754,N_3610,N_2947);
nand U11755 (N_11755,N_7795,N_3612);
nor U11756 (N_11756,N_8936,N_6731);
nand U11757 (N_11757,N_9291,N_6794);
and U11758 (N_11758,N_3214,N_4372);
nor U11759 (N_11759,N_120,N_8249);
or U11760 (N_11760,N_6937,N_7889);
and U11761 (N_11761,N_4838,N_5179);
nand U11762 (N_11762,N_8848,N_556);
nand U11763 (N_11763,N_3661,N_5901);
and U11764 (N_11764,N_6360,N_5978);
nand U11765 (N_11765,N_7299,N_7996);
xnor U11766 (N_11766,N_2910,N_5371);
and U11767 (N_11767,N_6191,N_910);
nand U11768 (N_11768,N_9344,N_664);
nand U11769 (N_11769,N_8610,N_4402);
nand U11770 (N_11770,N_1557,N_7714);
xor U11771 (N_11771,N_4106,N_9457);
nor U11772 (N_11772,N_6631,N_4855);
xnor U11773 (N_11773,N_7538,N_8022);
nor U11774 (N_11774,N_5600,N_4455);
or U11775 (N_11775,N_9044,N_1000);
nand U11776 (N_11776,N_3382,N_6090);
or U11777 (N_11777,N_6763,N_2522);
or U11778 (N_11778,N_7126,N_5404);
nor U11779 (N_11779,N_5262,N_2008);
nand U11780 (N_11780,N_7125,N_4739);
nor U11781 (N_11781,N_5709,N_6870);
nor U11782 (N_11782,N_407,N_9850);
nand U11783 (N_11783,N_2906,N_7413);
or U11784 (N_11784,N_1273,N_6307);
or U11785 (N_11785,N_2850,N_707);
or U11786 (N_11786,N_586,N_7899);
nand U11787 (N_11787,N_6120,N_4863);
or U11788 (N_11788,N_3339,N_3175);
and U11789 (N_11789,N_3432,N_5650);
nand U11790 (N_11790,N_2106,N_8563);
nand U11791 (N_11791,N_996,N_6109);
nand U11792 (N_11792,N_7499,N_3356);
nand U11793 (N_11793,N_7847,N_7824);
and U11794 (N_11794,N_5422,N_1870);
nand U11795 (N_11795,N_6161,N_9436);
and U11796 (N_11796,N_9363,N_8961);
nand U11797 (N_11797,N_8059,N_1667);
and U11798 (N_11798,N_8419,N_9618);
or U11799 (N_11799,N_311,N_8746);
or U11800 (N_11800,N_4043,N_857);
nor U11801 (N_11801,N_9662,N_5853);
nand U11802 (N_11802,N_23,N_3321);
nor U11803 (N_11803,N_7485,N_9286);
nand U11804 (N_11804,N_2147,N_1115);
nand U11805 (N_11805,N_3428,N_4649);
xnor U11806 (N_11806,N_6268,N_1774);
or U11807 (N_11807,N_465,N_8176);
or U11808 (N_11808,N_613,N_5899);
and U11809 (N_11809,N_4542,N_6520);
and U11810 (N_11810,N_5100,N_8896);
and U11811 (N_11811,N_2767,N_3714);
nand U11812 (N_11812,N_7006,N_9409);
or U11813 (N_11813,N_498,N_6076);
nor U11814 (N_11814,N_9978,N_4875);
nand U11815 (N_11815,N_1258,N_1843);
or U11816 (N_11816,N_4248,N_8652);
nor U11817 (N_11817,N_7522,N_2290);
and U11818 (N_11818,N_3673,N_6629);
nand U11819 (N_11819,N_4108,N_8270);
and U11820 (N_11820,N_2154,N_408);
nor U11821 (N_11821,N_1874,N_5867);
or U11822 (N_11822,N_1676,N_7264);
and U11823 (N_11823,N_4314,N_874);
nand U11824 (N_11824,N_5251,N_3929);
nand U11825 (N_11825,N_8100,N_72);
and U11826 (N_11826,N_5167,N_3512);
and U11827 (N_11827,N_6242,N_793);
xor U11828 (N_11828,N_6271,N_3809);
xor U11829 (N_11829,N_3695,N_5374);
and U11830 (N_11830,N_341,N_6083);
or U11831 (N_11831,N_5214,N_2941);
nand U11832 (N_11832,N_7060,N_3793);
or U11833 (N_11833,N_681,N_8269);
nor U11834 (N_11834,N_364,N_8284);
xnor U11835 (N_11835,N_9144,N_3337);
nor U11836 (N_11836,N_9337,N_9200);
xor U11837 (N_11837,N_59,N_7726);
or U11838 (N_11838,N_5346,N_7776);
xor U11839 (N_11839,N_6945,N_5925);
and U11840 (N_11840,N_6902,N_948);
nand U11841 (N_11841,N_861,N_4655);
nor U11842 (N_11842,N_284,N_5485);
nand U11843 (N_11843,N_52,N_9394);
nand U11844 (N_11844,N_4397,N_3966);
nand U11845 (N_11845,N_7463,N_2260);
and U11846 (N_11846,N_3709,N_4577);
and U11847 (N_11847,N_9800,N_6323);
nand U11848 (N_11848,N_192,N_3867);
xor U11849 (N_11849,N_7647,N_4794);
nand U11850 (N_11850,N_3308,N_8876);
nor U11851 (N_11851,N_4238,N_5918);
and U11852 (N_11852,N_2364,N_5008);
xor U11853 (N_11853,N_1662,N_1931);
and U11854 (N_11854,N_7151,N_8230);
nand U11855 (N_11855,N_5649,N_2314);
nand U11856 (N_11856,N_9990,N_2555);
nand U11857 (N_11857,N_7663,N_2049);
xnor U11858 (N_11858,N_5764,N_5391);
nor U11859 (N_11859,N_1191,N_3448);
nand U11860 (N_11860,N_8744,N_5613);
or U11861 (N_11861,N_5168,N_5311);
and U11862 (N_11862,N_345,N_884);
and U11863 (N_11863,N_7182,N_2063);
nor U11864 (N_11864,N_7211,N_5036);
nor U11865 (N_11865,N_7410,N_8492);
nor U11866 (N_11866,N_1343,N_4971);
xor U11867 (N_11867,N_7839,N_5989);
or U11868 (N_11868,N_4827,N_5634);
or U11869 (N_11869,N_8242,N_9772);
xor U11870 (N_11870,N_7703,N_7594);
nand U11871 (N_11871,N_3002,N_1974);
xor U11872 (N_11872,N_9251,N_1391);
or U11873 (N_11873,N_7422,N_4161);
nor U11874 (N_11874,N_3408,N_3533);
nor U11875 (N_11875,N_1684,N_8151);
and U11876 (N_11876,N_2541,N_8626);
or U11877 (N_11877,N_7937,N_7793);
nand U11878 (N_11878,N_456,N_7686);
nand U11879 (N_11879,N_1486,N_1413);
nand U11880 (N_11880,N_4059,N_3184);
nor U11881 (N_11881,N_6928,N_8251);
nand U11882 (N_11882,N_1390,N_7515);
or U11883 (N_11883,N_900,N_1885);
xor U11884 (N_11884,N_5972,N_2804);
xnor U11885 (N_11885,N_4300,N_9627);
or U11886 (N_11886,N_8495,N_3783);
nand U11887 (N_11887,N_2399,N_5550);
nor U11888 (N_11888,N_2263,N_686);
or U11889 (N_11889,N_9985,N_6129);
nand U11890 (N_11890,N_7613,N_3870);
nand U11891 (N_11891,N_4276,N_277);
xnor U11892 (N_11892,N_1329,N_1913);
xor U11893 (N_11893,N_9501,N_3090);
or U11894 (N_11894,N_3941,N_9714);
nor U11895 (N_11895,N_5915,N_201);
and U11896 (N_11896,N_8136,N_2697);
xor U11897 (N_11897,N_621,N_3817);
and U11898 (N_11898,N_1254,N_5851);
nor U11899 (N_11899,N_4012,N_3703);
nor U11900 (N_11900,N_3840,N_9477);
xnor U11901 (N_11901,N_1469,N_3498);
nor U11902 (N_11902,N_3286,N_6336);
nor U11903 (N_11903,N_5895,N_8511);
nor U11904 (N_11904,N_5728,N_5206);
nand U11905 (N_11905,N_4953,N_5855);
or U11906 (N_11906,N_6976,N_8403);
or U11907 (N_11907,N_6598,N_8518);
nor U11908 (N_11908,N_5012,N_6217);
nor U11909 (N_11909,N_5380,N_5298);
or U11910 (N_11910,N_3424,N_8537);
nor U11911 (N_11911,N_2051,N_5590);
or U11912 (N_11912,N_4537,N_9639);
and U11913 (N_11913,N_567,N_6826);
nand U11914 (N_11914,N_9921,N_3052);
nor U11915 (N_11915,N_5934,N_6758);
or U11916 (N_11916,N_423,N_5891);
nor U11917 (N_11917,N_6872,N_3729);
and U11918 (N_11918,N_7614,N_3163);
nand U11919 (N_11919,N_8903,N_1116);
or U11920 (N_11920,N_3083,N_7540);
xor U11921 (N_11921,N_4931,N_3765);
or U11922 (N_11922,N_4600,N_7216);
nor U11923 (N_11923,N_4405,N_2792);
and U11924 (N_11924,N_7323,N_737);
or U11925 (N_11925,N_9143,N_1036);
xnor U11926 (N_11926,N_9842,N_7599);
nor U11927 (N_11927,N_9525,N_6903);
xor U11928 (N_11928,N_6691,N_1791);
or U11929 (N_11929,N_1448,N_8065);
nor U11930 (N_11930,N_6785,N_7338);
nand U11931 (N_11931,N_2723,N_6637);
nand U11932 (N_11932,N_4903,N_2269);
and U11933 (N_11933,N_727,N_2725);
xor U11934 (N_11934,N_9443,N_8325);
nand U11935 (N_11935,N_3107,N_1303);
and U11936 (N_11936,N_1597,N_4158);
or U11937 (N_11937,N_1767,N_8749);
or U11938 (N_11938,N_262,N_7374);
xor U11939 (N_11939,N_9077,N_4811);
nand U11940 (N_11940,N_5440,N_5457);
nor U11941 (N_11941,N_8674,N_2996);
and U11942 (N_11942,N_2398,N_1526);
nand U11943 (N_11943,N_5059,N_9198);
or U11944 (N_11944,N_9465,N_4885);
nand U11945 (N_11945,N_7459,N_4830);
nor U11946 (N_11946,N_4825,N_7593);
or U11947 (N_11947,N_427,N_3325);
or U11948 (N_11948,N_8476,N_1947);
and U11949 (N_11949,N_2535,N_2511);
nand U11950 (N_11950,N_535,N_1742);
or U11951 (N_11951,N_6611,N_5598);
nand U11952 (N_11952,N_7803,N_3439);
nor U11953 (N_11953,N_6717,N_2765);
or U11954 (N_11954,N_2821,N_7707);
or U11955 (N_11955,N_9721,N_3788);
nor U11956 (N_11956,N_6117,N_5807);
or U11957 (N_11957,N_4777,N_4854);
nor U11958 (N_11958,N_6912,N_9524);
and U11959 (N_11959,N_6177,N_6034);
and U11960 (N_11960,N_4425,N_4721);
nor U11961 (N_11961,N_1094,N_9289);
nand U11962 (N_11962,N_2917,N_9485);
nand U11963 (N_11963,N_8374,N_2191);
nand U11964 (N_11964,N_4549,N_7526);
nand U11965 (N_11965,N_1731,N_5902);
nor U11966 (N_11966,N_2717,N_8441);
nor U11967 (N_11967,N_2365,N_9298);
xor U11968 (N_11968,N_4653,N_7595);
nor U11969 (N_11969,N_9819,N_2674);
and U11970 (N_11970,N_5320,N_4541);
nor U11971 (N_11971,N_8050,N_2460);
or U11972 (N_11972,N_1428,N_5501);
xnor U11973 (N_11973,N_9300,N_4666);
nand U11974 (N_11974,N_1241,N_2366);
nand U11975 (N_11975,N_9381,N_7685);
nor U11976 (N_11976,N_7155,N_4098);
xnor U11977 (N_11977,N_809,N_2621);
nand U11978 (N_11978,N_5864,N_6250);
nor U11979 (N_11979,N_7222,N_1150);
or U11980 (N_11980,N_4594,N_3797);
or U11981 (N_11981,N_7603,N_3407);
nand U11982 (N_11982,N_538,N_1965);
xor U11983 (N_11983,N_9030,N_5676);
and U11984 (N_11984,N_7432,N_107);
xnor U11985 (N_11985,N_9859,N_2640);
nor U11986 (N_11986,N_4718,N_441);
or U11987 (N_11987,N_2738,N_475);
or U11988 (N_11988,N_8895,N_933);
nand U11989 (N_11989,N_1797,N_1590);
nor U11990 (N_11990,N_8447,N_8712);
or U11991 (N_11991,N_2018,N_926);
or U11992 (N_11992,N_476,N_6272);
nand U11993 (N_11993,N_8015,N_3888);
nor U11994 (N_11994,N_3249,N_7625);
xor U11995 (N_11995,N_7181,N_2784);
nor U11996 (N_11996,N_9104,N_8238);
nor U11997 (N_11997,N_1876,N_8566);
nor U11998 (N_11998,N_1400,N_8918);
nand U11999 (N_11999,N_110,N_8831);
xnor U12000 (N_12000,N_3149,N_2488);
or U12001 (N_12001,N_5597,N_1525);
nand U12002 (N_12002,N_8571,N_4807);
or U12003 (N_12003,N_3131,N_7385);
and U12004 (N_12004,N_6516,N_1795);
or U12005 (N_12005,N_6441,N_7089);
and U12006 (N_12006,N_555,N_9864);
nand U12007 (N_12007,N_3042,N_3666);
xor U12008 (N_12008,N_682,N_1743);
nor U12009 (N_12009,N_5151,N_63);
or U12010 (N_12010,N_7361,N_7650);
nand U12011 (N_12011,N_9608,N_683);
and U12012 (N_12012,N_9328,N_9521);
nor U12013 (N_12013,N_4515,N_8782);
or U12014 (N_12014,N_4556,N_9966);
and U12015 (N_12015,N_1957,N_2648);
and U12016 (N_12016,N_887,N_6011);
nor U12017 (N_12017,N_599,N_2961);
nor U12018 (N_12018,N_8335,N_9959);
or U12019 (N_12019,N_4958,N_2747);
and U12020 (N_12020,N_4223,N_8851);
or U12021 (N_12021,N_416,N_4173);
nand U12022 (N_12022,N_8615,N_4829);
nor U12023 (N_12023,N_1334,N_9613);
or U12024 (N_12024,N_3446,N_6189);
or U12025 (N_12025,N_1409,N_8630);
nand U12026 (N_12026,N_6545,N_7084);
or U12027 (N_12027,N_1622,N_6690);
nor U12028 (N_12028,N_7588,N_5019);
or U12029 (N_12029,N_3457,N_3156);
nand U12030 (N_12030,N_7774,N_1529);
nand U12031 (N_12031,N_6297,N_2128);
or U12032 (N_12032,N_1720,N_153);
or U12033 (N_12033,N_8280,N_6212);
nor U12034 (N_12034,N_8680,N_562);
nor U12035 (N_12035,N_6310,N_3035);
xor U12036 (N_12036,N_4674,N_8897);
and U12037 (N_12037,N_2417,N_6325);
and U12038 (N_12038,N_9675,N_7473);
nor U12039 (N_12039,N_1041,N_9173);
or U12040 (N_12040,N_6432,N_184);
and U12041 (N_12041,N_2436,N_7789);
nor U12042 (N_12042,N_2776,N_9830);
and U12043 (N_12043,N_3626,N_4606);
xnor U12044 (N_12044,N_7501,N_1300);
nand U12045 (N_12045,N_4998,N_3162);
nor U12046 (N_12046,N_8922,N_97);
and U12047 (N_12047,N_187,N_6486);
nor U12048 (N_12048,N_6348,N_4812);
or U12049 (N_12049,N_956,N_4169);
xor U12050 (N_12050,N_6489,N_9666);
or U12051 (N_12051,N_175,N_1946);
or U12052 (N_12052,N_9725,N_5870);
nor U12053 (N_12053,N_6894,N_1862);
nand U12054 (N_12054,N_5939,N_2817);
nor U12055 (N_12055,N_1588,N_344);
nor U12056 (N_12056,N_2902,N_804);
and U12057 (N_12057,N_5383,N_9894);
and U12058 (N_12058,N_9563,N_7984);
nor U12059 (N_12059,N_649,N_2319);
nand U12060 (N_12060,N_2603,N_3685);
nand U12061 (N_12061,N_6883,N_5466);
nand U12062 (N_12062,N_2078,N_1978);
and U12063 (N_12063,N_2811,N_4502);
and U12064 (N_12064,N_8906,N_8548);
nand U12065 (N_12065,N_7347,N_8668);
nor U12066 (N_12066,N_5632,N_9417);
or U12067 (N_12067,N_941,N_8409);
and U12068 (N_12068,N_8115,N_9892);
and U12069 (N_12069,N_4752,N_5583);
nand U12070 (N_12070,N_1283,N_3541);
nand U12071 (N_12071,N_7167,N_9797);
nand U12072 (N_12072,N_883,N_9393);
nand U12073 (N_12073,N_806,N_1449);
nand U12074 (N_12074,N_7448,N_922);
nor U12075 (N_12075,N_2868,N_1641);
or U12076 (N_12076,N_4525,N_2326);
nand U12077 (N_12077,N_9452,N_3509);
and U12078 (N_12078,N_2607,N_2268);
nand U12079 (N_12079,N_1137,N_2446);
and U12080 (N_12080,N_270,N_7514);
and U12081 (N_12081,N_4946,N_4410);
and U12082 (N_12082,N_7187,N_5838);
nor U12083 (N_12083,N_274,N_703);
or U12084 (N_12084,N_1257,N_1835);
xor U12085 (N_12085,N_7771,N_729);
xnor U12086 (N_12086,N_5609,N_9808);
and U12087 (N_12087,N_2625,N_2561);
nor U12088 (N_12088,N_156,N_1863);
nor U12089 (N_12089,N_2752,N_1896);
xnor U12090 (N_12090,N_2464,N_7250);
or U12091 (N_12091,N_2309,N_7148);
nor U12092 (N_12092,N_5640,N_1264);
nand U12093 (N_12093,N_1377,N_4471);
nor U12094 (N_12094,N_9243,N_7071);
nand U12095 (N_12095,N_321,N_3154);
nand U12096 (N_12096,N_5638,N_5624);
and U12097 (N_12097,N_3501,N_1840);
and U12098 (N_12098,N_8644,N_7433);
and U12099 (N_12099,N_5696,N_3401);
nand U12100 (N_12100,N_3508,N_25);
and U12101 (N_12101,N_5232,N_5774);
and U12102 (N_12102,N_8165,N_7892);
and U12103 (N_12103,N_1394,N_4004);
nor U12104 (N_12104,N_1074,N_1485);
and U12105 (N_12105,N_2318,N_1153);
or U12106 (N_12106,N_171,N_5672);
or U12107 (N_12107,N_990,N_3352);
nor U12108 (N_12108,N_5317,N_6119);
nand U12109 (N_12109,N_3161,N_3109);
or U12110 (N_12110,N_178,N_5773);
or U12111 (N_12111,N_3955,N_3078);
and U12112 (N_12112,N_9315,N_865);
nand U12113 (N_12113,N_2455,N_7349);
nor U12114 (N_12114,N_128,N_4374);
and U12115 (N_12115,N_1554,N_2575);
nor U12116 (N_12116,N_4622,N_6645);
or U12117 (N_12117,N_3361,N_3618);
xor U12118 (N_12118,N_4480,N_6897);
and U12119 (N_12119,N_9241,N_4961);
nand U12120 (N_12120,N_8485,N_2580);
and U12121 (N_12121,N_442,N_6574);
or U12122 (N_12122,N_209,N_6040);
and U12123 (N_12123,N_6969,N_1860);
or U12124 (N_12124,N_3155,N_9861);
nor U12125 (N_12125,N_6828,N_5871);
nor U12126 (N_12126,N_2277,N_581);
xnor U12127 (N_12127,N_2259,N_7495);
or U12128 (N_12128,N_3328,N_2658);
xor U12129 (N_12129,N_6830,N_3063);
or U12130 (N_12130,N_3832,N_7191);
nand U12131 (N_12131,N_3587,N_6825);
or U12132 (N_12132,N_5636,N_5888);
and U12133 (N_12133,N_7503,N_343);
nand U12134 (N_12134,N_9228,N_3203);
nor U12135 (N_12135,N_4426,N_3568);
nor U12136 (N_12136,N_8465,N_2856);
nand U12137 (N_12137,N_9712,N_7505);
nor U12138 (N_12138,N_7342,N_6869);
and U12139 (N_12139,N_3637,N_8657);
and U12140 (N_12140,N_9415,N_6292);
or U12141 (N_12141,N_5898,N_3324);
xor U12142 (N_12142,N_4419,N_8766);
xor U12143 (N_12143,N_9744,N_2543);
or U12144 (N_12144,N_5794,N_7835);
xnor U12145 (N_12145,N_7875,N_7023);
or U12146 (N_12146,N_7924,N_2702);
nor U12147 (N_12147,N_6697,N_7419);
xor U12148 (N_12148,N_909,N_8484);
or U12149 (N_12149,N_8431,N_939);
nand U12150 (N_12150,N_508,N_6834);
and U12151 (N_12151,N_2295,N_1829);
and U12152 (N_12152,N_8312,N_1754);
nand U12153 (N_12153,N_3722,N_7472);
and U12154 (N_12154,N_6218,N_9389);
nor U12155 (N_12155,N_8183,N_7712);
nand U12156 (N_12156,N_3250,N_3423);
or U12157 (N_12157,N_6338,N_4804);
nor U12158 (N_12158,N_6453,N_5938);
and U12159 (N_12159,N_791,N_7976);
nand U12160 (N_12160,N_4887,N_1177);
nand U12161 (N_12161,N_8038,N_5290);
nand U12162 (N_12162,N_3347,N_8824);
and U12163 (N_12163,N_8544,N_3150);
or U12164 (N_12164,N_255,N_5104);
xnor U12165 (N_12165,N_7421,N_2175);
xor U12166 (N_12166,N_9807,N_8221);
or U12167 (N_12167,N_1749,N_4907);
xor U12168 (N_12168,N_5092,N_2210);
nor U12169 (N_12169,N_807,N_3376);
or U12170 (N_12170,N_3785,N_4447);
nor U12171 (N_12171,N_3455,N_6209);
or U12172 (N_12172,N_2586,N_5412);
and U12173 (N_12173,N_1371,N_7681);
and U12174 (N_12174,N_3417,N_7240);
or U12175 (N_12175,N_6368,N_6974);
xnor U12176 (N_12176,N_310,N_6556);
nand U12177 (N_12177,N_5345,N_3990);
nand U12178 (N_12178,N_319,N_231);
and U12179 (N_12179,N_9702,N_4546);
and U12180 (N_12180,N_240,N_4620);
nor U12181 (N_12181,N_5822,N_425);
nor U12182 (N_12182,N_4371,N_7576);
and U12183 (N_12183,N_8393,N_3345);
nor U12184 (N_12184,N_8545,N_5163);
or U12185 (N_12185,N_2512,N_3427);
and U12186 (N_12186,N_7993,N_254);
nor U12187 (N_12187,N_4293,N_2816);
nor U12188 (N_12188,N_9445,N_7110);
nand U12189 (N_12189,N_6688,N_6468);
nor U12190 (N_12190,N_2346,N_5400);
xor U12191 (N_12191,N_6665,N_1212);
and U12192 (N_12192,N_6425,N_1269);
nor U12193 (N_12193,N_5399,N_9576);
nor U12194 (N_12194,N_2847,N_7477);
nand U12195 (N_12195,N_9399,N_3874);
nand U12196 (N_12196,N_4006,N_2300);
nand U12197 (N_12197,N_6155,N_7429);
and U12198 (N_12198,N_3606,N_5248);
nor U12199 (N_12199,N_7636,N_3084);
or U12200 (N_12200,N_44,N_533);
nor U12201 (N_12201,N_8422,N_6092);
nand U12202 (N_12202,N_1814,N_402);
nand U12203 (N_12203,N_2900,N_2014);
or U12204 (N_12204,N_1368,N_8560);
or U12205 (N_12205,N_5326,N_6953);
and U12206 (N_12206,N_3692,N_5879);
nor U12207 (N_12207,N_655,N_2482);
or U12208 (N_12208,N_2430,N_1479);
or U12209 (N_12209,N_4416,N_9768);
xor U12210 (N_12210,N_4512,N_491);
nand U12211 (N_12211,N_3137,N_3211);
nand U12212 (N_12212,N_2844,N_6525);
nand U12213 (N_12213,N_2665,N_8808);
and U12214 (N_12214,N_180,N_7238);
or U12215 (N_12215,N_4592,N_3327);
nand U12216 (N_12216,N_1275,N_3792);
xnor U12217 (N_12217,N_2828,N_2782);
and U12218 (N_12218,N_2320,N_5031);
or U12219 (N_12219,N_9158,N_1527);
xnor U12220 (N_12220,N_8761,N_6823);
nor U12221 (N_12221,N_6138,N_1682);
xnor U12222 (N_12222,N_1939,N_915);
nand U12223 (N_12223,N_1243,N_3653);
and U12224 (N_12224,N_8645,N_8620);
nand U12225 (N_12225,N_1773,N_3353);
nor U12226 (N_12226,N_9858,N_9410);
and U12227 (N_12227,N_3752,N_7626);
nor U12228 (N_12228,N_5724,N_6981);
and U12229 (N_12229,N_7489,N_3103);
and U12230 (N_12230,N_9880,N_9872);
or U12231 (N_12231,N_6075,N_8152);
nor U12232 (N_12232,N_5548,N_6471);
nor U12233 (N_12233,N_704,N_7657);
nor U12234 (N_12234,N_8372,N_9532);
nor U12235 (N_12235,N_7474,N_5426);
and U12236 (N_12236,N_4087,N_2988);
and U12237 (N_12237,N_2477,N_1281);
and U12238 (N_12238,N_9607,N_6469);
nand U12239 (N_12239,N_6058,N_2498);
nor U12240 (N_12240,N_5861,N_3433);
or U12241 (N_12241,N_902,N_9518);
nor U12242 (N_12242,N_8225,N_8978);
or U12243 (N_12243,N_5747,N_6566);
nand U12244 (N_12244,N_3151,N_5201);
or U12245 (N_12245,N_8523,N_1599);
xnor U12246 (N_12246,N_8125,N_5063);
and U12247 (N_12247,N_2422,N_4882);
nand U12248 (N_12248,N_4540,N_1781);
and U12249 (N_12249,N_8415,N_7234);
or U12250 (N_12250,N_8745,N_8434);
nor U12251 (N_12251,N_5178,N_1653);
nor U12252 (N_12252,N_2159,N_7787);
and U12253 (N_12253,N_2254,N_3510);
nor U12254 (N_12254,N_4602,N_5020);
nand U12255 (N_12255,N_1277,N_4516);
nor U12256 (N_12256,N_1772,N_2957);
or U12257 (N_12257,N_7135,N_2466);
or U12258 (N_12258,N_1587,N_4976);
nor U12259 (N_12259,N_1445,N_9392);
and U12260 (N_12260,N_6178,N_2266);
and U12261 (N_12261,N_3481,N_4028);
nor U12262 (N_12262,N_1027,N_4401);
or U12263 (N_12263,N_3055,N_6245);
nor U12264 (N_12264,N_8765,N_9101);
or U12265 (N_12265,N_7015,N_253);
nand U12266 (N_12266,N_3836,N_4859);
nor U12267 (N_12267,N_7748,N_4156);
or U12268 (N_12268,N_7021,N_7840);
nor U12269 (N_12269,N_1125,N_5469);
or U12270 (N_12270,N_9268,N_5110);
nor U12271 (N_12271,N_2613,N_4312);
nor U12272 (N_12272,N_6492,N_5593);
and U12273 (N_12273,N_7194,N_3171);
nor U12274 (N_12274,N_6009,N_2999);
or U12275 (N_12275,N_4191,N_1476);
nand U12276 (N_12276,N_9988,N_2438);
nor U12277 (N_12277,N_2852,N_6397);
or U12278 (N_12278,N_7297,N_7334);
and U12279 (N_12279,N_2785,N_3843);
or U12280 (N_12280,N_6267,N_7161);
nor U12281 (N_12281,N_7069,N_8857);
nand U12282 (N_12282,N_6694,N_9340);
or U12283 (N_12283,N_1543,N_512);
nor U12284 (N_12284,N_2871,N_8233);
nor U12285 (N_12285,N_694,N_116);
nor U12286 (N_12286,N_9919,N_5556);
and U12287 (N_12287,N_9581,N_4663);
nand U12288 (N_12288,N_5565,N_9474);
and U12289 (N_12289,N_2387,N_1420);
xnor U12290 (N_12290,N_8396,N_5574);
nor U12291 (N_12291,N_2238,N_2786);
nor U12292 (N_12292,N_4249,N_8732);
nand U12293 (N_12293,N_4053,N_2251);
nand U12294 (N_12294,N_2881,N_982);
nand U12295 (N_12295,N_2685,N_9646);
nor U12296 (N_12296,N_6628,N_7170);
and U12297 (N_12297,N_3813,N_2183);
nor U12298 (N_12298,N_1535,N_1030);
and U12299 (N_12299,N_6431,N_4884);
nor U12300 (N_12300,N_330,N_9266);
nor U12301 (N_12301,N_7065,N_8339);
or U12302 (N_12302,N_9426,N_2766);
or U12303 (N_12303,N_7307,N_457);
and U12304 (N_12304,N_7668,N_2247);
and U12305 (N_12305,N_9194,N_7112);
xor U12306 (N_12306,N_6201,N_5874);
xor U12307 (N_12307,N_4544,N_1484);
xor U12308 (N_12308,N_2622,N_750);
xor U12309 (N_12309,N_1450,N_7186);
and U12310 (N_12310,N_3398,N_7171);
or U12311 (N_12311,N_9278,N_2820);
xor U12312 (N_12312,N_1660,N_2447);
nor U12313 (N_12313,N_8410,N_6730);
nand U12314 (N_12314,N_8816,N_8201);
nand U12315 (N_12315,N_648,N_9832);
nand U12316 (N_12316,N_2970,N_9980);
and U12317 (N_12317,N_1569,N_3173);
nor U12318 (N_12318,N_800,N_4878);
nand U12319 (N_12319,N_1121,N_8254);
nand U12320 (N_12320,N_6460,N_4495);
nor U12321 (N_12321,N_2403,N_9713);
or U12322 (N_12322,N_8625,N_4822);
or U12323 (N_12323,N_7345,N_8762);
and U12324 (N_12324,N_8262,N_8614);
nor U12325 (N_12325,N_2393,N_1819);
nor U12326 (N_12326,N_7266,N_6664);
or U12327 (N_12327,N_5027,N_7660);
nor U12328 (N_12328,N_1362,N_9708);
nor U12329 (N_12329,N_6653,N_4118);
and U12330 (N_12330,N_5768,N_4103);
nand U12331 (N_12331,N_9733,N_9112);
or U12332 (N_12332,N_8889,N_5733);
or U12333 (N_12333,N_6677,N_5701);
and U12334 (N_12334,N_1480,N_3247);
nand U12335 (N_12335,N_9327,N_6195);
nand U12336 (N_12336,N_6693,N_380);
and U12337 (N_12337,N_7027,N_3259);
nor U12338 (N_12338,N_2245,N_6314);
nand U12339 (N_12339,N_1048,N_2955);
or U12340 (N_12340,N_2653,N_8715);
nand U12341 (N_12341,N_4917,N_3769);
or U12342 (N_12342,N_1157,N_7715);
nor U12343 (N_12343,N_8320,N_4370);
or U12344 (N_12344,N_8958,N_1147);
nand U12345 (N_12345,N_7337,N_6714);
nand U12346 (N_12346,N_3635,N_5479);
xnor U12347 (N_12347,N_3011,N_9188);
or U12348 (N_12348,N_3297,N_1866);
and U12349 (N_12349,N_1122,N_1330);
and U12350 (N_12350,N_2929,N_3700);
and U12351 (N_12351,N_3234,N_8809);
nand U12352 (N_12352,N_9370,N_236);
xnor U12353 (N_12353,N_5030,N_7000);
or U12354 (N_12354,N_1794,N_5041);
nand U12355 (N_12355,N_6127,N_5428);
or U12356 (N_12356,N_7751,N_6303);
or U12357 (N_12357,N_5138,N_2645);
xnor U12358 (N_12358,N_4714,N_3009);
xnor U12359 (N_12359,N_2791,N_6319);
and U12360 (N_12360,N_9089,N_9647);
nand U12361 (N_12361,N_4291,N_8428);
and U12362 (N_12362,N_9726,N_1339);
or U12363 (N_12363,N_1577,N_4355);
and U12364 (N_12364,N_2442,N_1694);
or U12365 (N_12365,N_6093,N_1670);
and U12366 (N_12366,N_7059,N_6502);
nand U12367 (N_12367,N_7667,N_6130);
xor U12368 (N_12368,N_5324,N_6935);
or U12369 (N_12369,N_6136,N_2187);
or U12370 (N_12370,N_2841,N_5257);
and U12371 (N_12371,N_7570,N_1386);
nor U12372 (N_12372,N_3017,N_8105);
or U12373 (N_12373,N_3326,N_9447);
nor U12374 (N_12374,N_217,N_8870);
or U12375 (N_12375,N_5072,N_3231);
and U12376 (N_12376,N_934,N_622);
nand U12377 (N_12377,N_6686,N_5162);
nor U12378 (N_12378,N_4008,N_5230);
and U12379 (N_12379,N_6676,N_6612);
and U12380 (N_12380,N_8985,N_3577);
xor U12381 (N_12381,N_6230,N_3219);
nand U12382 (N_12382,N_2521,N_3147);
xor U12383 (N_12383,N_3970,N_6461);
nand U12384 (N_12384,N_6411,N_4010);
nor U12385 (N_12385,N_4244,N_4598);
or U12386 (N_12386,N_2412,N_5738);
or U12387 (N_12387,N_8993,N_412);
xnor U12388 (N_12388,N_9945,N_609);
or U12389 (N_12389,N_1668,N_3861);
and U12390 (N_12390,N_5481,N_6542);
nor U12391 (N_12391,N_5477,N_422);
xor U12392 (N_12392,N_1605,N_5419);
and U12393 (N_12393,N_8451,N_8951);
and U12394 (N_12394,N_3539,N_4669);
xor U12395 (N_12395,N_5064,N_5433);
nor U12396 (N_12396,N_1853,N_1471);
nor U12397 (N_12397,N_4458,N_5631);
nand U12398 (N_12398,N_3285,N_8597);
nand U12399 (N_12399,N_4284,N_3316);
or U12400 (N_12400,N_1415,N_4152);
and U12401 (N_12401,N_322,N_657);
or U12402 (N_12402,N_7986,N_5411);
nor U12403 (N_12403,N_740,N_1953);
nor U12404 (N_12404,N_1728,N_1845);
nand U12405 (N_12405,N_3036,N_1268);
and U12406 (N_12406,N_6557,N_6704);
and U12407 (N_12407,N_7827,N_9710);
nor U12408 (N_12408,N_2696,N_5530);
or U12409 (N_12409,N_6662,N_9636);
nor U12410 (N_12410,N_2706,N_8389);
or U12411 (N_12411,N_917,N_8540);
nor U12412 (N_12412,N_8552,N_9514);
nand U12413 (N_12413,N_1658,N_1280);
nor U12414 (N_12414,N_6831,N_7082);
or U12415 (N_12415,N_7435,N_33);
or U12416 (N_12416,N_8947,N_7094);
nand U12417 (N_12417,N_6839,N_7030);
nand U12418 (N_12418,N_6381,N_7933);
nand U12419 (N_12419,N_1636,N_167);
nor U12420 (N_12420,N_8432,N_9427);
or U12421 (N_12421,N_780,N_5943);
nor U12422 (N_12422,N_7243,N_6454);
or U12423 (N_12423,N_984,N_9979);
nor U12424 (N_12424,N_3265,N_2746);
nand U12425 (N_12425,N_3686,N_976);
and U12426 (N_12426,N_6874,N_5490);
xor U12427 (N_12427,N_1454,N_4135);
nor U12428 (N_12428,N_3940,N_8756);
or U12429 (N_12429,N_6829,N_2296);
nand U12430 (N_12430,N_7673,N_7719);
nand U12431 (N_12431,N_5474,N_1407);
nand U12432 (N_12432,N_842,N_22);
or U12433 (N_12433,N_3553,N_742);
nand U12434 (N_12434,N_3887,N_9247);
nor U12435 (N_12435,N_4921,N_4340);
or U12436 (N_12436,N_1446,N_4221);
nor U12437 (N_12437,N_9181,N_8909);
nor U12438 (N_12438,N_2407,N_6802);
nor U12439 (N_12439,N_9601,N_738);
or U12440 (N_12440,N_1804,N_3830);
nand U12441 (N_12441,N_5827,N_2034);
or U12442 (N_12442,N_2591,N_6873);
and U12443 (N_12443,N_147,N_1735);
and U12444 (N_12444,N_5460,N_4469);
and U12445 (N_12445,N_9693,N_3767);
or U12446 (N_12446,N_5667,N_1323);
and U12447 (N_12447,N_3478,N_4346);
and U12448 (N_12448,N_7861,N_5906);
and U12449 (N_12449,N_4091,N_6503);
nand U12450 (N_12450,N_2148,N_1873);
nor U12451 (N_12451,N_5580,N_1784);
and U12452 (N_12452,N_3965,N_9543);
nand U12453 (N_12453,N_1961,N_6875);
nor U12454 (N_12454,N_6722,N_7111);
or U12455 (N_12455,N_8884,N_1467);
and U12456 (N_12456,N_5668,N_5792);
nand U12457 (N_12457,N_3313,N_7319);
or U12458 (N_12458,N_6775,N_5291);
and U12459 (N_12459,N_4876,N_400);
nand U12460 (N_12460,N_1070,N_3160);
xnor U12461 (N_12461,N_7034,N_279);
nor U12462 (N_12462,N_591,N_1316);
and U12463 (N_12463,N_3049,N_2635);
and U12464 (N_12464,N_5987,N_1219);
and U12465 (N_12465,N_1403,N_5165);
xor U12466 (N_12466,N_2285,N_7925);
nand U12467 (N_12467,N_7710,N_7537);
or U12468 (N_12468,N_9222,N_7259);
or U12469 (N_12469,N_4077,N_3831);
nor U12470 (N_12470,N_5821,N_4232);
or U12471 (N_12471,N_7511,N_1824);
or U12472 (N_12472,N_8718,N_6440);
nor U12473 (N_12473,N_3270,N_4711);
nor U12474 (N_12474,N_7578,N_8590);
nand U12475 (N_12475,N_8420,N_8931);
nor U12476 (N_12476,N_8148,N_5894);
nand U12477 (N_12477,N_7500,N_6540);
nand U12478 (N_12478,N_1322,N_5995);
nand U12479 (N_12479,N_7509,N_4197);
and U12480 (N_12480,N_2517,N_359);
nand U12481 (N_12481,N_367,N_5889);
and U12482 (N_12482,N_6364,N_8983);
nor U12483 (N_12483,N_1262,N_3875);
and U12484 (N_12484,N_8047,N_6813);
nand U12485 (N_12485,N_4129,N_8535);
nand U12486 (N_12486,N_42,N_8913);
and U12487 (N_12487,N_3764,N_1596);
nand U12488 (N_12488,N_7490,N_9657);
and U12489 (N_12489,N_7952,N_5880);
or U12490 (N_12490,N_6012,N_4001);
or U12491 (N_12491,N_484,N_5760);
or U12492 (N_12492,N_2869,N_4437);
or U12493 (N_12493,N_3430,N_5011);
or U12494 (N_12494,N_8106,N_4277);
nor U12495 (N_12495,N_8649,N_8636);
xnor U12496 (N_12496,N_8390,N_4477);
nand U12497 (N_12497,N_6429,N_4800);
and U12498 (N_12498,N_1859,N_5810);
and U12499 (N_12499,N_3054,N_2169);
nand U12500 (N_12500,N_8341,N_4189);
or U12501 (N_12501,N_7919,N_5486);
nor U12502 (N_12502,N_8414,N_6655);
or U12503 (N_12503,N_5431,N_4044);
and U12504 (N_12504,N_2429,N_2610);
xnor U12505 (N_12505,N_1854,N_445);
nor U12506 (N_12506,N_7551,N_8595);
nor U12507 (N_12507,N_9171,N_9598);
and U12508 (N_12508,N_7706,N_4793);
and U12509 (N_12509,N_1547,N_3759);
nor U12510 (N_12510,N_5935,N_3453);
and U12511 (N_12511,N_8676,N_5200);
and U12512 (N_12512,N_3176,N_3805);
nor U12513 (N_12513,N_1114,N_9254);
or U12514 (N_12514,N_2682,N_3470);
nor U12515 (N_12515,N_5136,N_1261);
nor U12516 (N_12516,N_3814,N_4769);
xnor U12517 (N_12517,N_7882,N_5620);
nor U12518 (N_12518,N_8232,N_5438);
or U12519 (N_12519,N_6317,N_7180);
or U12520 (N_12520,N_5285,N_3991);
or U12521 (N_12521,N_3997,N_4133);
and U12522 (N_12522,N_721,N_8191);
xor U12523 (N_12523,N_1001,N_6448);
or U12524 (N_12524,N_4832,N_3496);
or U12525 (N_12525,N_5635,N_9932);
and U12526 (N_12526,N_2749,N_6315);
or U12527 (N_12527,N_7816,N_830);
and U12528 (N_12528,N_5354,N_7263);
xnor U12529 (N_12529,N_4558,N_5971);
or U12530 (N_12530,N_4131,N_881);
nor U12531 (N_12531,N_8964,N_2818);
or U12532 (N_12532,N_6782,N_2509);
nand U12533 (N_12533,N_6496,N_1762);
nand U12534 (N_12534,N_9217,N_8833);
xnor U12535 (N_12535,N_985,N_5014);
nor U12536 (N_12536,N_170,N_8066);
nand U12537 (N_12537,N_5347,N_2437);
or U12538 (N_12538,N_3388,N_5283);
nor U12539 (N_12539,N_2526,N_75);
nand U12540 (N_12540,N_3322,N_5659);
and U12541 (N_12541,N_7508,N_6518);
xor U12542 (N_12542,N_6091,N_4680);
and U12543 (N_12543,N_1513,N_1539);
or U12544 (N_12544,N_685,N_2345);
nand U12545 (N_12545,N_7281,N_4159);
nand U12546 (N_12546,N_5708,N_9);
nand U12547 (N_12547,N_5698,N_3774);
nand U12548 (N_12548,N_470,N_7870);
nand U12549 (N_12549,N_8248,N_730);
and U12550 (N_12550,N_6858,N_9009);
nor U12551 (N_12551,N_1224,N_6952);
nor U12552 (N_12552,N_6909,N_9570);
and U12553 (N_12553,N_6394,N_4654);
or U12554 (N_12554,N_6004,N_4689);
nand U12555 (N_12555,N_634,N_2486);
and U12556 (N_12556,N_6278,N_7005);
nor U12557 (N_12557,N_5582,N_4768);
and U12558 (N_12558,N_4778,N_5468);
or U12559 (N_12559,N_4264,N_5186);
or U12560 (N_12560,N_1960,N_2582);
nand U12561 (N_12561,N_348,N_9376);
and U12562 (N_12562,N_8307,N_3095);
nand U12563 (N_12563,N_2396,N_2950);
and U12564 (N_12564,N_9448,N_3821);
nand U12565 (N_12565,N_1536,N_3556);
or U12566 (N_12566,N_6284,N_429);
nor U12567 (N_12567,N_8051,N_8806);
nor U12568 (N_12568,N_3969,N_8487);
and U12569 (N_12569,N_6733,N_1820);
and U12570 (N_12570,N_756,N_3377);
nor U12571 (N_12571,N_2956,N_409);
and U12572 (N_12572,N_5999,N_714);
or U12573 (N_12573,N_8938,N_2692);
or U12574 (N_12574,N_215,N_774);
nand U12575 (N_12575,N_431,N_8345);
xnor U12576 (N_12576,N_9685,N_9747);
nor U12577 (N_12577,N_5601,N_2514);
nor U12578 (N_12578,N_3097,N_9620);
and U12579 (N_12579,N_864,N_4319);
xor U12580 (N_12580,N_8083,N_529);
or U12581 (N_12581,N_7303,N_7519);
nand U12582 (N_12582,N_2484,N_7017);
nand U12583 (N_12583,N_6533,N_312);
nor U12584 (N_12584,N_6081,N_4281);
nand U12585 (N_12585,N_8025,N_7902);
nor U12586 (N_12586,N_4926,N_5153);
xor U12587 (N_12587,N_243,N_9157);
nor U12588 (N_12588,N_414,N_4396);
or U12589 (N_12589,N_3323,N_9596);
nor U12590 (N_12590,N_6176,N_1063);
and U12591 (N_12591,N_9180,N_8342);
or U12592 (N_12592,N_1221,N_6277);
or U12593 (N_12593,N_6960,N_5651);
nor U12594 (N_12594,N_7731,N_4848);
xnor U12595 (N_12595,N_8822,N_7348);
and U12596 (N_12596,N_3349,N_3984);
or U12597 (N_12597,N_300,N_3878);
nor U12598 (N_12598,N_6788,N_2047);
nor U12599 (N_12599,N_8924,N_5423);
nor U12600 (N_12600,N_1255,N_4289);
or U12601 (N_12601,N_3139,N_1951);
or U12602 (N_12602,N_135,N_7178);
nand U12603 (N_12603,N_7968,N_6776);
or U12604 (N_12604,N_7253,N_4073);
xor U12605 (N_12605,N_7583,N_2439);
or U12606 (N_12606,N_2901,N_7516);
and U12607 (N_12607,N_2887,N_5196);
or U12608 (N_12608,N_7105,N_1061);
nor U12609 (N_12609,N_863,N_233);
nor U12610 (N_12610,N_3906,N_9302);
nand U12611 (N_12611,N_2710,N_547);
or U12612 (N_12612,N_797,N_3172);
nand U12613 (N_12613,N_6790,N_2395);
or U12614 (N_12614,N_4265,N_7415);
or U12615 (N_12615,N_4715,N_626);
and U12616 (N_12616,N_3196,N_8880);
and U12617 (N_12617,N_4304,N_8898);
nor U12618 (N_12618,N_3977,N_4631);
or U12619 (N_12619,N_7796,N_3607);
and U12620 (N_12620,N_1124,N_5976);
nand U12621 (N_12621,N_4687,N_6184);
and U12622 (N_12622,N_6456,N_8382);
and U12623 (N_12623,N_6424,N_7249);
nand U12624 (N_12624,N_4411,N_2059);
nor U12625 (N_12625,N_7738,N_8655);
or U12626 (N_12626,N_8006,N_8348);
nand U12627 (N_12627,N_7016,N_4511);
and U12628 (N_12628,N_3872,N_4309);
nand U12629 (N_12629,N_8660,N_9716);
nand U12630 (N_12630,N_1372,N_943);
xor U12631 (N_12631,N_6762,N_5829);
xor U12632 (N_12632,N_9397,N_7845);
and U12633 (N_12633,N_4435,N_2255);
nand U12634 (N_12634,N_891,N_7452);
and U12635 (N_12635,N_8793,N_7441);
and U12636 (N_12636,N_5183,N_1460);
and U12637 (N_12637,N_2715,N_3062);
and U12638 (N_12638,N_2381,N_1163);
nor U12639 (N_12639,N_9303,N_3506);
or U12640 (N_12640,N_7569,N_9107);
nor U12641 (N_12641,N_6367,N_9284);
nand U12642 (N_12642,N_8175,N_9346);
nand U12643 (N_12643,N_3516,N_7705);
nand U12644 (N_12644,N_3860,N_1242);
xor U12645 (N_12645,N_1801,N_1296);
or U12646 (N_12646,N_7935,N_6257);
xor U12647 (N_12647,N_6620,N_5990);
or U12648 (N_12648,N_8488,N_3711);
nand U12649 (N_12649,N_4154,N_6445);
and U12650 (N_12650,N_9134,N_8837);
or U12651 (N_12651,N_9949,N_7643);
or U12652 (N_12652,N_6464,N_6944);
nor U12653 (N_12653,N_3629,N_9479);
and U12654 (N_12654,N_4260,N_235);
and U12655 (N_12655,N_6026,N_7031);
xor U12656 (N_12656,N_8184,N_7879);
nor U12657 (N_12657,N_2324,N_8666);
and U12658 (N_12658,N_2071,N_1455);
nor U12659 (N_12659,N_6060,N_2989);
and U12660 (N_12660,N_9775,N_3742);
nor U12661 (N_12661,N_9349,N_8290);
or U12662 (N_12662,N_955,N_6595);
nor U12663 (N_12663,N_1360,N_9548);
nand U12664 (N_12664,N_8789,N_925);
nand U12665 (N_12665,N_1417,N_6059);
xnor U12666 (N_12666,N_5334,N_7745);
and U12667 (N_12667,N_6006,N_1425);
xnor U12668 (N_12668,N_6767,N_5941);
or U12669 (N_12669,N_1464,N_9609);
nand U12670 (N_12670,N_9480,N_2231);
nand U12671 (N_12671,N_8557,N_3212);
nor U12672 (N_12672,N_5071,N_9580);
and U12673 (N_12673,N_6270,N_8950);
or U12674 (N_12674,N_8456,N_7690);
and U12675 (N_12675,N_3555,N_3334);
nand U12676 (N_12676,N_7239,N_8753);
nand U12677 (N_12677,N_9827,N_3693);
nand U12678 (N_12678,N_6888,N_4432);
nor U12679 (N_12679,N_1522,N_165);
xnor U12680 (N_12680,N_8786,N_3798);
xnor U12681 (N_12681,N_4147,N_8253);
nor U12682 (N_12682,N_3928,N_7346);
nand U12683 (N_12683,N_7871,N_9338);
or U12684 (N_12684,N_3260,N_3006);
and U12685 (N_12685,N_8561,N_6695);
nand U12686 (N_12686,N_390,N_9582);
and U12687 (N_12687,N_3916,N_9149);
or U12688 (N_12688,N_1085,N_5047);
and U12689 (N_12689,N_9994,N_9414);
or U12690 (N_12690,N_1700,N_7888);
xor U12691 (N_12691,N_5944,N_2068);
nand U12692 (N_12692,N_6998,N_1558);
and U12693 (N_12693,N_6494,N_8271);
nor U12694 (N_12694,N_7810,N_7132);
nand U12695 (N_12695,N_2223,N_4417);
nor U12696 (N_12696,N_2031,N_7834);
and U12697 (N_12697,N_8302,N_1709);
nor U12698 (N_12698,N_9668,N_6610);
or U12699 (N_12699,N_2534,N_5862);
nand U12700 (N_12700,N_4507,N_3892);
nor U12701 (N_12701,N_3182,N_6343);
or U12702 (N_12702,N_7966,N_3643);
nor U12703 (N_12703,N_2824,N_2105);
or U12704 (N_12704,N_6859,N_1673);
and U12705 (N_12705,N_7072,N_4575);
nand U12706 (N_12706,N_7087,N_588);
nor U12707 (N_12707,N_8222,N_8952);
and U12708 (N_12708,N_6643,N_9099);
nor U12709 (N_12709,N_9453,N_3466);
or U12710 (N_12710,N_6174,N_3701);
or U12711 (N_12711,N_9503,N_8101);
or U12712 (N_12712,N_7841,N_5865);
and U12713 (N_12713,N_9999,N_6438);
nor U12714 (N_12714,N_4632,N_5842);
and U12715 (N_12715,N_4522,N_90);
nand U12716 (N_12716,N_1632,N_8362);
nor U12717 (N_12717,N_1142,N_625);
or U12718 (N_12718,N_9209,N_3101);
xnor U12719 (N_12719,N_8128,N_8469);
nor U12720 (N_12720,N_5498,N_9724);
and U12721 (N_12721,N_5068,N_2662);
or U12722 (N_12722,N_1528,N_3198);
and U12723 (N_12723,N_4274,N_5356);
nor U12724 (N_12724,N_545,N_86);
nor U12725 (N_12725,N_8308,N_5158);
or U12726 (N_12726,N_5147,N_8967);
nand U12727 (N_12727,N_9690,N_9849);
and U12728 (N_12728,N_7475,N_7383);
xor U12729 (N_12729,N_8364,N_5984);
and U12730 (N_12730,N_6049,N_7579);
or U12731 (N_12731,N_1929,N_6607);
or U12732 (N_12732,N_9684,N_2222);
and U12733 (N_12733,N_6252,N_6305);
and U12734 (N_12734,N_5832,N_1412);
and U12735 (N_12735,N_2596,N_8813);
or U12736 (N_12736,N_8835,N_5916);
nor U12737 (N_12737,N_8814,N_2952);
nor U12738 (N_12738,N_2862,N_7864);
nand U12739 (N_12739,N_4506,N_2595);
nand U12740 (N_12740,N_7718,N_1181);
nand U12741 (N_12741,N_8141,N_191);
nor U12742 (N_12742,N_11,N_3330);
and U12743 (N_12743,N_1120,N_2703);
and U12744 (N_12744,N_3047,N_8020);
and U12745 (N_12745,N_6564,N_1652);
nor U12746 (N_12746,N_8052,N_2007);
nand U12747 (N_12747,N_3003,N_4590);
or U12748 (N_12748,N_6805,N_31);
nor U12749 (N_12749,N_2248,N_8398);
nor U12750 (N_12750,N_3385,N_9615);
or U12751 (N_12751,N_1215,N_5780);
and U12752 (N_12752,N_6585,N_5216);
xnor U12753 (N_12753,N_5644,N_3146);
nor U12754 (N_12754,N_7412,N_2394);
nand U12755 (N_12755,N_6719,N_7592);
or U12756 (N_12756,N_2809,N_4413);
and U12757 (N_12757,N_6670,N_3467);
or U12758 (N_12758,N_8094,N_2305);
or U12759 (N_12759,N_2357,N_9814);
nor U12760 (N_12760,N_9838,N_5117);
or U12761 (N_12761,N_4660,N_4908);
nor U12762 (N_12762,N_7295,N_5981);
xnor U12763 (N_12763,N_2060,N_2092);
nand U12764 (N_12764,N_9441,N_2385);
nor U12765 (N_12765,N_3960,N_2831);
nor U12766 (N_12766,N_8953,N_6599);
and U12767 (N_12767,N_3389,N_3945);
xor U12768 (N_12768,N_8016,N_2916);
nand U12769 (N_12769,N_4280,N_9125);
nor U12770 (N_12770,N_8357,N_9248);
and U12771 (N_12771,N_7371,N_8209);
and U12772 (N_12772,N_6164,N_4145);
xor U12773 (N_12773,N_6997,N_7219);
nor U12774 (N_12774,N_612,N_7134);
nand U12775 (N_12775,N_3344,N_2386);
xnor U12776 (N_12776,N_8098,N_5021);
xor U12777 (N_12777,N_9900,N_4365);
and U12778 (N_12778,N_4202,N_3956);
or U12779 (N_12779,N_6718,N_8661);
or U12780 (N_12780,N_4464,N_2676);
nor U12781 (N_12781,N_1109,N_3699);
or U12782 (N_12782,N_3138,N_4219);
or U12783 (N_12783,N_906,N_256);
nor U12784 (N_12784,N_8844,N_3922);
or U12785 (N_12785,N_6401,N_7969);
nor U12786 (N_12786,N_9976,N_4121);
nand U12787 (N_12787,N_5288,N_145);
or U12788 (N_12788,N_5118,N_8670);
or U12789 (N_12789,N_4676,N_5156);
or U12790 (N_12790,N_6029,N_3071);
or U12791 (N_12791,N_9329,N_4798);
or U12792 (N_12792,N_4623,N_3768);
or U12793 (N_12793,N_4231,N_6710);
xnor U12794 (N_12794,N_6715,N_4438);
or U12795 (N_12795,N_7458,N_816);
xnor U12796 (N_12796,N_6370,N_5594);
nor U12797 (N_12797,N_7777,N_4734);
and U12798 (N_12798,N_5267,N_7874);
and U12799 (N_12799,N_8738,N_1848);
nand U12800 (N_12800,N_9837,N_3525);
and U12801 (N_12801,N_7807,N_2328);
or U12802 (N_12802,N_8466,N_1714);
nand U12803 (N_12803,N_9681,N_5327);
and U12804 (N_12804,N_2699,N_3596);
nor U12805 (N_12805,N_9567,N_4583);
xnor U12806 (N_12806,N_8074,N_3040);
nor U12807 (N_12807,N_4697,N_3642);
or U12808 (N_12808,N_4895,N_2846);
nor U12809 (N_12809,N_8180,N_5319);
nand U12810 (N_12810,N_8735,N_7284);
or U12811 (N_12811,N_6749,N_7147);
nor U12812 (N_12812,N_3076,N_8346);
and U12813 (N_12813,N_3072,N_3667);
and U12814 (N_12814,N_1338,N_9820);
or U12815 (N_12815,N_7742,N_2322);
nand U12816 (N_12816,N_3611,N_9275);
and U12817 (N_12817,N_4708,N_6113);
and U12818 (N_12818,N_3886,N_186);
xor U12819 (N_12819,N_1948,N_5520);
or U12820 (N_12820,N_6148,N_7648);
nor U12821 (N_12821,N_2351,N_8521);
nor U12822 (N_12822,N_7401,N_2449);
or U12823 (N_12823,N_3835,N_8068);
or U12824 (N_12824,N_8039,N_375);
or U12825 (N_12825,N_1310,N_2130);
nand U12826 (N_12826,N_5904,N_9049);
nor U12827 (N_12827,N_1090,N_3627);
or U12828 (N_12828,N_3750,N_5442);
or U12829 (N_12829,N_8032,N_7632);
and U12830 (N_12830,N_242,N_3153);
or U12831 (N_12831,N_8120,N_4833);
and U12832 (N_12832,N_636,N_6335);
nand U12833 (N_12833,N_539,N_391);
and U12834 (N_12834,N_5933,N_3126);
and U12835 (N_12835,N_9459,N_9815);
xor U12836 (N_12836,N_9866,N_2793);
or U12837 (N_12837,N_9365,N_4678);
nand U12838 (N_12838,N_163,N_1032);
nor U12839 (N_12839,N_4834,N_6115);
and U12840 (N_12840,N_803,N_5351);
nor U12841 (N_12841,N_3135,N_5799);
or U12842 (N_12842,N_1047,N_1073);
or U12843 (N_12843,N_7277,N_8473);
nand U12844 (N_12844,N_8213,N_9986);
nand U12845 (N_12845,N_7312,N_3241);
nand U12846 (N_12846,N_3039,N_7207);
nand U12847 (N_12847,N_4686,N_7367);
or U12848 (N_12848,N_8438,N_1188);
nand U12849 (N_12849,N_8714,N_1477);
nor U12850 (N_12850,N_3340,N_829);
and U12851 (N_12851,N_4897,N_1856);
or U12852 (N_12852,N_9197,N_5849);
or U12853 (N_12853,N_5222,N_6989);
nor U12854 (N_12854,N_4756,N_3027);
nor U12855 (N_12855,N_2310,N_4684);
and U12856 (N_12856,N_124,N_6592);
or U12857 (N_12857,N_6238,N_558);
and U12858 (N_12858,N_8008,N_1083);
or U12859 (N_12859,N_9736,N_6386);
or U12860 (N_12860,N_812,N_3197);
nor U12861 (N_12861,N_3441,N_2089);
nand U12862 (N_12862,N_3282,N_1604);
or U12863 (N_12863,N_7735,N_272);
and U12864 (N_12864,N_3919,N_3469);
xnor U12865 (N_12865,N_1151,N_4562);
and U12866 (N_12866,N_6074,N_244);
and U12867 (N_12867,N_6116,N_4242);
nand U12868 (N_12868,N_7995,N_6940);
nand U12869 (N_12869,N_230,N_6862);
nand U12870 (N_12870,N_5067,N_7898);
nor U12871 (N_12871,N_4881,N_5042);
or U12872 (N_12872,N_1785,N_2788);
or U12873 (N_12873,N_6135,N_782);
nand U12874 (N_12874,N_873,N_2379);
nand U12875 (N_12875,N_2981,N_8891);
nor U12876 (N_12876,N_9416,N_7365);
and U12877 (N_12877,N_9018,N_8551);
nand U12878 (N_12878,N_4114,N_7150);
or U12879 (N_12879,N_2614,N_9431);
nand U12880 (N_12880,N_4052,N_4938);
nor U12881 (N_12881,N_3520,N_1465);
nor U12882 (N_12882,N_4519,N_6882);
and U12883 (N_12883,N_9844,N_7833);
nand U12884 (N_12884,N_7045,N_1326);
and U12885 (N_12885,N_8311,N_4263);
nor U12886 (N_12886,N_5144,N_5652);
nor U12887 (N_12887,N_6995,N_4799);
or U12888 (N_12888,N_1837,N_373);
or U12889 (N_12889,N_1950,N_7304);
or U12890 (N_12890,N_8203,N_7054);
nand U12891 (N_12891,N_9191,N_8694);
nor U12892 (N_12892,N_6709,N_4945);
nand U12893 (N_12893,N_2719,N_5924);
xnor U12894 (N_12894,N_8196,N_8543);
or U12895 (N_12895,N_6377,N_3483);
nor U12896 (N_12896,N_2155,N_7313);
and U12897 (N_12897,N_9785,N_9812);
nand U12898 (N_12898,N_4192,N_1195);
and U12899 (N_12899,N_6743,N_5258);
nand U12900 (N_12900,N_100,N_2647);
nor U12901 (N_12901,N_4220,N_2490);
and U12902 (N_12902,N_324,N_6959);
or U12903 (N_12903,N_5043,N_9281);
nor U12904 (N_12904,N_9592,N_3140);
nand U12905 (N_12905,N_6039,N_7517);
or U12906 (N_12906,N_8423,N_4327);
nor U12907 (N_12907,N_7529,N_2507);
nand U12908 (N_12908,N_5314,N_866);
nor U12909 (N_12909,N_4995,N_6107);
nor U12910 (N_12910,N_3251,N_1945);
nand U12911 (N_12911,N_4728,N_5134);
or U12912 (N_12912,N_1354,N_189);
and U12913 (N_12913,N_1185,N_1664);
nand U12914 (N_12914,N_9853,N_6911);
nand U12915 (N_12915,N_3488,N_8892);
nor U12916 (N_12916,N_7192,N_8591);
and U12917 (N_12917,N_7972,N_4361);
or U12918 (N_12918,N_7085,N_9855);
and U12919 (N_12919,N_5410,N_6930);
and U12920 (N_12920,N_7267,N_5395);
xor U12921 (N_12921,N_9654,N_2356);
nand U12922 (N_12922,N_903,N_5711);
or U12923 (N_12923,N_772,N_2088);
nor U12924 (N_12924,N_1949,N_410);
nand U12925 (N_12925,N_8231,N_9783);
nor U12926 (N_12926,N_7653,N_4254);
nor U12927 (N_12927,N_3592,N_6239);
xor U12928 (N_12928,N_9321,N_9578);
and U12929 (N_12929,N_7616,N_8158);
and U12930 (N_12930,N_6963,N_3559);
nand U12931 (N_12931,N_8594,N_7741);
nor U12932 (N_12932,N_2654,N_8480);
or U12933 (N_12933,N_2550,N_4795);
nor U12934 (N_12934,N_232,N_8256);
nor U12935 (N_12935,N_4119,N_2772);
nand U12936 (N_12936,N_844,N_3604);
xnor U12937 (N_12937,N_4658,N_9679);
xnor U12938 (N_12938,N_1021,N_1972);
and U12939 (N_12939,N_4310,N_660);
and U12940 (N_12940,N_1193,N_6508);
or U12941 (N_12941,N_4579,N_7611);
and U12942 (N_12942,N_8853,N_7800);
nor U12943 (N_12943,N_7453,N_1402);
nor U12944 (N_12944,N_8702,N_1069);
or U12945 (N_12945,N_5128,N_6958);
nand U12946 (N_12946,N_7061,N_4442);
and U12947 (N_12947,N_4852,N_5212);
nor U12948 (N_12948,N_2626,N_83);
and U12949 (N_12949,N_1431,N_2142);
xnor U12950 (N_12950,N_6302,N_3105);
nand U12951 (N_12951,N_1872,N_4051);
nor U12952 (N_12952,N_3563,N_7539);
or U12953 (N_12953,N_8155,N_6415);
nor U12954 (N_12954,N_3460,N_8794);
nor U12955 (N_12955,N_5177,N_9992);
and U12956 (N_12956,N_9625,N_1175);
nor U12957 (N_12957,N_4986,N_9739);
or U12958 (N_12958,N_4041,N_1717);
xor U12959 (N_12959,N_1058,N_2876);
nand U12960 (N_12960,N_6488,N_6657);
nor U12961 (N_12961,N_2132,N_265);
xnor U12962 (N_12962,N_4628,N_216);
or U12963 (N_12963,N_4535,N_8268);
and U12964 (N_12964,N_7604,N_4572);
nor U12965 (N_12965,N_6258,N_675);
nor U12966 (N_12966,N_9611,N_1008);
and U12967 (N_12967,N_7945,N_2741);
or U12968 (N_12968,N_1713,N_9418);
and U12969 (N_12969,N_5506,N_6601);
or U12970 (N_12970,N_3591,N_2516);
and U12971 (N_12971,N_3873,N_5126);
and U12972 (N_12972,N_1161,N_4141);
or U12973 (N_12973,N_8516,N_2612);
or U12974 (N_12974,N_5207,N_7819);
nor U12975 (N_12975,N_9624,N_1846);
nor U12976 (N_12976,N_6741,N_8911);
and U12977 (N_12977,N_213,N_4751);
nor U12978 (N_12978,N_1610,N_7562);
nor U12979 (N_12979,N_6861,N_4070);
nor U12980 (N_12980,N_5048,N_4324);
or U12981 (N_12981,N_633,N_6157);
xor U12982 (N_12982,N_61,N_5060);
and U12983 (N_12983,N_2592,N_6025);
xnor U12984 (N_12984,N_5026,N_7525);
and U12985 (N_12985,N_7208,N_6583);
and U12986 (N_12986,N_6289,N_6519);
nor U12987 (N_12987,N_3477,N_91);
nand U12988 (N_12988,N_4716,N_6506);
nor U12989 (N_12989,N_1358,N_9823);
or U12990 (N_12990,N_3780,N_7215);
nor U12991 (N_12991,N_3931,N_4983);
nor U12992 (N_12992,N_7438,N_333);
nand U12993 (N_12993,N_7586,N_8905);
nand U12994 (N_12994,N_6632,N_9118);
nand U12995 (N_12995,N_101,N_7086);
and U12996 (N_12996,N_1324,N_7185);
or U12997 (N_12997,N_6185,N_9033);
nand U12998 (N_12998,N_3731,N_2211);
and U12999 (N_12999,N_7605,N_4250);
nor U13000 (N_13000,N_5608,N_5752);
nor U13001 (N_13001,N_2768,N_8693);
or U13002 (N_13002,N_7666,N_280);
and U13003 (N_13003,N_1227,N_6145);
nand U13004 (N_13004,N_9876,N_8199);
nor U13005 (N_13005,N_6792,N_1733);
nor U13006 (N_13006,N_2139,N_7634);
or U13007 (N_13007,N_576,N_6811);
or U13008 (N_13008,N_1297,N_9017);
or U13009 (N_13009,N_3465,N_6108);
nor U13010 (N_13010,N_8276,N_3246);
xnor U13011 (N_13011,N_5992,N_1011);
or U13012 (N_13012,N_1740,N_9765);
xnor U13013 (N_13013,N_3691,N_5401);
or U13014 (N_13014,N_5704,N_2659);
xnor U13015 (N_13015,N_9829,N_745);
nor U13016 (N_13016,N_9674,N_8322);
and U13017 (N_13017,N_7366,N_4032);
nand U13018 (N_13018,N_2744,N_9003);
and U13019 (N_13019,N_5893,N_1975);
nor U13020 (N_13020,N_6300,N_5615);
nor U13021 (N_13021,N_7659,N_1004);
nand U13022 (N_13022,N_6110,N_7507);
xor U13023 (N_13023,N_6957,N_1369);
nand U13024 (N_13024,N_3672,N_8954);
xor U13025 (N_13025,N_4861,N_4770);
or U13026 (N_13026,N_3189,N_4527);
nand U13027 (N_13027,N_4182,N_4104);
and U13028 (N_13028,N_4306,N_5231);
xnor U13029 (N_13029,N_9816,N_9989);
and U13030 (N_13030,N_7720,N_5332);
or U13031 (N_13031,N_7676,N_6101);
nand U13032 (N_13032,N_3583,N_3369);
nand U13033 (N_13033,N_2414,N_3295);
nor U13034 (N_13034,N_4266,N_1966);
nor U13035 (N_13035,N_9915,N_2865);
or U13036 (N_13036,N_4228,N_3186);
nand U13037 (N_13037,N_3957,N_7146);
and U13038 (N_13038,N_7285,N_8583);
nand U13039 (N_13039,N_2513,N_3557);
nand U13040 (N_13040,N_1671,N_7251);
nor U13041 (N_13041,N_3253,N_2615);
nor U13042 (N_13042,N_1299,N_1189);
nor U13043 (N_13043,N_766,N_698);
or U13044 (N_13044,N_6208,N_2349);
nand U13045 (N_13045,N_5023,N_1828);
xnor U13046 (N_13046,N_4567,N_3442);
nand U13047 (N_13047,N_5224,N_9316);
xor U13048 (N_13048,N_5509,N_4393);
or U13049 (N_13049,N_8087,N_8598);
and U13050 (N_13050,N_3443,N_6560);
xnor U13051 (N_13051,N_1164,N_6615);
nor U13052 (N_13052,N_718,N_2454);
or U13053 (N_13053,N_2527,N_7557);
nor U13054 (N_13054,N_4283,N_2280);
nor U13055 (N_13055,N_2472,N_5748);
and U13056 (N_13056,N_6430,N_9353);
nor U13057 (N_13057,N_2056,N_5734);
nand U13058 (N_13058,N_1291,N_3437);
and U13059 (N_13059,N_4524,N_1601);
or U13060 (N_13060,N_1973,N_3317);
and U13061 (N_13061,N_4115,N_8144);
xor U13062 (N_13062,N_644,N_1278);
and U13063 (N_13063,N_4573,N_8073);
and U13064 (N_13064,N_4215,N_7272);
or U13065 (N_13065,N_6479,N_3953);
nand U13066 (N_13066,N_1018,N_9533);
or U13067 (N_13067,N_3124,N_7662);
nor U13068 (N_13068,N_7129,N_2220);
nor U13069 (N_13069,N_3486,N_7044);
nand U13070 (N_13070,N_2735,N_377);
nand U13071 (N_13071,N_7022,N_7546);
nor U13072 (N_13072,N_8834,N_9750);
or U13073 (N_13073,N_8606,N_2350);
or U13074 (N_13074,N_582,N_3058);
nor U13075 (N_13075,N_1545,N_5663);
nand U13076 (N_13076,N_7700,N_2152);
nand U13077 (N_13077,N_4172,N_975);
xor U13078 (N_13078,N_2145,N_6283);
nand U13079 (N_13079,N_8667,N_3284);
nor U13080 (N_13080,N_8581,N_744);
nor U13081 (N_13081,N_9934,N_1461);
and U13082 (N_13082,N_3227,N_2904);
or U13083 (N_13083,N_146,N_8378);
nand U13084 (N_13084,N_9833,N_7286);
and U13085 (N_13085,N_5112,N_9996);
or U13086 (N_13086,N_1256,N_8506);
nand U13087 (N_13087,N_8663,N_4409);
nor U13088 (N_13088,N_4060,N_1247);
nand U13089 (N_13089,N_6183,N_7817);
nand U13090 (N_13090,N_4894,N_2691);
nor U13091 (N_13091,N_846,N_8218);
or U13092 (N_13092,N_1984,N_7831);
nor U13093 (N_13093,N_1076,N_6756);
or U13094 (N_13094,N_2997,N_4443);
nor U13095 (N_13095,N_4496,N_8075);
nand U13096 (N_13096,N_856,N_3992);
nand U13097 (N_13097,N_1210,N_1135);
and U13098 (N_13098,N_9287,N_258);
or U13099 (N_13099,N_2011,N_755);
or U13100 (N_13100,N_7038,N_4599);
or U13101 (N_13101,N_1779,N_1176);
nand U13102 (N_13102,N_580,N_1869);
and U13103 (N_13103,N_5922,N_2870);
xor U13104 (N_13104,N_1716,N_8323);
nand U13105 (N_13105,N_7761,N_8427);
and U13106 (N_13106,N_5910,N_9648);
nand U13107 (N_13107,N_471,N_9602);
or U13108 (N_13108,N_6308,N_1298);
and U13109 (N_13109,N_3862,N_7492);
nand U13110 (N_13110,N_9534,N_6951);
nor U13111 (N_13111,N_4596,N_7245);
nor U13112 (N_13112,N_30,N_3721);
or U13113 (N_13113,N_9776,N_550);
nand U13114 (N_13114,N_3087,N_815);
nand U13115 (N_13115,N_9901,N_2757);
or U13116 (N_13116,N_3206,N_7727);
or U13117 (N_13117,N_6509,N_5628);
or U13118 (N_13118,N_3989,N_8139);
nor U13119 (N_13119,N_6385,N_4652);
nor U13120 (N_13120,N_3517,N_9835);
and U13121 (N_13121,N_2839,N_9515);
nand U13122 (N_13122,N_6791,N_2830);
nand U13123 (N_13123,N_238,N_6476);
and U13124 (N_13124,N_3827,N_752);
and U13125 (N_13125,N_4157,N_4790);
and U13126 (N_13126,N_1541,N_6517);
nand U13127 (N_13127,N_5772,N_3978);
nor U13128 (N_13128,N_6398,N_9687);
and U13129 (N_13129,N_8160,N_1650);
nor U13130 (N_13130,N_8665,N_5090);
xor U13131 (N_13131,N_3422,N_307);
and U13132 (N_13132,N_9028,N_1512);
and U13133 (N_13133,N_601,N_6033);
or U13134 (N_13134,N_8758,N_530);
and U13135 (N_13135,N_1077,N_8920);
or U13136 (N_13136,N_8482,N_8981);
or U13137 (N_13137,N_9361,N_8701);
or U13138 (N_13138,N_3288,N_248);
or U13139 (N_13139,N_4394,N_5751);
and U13140 (N_13140,N_6863,N_8773);
nand U13141 (N_13141,N_522,N_5323);
and U13142 (N_13142,N_2722,N_3474);
nand U13143 (N_13143,N_5002,N_9752);
and U13144 (N_13144,N_6442,N_3031);
nand U13145 (N_13145,N_5213,N_2810);
or U13146 (N_13146,N_1634,N_5363);
nand U13147 (N_13147,N_3943,N_5261);
and U13148 (N_13148,N_1050,N_2762);
xnor U13149 (N_13149,N_1373,N_1898);
xnor U13150 (N_13150,N_989,N_4109);
or U13151 (N_13151,N_5589,N_8933);
xor U13152 (N_13152,N_9351,N_2400);
nand U13153 (N_13153,N_7584,N_1274);
nand U13154 (N_13154,N_9139,N_4014);
nor U13155 (N_13155,N_1040,N_41);
nand U13156 (N_13156,N_7375,N_8721);
xor U13157 (N_13157,N_3537,N_8752);
nor U13158 (N_13158,N_4040,N_2506);
and U13159 (N_13159,N_9041,N_5622);
or U13160 (N_13160,N_3760,N_5161);
nor U13161 (N_13161,N_6925,N_9405);
nand U13162 (N_13162,N_7450,N_2783);
or U13163 (N_13163,N_2731,N_860);
xor U13164 (N_13164,N_1759,N_385);
xnor U13165 (N_13165,N_531,N_6889);
or U13166 (N_13166,N_6663,N_4901);
nand U13167 (N_13167,N_9335,N_7753);
nand U13168 (N_13168,N_9632,N_9764);
and U13169 (N_13169,N_2923,N_399);
nor U13170 (N_13170,N_6122,N_9494);
or U13171 (N_13171,N_6070,N_4905);
or U13172 (N_13172,N_2080,N_2236);
nand U13173 (N_13173,N_5239,N_5614);
nor U13174 (N_13174,N_2568,N_4218);
nor U13175 (N_13175,N_5070,N_8547);
and U13176 (N_13176,N_4774,N_9379);
and U13177 (N_13177,N_5800,N_2860);
and U13178 (N_13178,N_3511,N_1626);
nor U13179 (N_13179,N_7498,N_8664);
nor U13180 (N_13180,N_9891,N_3499);
and U13181 (N_13181,N_9293,N_1703);
nand U13182 (N_13182,N_4990,N_1959);
nor U13183 (N_13183,N_1919,N_9895);
or U13184 (N_13184,N_6673,N_9458);
and U13185 (N_13185,N_4466,N_5160);
nor U13186 (N_13186,N_136,N_1171);
nand U13187 (N_13187,N_2570,N_3723);
and U13188 (N_13188,N_9085,N_8);
and U13189 (N_13189,N_9377,N_7606);
xnor U13190 (N_13190,N_9857,N_2001);
nor U13191 (N_13191,N_463,N_967);
nor U13192 (N_13192,N_4740,N_2930);
nand U13193 (N_13193,N_2905,N_6962);
nor U13194 (N_13194,N_7121,N_1500);
or U13195 (N_13195,N_7590,N_8586);
and U13196 (N_13196,N_6867,N_4873);
and U13197 (N_13197,N_6827,N_7554);
nand U13198 (N_13198,N_9238,N_3727);
nand U13199 (N_13199,N_3964,N_6692);
or U13200 (N_13200,N_9094,N_6294);
and U13201 (N_13201,N_7963,N_3232);
and U13202 (N_13202,N_8698,N_9843);
nand U13203 (N_13203,N_3662,N_679);
nor U13204 (N_13204,N_2209,N_3579);
nor U13205 (N_13205,N_6414,N_999);
xnor U13206 (N_13206,N_543,N_5655);
nand U13207 (N_13207,N_7384,N_656);
and U13208 (N_13208,N_7237,N_3527);
and U13209 (N_13209,N_6967,N_6727);
or U13210 (N_13210,N_5746,N_7884);
and U13211 (N_13211,N_2954,N_9817);
nand U13212 (N_13212,N_3293,N_318);
xnor U13213 (N_13213,N_5523,N_7142);
nor U13214 (N_13214,N_4481,N_8305);
nand U13215 (N_13215,N_7929,N_7783);
nor U13216 (N_13216,N_5302,N_8886);
nand U13217 (N_13217,N_5982,N_2842);
nor U13218 (N_13218,N_593,N_7179);
and U13219 (N_13219,N_1678,N_5475);
nand U13220 (N_13220,N_5722,N_3281);
nor U13221 (N_13221,N_8811,N_8377);
nor U13222 (N_13222,N_5569,N_4078);
and U13223 (N_13223,N_1155,N_834);
and U13224 (N_13224,N_5046,N_3971);
and U13225 (N_13225,N_1235,N_927);
or U13226 (N_13226,N_9554,N_7581);
nand U13227 (N_13227,N_7564,N_8352);
nor U13228 (N_13228,N_4279,N_308);
nand U13229 (N_13229,N_2107,N_7496);
nand U13230 (N_13230,N_4826,N_3923);
and U13231 (N_13231,N_1920,N_58);
nand U13232 (N_13232,N_5491,N_3652);
xor U13233 (N_13233,N_2834,N_4143);
and U13234 (N_13234,N_3804,N_6373);
xnor U13235 (N_13235,N_9234,N_4613);
nand U13236 (N_13236,N_2421,N_2192);
nor U13237 (N_13237,N_5993,N_6922);
nand U13238 (N_13238,N_1320,N_2537);
and U13239 (N_13239,N_6918,N_1158);
nor U13240 (N_13240,N_6359,N_9898);
and U13241 (N_13241,N_668,N_3434);
or U13242 (N_13242,N_9467,N_6675);
nand U13243 (N_13243,N_2790,N_6316);
and U13244 (N_13244,N_4729,N_4605);
nor U13245 (N_13245,N_7271,N_417);
nor U13246 (N_13246,N_630,N_9906);
or U13247 (N_13247,N_654,N_8449);
or U13248 (N_13248,N_5923,N_4063);
or U13249 (N_13249,N_1573,N_8097);
or U13250 (N_13250,N_6410,N_9794);
nor U13251 (N_13251,N_1508,N_876);
or U13252 (N_13252,N_3942,N_5252);
nand U13253 (N_13253,N_9406,N_7333);
xnor U13254 (N_13254,N_3988,N_2163);
nand U13255 (N_13255,N_9552,N_9558);
nand U13256 (N_13256,N_3726,N_2638);
nor U13257 (N_13257,N_8888,N_2935);
and U13258 (N_13258,N_9603,N_5462);
and U13259 (N_13259,N_9847,N_7822);
xor U13260 (N_13260,N_6575,N_5761);
and U13261 (N_13261,N_1075,N_5716);
or U13262 (N_13262,N_6577,N_3576);
or U13263 (N_13263,N_7818,N_3633);
nor U13264 (N_13264,N_9435,N_9569);
or U13265 (N_13265,N_266,N_4042);
or U13266 (N_13266,N_731,N_2754);
nor U13267 (N_13267,N_6936,N_129);
or U13268 (N_13268,N_3007,N_8740);
xor U13269 (N_13269,N_6801,N_123);
and U13270 (N_13270,N_5833,N_335);
or U13271 (N_13271,N_2520,N_9930);
nand U13272 (N_13272,N_5103,N_6327);
nand U13273 (N_13273,N_3116,N_9374);
nand U13274 (N_13274,N_1029,N_6901);
and U13275 (N_13275,N_7088,N_1661);
and U13276 (N_13276,N_8291,N_4528);
nand U13277 (N_13277,N_3303,N_2943);
nand U13278 (N_13278,N_965,N_8384);
or U13279 (N_13279,N_3848,N_2673);
nand U13280 (N_13280,N_3628,N_2331);
and U13281 (N_13281,N_2496,N_5210);
and U13282 (N_13282,N_9774,N_9498);
and U13283 (N_13283,N_4787,N_6821);
nand U13284 (N_13284,N_5497,N_6354);
or U13285 (N_13285,N_6420,N_5487);
nor U13286 (N_13286,N_6700,N_871);
or U13287 (N_13287,N_4031,N_9317);
nor U13288 (N_13288,N_1340,N_4989);
nor U13289 (N_13289,N_1198,N_1336);
nand U13290 (N_13290,N_4874,N_7642);
and U13291 (N_13291,N_6434,N_6774);
or U13292 (N_13292,N_3739,N_2153);
nand U13293 (N_13293,N_676,N_7279);
and U13294 (N_13294,N_4354,N_7702);
nand U13295 (N_13295,N_7641,N_5032);
nand U13296 (N_13296,N_667,N_77);
nor U13297 (N_13297,N_1230,N_1777);
or U13298 (N_13298,N_488,N_8700);
and U13299 (N_13299,N_9371,N_7983);
xnor U13300 (N_13300,N_1691,N_3037);
nor U13301 (N_13301,N_4603,N_9700);
nor U13302 (N_13302,N_868,N_2911);
nand U13303 (N_13303,N_2293,N_9454);
nor U13304 (N_13304,N_5106,N_747);
and U13305 (N_13305,N_6181,N_5278);
nor U13306 (N_13306,N_8949,N_6550);
xor U13307 (N_13307,N_6761,N_95);
and U13308 (N_13308,N_0,N_6523);
nor U13309 (N_13309,N_2329,N_6057);
or U13310 (N_13310,N_5182,N_4450);
nand U13311 (N_13311,N_8915,N_9048);
nor U13312 (N_13312,N_3893,N_3735);
or U13313 (N_13313,N_3066,N_4867);
xor U13314 (N_13314,N_2872,N_5575);
xnor U13315 (N_13315,N_3128,N_1861);
nor U13316 (N_13316,N_5513,N_3818);
and U13317 (N_13317,N_912,N_1127);
or U13318 (N_13318,N_4928,N_260);
nand U13319 (N_13319,N_5127,N_6222);
nand U13320 (N_13320,N_6764,N_5775);
nand U13321 (N_13321,N_6439,N_8770);
nand U13322 (N_13322,N_281,N_1065);
nand U13323 (N_13323,N_3900,N_1237);
xnor U13324 (N_13324,N_7574,N_9461);
nor U13325 (N_13325,N_5353,N_8167);
and U13326 (N_13326,N_5883,N_6366);
or U13327 (N_13327,N_3159,N_2404);
xor U13328 (N_13328,N_584,N_8613);
nor U13329 (N_13329,N_6961,N_2897);
nor U13330 (N_13330,N_1756,N_7678);
nand U13331 (N_13331,N_4703,N_2306);
nor U13332 (N_13332,N_9385,N_9096);
xor U13333 (N_13333,N_9314,N_8899);
nand U13334 (N_13334,N_8605,N_2276);
nand U13335 (N_13335,N_8801,N_7856);
and U13336 (N_13336,N_452,N_8781);
and U13337 (N_13337,N_5599,N_1910);
nor U13338 (N_13338,N_4935,N_7973);
or U13339 (N_13339,N_1542,N_3310);
and U13340 (N_13340,N_386,N_2532);
xor U13341 (N_13341,N_4295,N_1451);
and U13342 (N_13342,N_5340,N_5010);
and U13343 (N_13343,N_7542,N_5307);
nand U13344 (N_13344,N_2214,N_2050);
and U13345 (N_13345,N_578,N_2271);
nand U13346 (N_13346,N_6593,N_7317);
nor U13347 (N_13347,N_4058,N_162);
nor U13348 (N_13348,N_5986,N_8717);
nand U13349 (N_13349,N_6205,N_5942);
or U13350 (N_13350,N_4759,N_3812);
nand U13351 (N_13351,N_4247,N_4910);
or U13352 (N_13352,N_6254,N_392);
nand U13353 (N_13353,N_7255,N_6131);
or U13354 (N_13354,N_6030,N_2388);
xnor U13355 (N_13355,N_1134,N_8531);
and U13356 (N_13356,N_4682,N_3985);
or U13357 (N_13357,N_5220,N_164);
or U13358 (N_13358,N_1944,N_2577);
nor U13359 (N_13359,N_7917,N_9168);
xnor U13360 (N_13360,N_9053,N_7357);
nand U13361 (N_13361,N_9252,N_3185);
nand U13362 (N_13362,N_3877,N_337);
xor U13363 (N_13363,N_1708,N_8063);
or U13364 (N_13364,N_8240,N_241);
nor U13365 (N_13365,N_8972,N_6696);
and U13366 (N_13366,N_7160,N_9868);
and U13367 (N_13367,N_8301,N_5362);
and U13368 (N_13368,N_7434,N_3342);
nor U13369 (N_13369,N_9487,N_8009);
xnor U13370 (N_13370,N_7392,N_9889);
nor U13371 (N_13371,N_34,N_4919);
nand U13372 (N_13372,N_6244,N_4234);
and U13373 (N_13373,N_9034,N_7205);
or U13374 (N_13374,N_4701,N_5342);
nor U13375 (N_13375,N_6199,N_3005);
nand U13376 (N_13376,N_650,N_5352);
or U13377 (N_13377,N_722,N_8930);
nand U13378 (N_13378,N_5793,N_4858);
nand U13379 (N_13379,N_5619,N_2315);
and U13380 (N_13380,N_9982,N_9240);
and U13381 (N_13381,N_7417,N_2863);
or U13382 (N_13382,N_9065,N_155);
nor U13383 (N_13383,N_1905,N_6152);
nand U13384 (N_13384,N_7620,N_914);
nand U13385 (N_13385,N_8568,N_1503);
or U13386 (N_13386,N_7480,N_8494);
or U13387 (N_13387,N_898,N_1276);
nor U13388 (N_13388,N_5566,N_1231);
xnor U13389 (N_13389,N_2924,N_8279);
and U13390 (N_13390,N_9790,N_5854);
or U13391 (N_13391,N_7430,N_7815);
and U13392 (N_13392,N_2750,N_4201);
nand U13393 (N_13393,N_1209,N_2342);
or U13394 (N_13394,N_9605,N_4285);
and U13395 (N_13395,N_904,N_8508);
nand U13396 (N_13396,N_2538,N_6100);
nand U13397 (N_13397,N_7209,N_932);
or U13398 (N_13398,N_4061,N_6881);
nor U13399 (N_13399,N_796,N_4079);
or U13400 (N_13400,N_7341,N_8860);
nand U13401 (N_13401,N_2019,N_9628);
xnor U13402 (N_13402,N_3188,N_9792);
or U13403 (N_13403,N_6798,N_6600);
nor U13404 (N_13404,N_5610,N_7711);
or U13405 (N_13405,N_7930,N_4576);
nor U13406 (N_13406,N_1800,N_7633);
nor U13407 (N_13407,N_1380,N_6264);
nor U13408 (N_13408,N_468,N_2137);
and U13409 (N_13409,N_9019,N_5617);
nand U13410 (N_13410,N_351,N_6569);
nand U13411 (N_13411,N_3705,N_4100);
nand U13412 (N_13412,N_3122,N_8200);
or U13413 (N_13413,N_7026,N_1205);
nor U13414 (N_13414,N_5408,N_6648);
nand U13415 (N_13415,N_5875,N_6261);
and U13416 (N_13416,N_7305,N_4648);
and U13417 (N_13417,N_9408,N_4021);
and U13418 (N_13418,N_4473,N_4407);
nor U13419 (N_13419,N_4554,N_5260);
nor U13420 (N_13420,N_8129,N_1988);
nand U13421 (N_13421,N_6642,N_9255);
xor U13422 (N_13422,N_6173,N_6443);
nor U13423 (N_13423,N_6237,N_109);
nor U13424 (N_13424,N_9061,N_16);
nor U13425 (N_13425,N_4083,N_3784);
nor U13426 (N_13426,N_6810,N_9542);
and U13427 (N_13427,N_8127,N_7560);
and U13428 (N_13428,N_3370,N_1849);
nand U13429 (N_13429,N_7640,N_7923);
nand U13430 (N_13430,N_4390,N_2409);
and U13431 (N_13431,N_7362,N_8329);
or U13432 (N_13432,N_8117,N_9652);
nand U13433 (N_13433,N_2641,N_1940);
and U13434 (N_13434,N_4288,N_5960);
nor U13435 (N_13435,N_1757,N_1982);
and U13436 (N_13436,N_9439,N_5496);
xnor U13437 (N_13437,N_6417,N_6845);
nand U13438 (N_13438,N_7979,N_1755);
nor U13439 (N_13439,N_6971,N_5691);
nand U13440 (N_13440,N_4974,N_3374);
nor U13441 (N_13441,N_7876,N_1888);
nor U13442 (N_13442,N_4742,N_7697);
or U13443 (N_13443,N_1548,N_3061);
and U13444 (N_13444,N_8681,N_2118);
nand U13445 (N_13445,N_2492,N_3895);
and U13446 (N_13446,N_5202,N_732);
and U13447 (N_13447,N_8856,N_2814);
nor U13448 (N_13448,N_7794,N_7390);
nand U13449 (N_13449,N_8145,N_2669);
nand U13450 (N_13450,N_5586,N_2165);
xor U13451 (N_13451,N_1313,N_3896);
or U13452 (N_13452,N_9223,N_3174);
and U13453 (N_13453,N_9845,N_560);
or U13454 (N_13454,N_9732,N_4453);
and U13455 (N_13455,N_4494,N_5310);
nor U13456 (N_13456,N_5694,N_5788);
nand U13457 (N_13457,N_1442,N_8134);
or U13458 (N_13458,N_7808,N_320);
or U13459 (N_13459,N_8455,N_6306);
nor U13460 (N_13460,N_3620,N_8862);
or U13461 (N_13461,N_2336,N_3973);
and U13462 (N_13462,N_6046,N_1786);
nor U13463 (N_13463,N_3091,N_3092);
nor U13464 (N_13464,N_1815,N_149);
xnor U13465 (N_13465,N_9473,N_9939);
or U13466 (N_13466,N_6361,N_7577);
and U13467 (N_13467,N_1566,N_2452);
xnor U13468 (N_13468,N_5777,N_2427);
nand U13469 (N_13469,N_790,N_5682);
nand U13470 (N_13470,N_5330,N_5120);
and U13471 (N_13471,N_1381,N_7156);
nor U13472 (N_13472,N_851,N_590);
and U13473 (N_13473,N_802,N_112);
nand U13474 (N_13474,N_5914,N_2493);
nor U13475 (N_13475,N_9673,N_6045);
and U13476 (N_13476,N_5512,N_8028);
nand U13477 (N_13477,N_3743,N_114);
xor U13478 (N_13478,N_6661,N_8332);
xnor U13479 (N_13479,N_5187,N_5804);
xor U13480 (N_13480,N_8697,N_9881);
nor U13481 (N_13481,N_4423,N_7241);
xor U13482 (N_13482,N_6067,N_6077);
nor U13483 (N_13483,N_9184,N_3190);
nand U13484 (N_13484,N_1051,N_9387);
or U13485 (N_13485,N_4357,N_1152);
nand U13486 (N_13486,N_8534,N_1042);
or U13487 (N_13487,N_5484,N_557);
nand U13488 (N_13488,N_7649,N_3899);
or U13489 (N_13489,N_8109,N_827);
or U13490 (N_13490,N_6787,N_5471);
nand U13491 (N_13491,N_1347,N_9694);
and U13492 (N_13492,N_9941,N_4836);
nor U13493 (N_13493,N_7947,N_2975);
or U13494 (N_13494,N_8784,N_9908);
nand U13495 (N_13495,N_1194,N_9126);
and U13496 (N_13496,N_5052,N_589);
nor U13497 (N_13497,N_7553,N_7360);
nor U13498 (N_13498,N_3913,N_5825);
and U13499 (N_13499,N_2705,N_3924);
xnor U13500 (N_13500,N_2004,N_1404);
nor U13501 (N_13501,N_4384,N_7407);
nand U13502 (N_13502,N_4723,N_5429);
and U13503 (N_13503,N_2038,N_483);
nor U13504 (N_13504,N_1637,N_7302);
or U13505 (N_13505,N_3601,N_8659);
nor U13506 (N_13506,N_6779,N_7269);
or U13507 (N_13507,N_6807,N_9005);
or U13508 (N_13508,N_4586,N_8440);
and U13509 (N_13509,N_3414,N_8507);
xnor U13510 (N_13510,N_6623,N_39);
nor U13511 (N_13511,N_227,N_4476);
or U13512 (N_13512,N_9661,N_1434);
or U13513 (N_13513,N_3640,N_3471);
or U13514 (N_13514,N_6796,N_4278);
and U13515 (N_13515,N_1534,N_677);
nand U13516 (N_13516,N_7975,N_4391);
and U13517 (N_13517,N_603,N_2680);
and U13518 (N_13518,N_3225,N_2913);
and U13519 (N_13519,N_8785,N_2569);
and U13520 (N_13520,N_5784,N_1649);
xnor U13521 (N_13521,N_6537,N_8567);
or U13522 (N_13522,N_1760,N_1537);
and U13523 (N_13523,N_5693,N_6347);
nand U13524 (N_13524,N_6561,N_2390);
and U13525 (N_13525,N_7624,N_5979);
nor U13526 (N_13526,N_5478,N_5446);
or U13527 (N_13527,N_1317,N_962);
nor U13528 (N_13528,N_4840,N_4381);
nor U13529 (N_13529,N_4126,N_7336);
xor U13530 (N_13530,N_570,N_1753);
and U13531 (N_13531,N_2657,N_4985);
or U13532 (N_13532,N_7903,N_5198);
xnor U13533 (N_13533,N_6646,N_1899);
or U13534 (N_13534,N_4982,N_1284);
xor U13535 (N_13535,N_1217,N_2672);
and U13536 (N_13536,N_5567,N_9852);
nor U13537 (N_13537,N_9195,N_2982);
nand U13538 (N_13538,N_1440,N_2797);
nand U13539 (N_13539,N_3656,N_7327);
nor U13540 (N_13540,N_5703,N_5850);
or U13541 (N_13541,N_2958,N_2111);
nand U13542 (N_13542,N_7321,N_1977);
and U13543 (N_13543,N_3586,N_57);
or U13544 (N_13544,N_8132,N_509);
nor U13545 (N_13545,N_4137,N_5191);
xnor U13546 (N_13546,N_2445,N_4015);
nand U13547 (N_13547,N_5754,N_2360);
nand U13548 (N_13548,N_5483,N_5929);
and U13549 (N_13549,N_6803,N_9922);
nor U13550 (N_13550,N_9678,N_5413);
nor U13551 (N_13551,N_1196,N_4124);
xor U13552 (N_13552,N_4166,N_2141);
nand U13553 (N_13553,N_1739,N_5237);
nor U13554 (N_13554,N_5824,N_8046);
nand U13555 (N_13555,N_6815,N_4733);
nand U13556 (N_13556,N_1366,N_4913);
nor U13557 (N_13557,N_3634,N_5296);
or U13558 (N_13558,N_3375,N_2627);
or U13559 (N_13559,N_3707,N_5931);
nand U13560 (N_13560,N_9311,N_8026);
nand U13561 (N_13561,N_4353,N_7235);
nor U13562 (N_13562,N_3170,N_2208);
nand U13563 (N_13563,N_9557,N_5669);
nand U13564 (N_13564,N_6137,N_8699);
nand U13565 (N_13565,N_5017,N_8836);
and U13566 (N_13566,N_1884,N_687);
nand U13567 (N_13567,N_24,N_3962);
nor U13568 (N_13568,N_2129,N_5488);
nand U13569 (N_13569,N_3963,N_9574);
xor U13570 (N_13570,N_2055,N_5461);
nor U13571 (N_13571,N_6752,N_3200);
nand U13572 (N_13572,N_4007,N_5405);
nand U13573 (N_13573,N_8919,N_4930);
nand U13574 (N_13574,N_1521,N_3937);
xnor U13575 (N_13575,N_3775,N_1308);
nand U13576 (N_13576,N_1818,N_708);
nand U13577 (N_13577,N_8550,N_9796);
nor U13578 (N_13578,N_9806,N_566);
nor U13579 (N_13579,N_9871,N_8288);
nand U13580 (N_13580,N_1141,N_596);
nor U13581 (N_13581,N_9214,N_794);
or U13582 (N_13582,N_5602,N_5726);
or U13583 (N_13583,N_3779,N_4125);
and U13584 (N_13584,N_921,N_4702);
or U13585 (N_13585,N_7565,N_3697);
or U13586 (N_13586,N_7724,N_1389);
and U13587 (N_13587,N_108,N_3120);
or U13588 (N_13588,N_3671,N_430);
nand U13589 (N_13589,N_8871,N_1183);
nor U13590 (N_13590,N_7144,N_5476);
and U13591 (N_13591,N_513,N_9352);
or U13592 (N_13592,N_301,N_1994);
nor U13593 (N_13593,N_1473,N_8719);
and U13594 (N_13594,N_8573,N_371);
and U13595 (N_13595,N_8044,N_1594);
and U13596 (N_13596,N_8210,N_913);
and U13597 (N_13597,N_5522,N_4);
nand U13598 (N_13598,N_2919,N_8450);
nand U13599 (N_13599,N_4175,N_8587);
nor U13600 (N_13600,N_2729,N_2574);
nand U13601 (N_13601,N_8562,N_749);
nor U13602 (N_13602,N_783,N_7343);
or U13603 (N_13603,N_3228,N_5373);
and U13604 (N_13604,N_1864,N_624);
nor U13605 (N_13605,N_6635,N_5061);
nand U13606 (N_13606,N_3098,N_1253);
and U13607 (N_13607,N_1809,N_3134);
nor U13608 (N_13608,N_4763,N_4849);
and U13609 (N_13609,N_5578,N_8400);
and U13610 (N_13610,N_762,N_1955);
and U13611 (N_13611,N_2369,N_8048);
and U13612 (N_13612,N_7820,N_8375);
or U13613 (N_13613,N_3565,N_2216);
and U13614 (N_13614,N_7070,N_2020);
nand U13615 (N_13615,N_1013,N_4629);
nor U13616 (N_13616,N_7534,N_3903);
or U13617 (N_13617,N_2984,N_7545);
xor U13618 (N_13618,N_7652,N_5105);
nor U13619 (N_13619,N_5372,N_455);
xor U13620 (N_13620,N_3948,N_1680);
nand U13621 (N_13621,N_8003,N_8195);
nor U13622 (N_13622,N_3560,N_9279);
nor U13623 (N_13623,N_3256,N_4619);
or U13624 (N_13624,N_1037,N_5809);
or U13625 (N_13625,N_5740,N_997);
nand U13626 (N_13626,N_2780,N_7670);
or U13627 (N_13627,N_1202,N_5805);
and U13628 (N_13628,N_3938,N_8416);
nor U13629 (N_13629,N_9903,N_1507);
nand U13630 (N_13630,N_3534,N_6587);
or U13631 (N_13631,N_5872,N_8999);
nor U13632 (N_13632,N_5695,N_8582);
nor U13633 (N_13633,N_6017,N_8190);
and U13634 (N_13634,N_7254,N_1787);
nand U13635 (N_13635,N_9147,N_7575);
and U13636 (N_13636,N_2475,N_8250);
nor U13637 (N_13637,N_743,N_296);
nand U13638 (N_13638,N_6451,N_2593);
xnor U13639 (N_13639,N_4877,N_4102);
nand U13640 (N_13640,N_3694,N_4049);
nand U13641 (N_13641,N_8445,N_3542);
and U13642 (N_13642,N_6742,N_1088);
nor U13643 (N_13643,N_5715,N_4208);
and U13644 (N_13644,N_2643,N_9564);
and U13645 (N_13645,N_9400,N_9320);
nand U13646 (N_13646,N_4609,N_1439);
nor U13647 (N_13647,N_4347,N_9056);
nor U13648 (N_13648,N_4345,N_546);
and U13649 (N_13649,N_5348,N_9875);
nor U13650 (N_13650,N_6947,N_4072);
xor U13651 (N_13651,N_9186,N_5538);
nand U13652 (N_13652,N_7859,N_7645);
xor U13653 (N_13653,N_1350,N_1646);
nand U13654 (N_13654,N_1057,N_426);
nor U13655 (N_13655,N_1589,N_8296);
or U13656 (N_13656,N_2423,N_2944);
nand U13657 (N_13657,N_9488,N_9004);
and U13658 (N_13658,N_4865,N_2771);
xor U13659 (N_13659,N_3032,N_3791);
and U13660 (N_13660,N_4065,N_8990);
nor U13661 (N_13661,N_542,N_9836);
or U13662 (N_13662,N_8980,N_7940);
and U13663 (N_13663,N_5948,N_1911);
and U13664 (N_13664,N_7602,N_1805);
xnor U13665 (N_13665,N_134,N_3811);
or U13666 (N_13666,N_695,N_3449);
or U13667 (N_13667,N_3304,N_2392);
nand U13668 (N_13668,N_1627,N_292);
or U13669 (N_13669,N_9052,N_4788);
and U13670 (N_13670,N_2936,N_378);
nand U13671 (N_13671,N_9517,N_8879);
or U13672 (N_13672,N_8084,N_9973);
or U13673 (N_13673,N_4637,N_4614);
nor U13674 (N_13674,N_9202,N_907);
and U13675 (N_13675,N_5211,N_6536);
or U13676 (N_13676,N_6880,N_3311);
xor U13677 (N_13677,N_1489,N_2463);
nor U13678 (N_13678,N_17,N_8965);
and U13679 (N_13679,N_5732,N_9324);
xor U13680 (N_13680,N_3456,N_404);
nor U13681 (N_13681,N_9204,N_4941);
nand U13682 (N_13682,N_9546,N_3846);
or U13683 (N_13683,N_7067,N_7883);
nand U13684 (N_13684,N_2425,N_2833);
and U13685 (N_13685,N_7270,N_8483);
and U13686 (N_13686,N_3594,N_2219);
nor U13687 (N_13687,N_8872,N_3856);
and U13688 (N_13688,N_5705,N_1981);
nor U13689 (N_13689,N_2732,N_8446);
nor U13690 (N_13690,N_2131,N_1871);
xnor U13691 (N_13691,N_2980,N_1179);
or U13692 (N_13692,N_706,N_7535);
nand U13693 (N_13693,N_2067,N_6379);
xor U13694 (N_13694,N_6019,N_2397);
xor U13695 (N_13695,N_2332,N_7679);
nor U13696 (N_13696,N_7369,N_1927);
nand U13697 (N_13697,N_1758,N_5081);
nand U13698 (N_13698,N_6800,N_6538);
nor U13699 (N_13699,N_5796,N_7213);
and U13700 (N_13700,N_628,N_5000);
and U13701 (N_13701,N_150,N_3646);
nor U13702 (N_13702,N_838,N_524);
and U13703 (N_13703,N_712,N_4449);
or U13704 (N_13704,N_7862,N_5897);
or U13705 (N_13705,N_2940,N_437);
and U13706 (N_13706,N_4196,N_7262);
or U13707 (N_13707,N_489,N_2134);
nor U13708 (N_13708,N_930,N_4964);
nand U13709 (N_13709,N_3014,N_9210);
and U13710 (N_13710,N_9655,N_2781);
nand U13711 (N_13711,N_2597,N_7043);
and U13712 (N_13712,N_3266,N_3229);
and U13713 (N_13713,N_8328,N_6857);
or U13714 (N_13714,N_9253,N_7555);
or U13715 (N_13715,N_2524,N_5503);
nand U13716 (N_13716,N_8182,N_9308);
or U13717 (N_13717,N_4452,N_4297);
or U13718 (N_13718,N_6172,N_5680);
or U13719 (N_13719,N_3876,N_5953);
xnor U13720 (N_13720,N_7173,N_2334);
xor U13721 (N_13721,N_3479,N_2373);
nor U13722 (N_13722,N_5173,N_9382);
xnor U13723 (N_13723,N_1426,N_8310);
or U13724 (N_13724,N_1232,N_5949);
nor U13725 (N_13725,N_2389,N_7291);
and U13726 (N_13726,N_212,N_5056);
nand U13727 (N_13727,N_7154,N_8490);
and U13728 (N_13728,N_6404,N_2618);
or U13729 (N_13729,N_1307,N_7353);
nand U13730 (N_13730,N_8479,N_5843);
and U13731 (N_13731,N_4017,N_5964);
xnor U13732 (N_13732,N_1098,N_841);
nand U13733 (N_13733,N_5552,N_8359);
nand U13734 (N_13734,N_1640,N_4497);
or U13735 (N_13735,N_2299,N_6403);
nor U13736 (N_13736,N_1621,N_2497);
nor U13737 (N_13737,N_4375,N_1474);
nor U13738 (N_13738,N_952,N_2590);
nor U13739 (N_13739,N_4252,N_125);
nor U13740 (N_13740,N_7729,N_954);
nand U13741 (N_13741,N_6188,N_4424);
or U13742 (N_13742,N_2150,N_1617);
and U13743 (N_13743,N_9354,N_6168);
nor U13744 (N_13744,N_5660,N_2199);
nand U13745 (N_13745,N_5295,N_1490);
and U13746 (N_13746,N_5080,N_1239);
nand U13747 (N_13747,N_7767,N_5776);
nand U13748 (N_13748,N_6096,N_8805);
xnor U13749 (N_13749,N_3030,N_987);
or U13750 (N_13750,N_127,N_2133);
or U13751 (N_13751,N_8923,N_1138);
and U13752 (N_13752,N_7198,N_5859);
xor U13753 (N_13753,N_6339,N_2775);
and U13754 (N_13754,N_1867,N_7928);
nand U13755 (N_13755,N_7920,N_1361);
and U13756 (N_13756,N_1830,N_2918);
or U13757 (N_13757,N_401,N_608);
and U13758 (N_13758,N_4828,N_5240);
nor U13759 (N_13759,N_2634,N_3372);
nor U13760 (N_13760,N_986,N_7364);
nand U13761 (N_13761,N_2987,N_4067);
nand U13762 (N_13762,N_4816,N_3451);
nor U13763 (N_13763,N_3089,N_9575);
and U13764 (N_13764,N_4871,N_8629);
and U13765 (N_13765,N_1715,N_2374);
and U13766 (N_13766,N_5969,N_5113);
nand U13767 (N_13767,N_2753,N_5242);
or U13768 (N_13768,N_4766,N_7775);
nand U13769 (N_13769,N_7855,N_4842);
and U13770 (N_13770,N_4368,N_4333);
or U13771 (N_13771,N_2307,N_7200);
and U13772 (N_13772,N_5515,N_6904);
nand U13773 (N_13773,N_2156,N_8412);
or U13774 (N_13774,N_4459,N_7467);
or U13775 (N_13775,N_8092,N_5882);
nand U13776 (N_13776,N_2606,N_6390);
or U13777 (N_13777,N_651,N_3421);
xnor U13778 (N_13778,N_5289,N_8076);
nor U13779 (N_13779,N_9916,N_3669);
xor U13780 (N_13780,N_2405,N_5521);
and U13781 (N_13781,N_6984,N_2025);
xor U13782 (N_13782,N_2578,N_5921);
and U13783 (N_13783,N_7759,N_6572);
nor U13784 (N_13784,N_3631,N_4366);
nor U13785 (N_13785,N_5349,N_1748);
nor U13786 (N_13786,N_4997,N_7314);
nand U13787 (N_13787,N_8596,N_8054);
nand U13788 (N_13788,N_7943,N_5146);
nand U13789 (N_13789,N_2713,N_5286);
xnor U13790 (N_13790,N_1228,N_9016);
nand U13791 (N_13791,N_2663,N_5646);
or U13792 (N_13792,N_7330,N_3704);
or U13793 (N_13793,N_8632,N_890);
or U13794 (N_13794,N_1087,N_3536);
nand U13795 (N_13795,N_1644,N_1452);
or U13796 (N_13796,N_1799,N_6389);
and U13797 (N_13797,N_896,N_5097);
nand U13798 (N_13798,N_6405,N_2739);
nand U13799 (N_13799,N_2877,N_6548);
nor U13800 (N_13800,N_3545,N_9012);
or U13801 (N_13801,N_8126,N_6263);
nor U13802 (N_13802,N_5,N_5852);
or U13803 (N_13803,N_7062,N_2090);
nand U13804 (N_13804,N_9788,N_7701);
or U13805 (N_13805,N_7901,N_8245);
and U13806 (N_13806,N_4954,N_552);
or U13807 (N_13807,N_4122,N_5292);
nand U13808 (N_13808,N_8780,N_51);
or U13809 (N_13809,N_2851,N_8890);
or U13810 (N_13810,N_3208,N_3240);
nor U13811 (N_13811,N_9075,N_5339);
and U13812 (N_13812,N_1520,N_4633);
and U13813 (N_13813,N_8303,N_218);
and U13814 (N_13814,N_6493,N_1841);
nor U13815 (N_13815,N_8205,N_6783);
nor U13816 (N_13816,N_6994,N_3351);
or U13817 (N_13817,N_8173,N_4662);
nand U13818 (N_13818,N_821,N_6618);
or U13819 (N_13819,N_4725,N_4448);
nor U13820 (N_13820,N_4150,N_2661);
nor U13821 (N_13821,N_3386,N_12);
and U13822 (N_13822,N_8399,N_4704);
nand U13823 (N_13823,N_6221,N_5786);
nand U13824 (N_13824,N_8255,N_4305);
nand U13825 (N_13825,N_2563,N_220);
xnor U13826 (N_13826,N_8166,N_8265);
nand U13827 (N_13827,N_2518,N_9339);
nor U13828 (N_13828,N_6892,N_9388);
and U13829 (N_13829,N_2341,N_3415);
or U13830 (N_13830,N_6605,N_6907);
nor U13831 (N_13831,N_1655,N_4068);
or U13832 (N_13832,N_6334,N_14);
nor U13833 (N_13833,N_1710,N_640);
and U13834 (N_13834,N_3526,N_1712);
nor U13835 (N_13835,N_7829,N_6013);
and U13836 (N_13836,N_5381,N_9256);
or U13837 (N_13837,N_4239,N_2837);
or U13838 (N_13838,N_8716,N_808);
nand U13839 (N_13839,N_5725,N_8241);
xnor U13840 (N_13840,N_7896,N_1218);
nand U13841 (N_13841,N_1983,N_517);
and U13842 (N_13842,N_478,N_1693);
or U13843 (N_13843,N_9124,N_2963);
or U13844 (N_13844,N_9258,N_4155);
or U13845 (N_13845,N_528,N_7293);
nor U13846 (N_13846,N_6065,N_1169);
and U13847 (N_13847,N_6114,N_1595);
nand U13848 (N_13848,N_5621,N_7210);
xor U13849 (N_13849,N_1304,N_5911);
nand U13850 (N_13850,N_9063,N_2);
nand U13851 (N_13851,N_2892,N_573);
or U13852 (N_13852,N_1737,N_5887);
nor U13853 (N_13853,N_7052,N_6002);
or U13854 (N_13854,N_3933,N_1184);
nor U13855 (N_13855,N_9664,N_3223);
and U13856 (N_13856,N_6295,N_8376);
or U13857 (N_13857,N_3728,N_3060);
or U13858 (N_13858,N_4463,N_6658);
or U13859 (N_13859,N_1892,N_5603);
or U13860 (N_13860,N_4963,N_8121);
nand U13861 (N_13861,N_4363,N_1850);
nand U13862 (N_13862,N_2914,N_305);
or U13863 (N_13863,N_6604,N_4209);
nand U13864 (N_13864,N_4302,N_9037);
xor U13865 (N_13865,N_2633,N_6843);
nor U13866 (N_13866,N_7328,N_5811);
or U13867 (N_13867,N_4862,N_2932);
nor U13868 (N_13868,N_1751,N_7893);
nor U13869 (N_13869,N_7536,N_6211);
and U13870 (N_13870,N_7601,N_7189);
xor U13871 (N_13871,N_5749,N_6016);
or U13872 (N_13872,N_5227,N_7395);
xor U13873 (N_13873,N_1105,N_4909);
xor U13874 (N_13874,N_2451,N_8395);
and U13875 (N_13875,N_2859,N_7717);
nor U13876 (N_13876,N_7226,N_5396);
or U13877 (N_13877,N_6707,N_3655);
and U13878 (N_13878,N_198,N_3169);
xnor U13879 (N_13879,N_3399,N_2660);
or U13880 (N_13880,N_6372,N_9450);
nand U13881 (N_13881,N_1089,N_8723);
nand U13882 (N_13882,N_1600,N_5611);
or U13883 (N_13883,N_1220,N_7769);
nand U13884 (N_13884,N_9536,N_2053);
nor U13885 (N_13885,N_7406,N_3507);
nand U13886 (N_13886,N_2632,N_569);
xnor U13887 (N_13887,N_6126,N_2256);
or U13888 (N_13888,N_5368,N_221);
xor U13889 (N_13889,N_1117,N_4814);
nor U13890 (N_13890,N_4851,N_3762);
nor U13891 (N_13891,N_6048,N_572);
and U13892 (N_13892,N_9910,N_7911);
nor U13893 (N_13893,N_9151,N_3099);
or U13894 (N_13894,N_7301,N_9508);
or U13895 (N_13895,N_195,N_8996);
nand U13896 (N_13896,N_3575,N_9420);
or U13897 (N_13897,N_4796,N_119);
and U13898 (N_13898,N_9220,N_4403);
or U13899 (N_13899,N_2026,N_8498);
and U13900 (N_13900,N_919,N_7890);
xnor U13901 (N_13901,N_8601,N_1033);
and U13902 (N_13902,N_7959,N_6313);
nor U13903 (N_13903,N_4446,N_2937);
and U13904 (N_13904,N_4943,N_4171);
and U13905 (N_13905,N_776,N_2483);
or U13906 (N_13906,N_6852,N_2942);
or U13907 (N_13907,N_9203,N_1688);
nand U13908 (N_13908,N_9928,N_1764);
nor U13909 (N_13909,N_436,N_1156);
and U13910 (N_13910,N_7136,N_2301);
xnor U13911 (N_13911,N_2027,N_9367);
nand U13912 (N_13912,N_1505,N_8556);
or U13913 (N_13913,N_7197,N_1509);
and U13914 (N_13914,N_1793,N_6799);
nor U13915 (N_13915,N_6357,N_4003);
nor U13916 (N_13916,N_8090,N_8078);
and U13917 (N_13917,N_3546,N_8624);
nor U13918 (N_13918,N_3462,N_1376);
nand U13919 (N_13919,N_2920,N_204);
nor U13920 (N_13920,N_9299,N_1665);
or U13921 (N_13921,N_5674,N_1903);
nor U13922 (N_13922,N_2052,N_6112);
nor U13923 (N_13923,N_144,N_1443);
or U13924 (N_13924,N_4444,N_8237);
nor U13925 (N_13925,N_239,N_9430);
xor U13926 (N_13926,N_2855,N_8070);
or U13927 (N_13927,N_154,N_7865);
xor U13928 (N_13928,N_3621,N_4780);
xnor U13929 (N_13929,N_1741,N_6050);
nand U13930 (N_13930,N_4057,N_739);
nor U13931 (N_13931,N_5093,N_3413);
nor U13932 (N_13932,N_6215,N_3215);
and U13933 (N_13933,N_770,N_9108);
nand U13934 (N_13934,N_7172,N_9516);
nand U13935 (N_13935,N_482,N_7400);
xnor U13936 (N_13936,N_6491,N_5836);
nor U13937 (N_13937,N_7428,N_7743);
or U13938 (N_13938,N_1487,N_8576);
and U13939 (N_13939,N_8497,N_8875);
and U13940 (N_13940,N_602,N_5013);
or U13941 (N_13941,N_3967,N_6036);
and U13942 (N_13942,N_7849,N_813);
nor U13943 (N_13943,N_5604,N_3472);
xor U13944 (N_13944,N_7956,N_9170);
nand U13945 (N_13945,N_4883,N_4879);
and U13946 (N_13946,N_4638,N_1620);
nor U13947 (N_13947,N_3959,N_7791);
or U13948 (N_13948,N_2353,N_7083);
nand U13949 (N_13949,N_5528,N_7300);
nor U13950 (N_13950,N_1328,N_3708);
or U13951 (N_13951,N_6650,N_2012);
xnor U13952 (N_13952,N_4570,N_2552);
nor U13953 (N_13953,N_3802,N_2167);
nor U13954 (N_13954,N_7064,N_5847);
nor U13955 (N_13955,N_5035,N_7582);
and U13956 (N_13956,N_3894,N_6596);
and U13957 (N_13957,N_2708,N_9199);
and U13958 (N_13958,N_313,N_5050);
nand U13959 (N_13959,N_8295,N_781);
and U13960 (N_13960,N_3029,N_1679);
or U13961 (N_13961,N_6554,N_4584);
xor U13962 (N_13962,N_6472,N_7674);
or U13963 (N_13963,N_1802,N_7740);
nor U13964 (N_13964,N_7029,N_3807);
nand U13965 (N_13965,N_8509,N_972);
or U13966 (N_13966,N_6007,N_4048);
or U13967 (N_13967,N_5255,N_6353);
and U13968 (N_13968,N_8056,N_2281);
and U13969 (N_13969,N_8607,N_4214);
nand U13970 (N_13970,N_4835,N_2993);
and U13971 (N_13971,N_9904,N_9540);
nand U13972 (N_13972,N_2355,N_4722);
and U13973 (N_13973,N_3045,N_6249);
nand U13974 (N_13974,N_5741,N_7821);
and U13975 (N_13975,N_7644,N_2808);
xnor U13976 (N_13976,N_4561,N_4656);
and U13977 (N_13977,N_1752,N_264);
nor U13978 (N_13978,N_3584,N_9589);
and U13979 (N_13979,N_9931,N_228);
and U13980 (N_13980,N_1895,N_5107);
and U13981 (N_13981,N_2173,N_6287);
and U13982 (N_13982,N_1149,N_1110);
nand U13983 (N_13983,N_4737,N_6499);
or U13984 (N_13984,N_9977,N_4329);
or U13985 (N_13985,N_2478,N_4335);
xor U13986 (N_13986,N_6014,N_9062);
nand U13987 (N_13987,N_8986,N_2769);
nor U13988 (N_13988,N_6966,N_5455);
xnor U13989 (N_13989,N_450,N_2003);
or U13990 (N_13990,N_5089,N_6073);
and U13991 (N_13991,N_7063,N_9740);
nor U13992 (N_13992,N_8131,N_6187);
nor U13993 (N_13993,N_7247,N_4349);
and U13994 (N_13994,N_3998,N_9526);
nor U13995 (N_13995,N_1385,N_6522);
and U13996 (N_13996,N_4695,N_6382);
nand U13997 (N_13997,N_3000,N_9947);
nand U13998 (N_13998,N_9556,N_6571);
nand U13999 (N_13999,N_6983,N_7221);
nand U14000 (N_14000,N_6597,N_9130);
nand U14001 (N_14001,N_5322,N_5818);
nand U14002 (N_14002,N_2230,N_2874);
nand U14003 (N_14003,N_6224,N_6916);
and U14004 (N_14004,N_8628,N_9489);
nor U14005 (N_14005,N_79,N_6729);
or U14006 (N_14006,N_9249,N_5545);
or U14007 (N_14007,N_8800,N_8402);
and U14008 (N_14008,N_4922,N_9560);
xor U14009 (N_14009,N_466,N_1878);
or U14010 (N_14010,N_8861,N_464);
nor U14011 (N_14011,N_2474,N_5525);
or U14012 (N_14012,N_8705,N_6854);
and U14013 (N_14013,N_5245,N_2678);
and U14014 (N_14014,N_2951,N_4055);
and U14015 (N_14015,N_2032,N_6996);
nand U14016 (N_14016,N_7232,N_5409);
or U14017 (N_14017,N_9038,N_7637);
or U14018 (N_14018,N_6498,N_3418);
nand U14019 (N_14019,N_4977,N_3810);
and U14020 (N_14020,N_3004,N_2557);
or U14021 (N_14021,N_3815,N_1890);
and U14022 (N_14022,N_1166,N_7948);
and U14023 (N_14023,N_2240,N_6151);
xnor U14024 (N_14024,N_7244,N_7638);
xnor U14025 (N_14025,N_9970,N_7174);
nand U14026 (N_14026,N_5325,N_507);
and U14027 (N_14027,N_9026,N_8648);
and U14028 (N_14028,N_6769,N_4035);
nand U14029 (N_14029,N_8062,N_6146);
and U14030 (N_14030,N_7513,N_4301);
nor U14031 (N_14031,N_3658,N_7907);
or U14032 (N_14032,N_7830,N_1502);
nor U14033 (N_14033,N_5900,N_190);
and U14034 (N_14034,N_8845,N_3522);
or U14035 (N_14035,N_7493,N_294);
nor U14036 (N_14036,N_9176,N_67);
and U14037 (N_14037,N_2101,N_3022);
xnor U14038 (N_14038,N_9887,N_3712);
nor U14039 (N_14039,N_5336,N_5432);
nor U14040 (N_14040,N_825,N_420);
or U14041 (N_14041,N_5531,N_2233);
nand U14042 (N_14042,N_8246,N_5038);
xnor U14043 (N_14043,N_7288,N_9995);
or U14044 (N_14044,N_7552,N_7675);
nor U14045 (N_14045,N_8558,N_3346);
xnor U14046 (N_14046,N_6293,N_832);
xor U14047 (N_14047,N_7131,N_8130);
or U14048 (N_14048,N_6391,N_8914);
nand U14049 (N_14049,N_6228,N_4184);
nor U14050 (N_14050,N_7399,N_8037);
xnor U14051 (N_14051,N_4268,N_1834);
nor U14052 (N_14052,N_1421,N_7723);
nor U14053 (N_14053,N_3110,N_3566);
or U14054 (N_14054,N_2985,N_2164);
or U14055 (N_14055,N_1575,N_9021);
nor U14056 (N_14056,N_1891,N_56);
nand U14057 (N_14057,N_6128,N_1332);
and U14058 (N_14058,N_4267,N_8928);
nor U14059 (N_14059,N_4482,N_5139);
xnor U14060 (N_14060,N_9117,N_1701);
xor U14061 (N_14061,N_6530,N_8821);
nor U14062 (N_14062,N_5907,N_4839);
nor U14063 (N_14063,N_4313,N_4866);
nand U14064 (N_14064,N_6094,N_3869);
or U14065 (N_14065,N_4942,N_4612);
nor U14066 (N_14066,N_4081,N_9943);
and U14067 (N_14067,N_1609,N_6170);
or U14068 (N_14068,N_6501,N_5756);
nand U14069 (N_14069,N_5570,N_7765);
or U14070 (N_14070,N_5573,N_5194);
and U14071 (N_14071,N_8580,N_3306);
nand U14072 (N_14072,N_6027,N_346);
or U14073 (N_14073,N_140,N_3192);
and U14074 (N_14074,N_289,N_1356);
nand U14075 (N_14075,N_6018,N_5492);
nor U14076 (N_14076,N_3554,N_5828);
nor U14077 (N_14077,N_4831,N_6332);
nand U14078 (N_14078,N_7009,N_1964);
or U14079 (N_14079,N_1868,N_8071);
and U14080 (N_14080,N_6868,N_5069);
and U14081 (N_14081,N_9007,N_8863);
nand U14082 (N_14082,N_7246,N_2600);
nor U14083 (N_14083,N_1045,N_362);
or U14084 (N_14084,N_1663,N_5360);
or U14085 (N_14085,N_3698,N_8609);
and U14086 (N_14086,N_6156,N_9626);
nand U14087 (N_14087,N_3996,N_5892);
nor U14088 (N_14088,N_7805,N_3133);
and U14089 (N_14089,N_759,N_166);
and U14090 (N_14090,N_9882,N_6169);
and U14091 (N_14091,N_8684,N_6459);
and U14092 (N_14092,N_5930,N_1056);
and U14093 (N_14093,N_6576,N_5086);
nor U14094 (N_14094,N_3264,N_3141);
nor U14095 (N_14095,N_3426,N_2459);
and U14096 (N_14096,N_2583,N_5977);
or U14097 (N_14097,N_5518,N_7010);
nor U14098 (N_14098,N_6905,N_3736);
and U14099 (N_14099,N_342,N_7814);
nand U14100 (N_14100,N_2195,N_9964);
nor U14101 (N_14101,N_4082,N_7373);
nor U14102 (N_14102,N_877,N_5221);
and U14103 (N_14103,N_1598,N_6581);
xor U14104 (N_14104,N_6371,N_354);
nor U14105 (N_14105,N_6066,N_5585);
nor U14106 (N_14106,N_2157,N_6900);
nor U14107 (N_14107,N_9079,N_9572);
nor U14108 (N_14108,N_1302,N_3384);
and U14109 (N_14109,N_6512,N_2072);
nor U14110 (N_14110,N_5819,N_6991);
nand U14111 (N_14111,N_4726,N_9309);
and U14112 (N_14112,N_9599,N_5045);
nor U14113 (N_14113,N_8163,N_4657);
nand U14114 (N_14114,N_1803,N_5233);
nor U14115 (N_14115,N_6041,N_3958);
or U14116 (N_14116,N_3079,N_7449);
and U14117 (N_14117,N_446,N_897);
nand U14118 (N_14118,N_3269,N_8387);
or U14119 (N_14119,N_5510,N_9809);
and U14120 (N_14120,N_3675,N_8977);
xnor U14121 (N_14121,N_2995,N_9270);
nor U14122 (N_14122,N_1456,N_219);
nor U14123 (N_14123,N_5869,N_2619);
xnor U14124 (N_14124,N_619,N_331);
nand U14125 (N_14125,N_2721,N_4112);
or U14126 (N_14126,N_2927,N_4688);
nor U14127 (N_14127,N_7778,N_8294);
or U14128 (N_14128,N_2184,N_1941);
nand U14129 (N_14129,N_7282,N_5877);
and U14130 (N_14130,N_8259,N_7722);
nor U14131 (N_14131,N_2123,N_942);
nand U14132 (N_14132,N_4724,N_623);
and U14133 (N_14133,N_6481,N_8642);
nand U14134 (N_14134,N_773,N_6594);
or U14135 (N_14135,N_4235,N_486);
or U14136 (N_14136,N_3,N_4428);
or U14137 (N_14137,N_3570,N_5920);
nor U14138 (N_14138,N_2378,N_3505);
and U14139 (N_14139,N_9471,N_674);
and U14140 (N_14140,N_9192,N_886);
nor U14141 (N_14141,N_7212,N_7206);
nand U14142 (N_14142,N_3891,N_5903);
nor U14143 (N_14143,N_6478,N_4944);
nor U14144 (N_14144,N_1532,N_9332);
nor U14145 (N_14145,N_159,N_2800);
and U14146 (N_14146,N_6778,N_6082);
xor U14147 (N_14147,N_6340,N_7688);
nand U14148 (N_14148,N_374,N_8467);
and U14149 (N_14149,N_3291,N_3315);
nor U14150 (N_14150,N_5737,N_8641);
and U14151 (N_14151,N_3064,N_1991);
or U14152 (N_14152,N_8743,N_9159);
nand U14153 (N_14153,N_9464,N_4543);
and U14154 (N_14154,N_6737,N_1154);
and U14155 (N_14155,N_6968,N_6383);
and U14156 (N_14156,N_3993,N_5148);
nand U14157 (N_14157,N_60,N_3994);
nor U14158 (N_14158,N_8791,N_8043);
and U14159 (N_14159,N_6674,N_9064);
nor U14160 (N_14160,N_1009,N_4398);
nor U14161 (N_14161,N_8333,N_7363);
or U14162 (N_14162,N_5228,N_6409);
nor U14163 (N_14163,N_6754,N_46);
and U14164 (N_14164,N_1789,N_2264);
nand U14165 (N_14165,N_1986,N_6477);
nor U14166 (N_14166,N_2084,N_3320);
nand U14167 (N_14167,N_4385,N_6970);
nor U14168 (N_14168,N_5816,N_1200);
and U14169 (N_14169,N_8512,N_5831);
xor U14170 (N_14170,N_105,N_6504);
nor U14171 (N_14171,N_1321,N_8864);
nand U14172 (N_14172,N_5577,N_8926);
or U14173 (N_14173,N_4321,N_2588);
nand U14174 (N_14174,N_4781,N_2649);
or U14175 (N_14175,N_4270,N_631);
and U14176 (N_14176,N_7997,N_5908);
xnor U14177 (N_14177,N_7921,N_247);
or U14178 (N_14178,N_541,N_6251);
nand U14179 (N_14179,N_259,N_2037);
xnor U14180 (N_14180,N_6337,N_7268);
or U14181 (N_14181,N_8365,N_5472);
nor U14182 (N_14182,N_5612,N_4745);
nand U14183 (N_14183,N_3012,N_2716);
or U14184 (N_14184,N_885,N_3617);
or U14185 (N_14185,N_3863,N_6505);
nand U14186 (N_14186,N_9998,N_5988);
and U14187 (N_14187,N_9958,N_663);
or U14188 (N_14188,N_2023,N_9205);
nor U14189 (N_14189,N_7708,N_4563);
nor U14190 (N_14190,N_5040,N_8391);
nor U14191 (N_14191,N_5848,N_1747);
and U14192 (N_14192,N_6450,N_1223);
nor U14193 (N_14193,N_5434,N_250);
nand U14194 (N_14194,N_4224,N_4287);
nand U14195 (N_14195,N_7457,N_1319);
and U14196 (N_14196,N_4360,N_3409);
or U14197 (N_14197,N_3651,N_5666);
or U14198 (N_14198,N_7617,N_2567);
nand U14199 (N_14199,N_9555,N_8021);
xnor U14200 (N_14200,N_8912,N_2671);
nand U14201 (N_14201,N_5473,N_2361);
nand U14202 (N_14202,N_4186,N_3468);
and U14203 (N_14203,N_977,N_8153);
and U14204 (N_14204,N_604,N_7331);
and U14205 (N_14205,N_3057,N_271);
xnor U14206 (N_14206,N_9152,N_8460);
nor U14207 (N_14207,N_6923,N_8654);
xnor U14208 (N_14208,N_9032,N_8189);
and U14209 (N_14209,N_1017,N_514);
nor U14210 (N_14210,N_9229,N_2636);
or U14211 (N_14211,N_2945,N_9135);
nor U14212 (N_14212,N_8802,N_9333);
and U14213 (N_14213,N_4640,N_6893);
nand U14214 (N_14214,N_4180,N_2711);
nor U14215 (N_14215,N_4699,N_8634);
nand U14216 (N_14216,N_798,N_3082);
or U14217 (N_14217,N_3800,N_8177);
xor U14218 (N_14218,N_1971,N_2203);
xor U14219 (N_14219,N_7396,N_8520);
nor U14220 (N_14220,N_6780,N_617);
or U14221 (N_14221,N_4272,N_3183);
nor U14222 (N_14222,N_6819,N_627);
nor U14223 (N_14223,N_202,N_1043);
or U14224 (N_14224,N_1395,N_9545);
and U14225 (N_14225,N_2825,N_2677);
nand U14226 (N_14226,N_6760,N_302);
and U14227 (N_14227,N_7003,N_9923);
nor U14228 (N_14228,N_7749,N_3473);
nand U14229 (N_14229,N_6938,N_767);
and U14230 (N_14230,N_3113,N_118);
nand U14231 (N_14231,N_8040,N_8957);
and U14232 (N_14232,N_632,N_8317);
and U14233 (N_14233,N_7677,N_3440);
and U14234 (N_14234,N_9869,N_4328);
or U14235 (N_14235,N_3664,N_1399);
xor U14236 (N_14236,N_4980,N_810);
nor U14237 (N_14237,N_8336,N_1192);
or U14238 (N_14238,N_3395,N_1279);
xor U14239 (N_14239,N_1956,N_6265);
and U14240 (N_14240,N_3547,N_7868);
nand U14241 (N_14241,N_2560,N_4002);
or U14242 (N_14242,N_5730,N_3930);
and U14243 (N_14243,N_7113,N_1225);
nor U14244 (N_14244,N_8481,N_7350);
or U14245 (N_14245,N_4979,N_444);
or U14246 (N_14246,N_5770,N_4970);
or U14247 (N_14247,N_9728,N_8353);
and U14248 (N_14248,N_1968,N_2048);
nor U14249 (N_14249,N_4959,N_6124);
nor U14250 (N_14250,N_7988,N_6106);
and U14251 (N_14251,N_2903,N_4817);
nor U14252 (N_14252,N_3947,N_7802);
or U14253 (N_14253,N_8380,N_9971);
or U14254 (N_14254,N_882,N_7585);
or U14255 (N_14255,N_4705,N_1811);
and U14256 (N_14256,N_2267,N_4720);
and U14257 (N_14257,N_4075,N_7998);
nor U14258 (N_14258,N_6362,N_1066);
nand U14259 (N_14259,N_699,N_8067);
nor U14260 (N_14260,N_5706,N_8771);
and U14261 (N_14261,N_6555,N_6262);
and U14262 (N_14262,N_8192,N_8852);
or U14263 (N_14263,N_3411,N_1583);
or U14264 (N_14264,N_7423,N_1493);
nand U14265 (N_14265,N_6463,N_1732);
nor U14266 (N_14266,N_5645,N_8214);
xnor U14267 (N_14267,N_658,N_4591);
or U14268 (N_14268,N_9093,N_811);
and U14269 (N_14269,N_7825,N_9137);
xor U14270 (N_14270,N_5789,N_8679);
and U14271 (N_14271,N_4845,N_2542);
xor U14272 (N_14272,N_6038,N_8559);
or U14273 (N_14273,N_1436,N_5018);
nor U14274 (N_14274,N_5049,N_8424);
nand U14275 (N_14275,N_6231,N_9110);
xor U14276 (N_14276,N_4712,N_5009);
or U14277 (N_14277,N_2664,N_2174);
nand U14278 (N_14278,N_3416,N_4797);
nand U14279 (N_14279,N_3882,N_920);
nor U14280 (N_14280,N_8526,N_5385);
xor U14281 (N_14281,N_7153,N_9701);
nand U14282 (N_14282,N_7730,N_2457);
xnor U14283 (N_14283,N_9183,N_5235);
nand U14284 (N_14284,N_7386,N_6816);
nor U14285 (N_14285,N_9917,N_7378);
and U14286 (N_14286,N_7926,N_9031);
and U14287 (N_14287,N_9022,N_6985);
nand U14288 (N_14288,N_4636,N_2503);
and U14289 (N_14289,N_2751,N_9373);
or U14290 (N_14290,N_6329,N_7078);
nor U14291 (N_14291,N_960,N_3458);
and U14292 (N_14292,N_3476,N_4850);
or U14293 (N_14293,N_8349,N_8729);
or U14294 (N_14294,N_3915,N_2180);
nor U14295 (N_14295,N_2712,N_366);
and U14296 (N_14296,N_9781,N_7646);
xor U14297 (N_14297,N_2835,N_2420);
nor U14298 (N_14298,N_2207,N_1498);
nand U14299 (N_14299,N_2087,N_6910);
nand U14300 (N_14300,N_9029,N_1711);
xor U14301 (N_14301,N_3179,N_4940);
nand U14302 (N_14302,N_4389,N_7716);
and U14303 (N_14303,N_988,N_2819);
nor U14304 (N_14304,N_4508,N_2358);
nor U14305 (N_14305,N_3010,N_2182);
nor U14306 (N_14306,N_3318,N_9538);
and U14307 (N_14307,N_6419,N_1998);
xnor U14308 (N_14308,N_9705,N_3364);
nand U14309 (N_14309,N_4326,N_6274);
and U14310 (N_14310,N_7958,N_6573);
or U14311 (N_14311,N_6098,N_9318);
xor U14312 (N_14312,N_5116,N_9412);
nand U14313 (N_14313,N_7195,N_4951);
and U14314 (N_14314,N_4246,N_7661);
or U14315 (N_14315,N_2061,N_8338);
xor U14316 (N_14316,N_5720,N_411);
or U14317 (N_14317,N_4582,N_8226);
or U14318 (N_14318,N_4802,N_1943);
nand U14319 (N_14319,N_173,N_4630);
nor U14320 (N_14320,N_966,N_5607);
nor U14321 (N_14321,N_845,N_7007);
or U14322 (N_14322,N_5480,N_2536);
or U14323 (N_14323,N_7487,N_2962);
nand U14324 (N_14324,N_2096,N_724);
nand U14325 (N_14325,N_6063,N_4440);
xor U14326 (N_14326,N_8815,N_5164);
nor U14327 (N_14327,N_1180,N_2368);
and U14328 (N_14328,N_6946,N_7175);
or U14329 (N_14329,N_9313,N_7445);
nor U14330 (N_14330,N_7894,N_9787);
and U14331 (N_14331,N_9937,N_9960);
nand U14332 (N_14332,N_2435,N_5427);
or U14333 (N_14333,N_7872,N_3647);
nand U14334 (N_14334,N_5511,N_3514);
or U14335 (N_14335,N_7024,N_5338);
or U14336 (N_14336,N_2974,N_2287);
nor U14337 (N_14337,N_5975,N_5630);
nor U14338 (N_14338,N_8703,N_8355);
nand U14339 (N_14339,N_1173,N_8839);
and U14340 (N_14340,N_2058,N_3127);
and U14341 (N_14341,N_3495,N_9141);
xnor U14342 (N_14342,N_3730,N_3020);
nand U14343 (N_14343,N_1128,N_3077);
or U14344 (N_14344,N_9933,N_7224);
nor U14345 (N_14345,N_7853,N_1234);
or U14346 (N_14346,N_5189,N_4434);
and U14347 (N_14347,N_6331,N_6887);
nor U14348 (N_14348,N_4039,N_4992);
nand U14349 (N_14349,N_2467,N_5095);
xor U14350 (N_14350,N_2257,N_1540);
nand U14351 (N_14351,N_2376,N_5697);
nand U14352 (N_14352,N_705,N_2473);
and U14353 (N_14353,N_7596,N_9219);
or U14354 (N_14354,N_4621,N_8796);
or U14355 (N_14355,N_1,N_1091);
and U14356 (N_14356,N_8363,N_4713);
nand U14357 (N_14357,N_5055,N_3681);
nor U14358 (N_14358,N_949,N_1812);
or U14359 (N_14359,N_35,N_5007);
and U14360 (N_14360,N_8154,N_5946);
and U14361 (N_14361,N_7949,N_7456);
or U14362 (N_14362,N_6291,N_182);
or U14363 (N_14363,N_4493,N_826);
xor U14364 (N_14364,N_7571,N_3625);
nor U14365 (N_14365,N_4548,N_2202);
xnor U14366 (N_14366,N_8960,N_9216);
nand U14367 (N_14367,N_8682,N_9116);
nand U14368 (N_14368,N_3209,N_6328);
or U14369 (N_14369,N_64,N_7184);
nor U14370 (N_14370,N_3048,N_5623);
xnor U14371 (N_14371,N_5745,N_80);
and U14372 (N_14372,N_6842,N_4387);
and U14373 (N_14373,N_6840,N_3425);
xnor U14374 (N_14374,N_55,N_6726);
or U14375 (N_14375,N_9878,N_3136);
xor U14376 (N_14376,N_2655,N_9215);
nand U14377 (N_14377,N_5524,N_4259);
xnor U14378 (N_14378,N_8174,N_6973);
or U14379 (N_14379,N_8843,N_4226);
nor U14380 (N_14380,N_1206,N_9167);
nor U14381 (N_14381,N_4566,N_4618);
nor U14382 (N_14382,N_6047,N_6150);
or U14383 (N_14383,N_7418,N_3380);
and U14384 (N_14384,N_5801,N_2566);
or U14385 (N_14385,N_71,N_2416);
nor U14386 (N_14386,N_7630,N_3046);
or U14387 (N_14387,N_3016,N_4651);
or U14388 (N_14388,N_2121,N_8053);
nand U14389 (N_14389,N_1858,N_8161);
nor U14390 (N_14390,N_4996,N_5795);
nand U14391 (N_14391,N_9372,N_1229);
nor U14392 (N_14392,N_1562,N_2502);
nand U14393 (N_14393,N_963,N_8747);
nor U14394 (N_14394,N_2849,N_8941);
nand U14395 (N_14395,N_419,N_5626);
nor U14396 (N_14396,N_1510,N_1511);
nor U14397 (N_14397,N_20,N_9047);
or U14398 (N_14398,N_8962,N_8948);
or U14399 (N_14399,N_9658,N_2036);
and U14400 (N_14400,N_4776,N_5062);
nand U14401 (N_14401,N_1349,N_2558);
and U14402 (N_14402,N_454,N_5527);
nor U14403 (N_14403,N_1014,N_5341);
and U14404 (N_14404,N_6376,N_9786);
nor U14405 (N_14405,N_6833,N_9500);
and U14406 (N_14406,N_2594,N_3851);
nand U14407 (N_14407,N_6528,N_8963);
and U14408 (N_14408,N_9261,N_8023);
nand U14409 (N_14409,N_6392,N_4808);
xor U14410 (N_14410,N_1306,N_7158);
or U14411 (N_14411,N_8501,N_4824);
nand U14412 (N_14412,N_6055,N_4806);
or U14413 (N_14413,N_1883,N_3262);
xor U14414 (N_14414,N_728,N_5830);
nor U14415 (N_14415,N_393,N_89);
and U14416 (N_14416,N_4369,N_3593);
and U14417 (N_14417,N_5301,N_1314);
and U14418 (N_14418,N_4490,N_9653);
nand U14419 (N_14419,N_8319,N_3115);
and U14420 (N_14420,N_2908,N_7757);
xor U14421 (N_14421,N_69,N_1928);
nand U14422 (N_14422,N_8790,N_5470);
nand U14423 (N_14423,N_268,N_1623);
nor U14424 (N_14424,N_8907,N_8788);
or U14425 (N_14425,N_8868,N_323);
or U14426 (N_14426,N_3981,N_360);
and U14427 (N_14427,N_7359,N_8394);
nand U14428 (N_14428,N_8542,N_4005);
nor U14429 (N_14429,N_6061,N_9070);
nand U14430 (N_14430,N_4962,N_4331);
or U14431 (N_14431,N_8527,N_7035);
or U14432 (N_14432,N_3018,N_2733);
or U14433 (N_14433,N_2858,N_1882);
nor U14434 (N_14434,N_3961,N_6318);
and U14435 (N_14435,N_2896,N_2217);
or U14436 (N_14436,N_2523,N_8072);
or U14437 (N_14437,N_1958,N_8140);
nand U14438 (N_14438,N_2686,N_9081);
nand U14439 (N_14439,N_5727,N_1016);
and U14440 (N_14440,N_9927,N_4488);
nor U14441 (N_14441,N_1086,N_6558);
or U14442 (N_14442,N_5983,N_4675);
nand U14443 (N_14443,N_229,N_8792);
or U14444 (N_14444,N_6139,N_6275);
nor U14445 (N_14445,N_2093,N_9380);
nand U14446 (N_14446,N_5418,N_2934);
xor U14447 (N_14447,N_8969,N_6260);
nand U14448 (N_14448,N_7042,N_5554);
nor U14449 (N_14449,N_4273,N_5561);
and U14450 (N_14450,N_9544,N_2743);
or U14451 (N_14451,N_1782,N_6608);
nor U14452 (N_14452,N_6917,N_795);
nand U14453 (N_14453,N_8236,N_1357);
nand U14454 (N_14454,N_4580,N_2605);
and U14455 (N_14455,N_9493,N_9025);
nor U14456 (N_14456,N_6986,N_7145);
and U14457 (N_14457,N_9155,N_9926);
xnor U14458 (N_14458,N_4036,N_3857);
or U14459 (N_14459,N_3237,N_1783);
or U14460 (N_14460,N_2200,N_1078);
nand U14461 (N_14461,N_4392,N_6630);
and U14462 (N_14462,N_7798,N_7900);
nor U14463 (N_14463,N_9802,N_8147);
or U14464 (N_14464,N_768,N_5912);
xnor U14465 (N_14465,N_9697,N_9707);
nand U14466 (N_14466,N_693,N_6725);
and U14467 (N_14467,N_4170,N_2774);
nor U14468 (N_14468,N_5884,N_616);
nor U14469 (N_14469,N_3816,N_9098);
or U14470 (N_14470,N_5685,N_2273);
or U14471 (N_14471,N_9350,N_1023);
nand U14472 (N_14472,N_2894,N_1119);
and U14473 (N_14473,N_1106,N_4153);
nor U14474 (N_14474,N_2278,N_8208);
or U14475 (N_14475,N_1902,N_1586);
or U14476 (N_14476,N_2761,N_3889);
nand U14477 (N_14477,N_7970,N_9325);
nand U14478 (N_14478,N_2039,N_9499);
or U14479 (N_14479,N_7692,N_4383);
or U14480 (N_14480,N_9411,N_9634);
nand U14481 (N_14481,N_7309,N_1639);
or U14482 (N_14482,N_8202,N_1265);
xor U14483 (N_14483,N_6449,N_1374);
and U14484 (N_14484,N_8411,N_1780);
and U14485 (N_14485,N_709,N_568);
xor U14486 (N_14486,N_1060,N_8239);
and U14487 (N_14487,N_432,N_3338);
nor U14488 (N_14488,N_8468,N_4860);
or U14489 (N_14489,N_6089,N_1160);
xor U14490 (N_14490,N_6844,N_4643);
and U14491 (N_14491,N_9604,N_872);
nor U14492 (N_14492,N_2176,N_6955);
and U14493 (N_14493,N_3598,N_6143);
and U14494 (N_14494,N_5406,N_9795);
or U14495 (N_14495,N_5247,N_6568);
nand U14496 (N_14496,N_352,N_5962);
xnor U14497 (N_14497,N_4809,N_4578);
nand U14498 (N_14498,N_4529,N_6750);
or U14499 (N_14499,N_4818,N_7563);
or U14500 (N_14500,N_8257,N_3368);
or U14501 (N_14501,N_2237,N_2343);
nor U14502 (N_14502,N_5305,N_4146);
or U14503 (N_14503,N_1852,N_9770);
and U14504 (N_14504,N_6422,N_7541);
xnor U14505 (N_14505,N_4362,N_7779);
nor U14506 (N_14506,N_3702,N_9631);
or U14507 (N_14507,N_4230,N_2122);
and U14508 (N_14508,N_8157,N_1266);
and U14509 (N_14509,N_2494,N_7790);
nor U14510 (N_14510,N_1687,N_2559);
and U14511 (N_14511,N_3847,N_8024);
nor U14512 (N_14512,N_7257,N_4510);
nor U14513 (N_14513,N_8942,N_4538);
or U14514 (N_14514,N_3590,N_715);
nor U14515 (N_14515,N_6465,N_540);
xnor U14516 (N_14516,N_3833,N_8706);
and U14517 (N_14517,N_2718,N_304);
nand U14518 (N_14518,N_7559,N_6140);
and U14519 (N_14519,N_8927,N_1129);
nand U14520 (N_14520,N_2756,N_1909);
and U14521 (N_14521,N_3597,N_978);
nand U14522 (N_14522,N_9272,N_9111);
nand U14523 (N_14523,N_5328,N_3013);
and U14524 (N_14524,N_9165,N_1563);
nand U14525 (N_14525,N_8818,N_4521);
and U14526 (N_14526,N_314,N_2135);
and U14527 (N_14527,N_4229,N_3378);
nand U14528 (N_14528,N_2016,N_1082);
nand U14529 (N_14529,N_433,N_9042);
and U14530 (N_14530,N_1272,N_1582);
nand U14531 (N_14531,N_3670,N_5053);
and U14532 (N_14532,N_3276,N_2608);
or U14533 (N_14533,N_3564,N_8457);
and U14534 (N_14534,N_9565,N_480);
or U14535 (N_14535,N_4338,N_7409);
nor U14536 (N_14536,N_8453,N_1625);
xnor U14537 (N_14537,N_5782,N_7931);
nor U14538 (N_14538,N_9011,N_8939);
or U14539 (N_14539,N_501,N_3741);
nor U14540 (N_14540,N_4671,N_9665);
xnor U14541 (N_14541,N_8982,N_6621);
xnor U14542 (N_14542,N_7877,N_2533);
nor U14543 (N_14543,N_5275,N_8572);
xor U14544 (N_14544,N_8932,N_2726);
nor U14545 (N_14545,N_9345,N_47);
or U14546 (N_14546,N_2515,N_5605);
nand U14547 (N_14547,N_5028,N_4089);
or U14548 (N_14548,N_9446,N_4968);
nand U14549 (N_14549,N_5581,N_7225);
nand U14550 (N_14550,N_2650,N_2500);
nor U14551 (N_14551,N_6654,N_6285);
xnor U14552 (N_14552,N_2931,N_4016);
xnor U14553 (N_14553,N_1933,N_7204);
nor U14554 (N_14554,N_3051,N_4949);
xor U14555 (N_14555,N_4427,N_6446);
and U14556 (N_14556,N_4308,N_2495);
nor U14557 (N_14557,N_8370,N_8504);
or U14558 (N_14558,N_6999,N_973);
and U14559 (N_14559,N_7980,N_4367);
and U14560 (N_14560,N_2075,N_7014);
nand U14561 (N_14561,N_3639,N_1408);
nand U14562 (N_14562,N_1606,N_3026);
or U14563 (N_14563,N_8188,N_5579);
and U14564 (N_14564,N_1807,N_9020);
nor U14565 (N_14565,N_381,N_4927);
or U14566 (N_14566,N_6982,N_3524);
nor U14567 (N_14567,N_32,N_9211);
or U14568 (N_14568,N_5135,N_3725);
xnor U14569 (N_14569,N_7639,N_3954);
or U14570 (N_14570,N_5823,N_614);
nor U14571 (N_14571,N_4771,N_7739);
or U14572 (N_14572,N_5517,N_666);
nand U14573 (N_14573,N_7964,N_4148);
nand U14574 (N_14574,N_2948,N_6939);
xor U14575 (N_14575,N_3359,N_3019);
and U14576 (N_14576,N_3362,N_2431);
nor U14577 (N_14577,N_6005,N_6954);
or U14578 (N_14578,N_7848,N_5841);
and U14579 (N_14579,N_5264,N_4000);
xor U14580 (N_14580,N_214,N_6216);
nand U14581 (N_14581,N_7785,N_3796);
and U14582 (N_14582,N_8775,N_7684);
xnor U14583 (N_14583,N_3551,N_500);
and U14584 (N_14584,N_8426,N_5132);
or U14585 (N_14585,N_7075,N_6736);
nor U14586 (N_14586,N_4465,N_4257);
and U14587 (N_14587,N_2054,N_1145);
nor U14588 (N_14588,N_4472,N_993);
and U14589 (N_14589,N_5176,N_5787);
or U14590 (N_14590,N_329,N_3254);
or U14591 (N_14591,N_5300,N_1140);
nand U14592 (N_14592,N_1585,N_9010);
nand U14593 (N_14593,N_9455,N_8030);
nand U14594 (N_14594,N_6578,N_6914);
nor U14595 (N_14595,N_639,N_8736);
nand U14596 (N_14596,N_1618,N_2344);
nand U14597 (N_14597,N_1942,N_2898);
nand U14598 (N_14598,N_1806,N_9055);
nand U14599 (N_14599,N_3118,N_4553);
or U14600 (N_14600,N_4923,N_3158);
nor U14601 (N_14601,N_54,N_5790);
or U14602 (N_14602,N_908,N_4587);
nand U14603 (N_14603,N_143,N_10);
nand U14604 (N_14604,N_4029,N_467);
nand U14605 (N_14605,N_4743,N_5759);
or U14606 (N_14606,N_1842,N_469);
nand U14607 (N_14607,N_8741,N_5078);
or U14608 (N_14608,N_6406,N_6669);
and U14609 (N_14609,N_1226,N_172);
or U14610 (N_14610,N_847,N_2998);
or U14611 (N_14611,N_5266,N_4698);
and U14612 (N_14612,N_3044,N_2544);
and U14613 (N_14613,N_9839,N_6458);
or U14614 (N_14614,N_8538,N_6079);
or U14615 (N_14615,N_4261,N_7955);
and U14616 (N_14616,N_4916,N_8827);
nor U14617 (N_14617,N_7906,N_4880);
and U14618 (N_14618,N_3088,N_4188);
and U14619 (N_14619,N_9484,N_3275);
nor U14620 (N_14620,N_2333,N_325);
and U14621 (N_14621,N_7547,N_9672);
and U14622 (N_14622,N_775,N_269);
nor U14623 (N_14623,N_7289,N_4134);
nand U14624 (N_14624,N_8739,N_994);
xnor U14625 (N_14625,N_8841,N_5272);
nand U14626 (N_14626,N_9763,N_2151);
and U14627 (N_14627,N_7544,N_6751);
and U14628 (N_14628,N_4803,N_6544);
or U14629 (N_14629,N_4731,N_5502);
and U14630 (N_14630,N_7713,N_7437);
or U14631 (N_14631,N_5835,N_6795);
nand U14632 (N_14632,N_6032,N_4086);
nor U14633 (N_14633,N_7095,N_9390);
xnor U14634 (N_14634,N_37,N_3979);
and U14635 (N_14635,N_8283,N_4984);
and U14636 (N_14636,N_4047,N_905);
xor U14637 (N_14637,N_9911,N_7001);
nand U14638 (N_14638,N_2853,N_4085);
nor U14639 (N_14639,N_9095,N_7608);
xnor U14640 (N_14640,N_6678,N_2629);
and U14641 (N_14641,N_2302,N_5763);
nor U14642 (N_14642,N_1823,N_9175);
and U14643 (N_14643,N_7752,N_9743);
and U14644 (N_14644,N_521,N_439);
xor U14645 (N_14645,N_1002,N_537);
xor U14646 (N_14646,N_7573,N_2242);
or U14647 (N_14647,N_6304,N_8975);
nor U14648 (N_14648,N_8392,N_4659);
and U14649 (N_14649,N_2572,N_4805);
nor U14650 (N_14650,N_1531,N_8600);
or U14651 (N_14651,N_5909,N_583);
or U14652 (N_14652,N_3737,N_3307);
and U14653 (N_14653,N_6721,N_7325);
and U14654 (N_14654,N_2826,N_3638);
and U14655 (N_14655,N_8454,N_121);
nand U14656 (N_14656,N_3454,N_4475);
and U14657 (N_14657,N_1311,N_1093);
or U14658 (N_14658,N_9357,N_6687);
nor U14659 (N_14659,N_3021,N_5190);
or U14660 (N_14660,N_9650,N_7091);
or U14661 (N_14661,N_7941,N_7618);
nor U14662 (N_14662,N_8293,N_6570);
and U14663 (N_14663,N_4022,N_7394);
xnor U14664 (N_14664,N_2737,N_5535);
nor U14665 (N_14665,N_1233,N_5679);
nor U14666 (N_14666,N_9463,N_8458);
and U14667 (N_14667,N_5425,N_3677);
and U14668 (N_14668,N_2933,N_3688);
nand U14669 (N_14669,N_1704,N_6789);
nand U14670 (N_14670,N_2480,N_6921);
and U14671 (N_14671,N_692,N_5519);
xor U14672 (N_14672,N_1570,N_5856);
or U14673 (N_14673,N_9138,N_3358);
and U14674 (N_14674,N_2687,N_5686);
nand U14675 (N_14675,N_8760,N_1923);
and U14676 (N_14676,N_473,N_8095);
and U14677 (N_14677,N_2630,N_499);
or U14678 (N_14678,N_8925,N_7812);
and U14679 (N_14679,N_8461,N_4233);
nand U14680 (N_14680,N_9262,N_4168);
and U14681 (N_14681,N_7140,N_2690);
and U14682 (N_14682,N_8401,N_7041);
or U14683 (N_14683,N_2194,N_5684);
nor U14684 (N_14684,N_5642,N_3366);
nand U14685 (N_14685,N_4470,N_2158);
nand U14686 (N_14686,N_9355,N_5082);
and U14687 (N_14687,N_7141,N_3070);
nand U14688 (N_14688,N_3519,N_9334);
nand U14689 (N_14689,N_1642,N_7994);
nand U14690 (N_14690,N_4116,N_4195);
xor U14691 (N_14691,N_8277,N_2265);
nor U14692 (N_14692,N_9119,N_6160);
and U14693 (N_14693,N_5681,N_717);
or U14694 (N_14694,N_8417,N_1250);
nand U14695 (N_14695,N_5263,N_9825);
or U14696 (N_14696,N_9584,N_1457);
nand U14697 (N_14697,N_974,N_6234);
nor U14698 (N_14698,N_7521,N_1963);
or U14699 (N_14699,N_372,N_3852);
and U14700 (N_14700,N_7143,N_1411);
nand U14701 (N_14701,N_1674,N_8759);
and U14702 (N_14702,N_5802,N_9428);
or U14703 (N_14703,N_7380,N_8878);
and U14704 (N_14704,N_8616,N_8651);
nor U14705 (N_14705,N_4177,N_9023);
nor U14706 (N_14706,N_347,N_8934);
nand U14707 (N_14707,N_43,N_4920);
nand U14708 (N_14708,N_6043,N_8720);
or U14709 (N_14709,N_1887,N_2707);
nor U14710 (N_14710,N_3354,N_7885);
nand U14711 (N_14711,N_2693,N_1518);
xnor U14712 (N_14712,N_9437,N_2074);
and U14713 (N_14713,N_383,N_9559);
nand U14714 (N_14714,N_4641,N_5542);
and U14715 (N_14715,N_9651,N_5279);
nand U14716 (N_14716,N_6529,N_9288);
nand U14717 (N_14717,N_2562,N_1914);
nor U14718 (N_14718,N_2491,N_1108);
and U14719 (N_14719,N_2609,N_4318);
or U14720 (N_14720,N_3668,N_672);
xor U14721 (N_14721,N_6745,N_5370);
or U14722 (N_14722,N_3406,N_7188);
and U14723 (N_14723,N_8627,N_4210);
nor U14724 (N_14724,N_4111,N_7116);
and U14725 (N_14725,N_3497,N_3292);
or U14726 (N_14726,N_2688,N_8987);
nand U14727 (N_14727,N_4679,N_607);
and U14728 (N_14728,N_6699,N_4801);
and U14729 (N_14729,N_297,N_9132);
or U14730 (N_14730,N_4772,N_7960);
nand U14731 (N_14731,N_3829,N_6000);
nand U14732 (N_14732,N_5122,N_6421);
nor U14733 (N_14733,N_5205,N_3233);
xor U14734 (N_14734,N_4467,N_6860);
nand U14735 (N_14735,N_9476,N_7981);
or U14736 (N_14736,N_8164,N_9969);
and U14737 (N_14737,N_8973,N_8435);
or U14738 (N_14738,N_2510,N_2476);
nor U14739 (N_14739,N_5459,N_7107);
or U14740 (N_14740,N_78,N_3068);
or U14741 (N_14741,N_6052,N_6812);
nor U14742 (N_14742,N_49,N_6547);
or U14743 (N_14743,N_7316,N_8171);
nor U14744 (N_14744,N_4225,N_4064);
and U14745 (N_14745,N_5219,N_2602);
and U14746 (N_14746,N_6103,N_2109);
xnor U14747 (N_14747,N_1462,N_8866);
xor U14748 (N_14748,N_764,N_9244);
nor U14749 (N_14749,N_3689,N_131);
or U14750 (N_14750,N_8224,N_8768);
nand U14751 (N_14751,N_8418,N_9375);
and U14752 (N_14752,N_1211,N_6835);
and U14753 (N_14753,N_5967,N_4382);
or U14754 (N_14754,N_8979,N_6591);
nor U14755 (N_14755,N_1865,N_7750);
nand U14756 (N_14756,N_5172,N_9769);
nand U14757 (N_14757,N_7913,N_6078);
nand U14758 (N_14758,N_5937,N_8730);
nor U14759 (N_14759,N_7120,N_3920);
nor U14760 (N_14760,N_2883,N_3550);
nor U14761 (N_14761,N_4489,N_3732);
and U14762 (N_14762,N_3041,N_4581);
or U14763 (N_14763,N_575,N_5928);
or U14764 (N_14764,N_3909,N_365);
or U14765 (N_14765,N_4625,N_2969);
or U14766 (N_14766,N_7162,N_8443);
and U14767 (N_14767,N_1104,N_4320);
or U14768 (N_14768,N_8055,N_7737);
nor U14769 (N_14769,N_4336,N_9348);
or U14770 (N_14770,N_8217,N_9071);
nor U14771 (N_14771,N_7164,N_8795);
xor U14772 (N_14772,N_8206,N_1675);
nor U14773 (N_14773,N_6933,N_6781);
and U14774 (N_14774,N_1084,N_4981);
or U14775 (N_14775,N_1657,N_2623);
nor U14776 (N_14776,N_4162,N_9529);
nor U14777 (N_14777,N_605,N_3680);
nor U14778 (N_14778,N_5639,N_1252);
nand U14779 (N_14779,N_1197,N_2064);
xor U14780 (N_14780,N_8647,N_4483);
nor U14781 (N_14781,N_7754,N_4560);
nor U14782 (N_14782,N_2041,N_9069);
or U14783 (N_14783,N_6609,N_879);
and U14784 (N_14784,N_9897,N_7096);
nor U14785 (N_14785,N_7691,N_169);
or U14786 (N_14786,N_8842,N_5254);
or U14787 (N_14787,N_2261,N_7478);
nand U14788 (N_14788,N_9304,N_2867);
nor U14789 (N_14789,N_1482,N_1346);
nand U14790 (N_14790,N_4299,N_1936);
and U14791 (N_14791,N_8867,N_6447);
xor U14792 (N_14792,N_5142,N_5905);
and U14793 (N_14793,N_5037,N_4604);
nor U14794 (N_14794,N_206,N_2799);
nand U14795 (N_14795,N_6416,N_6462);
and U14796 (N_14796,N_5885,N_4019);
or U14797 (N_14797,N_6814,N_9449);
and U14798 (N_14798,N_7214,N_5562);
and U14799 (N_14799,N_4820,N_7965);
and U14800 (N_14800,N_1080,N_3263);
and U14801 (N_14801,N_5739,N_2046);
nor U14802 (N_14802,N_859,N_461);
nor U14803 (N_14803,N_4536,N_4056);
and U14804 (N_14804,N_8243,N_5537);
or U14805 (N_14805,N_8091,N_9595);
nor U14806 (N_14806,N_82,N_6144);
or U14807 (N_14807,N_3663,N_7227);
nand U14808 (N_14808,N_3747,N_3927);
or U14809 (N_14809,N_479,N_9929);
nand U14810 (N_14810,N_9091,N_7721);
nand U14811 (N_14811,N_888,N_9799);
nor U14812 (N_14812,N_5529,N_1705);
nand U14813 (N_14813,N_3776,N_8045);
nor U14814 (N_14814,N_6253,N_9403);
or U14815 (N_14815,N_7695,N_1019);
or U14816 (N_14816,N_5253,N_7781);
or U14817 (N_14817,N_3145,N_2465);
nor U14818 (N_14818,N_6088,N_2282);
nand U14819 (N_14819,N_4694,N_92);
nand U14820 (N_14820,N_3855,N_3715);
nand U14821 (N_14821,N_7916,N_523);
nor U14822 (N_14822,N_1987,N_4530);
nor U14823 (N_14823,N_5244,N_4518);
or U14824 (N_14824,N_9967,N_6149);
nor U14825 (N_14825,N_4821,N_1546);
nand U14826 (N_14826,N_396,N_3204);
nor U14827 (N_14827,N_448,N_9530);
nor U14828 (N_14828,N_3650,N_9616);
nand U14829 (N_14829,N_9128,N_9703);
and U14830 (N_14830,N_4779,N_610);
nand U14831 (N_14831,N_2291,N_5973);
nor U14832 (N_14832,N_5150,N_5952);
or U14833 (N_14833,N_2197,N_4132);
and U14834 (N_14834,N_1635,N_6086);
xnor U14835 (N_14835,N_1796,N_735);
nor U14836 (N_14836,N_2359,N_2714);
nor U14837 (N_14837,N_9008,N_1685);
and U14838 (N_14838,N_8968,N_2110);
and U14839 (N_14839,N_3679,N_5121);
nor U14840 (N_14840,N_5516,N_2279);
nor U14841 (N_14841,N_493,N_3053);
nand U14842 (N_14842,N_7600,N_3841);
or U14843 (N_14843,N_6054,N_2252);
nor U14844 (N_14844,N_7852,N_5066);
nand U14845 (N_14845,N_7379,N_5335);
nand U14846 (N_14846,N_8318,N_338);
and U14847 (N_14847,N_1379,N_9043);
nand U14848 (N_14848,N_3901,N_5670);
nor U14849 (N_14849,N_5689,N_4645);
or U14850 (N_14850,N_3493,N_2838);
nand U14851 (N_14851,N_4045,N_516);
nor U14852 (N_14852,N_3719,N_9877);
or U14853 (N_14853,N_4399,N_850);
nand U14854 (N_14854,N_9207,N_3239);
xnor U14855 (N_14855,N_9208,N_5765);
nor U14856 (N_14856,N_4937,N_7612);
nand U14857 (N_14857,N_9997,N_4207);
and U14858 (N_14858,N_303,N_553);
and U14859 (N_14859,N_6485,N_8908);
nor U14860 (N_14860,N_7598,N_9974);
or U14861 (N_14861,N_9594,N_7138);
or U14862 (N_14862,N_285,N_1855);
or U14863 (N_14863,N_5753,N_818);
and U14864 (N_14864,N_7533,N_8031);
and U14865 (N_14865,N_203,N_9260);
nand U14866 (N_14866,N_970,N_7117);
nand U14867 (N_14867,N_6735,N_9277);
nand U14868 (N_14868,N_4610,N_7115);
nor U14869 (N_14869,N_7427,N_1930);
nand U14870 (N_14870,N_7922,N_4241);
or U14871 (N_14871,N_6312,N_3379);
or U14872 (N_14872,N_6706,N_8823);
or U14873 (N_14873,N_6747,N_3986);
nand U14874 (N_14874,N_1095,N_7962);
nand U14875 (N_14875,N_3217,N_8385);
nor U14876 (N_14876,N_2372,N_7202);
nand U14877 (N_14877,N_1683,N_4418);
nand U14878 (N_14878,N_9468,N_2284);
xor U14879 (N_14879,N_9054,N_2812);
or U14880 (N_14880,N_1724,N_8263);
nand U14881 (N_14881,N_3393,N_2228);
nor U14882 (N_14882,N_1101,N_326);
or U14883 (N_14883,N_1616,N_510);
and U14884 (N_14884,N_5416,N_1245);
and U14885 (N_14885,N_8617,N_3245);
or U14886 (N_14886,N_5641,N_1706);
and U14887 (N_14887,N_9590,N_8347);
or U14888 (N_14888,N_2229,N_518);
xnor U14889 (N_14889,N_6204,N_8602);
nand U14890 (N_14890,N_1608,N_4691);
xor U14891 (N_14891,N_5379,N_8901);
nand U14892 (N_14892,N_7836,N_8274);
nand U14893 (N_14893,N_8579,N_6165);
xor U14894 (N_14894,N_6934,N_1305);
nand U14895 (N_14895,N_9791,N_7689);
nor U14896 (N_14896,N_2303,N_1010);
nand U14897 (N_14897,N_7905,N_2823);
nand U14898 (N_14898,N_7049,N_9527);
nor U14899 (N_14899,N_6320,N_8940);
nand U14900 (N_14900,N_961,N_7046);
or U14901 (N_14901,N_9510,N_3314);
nor U14902 (N_14902,N_9862,N_4505);
nor U14903 (N_14903,N_8013,N_405);
nand U14904 (N_14904,N_3795,N_4869);
nand U14905 (N_14905,N_4517,N_434);
and U14906 (N_14906,N_1111,N_6413);
nand U14907 (N_14907,N_3104,N_8779);
xnor U14908 (N_14908,N_9953,N_4251);
xnor U14909 (N_14909,N_4095,N_9059);
and U14910 (N_14910,N_7176,N_9097);
nand U14911 (N_14911,N_9310,N_8012);
and U14912 (N_14912,N_9585,N_6299);
xor U14913 (N_14913,N_5555,N_5441);
or U14914 (N_14914,N_5656,N_8124);
or U14915 (N_14915,N_5458,N_1288);
nor U14916 (N_14916,N_1576,N_8574);
or U14917 (N_14917,N_8172,N_1463);
and U14918 (N_14918,N_3951,N_8692);
and U14919 (N_14919,N_2270,N_9024);
nand U14920 (N_14920,N_3773,N_3838);
nand U14921 (N_14921,N_6280,N_40);
nand U14922 (N_14922,N_8991,N_2479);
or U14923 (N_14923,N_4955,N_5001);
nand U14924 (N_14924,N_7220,N_2549);
and U14925 (N_14925,N_3420,N_3100);
or U14926 (N_14926,N_7344,N_5541);
nand U14927 (N_14927,N_4571,N_839);
and U14928 (N_14928,N_646,N_8103);
xor U14929 (N_14929,N_5536,N_5840);
or U14930 (N_14930,N_8929,N_4378);
nor U14931 (N_14931,N_6908,N_4011);
nor U14932 (N_14932,N_1103,N_3884);
xnor U14933 (N_14933,N_7669,N_5654);
nand U14934 (N_14934,N_257,N_5671);
or U14935 (N_14935,N_9398,N_840);
or U14936 (N_14936,N_8041,N_8135);
and U14937 (N_14937,N_8337,N_188);
nand U14938 (N_14938,N_7506,N_1348);
or U14939 (N_14939,N_9606,N_9913);
or U14940 (N_14940,N_6639,N_8513);
or U14941 (N_14941,N_2730,N_160);
xnor U14942 (N_14942,N_9237,N_1808);
xnor U14943 (N_14943,N_799,N_1162);
nor U14944 (N_14944,N_3355,N_9924);
or U14945 (N_14945,N_944,N_5398);
nand U14946 (N_14946,N_4886,N_5771);
nor U14947 (N_14947,N_1131,N_7939);
and U14948 (N_14948,N_6744,N_9045);
nor U14949 (N_14949,N_7548,N_1497);
and U14950 (N_14950,N_1593,N_2126);
nand U14951 (N_14951,N_1697,N_579);
and U14952 (N_14952,N_1997,N_1049);
nor U14953 (N_14953,N_8683,N_7953);
xnor U14954 (N_14954,N_4013,N_3494);
nand U14955 (N_14955,N_26,N_4194);
nor U14956 (N_14956,N_5932,N_9523);
or U14957 (N_14957,N_7352,N_3287);
and U14958 (N_14958,N_6279,N_8519);
xor U14959 (N_14959,N_4485,N_4555);
and U14960 (N_14960,N_9378,N_8748);
xor U14961 (N_14961,N_6341,N_4693);
or U14962 (N_14962,N_1096,N_2587);
or U14963 (N_14963,N_4105,N_6824);
or U14964 (N_14964,N_1112,N_2893);
and U14965 (N_14965,N_4843,N_3226);
xor U14966 (N_14966,N_7566,N_9715);
or U14967 (N_14967,N_5238,N_6240);
nor U14968 (N_14968,N_4748,N_7531);
xor U14969 (N_14969,N_7294,N_9698);
nor U14970 (N_14970,N_9547,N_4762);
or U14971 (N_14971,N_4550,N_2347);
and U14972 (N_14972,N_8637,N_6408);
and U14973 (N_14973,N_7518,N_9166);
nand U14974 (N_14974,N_6521,N_4092);
or U14975 (N_14975,N_4841,N_5688);
or U14976 (N_14976,N_2177,N_5359);
nor U14977 (N_14977,N_7967,N_4574);
nor U14978 (N_14978,N_5377,N_9742);
nor U14979 (N_14979,N_4062,N_9640);
nand U14980 (N_14980,N_6487,N_5229);
nand U14981 (N_14981,N_2886,N_418);
and U14982 (N_14982,N_757,N_3569);
nand U14983 (N_14983,N_1216,N_6154);
or U14984 (N_14984,N_5563,N_2505);
nand U14985 (N_14985,N_6269,N_1113);
nand U14986 (N_14986,N_4627,N_6467);
nor U14987 (N_14987,N_1186,N_3205);
nor U14988 (N_14988,N_2922,N_4967);
or U14989 (N_14989,N_6990,N_7768);
nand U14990 (N_14990,N_4474,N_6123);
nor U14991 (N_14991,N_4601,N_5762);
or U14992 (N_14992,N_643,N_5111);
and U14993 (N_14993,N_3883,N_554);
or U14994 (N_14994,N_9621,N_6702);
nor U14995 (N_14995,N_4341,N_4237);
nand U14996 (N_14996,N_2964,N_852);
xor U14997 (N_14997,N_5004,N_2443);
and U14998 (N_14998,N_6495,N_85);
and U14999 (N_14999,N_8133,N_2579);
nor U15000 (N_15000,N_1208,N_9638);
nand U15001 (N_15001,N_5518,N_7826);
nand U15002 (N_15002,N_4183,N_3745);
nand U15003 (N_15003,N_5146,N_8824);
nand U15004 (N_15004,N_9676,N_788);
nor U15005 (N_15005,N_4847,N_131);
nor U15006 (N_15006,N_1615,N_4622);
xor U15007 (N_15007,N_2095,N_2656);
nand U15008 (N_15008,N_4134,N_9639);
or U15009 (N_15009,N_9703,N_4754);
and U15010 (N_15010,N_6831,N_8952);
nand U15011 (N_15011,N_1742,N_3081);
or U15012 (N_15012,N_9578,N_1904);
nor U15013 (N_15013,N_7344,N_1334);
or U15014 (N_15014,N_2625,N_7629);
or U15015 (N_15015,N_2208,N_1018);
nand U15016 (N_15016,N_5024,N_4430);
or U15017 (N_15017,N_3159,N_2844);
nand U15018 (N_15018,N_5865,N_1175);
and U15019 (N_15019,N_4331,N_8118);
or U15020 (N_15020,N_1299,N_5904);
xor U15021 (N_15021,N_1070,N_4204);
nand U15022 (N_15022,N_3397,N_5998);
and U15023 (N_15023,N_7357,N_6166);
nand U15024 (N_15024,N_6234,N_3700);
or U15025 (N_15025,N_2047,N_1098);
nor U15026 (N_15026,N_2073,N_2433);
or U15027 (N_15027,N_1384,N_5482);
nor U15028 (N_15028,N_8217,N_5131);
or U15029 (N_15029,N_7145,N_7923);
nand U15030 (N_15030,N_6478,N_9182);
nor U15031 (N_15031,N_3289,N_4147);
and U15032 (N_15032,N_137,N_2776);
nor U15033 (N_15033,N_7862,N_8017);
nor U15034 (N_15034,N_7273,N_6521);
or U15035 (N_15035,N_1571,N_2693);
nor U15036 (N_15036,N_7613,N_7910);
nand U15037 (N_15037,N_1651,N_6375);
nand U15038 (N_15038,N_3433,N_2269);
and U15039 (N_15039,N_8372,N_5216);
nand U15040 (N_15040,N_1644,N_3629);
nand U15041 (N_15041,N_9515,N_1219);
nand U15042 (N_15042,N_8671,N_6101);
and U15043 (N_15043,N_4255,N_4697);
nor U15044 (N_15044,N_5980,N_2677);
nor U15045 (N_15045,N_5030,N_9792);
and U15046 (N_15046,N_2735,N_9098);
nor U15047 (N_15047,N_3741,N_7583);
and U15048 (N_15048,N_3276,N_4791);
nor U15049 (N_15049,N_7779,N_7362);
or U15050 (N_15050,N_1163,N_4113);
and U15051 (N_15051,N_6826,N_9991);
nand U15052 (N_15052,N_7408,N_2164);
nor U15053 (N_15053,N_2142,N_4026);
or U15054 (N_15054,N_2974,N_2529);
nor U15055 (N_15055,N_8671,N_328);
xor U15056 (N_15056,N_901,N_4192);
nor U15057 (N_15057,N_6311,N_326);
and U15058 (N_15058,N_7351,N_6161);
nor U15059 (N_15059,N_1648,N_6393);
xnor U15060 (N_15060,N_7619,N_1780);
xnor U15061 (N_15061,N_2793,N_5119);
or U15062 (N_15062,N_1691,N_1808);
nand U15063 (N_15063,N_5844,N_3830);
and U15064 (N_15064,N_4540,N_4143);
and U15065 (N_15065,N_797,N_8476);
nor U15066 (N_15066,N_3896,N_4068);
nor U15067 (N_15067,N_5714,N_8390);
and U15068 (N_15068,N_7157,N_1028);
and U15069 (N_15069,N_3911,N_6008);
or U15070 (N_15070,N_8460,N_994);
or U15071 (N_15071,N_7798,N_1687);
or U15072 (N_15072,N_9645,N_2321);
nand U15073 (N_15073,N_5905,N_6466);
and U15074 (N_15074,N_7739,N_3487);
nand U15075 (N_15075,N_3843,N_9332);
or U15076 (N_15076,N_9052,N_719);
nand U15077 (N_15077,N_1935,N_7122);
xor U15078 (N_15078,N_8392,N_2259);
and U15079 (N_15079,N_3040,N_3247);
nand U15080 (N_15080,N_1199,N_2319);
nor U15081 (N_15081,N_7660,N_7779);
xnor U15082 (N_15082,N_5243,N_6946);
nor U15083 (N_15083,N_4042,N_5870);
nor U15084 (N_15084,N_3147,N_8933);
or U15085 (N_15085,N_1653,N_9946);
xor U15086 (N_15086,N_953,N_1860);
nand U15087 (N_15087,N_5062,N_9616);
or U15088 (N_15088,N_8150,N_9644);
nor U15089 (N_15089,N_4001,N_8015);
and U15090 (N_15090,N_6796,N_7643);
nand U15091 (N_15091,N_3124,N_1027);
xor U15092 (N_15092,N_3763,N_8458);
and U15093 (N_15093,N_2784,N_9058);
or U15094 (N_15094,N_4112,N_7096);
nand U15095 (N_15095,N_8541,N_5567);
or U15096 (N_15096,N_590,N_2380);
nand U15097 (N_15097,N_3587,N_1409);
nand U15098 (N_15098,N_1850,N_2115);
nor U15099 (N_15099,N_9033,N_5608);
and U15100 (N_15100,N_5590,N_3480);
nand U15101 (N_15101,N_9988,N_4750);
nor U15102 (N_15102,N_7193,N_304);
xnor U15103 (N_15103,N_238,N_4239);
or U15104 (N_15104,N_7602,N_8);
and U15105 (N_15105,N_8854,N_9104);
nand U15106 (N_15106,N_7788,N_658);
xnor U15107 (N_15107,N_2424,N_400);
nand U15108 (N_15108,N_2019,N_2709);
nand U15109 (N_15109,N_3005,N_1891);
xnor U15110 (N_15110,N_2236,N_8403);
nor U15111 (N_15111,N_0,N_9325);
or U15112 (N_15112,N_9476,N_2383);
nand U15113 (N_15113,N_1261,N_4443);
nand U15114 (N_15114,N_3960,N_1493);
and U15115 (N_15115,N_4307,N_3708);
or U15116 (N_15116,N_2552,N_8413);
xnor U15117 (N_15117,N_447,N_1507);
nand U15118 (N_15118,N_246,N_6734);
or U15119 (N_15119,N_5118,N_9878);
and U15120 (N_15120,N_2037,N_4876);
and U15121 (N_15121,N_9187,N_6415);
nor U15122 (N_15122,N_1207,N_6117);
nor U15123 (N_15123,N_7601,N_249);
xnor U15124 (N_15124,N_7734,N_8851);
and U15125 (N_15125,N_6682,N_6603);
or U15126 (N_15126,N_8356,N_607);
xnor U15127 (N_15127,N_3525,N_7250);
and U15128 (N_15128,N_2861,N_661);
and U15129 (N_15129,N_5502,N_3067);
and U15130 (N_15130,N_8659,N_3902);
xor U15131 (N_15131,N_5598,N_3459);
or U15132 (N_15132,N_3539,N_3231);
nand U15133 (N_15133,N_1656,N_3744);
and U15134 (N_15134,N_3435,N_4270);
nor U15135 (N_15135,N_5530,N_9798);
or U15136 (N_15136,N_7888,N_9389);
nor U15137 (N_15137,N_118,N_8138);
nand U15138 (N_15138,N_4442,N_3885);
or U15139 (N_15139,N_7030,N_9239);
nor U15140 (N_15140,N_5932,N_4692);
or U15141 (N_15141,N_2793,N_4889);
nor U15142 (N_15142,N_1490,N_386);
nor U15143 (N_15143,N_299,N_4304);
or U15144 (N_15144,N_4584,N_6167);
nand U15145 (N_15145,N_9094,N_1189);
nor U15146 (N_15146,N_6010,N_7634);
nand U15147 (N_15147,N_5633,N_8108);
or U15148 (N_15148,N_2706,N_473);
nand U15149 (N_15149,N_7680,N_8781);
nand U15150 (N_15150,N_3289,N_1832);
and U15151 (N_15151,N_6932,N_126);
and U15152 (N_15152,N_94,N_196);
nand U15153 (N_15153,N_24,N_5791);
nor U15154 (N_15154,N_5531,N_8548);
nand U15155 (N_15155,N_8152,N_7889);
nor U15156 (N_15156,N_2788,N_5433);
and U15157 (N_15157,N_7607,N_3221);
and U15158 (N_15158,N_1630,N_8461);
or U15159 (N_15159,N_9249,N_8488);
and U15160 (N_15160,N_7322,N_4489);
nand U15161 (N_15161,N_8028,N_1558);
nand U15162 (N_15162,N_4456,N_8039);
nor U15163 (N_15163,N_8353,N_8135);
nor U15164 (N_15164,N_3528,N_2081);
xnor U15165 (N_15165,N_148,N_6524);
nor U15166 (N_15166,N_8322,N_2854);
nor U15167 (N_15167,N_6886,N_7291);
nor U15168 (N_15168,N_1,N_4191);
and U15169 (N_15169,N_3286,N_5643);
and U15170 (N_15170,N_4649,N_4779);
nor U15171 (N_15171,N_5227,N_2090);
and U15172 (N_15172,N_9212,N_1103);
nor U15173 (N_15173,N_9164,N_6442);
and U15174 (N_15174,N_2225,N_6424);
and U15175 (N_15175,N_7934,N_3366);
nand U15176 (N_15176,N_8410,N_5644);
nand U15177 (N_15177,N_822,N_7883);
nor U15178 (N_15178,N_998,N_9652);
nor U15179 (N_15179,N_1611,N_3805);
or U15180 (N_15180,N_8823,N_3282);
or U15181 (N_15181,N_8624,N_3971);
nand U15182 (N_15182,N_4589,N_9847);
nand U15183 (N_15183,N_7811,N_247);
and U15184 (N_15184,N_6827,N_7381);
nand U15185 (N_15185,N_5913,N_5584);
xor U15186 (N_15186,N_4305,N_5816);
nor U15187 (N_15187,N_3027,N_1029);
nor U15188 (N_15188,N_4710,N_7454);
or U15189 (N_15189,N_7801,N_4667);
nand U15190 (N_15190,N_7742,N_6502);
nor U15191 (N_15191,N_9725,N_9942);
and U15192 (N_15192,N_8026,N_5885);
nand U15193 (N_15193,N_8727,N_8248);
xnor U15194 (N_15194,N_913,N_2047);
or U15195 (N_15195,N_3590,N_6843);
or U15196 (N_15196,N_931,N_1202);
nor U15197 (N_15197,N_3534,N_1792);
nand U15198 (N_15198,N_4212,N_3488);
or U15199 (N_15199,N_5969,N_4913);
nor U15200 (N_15200,N_9897,N_7815);
nand U15201 (N_15201,N_7281,N_9734);
and U15202 (N_15202,N_8743,N_3474);
or U15203 (N_15203,N_7944,N_9504);
nor U15204 (N_15204,N_8524,N_4060);
nand U15205 (N_15205,N_6388,N_2566);
nand U15206 (N_15206,N_8449,N_6299);
nand U15207 (N_15207,N_9038,N_3650);
and U15208 (N_15208,N_2654,N_4919);
and U15209 (N_15209,N_5304,N_5281);
xor U15210 (N_15210,N_9033,N_2132);
nor U15211 (N_15211,N_842,N_1711);
nand U15212 (N_15212,N_7757,N_8657);
nor U15213 (N_15213,N_6941,N_8736);
or U15214 (N_15214,N_4953,N_423);
and U15215 (N_15215,N_5458,N_285);
xor U15216 (N_15216,N_9577,N_5232);
nand U15217 (N_15217,N_7334,N_5010);
and U15218 (N_15218,N_2627,N_761);
and U15219 (N_15219,N_8508,N_5748);
nand U15220 (N_15220,N_3279,N_3624);
nor U15221 (N_15221,N_3599,N_2828);
and U15222 (N_15222,N_8491,N_8654);
xor U15223 (N_15223,N_4768,N_1935);
nand U15224 (N_15224,N_3723,N_129);
nand U15225 (N_15225,N_9627,N_2252);
nor U15226 (N_15226,N_8587,N_672);
nand U15227 (N_15227,N_1652,N_262);
nand U15228 (N_15228,N_6613,N_7273);
nand U15229 (N_15229,N_1236,N_4012);
nand U15230 (N_15230,N_4976,N_9742);
xnor U15231 (N_15231,N_2127,N_905);
or U15232 (N_15232,N_9784,N_1341);
nand U15233 (N_15233,N_107,N_4399);
nor U15234 (N_15234,N_5725,N_9598);
and U15235 (N_15235,N_3410,N_3516);
and U15236 (N_15236,N_4864,N_6081);
and U15237 (N_15237,N_4099,N_8037);
xor U15238 (N_15238,N_7210,N_1860);
and U15239 (N_15239,N_2326,N_9614);
nand U15240 (N_15240,N_6807,N_9962);
nand U15241 (N_15241,N_9726,N_7450);
nor U15242 (N_15242,N_4697,N_5895);
nor U15243 (N_15243,N_729,N_9507);
or U15244 (N_15244,N_3208,N_6858);
and U15245 (N_15245,N_6875,N_6858);
or U15246 (N_15246,N_4449,N_5807);
nor U15247 (N_15247,N_9312,N_6014);
nand U15248 (N_15248,N_123,N_5190);
nor U15249 (N_15249,N_1349,N_3037);
or U15250 (N_15250,N_3402,N_9604);
nand U15251 (N_15251,N_4549,N_2445);
nand U15252 (N_15252,N_8427,N_4444);
nor U15253 (N_15253,N_4026,N_5066);
and U15254 (N_15254,N_9155,N_6149);
or U15255 (N_15255,N_9748,N_7704);
and U15256 (N_15256,N_2318,N_2963);
or U15257 (N_15257,N_1648,N_5466);
nor U15258 (N_15258,N_7893,N_9310);
and U15259 (N_15259,N_9619,N_967);
and U15260 (N_15260,N_450,N_8093);
nand U15261 (N_15261,N_8822,N_9981);
nor U15262 (N_15262,N_6030,N_6273);
or U15263 (N_15263,N_2862,N_7625);
or U15264 (N_15264,N_3846,N_6421);
or U15265 (N_15265,N_4070,N_483);
or U15266 (N_15266,N_1597,N_3592);
and U15267 (N_15267,N_9547,N_8514);
or U15268 (N_15268,N_5089,N_6511);
or U15269 (N_15269,N_7893,N_4073);
nand U15270 (N_15270,N_4019,N_1374);
or U15271 (N_15271,N_3828,N_9322);
nor U15272 (N_15272,N_572,N_8375);
and U15273 (N_15273,N_1860,N_367);
nand U15274 (N_15274,N_8398,N_458);
or U15275 (N_15275,N_5788,N_8721);
or U15276 (N_15276,N_6676,N_3312);
nand U15277 (N_15277,N_2901,N_5689);
and U15278 (N_15278,N_8623,N_6732);
nand U15279 (N_15279,N_3490,N_6594);
or U15280 (N_15280,N_2463,N_3869);
xor U15281 (N_15281,N_7638,N_5322);
or U15282 (N_15282,N_486,N_3394);
nand U15283 (N_15283,N_3718,N_5563);
nor U15284 (N_15284,N_6002,N_9993);
and U15285 (N_15285,N_4074,N_9213);
nand U15286 (N_15286,N_8081,N_1982);
nand U15287 (N_15287,N_5263,N_8121);
nor U15288 (N_15288,N_3627,N_4827);
xnor U15289 (N_15289,N_328,N_6133);
and U15290 (N_15290,N_3034,N_7271);
nor U15291 (N_15291,N_4196,N_6628);
nor U15292 (N_15292,N_4491,N_9418);
nor U15293 (N_15293,N_5604,N_9152);
nand U15294 (N_15294,N_991,N_6987);
xor U15295 (N_15295,N_2631,N_8779);
nand U15296 (N_15296,N_2509,N_4210);
nand U15297 (N_15297,N_743,N_7755);
or U15298 (N_15298,N_235,N_9069);
nand U15299 (N_15299,N_3550,N_1065);
nor U15300 (N_15300,N_3966,N_5063);
and U15301 (N_15301,N_2650,N_4933);
nor U15302 (N_15302,N_1024,N_4276);
and U15303 (N_15303,N_8392,N_6857);
or U15304 (N_15304,N_4020,N_1109);
nand U15305 (N_15305,N_2781,N_119);
nand U15306 (N_15306,N_3995,N_4557);
or U15307 (N_15307,N_8020,N_2250);
nand U15308 (N_15308,N_4295,N_1554);
or U15309 (N_15309,N_2324,N_2475);
nand U15310 (N_15310,N_7224,N_1769);
or U15311 (N_15311,N_1182,N_1794);
xnor U15312 (N_15312,N_2337,N_9555);
and U15313 (N_15313,N_184,N_8723);
or U15314 (N_15314,N_4289,N_3678);
nand U15315 (N_15315,N_6400,N_451);
and U15316 (N_15316,N_739,N_7982);
xor U15317 (N_15317,N_6312,N_4225);
and U15318 (N_15318,N_7603,N_6413);
nand U15319 (N_15319,N_5498,N_3457);
nor U15320 (N_15320,N_8940,N_6415);
and U15321 (N_15321,N_5716,N_1275);
and U15322 (N_15322,N_418,N_633);
or U15323 (N_15323,N_3295,N_8520);
nand U15324 (N_15324,N_4653,N_1158);
nand U15325 (N_15325,N_5917,N_9670);
nor U15326 (N_15326,N_378,N_9654);
and U15327 (N_15327,N_4068,N_8760);
or U15328 (N_15328,N_338,N_7319);
xnor U15329 (N_15329,N_9793,N_8877);
or U15330 (N_15330,N_917,N_6083);
or U15331 (N_15331,N_7210,N_7044);
and U15332 (N_15332,N_3043,N_7962);
or U15333 (N_15333,N_3463,N_4593);
nand U15334 (N_15334,N_4919,N_7406);
xor U15335 (N_15335,N_2185,N_8618);
and U15336 (N_15336,N_1254,N_5119);
or U15337 (N_15337,N_5605,N_257);
nand U15338 (N_15338,N_3110,N_5163);
or U15339 (N_15339,N_7280,N_5283);
xor U15340 (N_15340,N_5434,N_2151);
xor U15341 (N_15341,N_9141,N_9324);
nor U15342 (N_15342,N_7009,N_4516);
and U15343 (N_15343,N_1604,N_2930);
or U15344 (N_15344,N_7301,N_5361);
or U15345 (N_15345,N_3346,N_6389);
nor U15346 (N_15346,N_904,N_1295);
and U15347 (N_15347,N_549,N_4947);
or U15348 (N_15348,N_1669,N_547);
xnor U15349 (N_15349,N_25,N_3343);
nor U15350 (N_15350,N_1656,N_7120);
nand U15351 (N_15351,N_5798,N_6763);
or U15352 (N_15352,N_4281,N_4074);
and U15353 (N_15353,N_3713,N_3515);
nor U15354 (N_15354,N_4228,N_7896);
or U15355 (N_15355,N_312,N_5341);
nor U15356 (N_15356,N_6920,N_9255);
or U15357 (N_15357,N_3615,N_3879);
nor U15358 (N_15358,N_2887,N_964);
nor U15359 (N_15359,N_4080,N_6238);
xor U15360 (N_15360,N_5912,N_9254);
or U15361 (N_15361,N_7208,N_8418);
and U15362 (N_15362,N_8327,N_1188);
nand U15363 (N_15363,N_2642,N_5132);
and U15364 (N_15364,N_8600,N_2337);
nor U15365 (N_15365,N_5047,N_3548);
nand U15366 (N_15366,N_9700,N_1144);
and U15367 (N_15367,N_9515,N_7888);
or U15368 (N_15368,N_8548,N_8170);
and U15369 (N_15369,N_2625,N_6745);
nand U15370 (N_15370,N_5799,N_3758);
and U15371 (N_15371,N_9548,N_7473);
and U15372 (N_15372,N_1966,N_414);
nor U15373 (N_15373,N_1743,N_7200);
nor U15374 (N_15374,N_6711,N_6551);
and U15375 (N_15375,N_5844,N_5506);
xnor U15376 (N_15376,N_7410,N_5563);
nand U15377 (N_15377,N_8605,N_2977);
xnor U15378 (N_15378,N_8235,N_4885);
and U15379 (N_15379,N_813,N_1737);
nor U15380 (N_15380,N_3195,N_3453);
nand U15381 (N_15381,N_7303,N_9084);
and U15382 (N_15382,N_6189,N_4198);
nand U15383 (N_15383,N_1242,N_5759);
or U15384 (N_15384,N_282,N_7182);
nand U15385 (N_15385,N_6638,N_1405);
xnor U15386 (N_15386,N_4350,N_4059);
nor U15387 (N_15387,N_9784,N_2876);
nand U15388 (N_15388,N_842,N_5722);
or U15389 (N_15389,N_4330,N_4917);
or U15390 (N_15390,N_1601,N_5317);
and U15391 (N_15391,N_9174,N_9888);
nor U15392 (N_15392,N_8323,N_9764);
and U15393 (N_15393,N_821,N_1856);
nor U15394 (N_15394,N_4047,N_6037);
xnor U15395 (N_15395,N_2782,N_6219);
nor U15396 (N_15396,N_7189,N_239);
nand U15397 (N_15397,N_7922,N_5578);
and U15398 (N_15398,N_7780,N_829);
and U15399 (N_15399,N_1719,N_7462);
nor U15400 (N_15400,N_6310,N_8549);
or U15401 (N_15401,N_4726,N_3307);
nor U15402 (N_15402,N_4704,N_1878);
nor U15403 (N_15403,N_2615,N_3774);
and U15404 (N_15404,N_1572,N_9338);
and U15405 (N_15405,N_811,N_5866);
or U15406 (N_15406,N_3823,N_2580);
and U15407 (N_15407,N_3631,N_5344);
or U15408 (N_15408,N_9308,N_1269);
xnor U15409 (N_15409,N_7818,N_1877);
and U15410 (N_15410,N_1460,N_4199);
nand U15411 (N_15411,N_3760,N_4895);
nor U15412 (N_15412,N_8963,N_344);
nand U15413 (N_15413,N_613,N_9904);
and U15414 (N_15414,N_6502,N_3940);
nor U15415 (N_15415,N_2357,N_9276);
or U15416 (N_15416,N_1625,N_1081);
or U15417 (N_15417,N_3408,N_4242);
nand U15418 (N_15418,N_3672,N_9414);
nand U15419 (N_15419,N_1889,N_4859);
and U15420 (N_15420,N_1160,N_1741);
nand U15421 (N_15421,N_4491,N_3235);
and U15422 (N_15422,N_3345,N_7587);
xor U15423 (N_15423,N_3411,N_9077);
and U15424 (N_15424,N_5928,N_7573);
and U15425 (N_15425,N_1638,N_3128);
and U15426 (N_15426,N_6298,N_3989);
nand U15427 (N_15427,N_3249,N_8690);
and U15428 (N_15428,N_1847,N_1011);
nand U15429 (N_15429,N_6702,N_3301);
and U15430 (N_15430,N_4918,N_3003);
and U15431 (N_15431,N_8828,N_2329);
nand U15432 (N_15432,N_7929,N_3244);
or U15433 (N_15433,N_714,N_4238);
nor U15434 (N_15434,N_905,N_1817);
or U15435 (N_15435,N_1305,N_3229);
nand U15436 (N_15436,N_3446,N_6456);
nand U15437 (N_15437,N_7154,N_3021);
nor U15438 (N_15438,N_7601,N_779);
nand U15439 (N_15439,N_6315,N_7810);
nand U15440 (N_15440,N_2400,N_3962);
or U15441 (N_15441,N_5544,N_7137);
and U15442 (N_15442,N_4147,N_604);
nand U15443 (N_15443,N_4537,N_9234);
or U15444 (N_15444,N_9759,N_5179);
xor U15445 (N_15445,N_936,N_9352);
nand U15446 (N_15446,N_4579,N_2887);
and U15447 (N_15447,N_6179,N_3713);
or U15448 (N_15448,N_7084,N_63);
or U15449 (N_15449,N_9229,N_6107);
nand U15450 (N_15450,N_1101,N_7611);
xnor U15451 (N_15451,N_5,N_9669);
xnor U15452 (N_15452,N_2324,N_4345);
or U15453 (N_15453,N_3093,N_6166);
nor U15454 (N_15454,N_8034,N_6560);
nor U15455 (N_15455,N_3896,N_7101);
nor U15456 (N_15456,N_7065,N_7388);
or U15457 (N_15457,N_6578,N_1157);
and U15458 (N_15458,N_9623,N_9458);
or U15459 (N_15459,N_2287,N_1549);
or U15460 (N_15460,N_802,N_8698);
nand U15461 (N_15461,N_5084,N_9245);
or U15462 (N_15462,N_9865,N_1253);
and U15463 (N_15463,N_8497,N_7181);
and U15464 (N_15464,N_8089,N_5405);
xor U15465 (N_15465,N_7961,N_6854);
or U15466 (N_15466,N_3500,N_6891);
and U15467 (N_15467,N_7330,N_9336);
nor U15468 (N_15468,N_5024,N_8737);
or U15469 (N_15469,N_1992,N_6966);
nor U15470 (N_15470,N_7730,N_506);
nand U15471 (N_15471,N_5176,N_3393);
xor U15472 (N_15472,N_7897,N_6900);
or U15473 (N_15473,N_4263,N_2214);
xor U15474 (N_15474,N_4665,N_4337);
nor U15475 (N_15475,N_4645,N_5176);
nor U15476 (N_15476,N_925,N_5309);
nand U15477 (N_15477,N_8477,N_8372);
nor U15478 (N_15478,N_2380,N_7904);
and U15479 (N_15479,N_6684,N_4453);
nor U15480 (N_15480,N_3665,N_3978);
or U15481 (N_15481,N_9118,N_5110);
nor U15482 (N_15482,N_194,N_2548);
nor U15483 (N_15483,N_1092,N_1436);
or U15484 (N_15484,N_5824,N_3221);
or U15485 (N_15485,N_6273,N_6565);
nand U15486 (N_15486,N_3245,N_9013);
nand U15487 (N_15487,N_1674,N_4234);
nor U15488 (N_15488,N_7590,N_5743);
nor U15489 (N_15489,N_3460,N_2264);
or U15490 (N_15490,N_9399,N_3509);
and U15491 (N_15491,N_2487,N_3389);
nor U15492 (N_15492,N_2884,N_7360);
nand U15493 (N_15493,N_7005,N_8023);
nand U15494 (N_15494,N_5294,N_4925);
nor U15495 (N_15495,N_7420,N_8972);
and U15496 (N_15496,N_3081,N_3641);
xnor U15497 (N_15497,N_510,N_6751);
nor U15498 (N_15498,N_3956,N_3369);
nand U15499 (N_15499,N_8575,N_2267);
nor U15500 (N_15500,N_7674,N_5909);
or U15501 (N_15501,N_4376,N_7415);
and U15502 (N_15502,N_1995,N_164);
nand U15503 (N_15503,N_4802,N_3532);
nor U15504 (N_15504,N_3653,N_4655);
nand U15505 (N_15505,N_1216,N_3624);
nand U15506 (N_15506,N_5327,N_1820);
nor U15507 (N_15507,N_3074,N_2658);
nand U15508 (N_15508,N_3652,N_4647);
nor U15509 (N_15509,N_5866,N_215);
nor U15510 (N_15510,N_7499,N_4276);
nand U15511 (N_15511,N_8922,N_142);
nor U15512 (N_15512,N_8933,N_8542);
or U15513 (N_15513,N_9699,N_4799);
or U15514 (N_15514,N_8392,N_9884);
or U15515 (N_15515,N_9220,N_7179);
nor U15516 (N_15516,N_6613,N_2149);
nor U15517 (N_15517,N_6409,N_4032);
and U15518 (N_15518,N_541,N_7026);
xnor U15519 (N_15519,N_2163,N_9802);
and U15520 (N_15520,N_2109,N_1885);
xor U15521 (N_15521,N_8187,N_8070);
nor U15522 (N_15522,N_2082,N_6667);
or U15523 (N_15523,N_2429,N_3760);
and U15524 (N_15524,N_9657,N_3092);
nand U15525 (N_15525,N_1747,N_3981);
nor U15526 (N_15526,N_5753,N_1348);
nor U15527 (N_15527,N_7359,N_4218);
and U15528 (N_15528,N_3222,N_3832);
nand U15529 (N_15529,N_8233,N_9338);
nand U15530 (N_15530,N_3327,N_6880);
nand U15531 (N_15531,N_7366,N_6394);
nor U15532 (N_15532,N_4435,N_6428);
or U15533 (N_15533,N_71,N_1194);
and U15534 (N_15534,N_1895,N_4015);
nand U15535 (N_15535,N_3656,N_1911);
or U15536 (N_15536,N_3152,N_6451);
nand U15537 (N_15537,N_2885,N_6539);
nor U15538 (N_15538,N_3059,N_6669);
xor U15539 (N_15539,N_3879,N_2638);
nand U15540 (N_15540,N_2871,N_9700);
nor U15541 (N_15541,N_5562,N_6494);
and U15542 (N_15542,N_5709,N_4263);
and U15543 (N_15543,N_5202,N_1722);
nand U15544 (N_15544,N_9833,N_3970);
nor U15545 (N_15545,N_7100,N_1180);
nand U15546 (N_15546,N_7688,N_9684);
or U15547 (N_15547,N_7344,N_832);
or U15548 (N_15548,N_1502,N_9465);
or U15549 (N_15549,N_9571,N_6563);
xor U15550 (N_15550,N_7193,N_7369);
and U15551 (N_15551,N_2522,N_3155);
and U15552 (N_15552,N_6027,N_8196);
and U15553 (N_15553,N_390,N_1007);
or U15554 (N_15554,N_5136,N_2869);
and U15555 (N_15555,N_7169,N_5420);
nand U15556 (N_15556,N_7665,N_5820);
nor U15557 (N_15557,N_2609,N_6735);
or U15558 (N_15558,N_9553,N_946);
and U15559 (N_15559,N_858,N_2611);
or U15560 (N_15560,N_5106,N_6821);
and U15561 (N_15561,N_7321,N_6521);
nor U15562 (N_15562,N_6130,N_8011);
or U15563 (N_15563,N_9741,N_5854);
xor U15564 (N_15564,N_2263,N_5779);
nand U15565 (N_15565,N_6785,N_4542);
nand U15566 (N_15566,N_9372,N_5117);
or U15567 (N_15567,N_8671,N_9135);
or U15568 (N_15568,N_4699,N_275);
nand U15569 (N_15569,N_9798,N_9165);
and U15570 (N_15570,N_6285,N_6843);
nor U15571 (N_15571,N_6301,N_4057);
xnor U15572 (N_15572,N_9232,N_7888);
or U15573 (N_15573,N_5942,N_3607);
and U15574 (N_15574,N_8473,N_4773);
or U15575 (N_15575,N_770,N_169);
xor U15576 (N_15576,N_7129,N_4028);
nor U15577 (N_15577,N_3697,N_4514);
nor U15578 (N_15578,N_1297,N_6018);
nand U15579 (N_15579,N_4053,N_2506);
nor U15580 (N_15580,N_8363,N_1789);
nand U15581 (N_15581,N_5432,N_4444);
nor U15582 (N_15582,N_1233,N_8044);
xnor U15583 (N_15583,N_9571,N_9626);
nor U15584 (N_15584,N_7474,N_4919);
or U15585 (N_15585,N_7124,N_37);
nor U15586 (N_15586,N_8738,N_958);
and U15587 (N_15587,N_4105,N_1427);
nor U15588 (N_15588,N_8822,N_3433);
and U15589 (N_15589,N_4552,N_2244);
and U15590 (N_15590,N_898,N_711);
xnor U15591 (N_15591,N_4257,N_144);
and U15592 (N_15592,N_8821,N_3954);
nand U15593 (N_15593,N_3790,N_2071);
nor U15594 (N_15594,N_7320,N_5946);
nor U15595 (N_15595,N_5337,N_9382);
nor U15596 (N_15596,N_9475,N_2522);
and U15597 (N_15597,N_9258,N_7209);
nor U15598 (N_15598,N_4547,N_7892);
and U15599 (N_15599,N_6529,N_8634);
and U15600 (N_15600,N_8839,N_4459);
nor U15601 (N_15601,N_3522,N_377);
nand U15602 (N_15602,N_8827,N_3116);
xnor U15603 (N_15603,N_6550,N_5248);
or U15604 (N_15604,N_9613,N_332);
and U15605 (N_15605,N_4982,N_3514);
nand U15606 (N_15606,N_5671,N_3206);
and U15607 (N_15607,N_3335,N_2493);
nand U15608 (N_15608,N_4736,N_6276);
or U15609 (N_15609,N_3178,N_8997);
nor U15610 (N_15610,N_4549,N_6951);
or U15611 (N_15611,N_9053,N_1521);
or U15612 (N_15612,N_4279,N_9699);
nand U15613 (N_15613,N_604,N_4703);
nor U15614 (N_15614,N_5144,N_9006);
nand U15615 (N_15615,N_4772,N_5374);
xor U15616 (N_15616,N_3101,N_6078);
and U15617 (N_15617,N_5400,N_9240);
nand U15618 (N_15618,N_387,N_5209);
and U15619 (N_15619,N_9020,N_2269);
and U15620 (N_15620,N_2335,N_8210);
nand U15621 (N_15621,N_5638,N_3446);
nand U15622 (N_15622,N_5230,N_4853);
nor U15623 (N_15623,N_1521,N_1552);
nor U15624 (N_15624,N_9123,N_9896);
or U15625 (N_15625,N_5781,N_3679);
and U15626 (N_15626,N_8631,N_3938);
nand U15627 (N_15627,N_161,N_2112);
nand U15628 (N_15628,N_1724,N_3132);
nand U15629 (N_15629,N_97,N_5196);
and U15630 (N_15630,N_7156,N_5286);
or U15631 (N_15631,N_5317,N_2670);
or U15632 (N_15632,N_5827,N_3723);
and U15633 (N_15633,N_8735,N_9476);
and U15634 (N_15634,N_3336,N_4946);
or U15635 (N_15635,N_1959,N_5946);
xor U15636 (N_15636,N_6866,N_4573);
and U15637 (N_15637,N_5406,N_1642);
or U15638 (N_15638,N_3374,N_542);
nand U15639 (N_15639,N_529,N_8130);
nand U15640 (N_15640,N_948,N_2740);
nor U15641 (N_15641,N_2014,N_9250);
or U15642 (N_15642,N_6463,N_2796);
nor U15643 (N_15643,N_9378,N_651);
nand U15644 (N_15644,N_4296,N_9448);
nand U15645 (N_15645,N_3820,N_498);
or U15646 (N_15646,N_7027,N_5861);
or U15647 (N_15647,N_2619,N_5756);
xor U15648 (N_15648,N_108,N_6510);
nand U15649 (N_15649,N_2668,N_4958);
and U15650 (N_15650,N_1750,N_4365);
nand U15651 (N_15651,N_1595,N_1132);
nor U15652 (N_15652,N_19,N_5269);
nand U15653 (N_15653,N_7059,N_5650);
xnor U15654 (N_15654,N_2651,N_6018);
nor U15655 (N_15655,N_7365,N_4947);
xor U15656 (N_15656,N_6119,N_9778);
nand U15657 (N_15657,N_2551,N_3123);
xnor U15658 (N_15658,N_6312,N_5530);
nor U15659 (N_15659,N_9289,N_7338);
nand U15660 (N_15660,N_3964,N_7074);
nand U15661 (N_15661,N_5422,N_8499);
nor U15662 (N_15662,N_1073,N_2550);
nor U15663 (N_15663,N_4951,N_6544);
nand U15664 (N_15664,N_1362,N_343);
nand U15665 (N_15665,N_3322,N_693);
or U15666 (N_15666,N_1921,N_4775);
and U15667 (N_15667,N_1812,N_6877);
xor U15668 (N_15668,N_3172,N_3030);
nand U15669 (N_15669,N_3110,N_3706);
nand U15670 (N_15670,N_761,N_8053);
or U15671 (N_15671,N_5691,N_9416);
nand U15672 (N_15672,N_668,N_9915);
or U15673 (N_15673,N_1405,N_658);
nand U15674 (N_15674,N_529,N_9156);
nand U15675 (N_15675,N_1556,N_1299);
or U15676 (N_15676,N_5873,N_7675);
nor U15677 (N_15677,N_6924,N_7228);
nand U15678 (N_15678,N_8574,N_5217);
and U15679 (N_15679,N_4866,N_7033);
nor U15680 (N_15680,N_1005,N_2623);
or U15681 (N_15681,N_7222,N_809);
and U15682 (N_15682,N_6798,N_7528);
and U15683 (N_15683,N_9050,N_3581);
xnor U15684 (N_15684,N_2041,N_7933);
nor U15685 (N_15685,N_3952,N_532);
xnor U15686 (N_15686,N_347,N_1804);
nand U15687 (N_15687,N_7278,N_7165);
nor U15688 (N_15688,N_250,N_1701);
or U15689 (N_15689,N_1724,N_3941);
nand U15690 (N_15690,N_9598,N_85);
nand U15691 (N_15691,N_3809,N_4155);
and U15692 (N_15692,N_5152,N_926);
nand U15693 (N_15693,N_2001,N_5784);
or U15694 (N_15694,N_1672,N_3513);
nor U15695 (N_15695,N_4701,N_9634);
and U15696 (N_15696,N_7199,N_3158);
and U15697 (N_15697,N_9047,N_5311);
nand U15698 (N_15698,N_2939,N_7698);
or U15699 (N_15699,N_9138,N_1520);
nor U15700 (N_15700,N_8133,N_5202);
xor U15701 (N_15701,N_4056,N_4749);
or U15702 (N_15702,N_4770,N_8813);
nor U15703 (N_15703,N_3554,N_794);
nand U15704 (N_15704,N_1780,N_3587);
and U15705 (N_15705,N_5895,N_9350);
nand U15706 (N_15706,N_3167,N_2758);
and U15707 (N_15707,N_5708,N_7099);
and U15708 (N_15708,N_6397,N_5931);
or U15709 (N_15709,N_412,N_610);
and U15710 (N_15710,N_838,N_4080);
and U15711 (N_15711,N_1591,N_4682);
or U15712 (N_15712,N_6468,N_4786);
nor U15713 (N_15713,N_4477,N_5358);
nor U15714 (N_15714,N_4849,N_4962);
or U15715 (N_15715,N_4988,N_1457);
xnor U15716 (N_15716,N_2849,N_1498);
and U15717 (N_15717,N_3929,N_8010);
nand U15718 (N_15718,N_9313,N_611);
nor U15719 (N_15719,N_4881,N_5411);
and U15720 (N_15720,N_4900,N_6960);
or U15721 (N_15721,N_2463,N_4803);
nand U15722 (N_15722,N_5838,N_1610);
xnor U15723 (N_15723,N_4415,N_6295);
or U15724 (N_15724,N_1711,N_8942);
nor U15725 (N_15725,N_8124,N_5829);
and U15726 (N_15726,N_6032,N_5125);
nand U15727 (N_15727,N_3873,N_5365);
and U15728 (N_15728,N_6345,N_243);
nor U15729 (N_15729,N_973,N_3998);
and U15730 (N_15730,N_3260,N_2672);
and U15731 (N_15731,N_7848,N_1637);
or U15732 (N_15732,N_4015,N_7704);
or U15733 (N_15733,N_4819,N_7743);
and U15734 (N_15734,N_5431,N_8186);
xnor U15735 (N_15735,N_8313,N_7284);
and U15736 (N_15736,N_3225,N_3180);
nor U15737 (N_15737,N_4481,N_8597);
and U15738 (N_15738,N_2058,N_1514);
nor U15739 (N_15739,N_6213,N_2668);
and U15740 (N_15740,N_1241,N_2824);
nand U15741 (N_15741,N_7373,N_9372);
nand U15742 (N_15742,N_5019,N_1924);
nand U15743 (N_15743,N_5207,N_9417);
or U15744 (N_15744,N_3904,N_2360);
nor U15745 (N_15745,N_9621,N_8669);
and U15746 (N_15746,N_1655,N_5683);
nor U15747 (N_15747,N_6232,N_6519);
nand U15748 (N_15748,N_2712,N_5319);
nor U15749 (N_15749,N_4949,N_9602);
xnor U15750 (N_15750,N_6670,N_9469);
nand U15751 (N_15751,N_6099,N_8220);
or U15752 (N_15752,N_1063,N_4680);
or U15753 (N_15753,N_9982,N_4149);
or U15754 (N_15754,N_956,N_9066);
and U15755 (N_15755,N_6230,N_7706);
or U15756 (N_15756,N_9860,N_2204);
and U15757 (N_15757,N_7873,N_8672);
or U15758 (N_15758,N_2004,N_6437);
and U15759 (N_15759,N_3227,N_7912);
nand U15760 (N_15760,N_5570,N_7020);
nor U15761 (N_15761,N_6450,N_3145);
nor U15762 (N_15762,N_7372,N_5308);
and U15763 (N_15763,N_245,N_522);
xor U15764 (N_15764,N_1373,N_5375);
or U15765 (N_15765,N_811,N_9995);
nor U15766 (N_15766,N_4539,N_6989);
nand U15767 (N_15767,N_1808,N_341);
and U15768 (N_15768,N_9687,N_2812);
nand U15769 (N_15769,N_4254,N_9503);
or U15770 (N_15770,N_3003,N_5284);
or U15771 (N_15771,N_3476,N_8492);
nor U15772 (N_15772,N_891,N_8352);
and U15773 (N_15773,N_5780,N_5653);
nand U15774 (N_15774,N_6590,N_2298);
or U15775 (N_15775,N_7527,N_7159);
and U15776 (N_15776,N_1559,N_7255);
nand U15777 (N_15777,N_672,N_8592);
or U15778 (N_15778,N_3970,N_3522);
and U15779 (N_15779,N_2273,N_8803);
and U15780 (N_15780,N_8267,N_8790);
xnor U15781 (N_15781,N_9487,N_7256);
nor U15782 (N_15782,N_8534,N_7110);
nor U15783 (N_15783,N_4361,N_8093);
nand U15784 (N_15784,N_399,N_1199);
and U15785 (N_15785,N_1247,N_9818);
xnor U15786 (N_15786,N_7896,N_1746);
and U15787 (N_15787,N_4240,N_2542);
nor U15788 (N_15788,N_8706,N_4171);
and U15789 (N_15789,N_1411,N_2370);
nor U15790 (N_15790,N_4047,N_8122);
xor U15791 (N_15791,N_2803,N_1636);
and U15792 (N_15792,N_6875,N_5887);
and U15793 (N_15793,N_3354,N_6786);
nor U15794 (N_15794,N_1978,N_7557);
nand U15795 (N_15795,N_2628,N_8436);
or U15796 (N_15796,N_7280,N_2127);
and U15797 (N_15797,N_5463,N_894);
xor U15798 (N_15798,N_7228,N_77);
xor U15799 (N_15799,N_6558,N_5431);
nor U15800 (N_15800,N_3152,N_7836);
and U15801 (N_15801,N_987,N_1772);
and U15802 (N_15802,N_7393,N_4494);
nand U15803 (N_15803,N_3105,N_7291);
nor U15804 (N_15804,N_1881,N_9718);
and U15805 (N_15805,N_9475,N_2421);
or U15806 (N_15806,N_3863,N_5240);
nor U15807 (N_15807,N_1358,N_4960);
and U15808 (N_15808,N_9621,N_8703);
nand U15809 (N_15809,N_7655,N_7872);
or U15810 (N_15810,N_4516,N_8537);
nor U15811 (N_15811,N_6136,N_6436);
or U15812 (N_15812,N_3018,N_1271);
nor U15813 (N_15813,N_3491,N_7003);
nor U15814 (N_15814,N_2636,N_8843);
nand U15815 (N_15815,N_4663,N_5802);
nor U15816 (N_15816,N_8093,N_3497);
or U15817 (N_15817,N_9933,N_990);
xnor U15818 (N_15818,N_8491,N_2861);
nor U15819 (N_15819,N_630,N_9504);
nand U15820 (N_15820,N_1308,N_284);
nor U15821 (N_15821,N_6664,N_7126);
xnor U15822 (N_15822,N_9236,N_6599);
and U15823 (N_15823,N_3705,N_2278);
nand U15824 (N_15824,N_1440,N_838);
nand U15825 (N_15825,N_2478,N_8373);
and U15826 (N_15826,N_6575,N_9895);
nor U15827 (N_15827,N_4143,N_4821);
nor U15828 (N_15828,N_3661,N_5867);
nor U15829 (N_15829,N_4370,N_1755);
nor U15830 (N_15830,N_7308,N_8288);
and U15831 (N_15831,N_121,N_6252);
nor U15832 (N_15832,N_4784,N_1106);
nand U15833 (N_15833,N_5324,N_4713);
nand U15834 (N_15834,N_847,N_2663);
nor U15835 (N_15835,N_6552,N_3887);
or U15836 (N_15836,N_8955,N_2694);
nand U15837 (N_15837,N_1888,N_1221);
nand U15838 (N_15838,N_6779,N_310);
and U15839 (N_15839,N_554,N_9711);
and U15840 (N_15840,N_5787,N_9128);
and U15841 (N_15841,N_5273,N_3616);
and U15842 (N_15842,N_6567,N_744);
nor U15843 (N_15843,N_6452,N_3020);
or U15844 (N_15844,N_7407,N_5097);
or U15845 (N_15845,N_2280,N_4431);
and U15846 (N_15846,N_888,N_5955);
xnor U15847 (N_15847,N_1805,N_6094);
and U15848 (N_15848,N_4934,N_6262);
nand U15849 (N_15849,N_597,N_6763);
and U15850 (N_15850,N_7886,N_7755);
and U15851 (N_15851,N_8814,N_3555);
or U15852 (N_15852,N_2571,N_4970);
or U15853 (N_15853,N_7435,N_8778);
or U15854 (N_15854,N_5551,N_2572);
or U15855 (N_15855,N_6016,N_9112);
or U15856 (N_15856,N_4957,N_2923);
nor U15857 (N_15857,N_5257,N_3352);
or U15858 (N_15858,N_2021,N_6380);
xor U15859 (N_15859,N_9445,N_9773);
or U15860 (N_15860,N_2964,N_7436);
and U15861 (N_15861,N_7955,N_2959);
and U15862 (N_15862,N_870,N_293);
or U15863 (N_15863,N_7543,N_1588);
nand U15864 (N_15864,N_7696,N_653);
or U15865 (N_15865,N_4175,N_5525);
and U15866 (N_15866,N_4608,N_3190);
nor U15867 (N_15867,N_2769,N_3891);
nand U15868 (N_15868,N_4763,N_3218);
or U15869 (N_15869,N_2113,N_8680);
nand U15870 (N_15870,N_3139,N_628);
and U15871 (N_15871,N_2969,N_5624);
or U15872 (N_15872,N_4770,N_5483);
or U15873 (N_15873,N_9183,N_3351);
nand U15874 (N_15874,N_9102,N_8193);
or U15875 (N_15875,N_7140,N_6226);
or U15876 (N_15876,N_1280,N_7315);
nand U15877 (N_15877,N_4507,N_5007);
nand U15878 (N_15878,N_8617,N_5904);
nor U15879 (N_15879,N_2248,N_4235);
or U15880 (N_15880,N_1140,N_3945);
nand U15881 (N_15881,N_4254,N_3739);
nor U15882 (N_15882,N_4453,N_4794);
or U15883 (N_15883,N_66,N_3219);
nor U15884 (N_15884,N_1606,N_91);
or U15885 (N_15885,N_5198,N_1485);
and U15886 (N_15886,N_4245,N_6220);
and U15887 (N_15887,N_3662,N_5291);
nor U15888 (N_15888,N_8982,N_764);
nor U15889 (N_15889,N_759,N_6385);
xor U15890 (N_15890,N_934,N_6600);
nor U15891 (N_15891,N_9227,N_1538);
or U15892 (N_15892,N_6909,N_3611);
and U15893 (N_15893,N_3534,N_7550);
nor U15894 (N_15894,N_5517,N_1421);
or U15895 (N_15895,N_4886,N_9126);
and U15896 (N_15896,N_2402,N_7091);
and U15897 (N_15897,N_5125,N_2469);
or U15898 (N_15898,N_2880,N_2654);
nand U15899 (N_15899,N_9942,N_9570);
nor U15900 (N_15900,N_1772,N_3341);
or U15901 (N_15901,N_7558,N_8088);
or U15902 (N_15902,N_2668,N_9646);
nor U15903 (N_15903,N_2599,N_2516);
xor U15904 (N_15904,N_6309,N_8830);
and U15905 (N_15905,N_5099,N_9326);
and U15906 (N_15906,N_9308,N_1183);
and U15907 (N_15907,N_5566,N_3525);
nand U15908 (N_15908,N_8438,N_105);
xor U15909 (N_15909,N_9164,N_6489);
or U15910 (N_15910,N_4361,N_5150);
or U15911 (N_15911,N_3587,N_3762);
nand U15912 (N_15912,N_864,N_4533);
and U15913 (N_15913,N_5071,N_4508);
xor U15914 (N_15914,N_2682,N_9299);
xnor U15915 (N_15915,N_362,N_869);
nand U15916 (N_15916,N_4634,N_6424);
or U15917 (N_15917,N_7005,N_9024);
nand U15918 (N_15918,N_6065,N_263);
and U15919 (N_15919,N_5785,N_9549);
nor U15920 (N_15920,N_7993,N_3136);
nor U15921 (N_15921,N_5402,N_8560);
or U15922 (N_15922,N_3349,N_2958);
and U15923 (N_15923,N_8073,N_4105);
or U15924 (N_15924,N_7622,N_8054);
and U15925 (N_15925,N_4012,N_2713);
xnor U15926 (N_15926,N_3726,N_2450);
nor U15927 (N_15927,N_4374,N_111);
or U15928 (N_15928,N_7779,N_5545);
or U15929 (N_15929,N_4534,N_1575);
nand U15930 (N_15930,N_2296,N_4380);
and U15931 (N_15931,N_1532,N_9648);
xnor U15932 (N_15932,N_7978,N_9778);
and U15933 (N_15933,N_109,N_3886);
nand U15934 (N_15934,N_4355,N_6022);
nand U15935 (N_15935,N_2258,N_3759);
nor U15936 (N_15936,N_697,N_1377);
xnor U15937 (N_15937,N_8370,N_3214);
xnor U15938 (N_15938,N_6672,N_7676);
nand U15939 (N_15939,N_8199,N_8289);
nor U15940 (N_15940,N_2736,N_8220);
and U15941 (N_15941,N_7957,N_3227);
or U15942 (N_15942,N_9422,N_2601);
and U15943 (N_15943,N_9154,N_6238);
nand U15944 (N_15944,N_8117,N_9027);
nor U15945 (N_15945,N_7097,N_6848);
or U15946 (N_15946,N_9692,N_2004);
nor U15947 (N_15947,N_7049,N_5123);
nor U15948 (N_15948,N_6272,N_6337);
and U15949 (N_15949,N_357,N_4173);
nor U15950 (N_15950,N_2294,N_5112);
xor U15951 (N_15951,N_7088,N_8511);
nor U15952 (N_15952,N_7000,N_5629);
xnor U15953 (N_15953,N_4401,N_4422);
and U15954 (N_15954,N_3180,N_5660);
and U15955 (N_15955,N_3112,N_338);
xor U15956 (N_15956,N_4972,N_6246);
and U15957 (N_15957,N_5437,N_9853);
and U15958 (N_15958,N_1341,N_3613);
or U15959 (N_15959,N_5277,N_3089);
nor U15960 (N_15960,N_1099,N_327);
nand U15961 (N_15961,N_5108,N_8255);
and U15962 (N_15962,N_5251,N_9551);
and U15963 (N_15963,N_1660,N_8010);
nor U15964 (N_15964,N_8775,N_8711);
and U15965 (N_15965,N_3388,N_9544);
nand U15966 (N_15966,N_778,N_7161);
nand U15967 (N_15967,N_792,N_4000);
or U15968 (N_15968,N_5235,N_8383);
or U15969 (N_15969,N_7651,N_2894);
nor U15970 (N_15970,N_3675,N_3404);
nand U15971 (N_15971,N_9551,N_6887);
or U15972 (N_15972,N_1973,N_5114);
nand U15973 (N_15973,N_3400,N_6991);
or U15974 (N_15974,N_1620,N_1974);
and U15975 (N_15975,N_7952,N_5022);
and U15976 (N_15976,N_4270,N_9699);
nand U15977 (N_15977,N_5470,N_6943);
and U15978 (N_15978,N_6963,N_4865);
nor U15979 (N_15979,N_5213,N_6541);
and U15980 (N_15980,N_747,N_2220);
nand U15981 (N_15981,N_55,N_1519);
nor U15982 (N_15982,N_6008,N_8171);
nand U15983 (N_15983,N_766,N_2925);
or U15984 (N_15984,N_7805,N_998);
and U15985 (N_15985,N_2701,N_7093);
nor U15986 (N_15986,N_5072,N_5494);
nor U15987 (N_15987,N_4628,N_6384);
and U15988 (N_15988,N_3494,N_3886);
and U15989 (N_15989,N_1081,N_3893);
or U15990 (N_15990,N_3517,N_8712);
nor U15991 (N_15991,N_7323,N_812);
xnor U15992 (N_15992,N_8976,N_6694);
and U15993 (N_15993,N_7282,N_2587);
nor U15994 (N_15994,N_5604,N_1018);
or U15995 (N_15995,N_8199,N_6941);
nor U15996 (N_15996,N_6982,N_9537);
nor U15997 (N_15997,N_7638,N_6874);
nand U15998 (N_15998,N_8544,N_8330);
nor U15999 (N_15999,N_8721,N_466);
xnor U16000 (N_16000,N_718,N_5477);
and U16001 (N_16001,N_3709,N_3976);
or U16002 (N_16002,N_6227,N_4449);
nand U16003 (N_16003,N_1623,N_9595);
nand U16004 (N_16004,N_2663,N_5761);
and U16005 (N_16005,N_3503,N_3073);
nand U16006 (N_16006,N_5244,N_2176);
nor U16007 (N_16007,N_8566,N_7341);
xnor U16008 (N_16008,N_6032,N_779);
or U16009 (N_16009,N_9675,N_839);
nor U16010 (N_16010,N_1243,N_5534);
nand U16011 (N_16011,N_3668,N_7740);
nand U16012 (N_16012,N_8200,N_9168);
nor U16013 (N_16013,N_8793,N_5444);
xnor U16014 (N_16014,N_5367,N_5452);
nor U16015 (N_16015,N_7065,N_8723);
nand U16016 (N_16016,N_6041,N_1726);
or U16017 (N_16017,N_4698,N_2600);
nor U16018 (N_16018,N_5465,N_361);
and U16019 (N_16019,N_7439,N_1500);
xnor U16020 (N_16020,N_5242,N_664);
or U16021 (N_16021,N_3310,N_2341);
or U16022 (N_16022,N_5020,N_8047);
nand U16023 (N_16023,N_8624,N_2854);
and U16024 (N_16024,N_4270,N_9037);
nor U16025 (N_16025,N_7879,N_5742);
and U16026 (N_16026,N_8310,N_5221);
nand U16027 (N_16027,N_3904,N_2953);
nand U16028 (N_16028,N_12,N_5613);
nor U16029 (N_16029,N_4439,N_4450);
or U16030 (N_16030,N_2743,N_3660);
and U16031 (N_16031,N_2195,N_127);
xor U16032 (N_16032,N_5560,N_7604);
nand U16033 (N_16033,N_5715,N_2185);
and U16034 (N_16034,N_2422,N_2706);
or U16035 (N_16035,N_1412,N_6505);
nand U16036 (N_16036,N_5110,N_3310);
nor U16037 (N_16037,N_6353,N_3704);
nand U16038 (N_16038,N_6379,N_5803);
nor U16039 (N_16039,N_2300,N_8606);
nor U16040 (N_16040,N_4755,N_8828);
nand U16041 (N_16041,N_3170,N_2140);
nand U16042 (N_16042,N_8218,N_3807);
nor U16043 (N_16043,N_5948,N_3445);
nand U16044 (N_16044,N_3932,N_9706);
and U16045 (N_16045,N_9668,N_8529);
or U16046 (N_16046,N_9644,N_8807);
nand U16047 (N_16047,N_4158,N_1526);
or U16048 (N_16048,N_6129,N_878);
nand U16049 (N_16049,N_2024,N_2784);
nor U16050 (N_16050,N_5872,N_772);
or U16051 (N_16051,N_4333,N_3785);
or U16052 (N_16052,N_5200,N_9220);
nor U16053 (N_16053,N_8056,N_8471);
or U16054 (N_16054,N_8100,N_8150);
xor U16055 (N_16055,N_8007,N_1204);
xnor U16056 (N_16056,N_6088,N_8861);
or U16057 (N_16057,N_5624,N_8171);
and U16058 (N_16058,N_2611,N_2226);
nand U16059 (N_16059,N_5947,N_1684);
or U16060 (N_16060,N_6515,N_1604);
and U16061 (N_16061,N_8915,N_1929);
and U16062 (N_16062,N_1057,N_2847);
nand U16063 (N_16063,N_1515,N_9283);
or U16064 (N_16064,N_4241,N_4778);
or U16065 (N_16065,N_6687,N_5931);
and U16066 (N_16066,N_8115,N_3757);
nor U16067 (N_16067,N_2045,N_7527);
and U16068 (N_16068,N_7432,N_5215);
nor U16069 (N_16069,N_3386,N_5693);
nor U16070 (N_16070,N_6974,N_9040);
nor U16071 (N_16071,N_1993,N_338);
and U16072 (N_16072,N_8815,N_6859);
nand U16073 (N_16073,N_7554,N_1233);
or U16074 (N_16074,N_6880,N_7690);
nand U16075 (N_16075,N_8226,N_4476);
and U16076 (N_16076,N_3346,N_4186);
and U16077 (N_16077,N_9053,N_8600);
xor U16078 (N_16078,N_10,N_5458);
nand U16079 (N_16079,N_4888,N_7907);
nand U16080 (N_16080,N_518,N_7092);
and U16081 (N_16081,N_5522,N_6420);
and U16082 (N_16082,N_4728,N_5903);
or U16083 (N_16083,N_2479,N_7890);
nand U16084 (N_16084,N_8961,N_1166);
xor U16085 (N_16085,N_9680,N_3352);
nand U16086 (N_16086,N_9021,N_3876);
nand U16087 (N_16087,N_3179,N_1917);
nor U16088 (N_16088,N_3855,N_7080);
or U16089 (N_16089,N_7597,N_2379);
or U16090 (N_16090,N_967,N_8370);
or U16091 (N_16091,N_569,N_2560);
or U16092 (N_16092,N_6532,N_8099);
nand U16093 (N_16093,N_2283,N_7825);
nor U16094 (N_16094,N_8181,N_9844);
nand U16095 (N_16095,N_3989,N_8818);
and U16096 (N_16096,N_2069,N_1152);
nor U16097 (N_16097,N_6840,N_3415);
nor U16098 (N_16098,N_571,N_4249);
xnor U16099 (N_16099,N_3608,N_1302);
nand U16100 (N_16100,N_3534,N_1359);
nor U16101 (N_16101,N_9140,N_3654);
nand U16102 (N_16102,N_1503,N_4653);
or U16103 (N_16103,N_6026,N_1535);
nand U16104 (N_16104,N_5780,N_8123);
nand U16105 (N_16105,N_8431,N_5189);
xnor U16106 (N_16106,N_2112,N_2525);
nand U16107 (N_16107,N_9057,N_6986);
nor U16108 (N_16108,N_6980,N_985);
nor U16109 (N_16109,N_5218,N_9042);
or U16110 (N_16110,N_7831,N_764);
or U16111 (N_16111,N_3724,N_1984);
and U16112 (N_16112,N_4310,N_7888);
or U16113 (N_16113,N_9592,N_8463);
xor U16114 (N_16114,N_7945,N_4630);
or U16115 (N_16115,N_3737,N_7778);
and U16116 (N_16116,N_4361,N_426);
nor U16117 (N_16117,N_1677,N_8415);
nor U16118 (N_16118,N_2747,N_3358);
or U16119 (N_16119,N_7439,N_337);
nor U16120 (N_16120,N_1793,N_2107);
and U16121 (N_16121,N_6167,N_1030);
nand U16122 (N_16122,N_1434,N_8048);
xnor U16123 (N_16123,N_5201,N_9813);
nand U16124 (N_16124,N_2732,N_2616);
nand U16125 (N_16125,N_4981,N_7142);
or U16126 (N_16126,N_5760,N_817);
nand U16127 (N_16127,N_3173,N_9525);
xor U16128 (N_16128,N_7531,N_4310);
nand U16129 (N_16129,N_5295,N_3725);
nand U16130 (N_16130,N_2844,N_4016);
xnor U16131 (N_16131,N_9666,N_7081);
and U16132 (N_16132,N_2459,N_7311);
nor U16133 (N_16133,N_4584,N_5146);
nor U16134 (N_16134,N_8671,N_102);
nor U16135 (N_16135,N_4149,N_6085);
and U16136 (N_16136,N_5877,N_9678);
xor U16137 (N_16137,N_8785,N_814);
and U16138 (N_16138,N_9793,N_1870);
and U16139 (N_16139,N_344,N_8134);
xnor U16140 (N_16140,N_3715,N_1096);
or U16141 (N_16141,N_3768,N_8814);
nand U16142 (N_16142,N_6377,N_7125);
or U16143 (N_16143,N_6048,N_2686);
or U16144 (N_16144,N_8651,N_7575);
and U16145 (N_16145,N_7456,N_6313);
nor U16146 (N_16146,N_7755,N_5121);
nor U16147 (N_16147,N_3621,N_6544);
nor U16148 (N_16148,N_2963,N_9147);
nand U16149 (N_16149,N_2666,N_7169);
xnor U16150 (N_16150,N_1398,N_249);
nor U16151 (N_16151,N_6292,N_5603);
nand U16152 (N_16152,N_6390,N_8105);
nand U16153 (N_16153,N_4043,N_5351);
nor U16154 (N_16154,N_7304,N_2471);
nand U16155 (N_16155,N_8113,N_6990);
and U16156 (N_16156,N_7762,N_2021);
and U16157 (N_16157,N_800,N_1363);
or U16158 (N_16158,N_6381,N_3880);
and U16159 (N_16159,N_2011,N_9303);
nor U16160 (N_16160,N_7972,N_7927);
nand U16161 (N_16161,N_7928,N_1172);
and U16162 (N_16162,N_9186,N_9744);
and U16163 (N_16163,N_6184,N_4220);
nor U16164 (N_16164,N_3628,N_3270);
nand U16165 (N_16165,N_2238,N_2245);
nand U16166 (N_16166,N_7470,N_1673);
nor U16167 (N_16167,N_2920,N_2987);
nand U16168 (N_16168,N_6595,N_8989);
and U16169 (N_16169,N_2724,N_9981);
nand U16170 (N_16170,N_5264,N_5189);
nand U16171 (N_16171,N_5389,N_6608);
or U16172 (N_16172,N_7825,N_7966);
nand U16173 (N_16173,N_7601,N_2092);
or U16174 (N_16174,N_2794,N_2306);
and U16175 (N_16175,N_2640,N_2036);
nand U16176 (N_16176,N_1410,N_7358);
and U16177 (N_16177,N_1232,N_9161);
nand U16178 (N_16178,N_5041,N_7221);
or U16179 (N_16179,N_6132,N_5173);
nor U16180 (N_16180,N_1478,N_3888);
nand U16181 (N_16181,N_8426,N_1462);
or U16182 (N_16182,N_94,N_939);
or U16183 (N_16183,N_9851,N_658);
or U16184 (N_16184,N_7540,N_2004);
nor U16185 (N_16185,N_8798,N_7375);
and U16186 (N_16186,N_6057,N_4234);
nand U16187 (N_16187,N_196,N_2630);
nand U16188 (N_16188,N_7133,N_4867);
and U16189 (N_16189,N_8777,N_176);
or U16190 (N_16190,N_9378,N_8982);
and U16191 (N_16191,N_5929,N_9774);
nor U16192 (N_16192,N_3993,N_8320);
and U16193 (N_16193,N_38,N_3615);
and U16194 (N_16194,N_9483,N_8086);
nor U16195 (N_16195,N_2948,N_4375);
nand U16196 (N_16196,N_6230,N_4838);
nor U16197 (N_16197,N_8309,N_947);
nand U16198 (N_16198,N_4305,N_1497);
nor U16199 (N_16199,N_430,N_8699);
or U16200 (N_16200,N_472,N_21);
and U16201 (N_16201,N_6515,N_3551);
nand U16202 (N_16202,N_9309,N_3366);
or U16203 (N_16203,N_6234,N_4542);
or U16204 (N_16204,N_7400,N_8203);
nor U16205 (N_16205,N_4517,N_5087);
nor U16206 (N_16206,N_5342,N_23);
or U16207 (N_16207,N_5062,N_4537);
or U16208 (N_16208,N_9679,N_6082);
nor U16209 (N_16209,N_2339,N_5616);
nand U16210 (N_16210,N_9263,N_3191);
and U16211 (N_16211,N_6833,N_7759);
xor U16212 (N_16212,N_1064,N_4219);
and U16213 (N_16213,N_9972,N_537);
nor U16214 (N_16214,N_3865,N_2114);
and U16215 (N_16215,N_9312,N_6234);
nand U16216 (N_16216,N_4928,N_3532);
nor U16217 (N_16217,N_3973,N_195);
nor U16218 (N_16218,N_5865,N_8422);
nand U16219 (N_16219,N_1956,N_8938);
and U16220 (N_16220,N_5835,N_9628);
or U16221 (N_16221,N_3828,N_7696);
nor U16222 (N_16222,N_890,N_9404);
and U16223 (N_16223,N_6107,N_1189);
nand U16224 (N_16224,N_9683,N_2764);
xnor U16225 (N_16225,N_9337,N_2675);
or U16226 (N_16226,N_6586,N_341);
or U16227 (N_16227,N_7045,N_4420);
or U16228 (N_16228,N_9504,N_1534);
nand U16229 (N_16229,N_8846,N_2596);
or U16230 (N_16230,N_4671,N_4253);
nand U16231 (N_16231,N_7488,N_3367);
or U16232 (N_16232,N_5342,N_3316);
nand U16233 (N_16233,N_8004,N_7697);
nand U16234 (N_16234,N_901,N_2625);
or U16235 (N_16235,N_1126,N_2068);
nand U16236 (N_16236,N_9617,N_263);
or U16237 (N_16237,N_4852,N_4346);
or U16238 (N_16238,N_8204,N_9502);
and U16239 (N_16239,N_7945,N_2315);
nor U16240 (N_16240,N_7657,N_2531);
and U16241 (N_16241,N_7294,N_1157);
nor U16242 (N_16242,N_9602,N_8220);
nor U16243 (N_16243,N_6791,N_3608);
nand U16244 (N_16244,N_9438,N_7291);
nand U16245 (N_16245,N_8144,N_425);
and U16246 (N_16246,N_9494,N_1784);
nand U16247 (N_16247,N_5721,N_4905);
and U16248 (N_16248,N_4740,N_946);
nor U16249 (N_16249,N_7236,N_273);
nand U16250 (N_16250,N_9978,N_5279);
nand U16251 (N_16251,N_4574,N_153);
nor U16252 (N_16252,N_7863,N_6185);
and U16253 (N_16253,N_7541,N_329);
nor U16254 (N_16254,N_8385,N_7086);
nand U16255 (N_16255,N_8872,N_2449);
nor U16256 (N_16256,N_6079,N_7546);
or U16257 (N_16257,N_1079,N_6202);
nor U16258 (N_16258,N_8742,N_6801);
and U16259 (N_16259,N_1330,N_6577);
and U16260 (N_16260,N_6669,N_1028);
nand U16261 (N_16261,N_4563,N_9627);
and U16262 (N_16262,N_6030,N_6356);
nand U16263 (N_16263,N_9360,N_8727);
nand U16264 (N_16264,N_8805,N_827);
nor U16265 (N_16265,N_6415,N_4331);
xor U16266 (N_16266,N_8988,N_800);
and U16267 (N_16267,N_9574,N_7538);
xor U16268 (N_16268,N_6705,N_7234);
xnor U16269 (N_16269,N_7500,N_4719);
and U16270 (N_16270,N_3601,N_1124);
nor U16271 (N_16271,N_5026,N_1596);
nand U16272 (N_16272,N_3377,N_3325);
or U16273 (N_16273,N_2044,N_5624);
nor U16274 (N_16274,N_4302,N_7112);
nor U16275 (N_16275,N_4907,N_6255);
and U16276 (N_16276,N_8694,N_5458);
and U16277 (N_16277,N_1280,N_5425);
nand U16278 (N_16278,N_5791,N_1240);
and U16279 (N_16279,N_434,N_4077);
and U16280 (N_16280,N_4590,N_7670);
nand U16281 (N_16281,N_8892,N_8135);
and U16282 (N_16282,N_6784,N_2379);
or U16283 (N_16283,N_8130,N_7495);
nand U16284 (N_16284,N_5410,N_1062);
or U16285 (N_16285,N_3459,N_7655);
and U16286 (N_16286,N_3558,N_3716);
nand U16287 (N_16287,N_7459,N_4244);
nor U16288 (N_16288,N_5783,N_6637);
and U16289 (N_16289,N_1482,N_8369);
nor U16290 (N_16290,N_1599,N_2452);
or U16291 (N_16291,N_7755,N_1480);
and U16292 (N_16292,N_8659,N_5669);
or U16293 (N_16293,N_8921,N_9142);
nand U16294 (N_16294,N_6087,N_4051);
nand U16295 (N_16295,N_1612,N_345);
and U16296 (N_16296,N_4078,N_7870);
nand U16297 (N_16297,N_365,N_2603);
and U16298 (N_16298,N_5712,N_6974);
or U16299 (N_16299,N_788,N_6843);
and U16300 (N_16300,N_9581,N_9453);
nor U16301 (N_16301,N_487,N_9834);
or U16302 (N_16302,N_1369,N_9252);
xnor U16303 (N_16303,N_866,N_909);
or U16304 (N_16304,N_8616,N_2383);
or U16305 (N_16305,N_2740,N_7301);
nor U16306 (N_16306,N_6432,N_5922);
and U16307 (N_16307,N_4878,N_6115);
and U16308 (N_16308,N_4301,N_3559);
nand U16309 (N_16309,N_1183,N_5464);
xnor U16310 (N_16310,N_2420,N_8856);
and U16311 (N_16311,N_9121,N_3385);
nand U16312 (N_16312,N_9927,N_7363);
nand U16313 (N_16313,N_1918,N_2529);
nor U16314 (N_16314,N_1733,N_5524);
xnor U16315 (N_16315,N_2750,N_677);
or U16316 (N_16316,N_3505,N_9503);
xor U16317 (N_16317,N_3296,N_1290);
nand U16318 (N_16318,N_9806,N_3083);
nor U16319 (N_16319,N_7783,N_1080);
or U16320 (N_16320,N_7246,N_320);
and U16321 (N_16321,N_3809,N_4973);
and U16322 (N_16322,N_9305,N_1568);
nor U16323 (N_16323,N_3589,N_8919);
or U16324 (N_16324,N_8493,N_4726);
nand U16325 (N_16325,N_8572,N_2561);
nor U16326 (N_16326,N_2975,N_5481);
nor U16327 (N_16327,N_263,N_2350);
or U16328 (N_16328,N_7379,N_9473);
and U16329 (N_16329,N_8065,N_1714);
nand U16330 (N_16330,N_2650,N_128);
nor U16331 (N_16331,N_8481,N_3045);
or U16332 (N_16332,N_2256,N_9937);
nor U16333 (N_16333,N_128,N_4881);
xnor U16334 (N_16334,N_2012,N_8137);
or U16335 (N_16335,N_6789,N_456);
and U16336 (N_16336,N_5161,N_9936);
and U16337 (N_16337,N_894,N_1799);
nand U16338 (N_16338,N_336,N_1949);
nor U16339 (N_16339,N_4048,N_5851);
nor U16340 (N_16340,N_3144,N_268);
nor U16341 (N_16341,N_7843,N_6733);
or U16342 (N_16342,N_3433,N_6457);
or U16343 (N_16343,N_4013,N_8816);
nor U16344 (N_16344,N_5097,N_1818);
and U16345 (N_16345,N_1823,N_9660);
xnor U16346 (N_16346,N_3733,N_8335);
nor U16347 (N_16347,N_5573,N_5087);
nor U16348 (N_16348,N_9245,N_1965);
nand U16349 (N_16349,N_1787,N_3340);
or U16350 (N_16350,N_6749,N_5727);
and U16351 (N_16351,N_1994,N_591);
nand U16352 (N_16352,N_1837,N_252);
nor U16353 (N_16353,N_9226,N_6480);
or U16354 (N_16354,N_2016,N_5418);
or U16355 (N_16355,N_2813,N_250);
or U16356 (N_16356,N_7937,N_8359);
and U16357 (N_16357,N_1199,N_9017);
and U16358 (N_16358,N_8558,N_6664);
or U16359 (N_16359,N_5006,N_348);
nand U16360 (N_16360,N_4270,N_8848);
nor U16361 (N_16361,N_4824,N_2770);
nor U16362 (N_16362,N_6470,N_9614);
nand U16363 (N_16363,N_82,N_2681);
or U16364 (N_16364,N_5407,N_5785);
xnor U16365 (N_16365,N_884,N_553);
nor U16366 (N_16366,N_1645,N_7481);
and U16367 (N_16367,N_9288,N_4980);
and U16368 (N_16368,N_4126,N_8975);
nand U16369 (N_16369,N_1486,N_450);
nand U16370 (N_16370,N_5021,N_6226);
or U16371 (N_16371,N_7124,N_9881);
or U16372 (N_16372,N_8308,N_2470);
nand U16373 (N_16373,N_966,N_9939);
and U16374 (N_16374,N_1200,N_1967);
or U16375 (N_16375,N_7730,N_1180);
nor U16376 (N_16376,N_7204,N_6578);
and U16377 (N_16377,N_257,N_6881);
nor U16378 (N_16378,N_2040,N_3441);
nor U16379 (N_16379,N_449,N_5641);
nand U16380 (N_16380,N_600,N_5854);
or U16381 (N_16381,N_8855,N_8440);
nor U16382 (N_16382,N_9259,N_6842);
nor U16383 (N_16383,N_9444,N_9288);
nand U16384 (N_16384,N_849,N_7488);
nor U16385 (N_16385,N_9414,N_3060);
or U16386 (N_16386,N_9892,N_7443);
nor U16387 (N_16387,N_5392,N_838);
or U16388 (N_16388,N_8645,N_8321);
and U16389 (N_16389,N_9390,N_7066);
nor U16390 (N_16390,N_5462,N_1212);
and U16391 (N_16391,N_3105,N_7731);
or U16392 (N_16392,N_3292,N_556);
nand U16393 (N_16393,N_9655,N_5173);
nand U16394 (N_16394,N_7522,N_1671);
and U16395 (N_16395,N_2691,N_6493);
and U16396 (N_16396,N_9982,N_5372);
and U16397 (N_16397,N_9594,N_6169);
nor U16398 (N_16398,N_2166,N_7424);
or U16399 (N_16399,N_6987,N_2246);
xnor U16400 (N_16400,N_5360,N_7484);
and U16401 (N_16401,N_6525,N_684);
and U16402 (N_16402,N_6237,N_1753);
nand U16403 (N_16403,N_9343,N_9166);
or U16404 (N_16404,N_1041,N_4356);
and U16405 (N_16405,N_4721,N_9860);
nor U16406 (N_16406,N_3062,N_6951);
xor U16407 (N_16407,N_2164,N_8265);
nand U16408 (N_16408,N_9985,N_8749);
nand U16409 (N_16409,N_8818,N_2655);
or U16410 (N_16410,N_9766,N_4035);
nand U16411 (N_16411,N_4456,N_2956);
nand U16412 (N_16412,N_9062,N_3235);
nor U16413 (N_16413,N_2607,N_5100);
or U16414 (N_16414,N_7334,N_1648);
nor U16415 (N_16415,N_6451,N_4084);
or U16416 (N_16416,N_2184,N_6437);
and U16417 (N_16417,N_9575,N_6291);
or U16418 (N_16418,N_7714,N_4244);
nand U16419 (N_16419,N_7067,N_4834);
nor U16420 (N_16420,N_8397,N_8071);
or U16421 (N_16421,N_4198,N_2992);
and U16422 (N_16422,N_3937,N_5896);
or U16423 (N_16423,N_3569,N_6134);
or U16424 (N_16424,N_1056,N_2105);
and U16425 (N_16425,N_6585,N_9584);
or U16426 (N_16426,N_1160,N_4864);
and U16427 (N_16427,N_5564,N_3278);
xor U16428 (N_16428,N_4845,N_2801);
nor U16429 (N_16429,N_1593,N_6251);
nor U16430 (N_16430,N_3586,N_7679);
nor U16431 (N_16431,N_7479,N_6553);
and U16432 (N_16432,N_6842,N_6785);
or U16433 (N_16433,N_444,N_845);
nor U16434 (N_16434,N_835,N_635);
xor U16435 (N_16435,N_5597,N_8170);
nand U16436 (N_16436,N_2876,N_7264);
and U16437 (N_16437,N_7096,N_1403);
nor U16438 (N_16438,N_2765,N_1544);
nand U16439 (N_16439,N_1819,N_7984);
and U16440 (N_16440,N_9350,N_7312);
xor U16441 (N_16441,N_7355,N_8298);
or U16442 (N_16442,N_3158,N_4268);
nand U16443 (N_16443,N_8281,N_6230);
or U16444 (N_16444,N_4279,N_9803);
and U16445 (N_16445,N_2789,N_5391);
nor U16446 (N_16446,N_3181,N_9841);
nand U16447 (N_16447,N_7760,N_7958);
or U16448 (N_16448,N_3343,N_2742);
nand U16449 (N_16449,N_6477,N_5441);
nand U16450 (N_16450,N_9956,N_8622);
nand U16451 (N_16451,N_3213,N_4784);
nand U16452 (N_16452,N_748,N_7212);
nor U16453 (N_16453,N_3595,N_44);
and U16454 (N_16454,N_5454,N_552);
nor U16455 (N_16455,N_52,N_1008);
or U16456 (N_16456,N_6771,N_1111);
and U16457 (N_16457,N_6633,N_2989);
nor U16458 (N_16458,N_1850,N_3126);
or U16459 (N_16459,N_7397,N_2599);
and U16460 (N_16460,N_8821,N_9391);
nor U16461 (N_16461,N_1619,N_7803);
and U16462 (N_16462,N_1321,N_9191);
xnor U16463 (N_16463,N_54,N_6295);
or U16464 (N_16464,N_3062,N_5998);
nor U16465 (N_16465,N_4041,N_2150);
nor U16466 (N_16466,N_1247,N_875);
and U16467 (N_16467,N_5429,N_4141);
or U16468 (N_16468,N_1467,N_7034);
or U16469 (N_16469,N_1193,N_5601);
nand U16470 (N_16470,N_5477,N_2146);
nor U16471 (N_16471,N_6450,N_5918);
nand U16472 (N_16472,N_4635,N_2726);
xor U16473 (N_16473,N_6537,N_9047);
and U16474 (N_16474,N_6081,N_6116);
nand U16475 (N_16475,N_1715,N_2841);
or U16476 (N_16476,N_5619,N_3247);
nand U16477 (N_16477,N_1665,N_7464);
or U16478 (N_16478,N_6383,N_2002);
nor U16479 (N_16479,N_3953,N_7719);
nor U16480 (N_16480,N_4271,N_1414);
and U16481 (N_16481,N_8177,N_6128);
and U16482 (N_16482,N_360,N_8350);
and U16483 (N_16483,N_4479,N_8965);
and U16484 (N_16484,N_1361,N_3695);
nor U16485 (N_16485,N_2838,N_3571);
or U16486 (N_16486,N_7183,N_3320);
xor U16487 (N_16487,N_667,N_9428);
xor U16488 (N_16488,N_4388,N_9492);
nor U16489 (N_16489,N_7876,N_3790);
or U16490 (N_16490,N_4813,N_3537);
nand U16491 (N_16491,N_5659,N_8862);
and U16492 (N_16492,N_2796,N_1536);
xnor U16493 (N_16493,N_3100,N_4343);
and U16494 (N_16494,N_9767,N_666);
and U16495 (N_16495,N_9067,N_9490);
nor U16496 (N_16496,N_4256,N_7527);
and U16497 (N_16497,N_5192,N_7195);
xnor U16498 (N_16498,N_6147,N_2382);
nand U16499 (N_16499,N_9983,N_6833);
or U16500 (N_16500,N_8127,N_6779);
nor U16501 (N_16501,N_6293,N_1937);
or U16502 (N_16502,N_688,N_4109);
and U16503 (N_16503,N_1557,N_4466);
nor U16504 (N_16504,N_96,N_1197);
nand U16505 (N_16505,N_4586,N_6502);
nand U16506 (N_16506,N_4908,N_7647);
or U16507 (N_16507,N_651,N_8402);
nand U16508 (N_16508,N_7333,N_8858);
and U16509 (N_16509,N_1787,N_1003);
nand U16510 (N_16510,N_9724,N_7103);
nor U16511 (N_16511,N_6406,N_5715);
or U16512 (N_16512,N_9203,N_3071);
xor U16513 (N_16513,N_3333,N_7020);
nor U16514 (N_16514,N_5443,N_773);
and U16515 (N_16515,N_5222,N_3907);
nor U16516 (N_16516,N_1918,N_4844);
xnor U16517 (N_16517,N_8535,N_2959);
or U16518 (N_16518,N_5591,N_2715);
nand U16519 (N_16519,N_5732,N_3868);
and U16520 (N_16520,N_6119,N_1222);
nor U16521 (N_16521,N_7475,N_9115);
nor U16522 (N_16522,N_5009,N_524);
or U16523 (N_16523,N_4342,N_5556);
xor U16524 (N_16524,N_6350,N_8054);
nor U16525 (N_16525,N_2217,N_6910);
nand U16526 (N_16526,N_4669,N_1912);
nand U16527 (N_16527,N_3663,N_8661);
xnor U16528 (N_16528,N_1824,N_6207);
and U16529 (N_16529,N_5714,N_1096);
and U16530 (N_16530,N_2686,N_2127);
and U16531 (N_16531,N_7570,N_253);
nor U16532 (N_16532,N_7991,N_4273);
or U16533 (N_16533,N_8603,N_887);
nor U16534 (N_16534,N_3699,N_8656);
or U16535 (N_16535,N_1276,N_4799);
nor U16536 (N_16536,N_2292,N_5652);
or U16537 (N_16537,N_3581,N_9276);
nand U16538 (N_16538,N_187,N_581);
nor U16539 (N_16539,N_810,N_727);
nor U16540 (N_16540,N_4905,N_4996);
nor U16541 (N_16541,N_5579,N_3278);
or U16542 (N_16542,N_4071,N_4672);
xor U16543 (N_16543,N_202,N_3364);
nand U16544 (N_16544,N_4026,N_8075);
nor U16545 (N_16545,N_9580,N_3958);
and U16546 (N_16546,N_1447,N_1445);
nor U16547 (N_16547,N_7349,N_8436);
nand U16548 (N_16548,N_6213,N_5636);
nor U16549 (N_16549,N_8708,N_3220);
or U16550 (N_16550,N_6755,N_2770);
or U16551 (N_16551,N_8953,N_5249);
nor U16552 (N_16552,N_2143,N_6084);
nand U16553 (N_16553,N_1482,N_8790);
xnor U16554 (N_16554,N_3251,N_1304);
nor U16555 (N_16555,N_2226,N_7356);
nor U16556 (N_16556,N_2890,N_6233);
nor U16557 (N_16557,N_7318,N_675);
xnor U16558 (N_16558,N_1418,N_3130);
xnor U16559 (N_16559,N_1860,N_2657);
or U16560 (N_16560,N_1671,N_5943);
nor U16561 (N_16561,N_6373,N_9948);
or U16562 (N_16562,N_9210,N_865);
xnor U16563 (N_16563,N_96,N_3909);
and U16564 (N_16564,N_4023,N_4479);
or U16565 (N_16565,N_8921,N_1859);
and U16566 (N_16566,N_4271,N_2421);
or U16567 (N_16567,N_4394,N_4612);
nor U16568 (N_16568,N_523,N_5671);
or U16569 (N_16569,N_3247,N_4194);
nand U16570 (N_16570,N_8106,N_4457);
and U16571 (N_16571,N_3271,N_6793);
or U16572 (N_16572,N_1805,N_6864);
and U16573 (N_16573,N_9293,N_9737);
nor U16574 (N_16574,N_3240,N_4003);
and U16575 (N_16575,N_4867,N_1830);
nand U16576 (N_16576,N_9430,N_6899);
xor U16577 (N_16577,N_9917,N_929);
nor U16578 (N_16578,N_4944,N_2192);
or U16579 (N_16579,N_2081,N_9510);
nand U16580 (N_16580,N_1071,N_8565);
nor U16581 (N_16581,N_2155,N_5009);
nand U16582 (N_16582,N_2334,N_441);
nor U16583 (N_16583,N_4236,N_7919);
and U16584 (N_16584,N_9736,N_926);
nor U16585 (N_16585,N_7168,N_3369);
or U16586 (N_16586,N_6689,N_2836);
xor U16587 (N_16587,N_8823,N_3628);
and U16588 (N_16588,N_6576,N_9414);
or U16589 (N_16589,N_5442,N_8381);
xor U16590 (N_16590,N_5584,N_3318);
nand U16591 (N_16591,N_4646,N_1221);
nand U16592 (N_16592,N_7756,N_1256);
or U16593 (N_16593,N_2828,N_7181);
and U16594 (N_16594,N_7725,N_6040);
nor U16595 (N_16595,N_2924,N_4764);
nand U16596 (N_16596,N_8288,N_30);
or U16597 (N_16597,N_7628,N_209);
nand U16598 (N_16598,N_3146,N_7869);
nor U16599 (N_16599,N_4750,N_8480);
nand U16600 (N_16600,N_7704,N_4139);
nor U16601 (N_16601,N_1090,N_4857);
or U16602 (N_16602,N_2733,N_8841);
nor U16603 (N_16603,N_5087,N_2022);
or U16604 (N_16604,N_5813,N_4938);
xnor U16605 (N_16605,N_4392,N_7556);
and U16606 (N_16606,N_2831,N_9814);
nor U16607 (N_16607,N_5093,N_8361);
and U16608 (N_16608,N_7878,N_3748);
nand U16609 (N_16609,N_7207,N_1845);
nor U16610 (N_16610,N_5190,N_3527);
nand U16611 (N_16611,N_2257,N_7007);
or U16612 (N_16612,N_726,N_9474);
xor U16613 (N_16613,N_5368,N_7136);
xor U16614 (N_16614,N_8249,N_2586);
nand U16615 (N_16615,N_3915,N_7747);
nor U16616 (N_16616,N_6202,N_4492);
or U16617 (N_16617,N_928,N_3287);
or U16618 (N_16618,N_9741,N_8339);
and U16619 (N_16619,N_1680,N_4223);
nand U16620 (N_16620,N_680,N_4223);
xnor U16621 (N_16621,N_1307,N_8938);
and U16622 (N_16622,N_5317,N_6590);
or U16623 (N_16623,N_6378,N_1666);
or U16624 (N_16624,N_8125,N_7295);
xnor U16625 (N_16625,N_1241,N_7422);
nand U16626 (N_16626,N_1415,N_9621);
or U16627 (N_16627,N_9495,N_341);
nand U16628 (N_16628,N_4869,N_9869);
and U16629 (N_16629,N_578,N_1344);
xnor U16630 (N_16630,N_8978,N_3996);
nand U16631 (N_16631,N_5804,N_2676);
nor U16632 (N_16632,N_1200,N_6139);
xnor U16633 (N_16633,N_6230,N_8984);
or U16634 (N_16634,N_170,N_5445);
nor U16635 (N_16635,N_779,N_9760);
or U16636 (N_16636,N_8249,N_9516);
xnor U16637 (N_16637,N_202,N_6274);
or U16638 (N_16638,N_3093,N_2350);
or U16639 (N_16639,N_8503,N_6206);
or U16640 (N_16640,N_9463,N_3745);
xor U16641 (N_16641,N_9888,N_21);
and U16642 (N_16642,N_1439,N_6819);
and U16643 (N_16643,N_4376,N_8192);
and U16644 (N_16644,N_5928,N_724);
nor U16645 (N_16645,N_7101,N_5203);
nor U16646 (N_16646,N_1831,N_3918);
nor U16647 (N_16647,N_2552,N_2933);
and U16648 (N_16648,N_7311,N_9167);
or U16649 (N_16649,N_136,N_9702);
or U16650 (N_16650,N_9625,N_4445);
or U16651 (N_16651,N_6896,N_2032);
nand U16652 (N_16652,N_7330,N_1067);
or U16653 (N_16653,N_7007,N_9326);
nand U16654 (N_16654,N_1504,N_2394);
or U16655 (N_16655,N_4074,N_7981);
nor U16656 (N_16656,N_5111,N_3452);
and U16657 (N_16657,N_1135,N_479);
or U16658 (N_16658,N_8761,N_5265);
nor U16659 (N_16659,N_6845,N_3197);
nor U16660 (N_16660,N_5380,N_7529);
and U16661 (N_16661,N_1316,N_6352);
or U16662 (N_16662,N_9939,N_1078);
xor U16663 (N_16663,N_8310,N_192);
or U16664 (N_16664,N_782,N_3036);
nand U16665 (N_16665,N_1647,N_4418);
or U16666 (N_16666,N_4976,N_5179);
nor U16667 (N_16667,N_3529,N_8370);
and U16668 (N_16668,N_2405,N_4869);
or U16669 (N_16669,N_7263,N_1570);
and U16670 (N_16670,N_5765,N_1261);
xnor U16671 (N_16671,N_2770,N_4119);
or U16672 (N_16672,N_750,N_5687);
nand U16673 (N_16673,N_8315,N_4551);
or U16674 (N_16674,N_637,N_1339);
xnor U16675 (N_16675,N_5613,N_5766);
and U16676 (N_16676,N_7809,N_7364);
or U16677 (N_16677,N_6293,N_9069);
nor U16678 (N_16678,N_6506,N_7292);
or U16679 (N_16679,N_701,N_4742);
xor U16680 (N_16680,N_8993,N_2415);
and U16681 (N_16681,N_9220,N_2127);
nand U16682 (N_16682,N_4263,N_1498);
nor U16683 (N_16683,N_1991,N_737);
nand U16684 (N_16684,N_634,N_1146);
or U16685 (N_16685,N_3608,N_9678);
xor U16686 (N_16686,N_4185,N_7054);
xor U16687 (N_16687,N_693,N_7785);
or U16688 (N_16688,N_3273,N_8769);
or U16689 (N_16689,N_6602,N_8061);
nor U16690 (N_16690,N_5804,N_6966);
or U16691 (N_16691,N_5161,N_2219);
or U16692 (N_16692,N_8849,N_4500);
and U16693 (N_16693,N_1832,N_113);
nor U16694 (N_16694,N_7534,N_1498);
xor U16695 (N_16695,N_7100,N_2738);
and U16696 (N_16696,N_6940,N_9781);
nand U16697 (N_16697,N_7105,N_6248);
nor U16698 (N_16698,N_1219,N_9235);
or U16699 (N_16699,N_5014,N_3589);
and U16700 (N_16700,N_3369,N_4671);
or U16701 (N_16701,N_2768,N_7667);
xnor U16702 (N_16702,N_9241,N_9183);
nor U16703 (N_16703,N_205,N_5379);
nor U16704 (N_16704,N_9874,N_7941);
nor U16705 (N_16705,N_6621,N_4600);
nor U16706 (N_16706,N_8801,N_4342);
xnor U16707 (N_16707,N_9706,N_5262);
or U16708 (N_16708,N_5430,N_5302);
or U16709 (N_16709,N_881,N_2645);
nor U16710 (N_16710,N_2703,N_1171);
or U16711 (N_16711,N_9231,N_4119);
nor U16712 (N_16712,N_5780,N_319);
and U16713 (N_16713,N_6276,N_5300);
nand U16714 (N_16714,N_3792,N_815);
nand U16715 (N_16715,N_8896,N_5853);
nand U16716 (N_16716,N_7879,N_9300);
and U16717 (N_16717,N_2625,N_3012);
nor U16718 (N_16718,N_5068,N_7249);
nand U16719 (N_16719,N_9480,N_2147);
nor U16720 (N_16720,N_3090,N_8442);
nor U16721 (N_16721,N_2909,N_6479);
and U16722 (N_16722,N_1621,N_6863);
nand U16723 (N_16723,N_8079,N_2949);
or U16724 (N_16724,N_6875,N_7126);
or U16725 (N_16725,N_8597,N_4936);
nand U16726 (N_16726,N_8236,N_2142);
nand U16727 (N_16727,N_2593,N_3819);
xor U16728 (N_16728,N_2489,N_5000);
nor U16729 (N_16729,N_1130,N_2562);
nand U16730 (N_16730,N_7396,N_6744);
nor U16731 (N_16731,N_4480,N_3236);
xor U16732 (N_16732,N_63,N_3917);
or U16733 (N_16733,N_4988,N_9748);
and U16734 (N_16734,N_4852,N_9553);
nand U16735 (N_16735,N_6322,N_6512);
or U16736 (N_16736,N_3653,N_9477);
and U16737 (N_16737,N_3185,N_4885);
nor U16738 (N_16738,N_8790,N_7801);
nand U16739 (N_16739,N_7290,N_6393);
nor U16740 (N_16740,N_7713,N_9291);
xor U16741 (N_16741,N_4002,N_1636);
nand U16742 (N_16742,N_9647,N_5468);
xor U16743 (N_16743,N_2203,N_7502);
and U16744 (N_16744,N_7643,N_5267);
and U16745 (N_16745,N_6106,N_8705);
nor U16746 (N_16746,N_4394,N_8625);
nor U16747 (N_16747,N_7002,N_1329);
nor U16748 (N_16748,N_3862,N_3645);
or U16749 (N_16749,N_1793,N_9877);
and U16750 (N_16750,N_7735,N_4404);
and U16751 (N_16751,N_2931,N_3053);
or U16752 (N_16752,N_3155,N_8205);
nand U16753 (N_16753,N_5337,N_1067);
nor U16754 (N_16754,N_8675,N_2678);
and U16755 (N_16755,N_614,N_9949);
nor U16756 (N_16756,N_4384,N_2725);
or U16757 (N_16757,N_7102,N_7675);
nor U16758 (N_16758,N_3024,N_3995);
or U16759 (N_16759,N_7990,N_1263);
and U16760 (N_16760,N_3646,N_2884);
xor U16761 (N_16761,N_6723,N_2928);
nor U16762 (N_16762,N_1614,N_2169);
or U16763 (N_16763,N_7820,N_5964);
xor U16764 (N_16764,N_3851,N_6873);
nand U16765 (N_16765,N_2259,N_8806);
or U16766 (N_16766,N_6639,N_3630);
nand U16767 (N_16767,N_540,N_6823);
nor U16768 (N_16768,N_6660,N_5385);
nor U16769 (N_16769,N_619,N_1062);
or U16770 (N_16770,N_9171,N_1437);
nand U16771 (N_16771,N_8376,N_4002);
nor U16772 (N_16772,N_7528,N_8403);
xor U16773 (N_16773,N_3624,N_9868);
and U16774 (N_16774,N_3953,N_4766);
or U16775 (N_16775,N_6711,N_7284);
or U16776 (N_16776,N_1580,N_7769);
nand U16777 (N_16777,N_3857,N_8119);
nor U16778 (N_16778,N_1874,N_8105);
nor U16779 (N_16779,N_3893,N_8957);
and U16780 (N_16780,N_7060,N_659);
nand U16781 (N_16781,N_5269,N_2046);
or U16782 (N_16782,N_6073,N_4691);
and U16783 (N_16783,N_9925,N_3085);
or U16784 (N_16784,N_4595,N_6670);
nand U16785 (N_16785,N_2580,N_9333);
xor U16786 (N_16786,N_9195,N_5616);
nor U16787 (N_16787,N_8984,N_7037);
nor U16788 (N_16788,N_7800,N_4868);
and U16789 (N_16789,N_2077,N_1714);
nand U16790 (N_16790,N_6318,N_5036);
and U16791 (N_16791,N_3527,N_4187);
nand U16792 (N_16792,N_8359,N_6415);
or U16793 (N_16793,N_8673,N_6884);
and U16794 (N_16794,N_6250,N_3041);
or U16795 (N_16795,N_9153,N_44);
or U16796 (N_16796,N_9968,N_2669);
nand U16797 (N_16797,N_1908,N_2533);
nor U16798 (N_16798,N_4619,N_6379);
or U16799 (N_16799,N_168,N_2869);
nand U16800 (N_16800,N_4634,N_6947);
nand U16801 (N_16801,N_1511,N_9564);
nand U16802 (N_16802,N_6760,N_5798);
nand U16803 (N_16803,N_1020,N_6975);
and U16804 (N_16804,N_3199,N_3794);
or U16805 (N_16805,N_8407,N_3817);
and U16806 (N_16806,N_2049,N_2180);
nor U16807 (N_16807,N_9515,N_3899);
and U16808 (N_16808,N_1704,N_5865);
or U16809 (N_16809,N_8044,N_9484);
nand U16810 (N_16810,N_1524,N_7152);
or U16811 (N_16811,N_3201,N_4498);
nand U16812 (N_16812,N_881,N_5483);
or U16813 (N_16813,N_3849,N_7479);
or U16814 (N_16814,N_2802,N_4786);
and U16815 (N_16815,N_8452,N_1766);
nand U16816 (N_16816,N_5414,N_3512);
and U16817 (N_16817,N_3497,N_2226);
and U16818 (N_16818,N_1392,N_1892);
xor U16819 (N_16819,N_11,N_9148);
and U16820 (N_16820,N_3572,N_2282);
nand U16821 (N_16821,N_3493,N_4983);
or U16822 (N_16822,N_8756,N_6667);
nand U16823 (N_16823,N_6157,N_3664);
nor U16824 (N_16824,N_2635,N_5433);
and U16825 (N_16825,N_6394,N_1593);
nand U16826 (N_16826,N_7141,N_2520);
nand U16827 (N_16827,N_3873,N_6295);
nor U16828 (N_16828,N_8187,N_4802);
nand U16829 (N_16829,N_3772,N_945);
nor U16830 (N_16830,N_9178,N_5663);
nand U16831 (N_16831,N_1412,N_4280);
or U16832 (N_16832,N_9744,N_148);
or U16833 (N_16833,N_4222,N_2686);
xor U16834 (N_16834,N_6831,N_7302);
xnor U16835 (N_16835,N_8182,N_5428);
nor U16836 (N_16836,N_9133,N_8066);
nor U16837 (N_16837,N_1092,N_1725);
nand U16838 (N_16838,N_5952,N_6049);
xor U16839 (N_16839,N_5491,N_8524);
nor U16840 (N_16840,N_701,N_2784);
nor U16841 (N_16841,N_3815,N_5346);
and U16842 (N_16842,N_4216,N_1132);
or U16843 (N_16843,N_5456,N_4620);
nand U16844 (N_16844,N_8016,N_1641);
nand U16845 (N_16845,N_794,N_2203);
and U16846 (N_16846,N_7260,N_7566);
or U16847 (N_16847,N_354,N_5853);
and U16848 (N_16848,N_5204,N_3860);
or U16849 (N_16849,N_4998,N_5958);
and U16850 (N_16850,N_5706,N_3020);
nor U16851 (N_16851,N_5385,N_372);
nand U16852 (N_16852,N_5757,N_6159);
or U16853 (N_16853,N_4522,N_3559);
nor U16854 (N_16854,N_7595,N_6887);
or U16855 (N_16855,N_8077,N_8784);
nand U16856 (N_16856,N_2583,N_3957);
nor U16857 (N_16857,N_4781,N_6758);
nand U16858 (N_16858,N_5865,N_4079);
nor U16859 (N_16859,N_166,N_7447);
nand U16860 (N_16860,N_3837,N_8160);
nand U16861 (N_16861,N_3966,N_12);
nor U16862 (N_16862,N_532,N_4542);
nor U16863 (N_16863,N_6343,N_9839);
nand U16864 (N_16864,N_5050,N_2515);
nand U16865 (N_16865,N_2735,N_108);
nor U16866 (N_16866,N_2335,N_9255);
and U16867 (N_16867,N_3090,N_8078);
nand U16868 (N_16868,N_197,N_3083);
or U16869 (N_16869,N_9326,N_7899);
nand U16870 (N_16870,N_3587,N_1809);
nor U16871 (N_16871,N_3405,N_256);
and U16872 (N_16872,N_3843,N_2469);
nand U16873 (N_16873,N_9005,N_9573);
nand U16874 (N_16874,N_8223,N_3125);
nand U16875 (N_16875,N_5688,N_5121);
xor U16876 (N_16876,N_1818,N_3231);
and U16877 (N_16877,N_3988,N_4963);
nand U16878 (N_16878,N_9313,N_9152);
and U16879 (N_16879,N_4280,N_349);
or U16880 (N_16880,N_4542,N_8379);
or U16881 (N_16881,N_9089,N_4268);
xor U16882 (N_16882,N_7010,N_1510);
nor U16883 (N_16883,N_5954,N_9053);
nor U16884 (N_16884,N_9801,N_3104);
nor U16885 (N_16885,N_8046,N_6113);
and U16886 (N_16886,N_9481,N_7770);
xnor U16887 (N_16887,N_6303,N_8184);
nor U16888 (N_16888,N_6451,N_4432);
xnor U16889 (N_16889,N_4949,N_6027);
or U16890 (N_16890,N_2019,N_4640);
and U16891 (N_16891,N_9175,N_8423);
and U16892 (N_16892,N_382,N_5295);
and U16893 (N_16893,N_8601,N_402);
and U16894 (N_16894,N_1038,N_5744);
and U16895 (N_16895,N_288,N_696);
or U16896 (N_16896,N_1077,N_9530);
nor U16897 (N_16897,N_2314,N_2694);
nand U16898 (N_16898,N_652,N_5874);
nor U16899 (N_16899,N_2113,N_7303);
nor U16900 (N_16900,N_4580,N_3117);
or U16901 (N_16901,N_3739,N_79);
and U16902 (N_16902,N_1147,N_8891);
nor U16903 (N_16903,N_8963,N_1279);
nand U16904 (N_16904,N_6027,N_4682);
and U16905 (N_16905,N_735,N_9019);
and U16906 (N_16906,N_4883,N_9553);
nor U16907 (N_16907,N_1142,N_1869);
xnor U16908 (N_16908,N_4252,N_6544);
nand U16909 (N_16909,N_2018,N_1523);
and U16910 (N_16910,N_8415,N_5970);
and U16911 (N_16911,N_4841,N_2968);
nand U16912 (N_16912,N_3333,N_9128);
and U16913 (N_16913,N_4965,N_2618);
or U16914 (N_16914,N_5934,N_9660);
xor U16915 (N_16915,N_7303,N_2559);
or U16916 (N_16916,N_2530,N_9737);
nand U16917 (N_16917,N_141,N_9813);
nor U16918 (N_16918,N_7162,N_2142);
nor U16919 (N_16919,N_3555,N_4776);
or U16920 (N_16920,N_4567,N_6959);
and U16921 (N_16921,N_5172,N_9662);
or U16922 (N_16922,N_9528,N_6862);
xnor U16923 (N_16923,N_5823,N_4184);
nor U16924 (N_16924,N_9512,N_2767);
or U16925 (N_16925,N_9051,N_4992);
or U16926 (N_16926,N_5768,N_9229);
nor U16927 (N_16927,N_4792,N_9054);
nand U16928 (N_16928,N_5322,N_4250);
and U16929 (N_16929,N_6765,N_23);
nor U16930 (N_16930,N_9215,N_1215);
nand U16931 (N_16931,N_4088,N_8523);
nor U16932 (N_16932,N_5709,N_2848);
nand U16933 (N_16933,N_4914,N_1844);
nor U16934 (N_16934,N_1697,N_4162);
or U16935 (N_16935,N_9611,N_6623);
nand U16936 (N_16936,N_5487,N_4332);
nor U16937 (N_16937,N_9834,N_1328);
or U16938 (N_16938,N_662,N_640);
or U16939 (N_16939,N_1691,N_7642);
nor U16940 (N_16940,N_7108,N_1120);
nand U16941 (N_16941,N_2873,N_4435);
nand U16942 (N_16942,N_3809,N_4801);
and U16943 (N_16943,N_3622,N_6290);
or U16944 (N_16944,N_5668,N_598);
xor U16945 (N_16945,N_7409,N_4340);
nor U16946 (N_16946,N_6983,N_6096);
nor U16947 (N_16947,N_1782,N_1582);
nor U16948 (N_16948,N_8835,N_5868);
nand U16949 (N_16949,N_8842,N_4754);
xor U16950 (N_16950,N_4477,N_7082);
nand U16951 (N_16951,N_5237,N_7915);
xnor U16952 (N_16952,N_8242,N_366);
nand U16953 (N_16953,N_9058,N_3045);
nor U16954 (N_16954,N_5434,N_8448);
or U16955 (N_16955,N_7927,N_5730);
xnor U16956 (N_16956,N_9596,N_8592);
and U16957 (N_16957,N_7519,N_8688);
nor U16958 (N_16958,N_570,N_596);
or U16959 (N_16959,N_5275,N_921);
or U16960 (N_16960,N_5005,N_197);
or U16961 (N_16961,N_8261,N_7245);
nor U16962 (N_16962,N_2195,N_1428);
and U16963 (N_16963,N_1830,N_7061);
nand U16964 (N_16964,N_9582,N_5872);
and U16965 (N_16965,N_2288,N_2020);
and U16966 (N_16966,N_7947,N_5490);
or U16967 (N_16967,N_8578,N_2311);
and U16968 (N_16968,N_160,N_9491);
or U16969 (N_16969,N_7211,N_8421);
xor U16970 (N_16970,N_5569,N_695);
nor U16971 (N_16971,N_4543,N_9013);
nand U16972 (N_16972,N_8693,N_6404);
xor U16973 (N_16973,N_6819,N_390);
and U16974 (N_16974,N_7593,N_2686);
nand U16975 (N_16975,N_902,N_7028);
and U16976 (N_16976,N_1859,N_896);
nor U16977 (N_16977,N_1291,N_1596);
or U16978 (N_16978,N_9354,N_3872);
or U16979 (N_16979,N_6915,N_2130);
nand U16980 (N_16980,N_2408,N_4030);
and U16981 (N_16981,N_4694,N_5431);
xnor U16982 (N_16982,N_8845,N_8760);
nand U16983 (N_16983,N_5136,N_7362);
nand U16984 (N_16984,N_7534,N_3099);
and U16985 (N_16985,N_7330,N_2647);
nor U16986 (N_16986,N_8875,N_3046);
and U16987 (N_16987,N_8053,N_905);
or U16988 (N_16988,N_5800,N_5810);
xnor U16989 (N_16989,N_8588,N_505);
nand U16990 (N_16990,N_3898,N_6651);
and U16991 (N_16991,N_338,N_920);
nand U16992 (N_16992,N_7712,N_9431);
nand U16993 (N_16993,N_5267,N_2315);
nor U16994 (N_16994,N_3633,N_9357);
or U16995 (N_16995,N_6933,N_7398);
xor U16996 (N_16996,N_3287,N_4387);
xnor U16997 (N_16997,N_8157,N_4434);
or U16998 (N_16998,N_1147,N_7590);
xnor U16999 (N_16999,N_936,N_1434);
xnor U17000 (N_17000,N_3930,N_7507);
nor U17001 (N_17001,N_8184,N_3645);
and U17002 (N_17002,N_8730,N_6969);
and U17003 (N_17003,N_1790,N_5871);
nor U17004 (N_17004,N_6380,N_803);
or U17005 (N_17005,N_5728,N_9214);
or U17006 (N_17006,N_7124,N_2543);
and U17007 (N_17007,N_2961,N_6351);
nand U17008 (N_17008,N_472,N_1952);
and U17009 (N_17009,N_9142,N_7016);
nand U17010 (N_17010,N_3858,N_9434);
nor U17011 (N_17011,N_568,N_3923);
nor U17012 (N_17012,N_6681,N_3492);
xnor U17013 (N_17013,N_7420,N_4253);
or U17014 (N_17014,N_8201,N_457);
nor U17015 (N_17015,N_2836,N_2602);
and U17016 (N_17016,N_5847,N_3424);
and U17017 (N_17017,N_4676,N_26);
or U17018 (N_17018,N_9414,N_6767);
nor U17019 (N_17019,N_41,N_8964);
nor U17020 (N_17020,N_1036,N_3114);
nor U17021 (N_17021,N_9600,N_8288);
and U17022 (N_17022,N_5660,N_9631);
or U17023 (N_17023,N_2701,N_7468);
and U17024 (N_17024,N_3263,N_1958);
and U17025 (N_17025,N_3911,N_8839);
or U17026 (N_17026,N_8397,N_3775);
or U17027 (N_17027,N_4152,N_6905);
and U17028 (N_17028,N_9241,N_9673);
nor U17029 (N_17029,N_4319,N_3679);
and U17030 (N_17030,N_2558,N_3685);
xnor U17031 (N_17031,N_3764,N_3987);
nand U17032 (N_17032,N_8222,N_4427);
or U17033 (N_17033,N_8684,N_3545);
and U17034 (N_17034,N_1240,N_5025);
nor U17035 (N_17035,N_3707,N_7138);
and U17036 (N_17036,N_8261,N_7029);
nor U17037 (N_17037,N_3422,N_850);
or U17038 (N_17038,N_3060,N_9189);
and U17039 (N_17039,N_898,N_8659);
and U17040 (N_17040,N_6191,N_526);
nand U17041 (N_17041,N_2026,N_1957);
nor U17042 (N_17042,N_3728,N_1705);
nor U17043 (N_17043,N_1218,N_2402);
nor U17044 (N_17044,N_2432,N_9837);
nand U17045 (N_17045,N_6201,N_62);
or U17046 (N_17046,N_9621,N_3882);
nand U17047 (N_17047,N_862,N_9804);
or U17048 (N_17048,N_3757,N_992);
or U17049 (N_17049,N_7492,N_3677);
nand U17050 (N_17050,N_6631,N_8676);
nor U17051 (N_17051,N_4093,N_789);
nand U17052 (N_17052,N_8615,N_5254);
nor U17053 (N_17053,N_8880,N_5079);
xor U17054 (N_17054,N_8330,N_119);
nor U17055 (N_17055,N_7844,N_1815);
nor U17056 (N_17056,N_4948,N_4887);
nor U17057 (N_17057,N_1772,N_7269);
nor U17058 (N_17058,N_7850,N_5123);
nor U17059 (N_17059,N_8541,N_4780);
and U17060 (N_17060,N_8424,N_9301);
xnor U17061 (N_17061,N_7164,N_8114);
or U17062 (N_17062,N_3126,N_8478);
nand U17063 (N_17063,N_806,N_7968);
and U17064 (N_17064,N_9621,N_9013);
or U17065 (N_17065,N_6704,N_4758);
and U17066 (N_17066,N_5524,N_7110);
and U17067 (N_17067,N_8737,N_8331);
nor U17068 (N_17068,N_1616,N_8438);
nor U17069 (N_17069,N_3758,N_2923);
nand U17070 (N_17070,N_36,N_9090);
and U17071 (N_17071,N_3445,N_7642);
nor U17072 (N_17072,N_8701,N_7367);
nand U17073 (N_17073,N_4205,N_5267);
nor U17074 (N_17074,N_4292,N_4813);
nor U17075 (N_17075,N_6881,N_261);
nand U17076 (N_17076,N_825,N_1705);
and U17077 (N_17077,N_6744,N_7320);
nand U17078 (N_17078,N_6051,N_2421);
xnor U17079 (N_17079,N_3661,N_6921);
nor U17080 (N_17080,N_7537,N_4222);
nand U17081 (N_17081,N_3697,N_4955);
nand U17082 (N_17082,N_4035,N_6435);
nand U17083 (N_17083,N_4086,N_6363);
or U17084 (N_17084,N_6999,N_4263);
and U17085 (N_17085,N_3473,N_2410);
and U17086 (N_17086,N_217,N_9073);
and U17087 (N_17087,N_5711,N_8047);
or U17088 (N_17088,N_9881,N_7018);
nand U17089 (N_17089,N_1289,N_4083);
xor U17090 (N_17090,N_4026,N_5756);
or U17091 (N_17091,N_4376,N_6115);
nor U17092 (N_17092,N_7196,N_7338);
nor U17093 (N_17093,N_188,N_8532);
nor U17094 (N_17094,N_5207,N_8513);
and U17095 (N_17095,N_3876,N_9733);
nand U17096 (N_17096,N_7595,N_2787);
or U17097 (N_17097,N_8372,N_1918);
or U17098 (N_17098,N_5699,N_2565);
nand U17099 (N_17099,N_4801,N_5351);
nand U17100 (N_17100,N_5837,N_1618);
nor U17101 (N_17101,N_4243,N_9414);
nor U17102 (N_17102,N_2465,N_1164);
nor U17103 (N_17103,N_6079,N_6067);
and U17104 (N_17104,N_2090,N_2160);
or U17105 (N_17105,N_8121,N_4864);
nand U17106 (N_17106,N_9598,N_1614);
or U17107 (N_17107,N_2761,N_5020);
and U17108 (N_17108,N_1488,N_7643);
nand U17109 (N_17109,N_715,N_6202);
or U17110 (N_17110,N_1693,N_7354);
and U17111 (N_17111,N_3332,N_5564);
nor U17112 (N_17112,N_6143,N_3126);
nor U17113 (N_17113,N_2390,N_9595);
xor U17114 (N_17114,N_1573,N_5054);
and U17115 (N_17115,N_4062,N_7750);
nor U17116 (N_17116,N_9258,N_142);
or U17117 (N_17117,N_5839,N_9014);
nor U17118 (N_17118,N_2388,N_1745);
nor U17119 (N_17119,N_4305,N_2417);
nor U17120 (N_17120,N_2717,N_5647);
nand U17121 (N_17121,N_762,N_1977);
and U17122 (N_17122,N_3494,N_7103);
or U17123 (N_17123,N_5253,N_1840);
and U17124 (N_17124,N_3640,N_9381);
nor U17125 (N_17125,N_9615,N_4161);
nor U17126 (N_17126,N_6600,N_7502);
nand U17127 (N_17127,N_5279,N_1064);
nand U17128 (N_17128,N_831,N_527);
nor U17129 (N_17129,N_8295,N_6581);
or U17130 (N_17130,N_6541,N_7891);
nor U17131 (N_17131,N_834,N_690);
and U17132 (N_17132,N_1671,N_9750);
or U17133 (N_17133,N_5108,N_1948);
nor U17134 (N_17134,N_9907,N_6145);
and U17135 (N_17135,N_4226,N_2283);
nor U17136 (N_17136,N_9485,N_484);
and U17137 (N_17137,N_759,N_1316);
and U17138 (N_17138,N_2184,N_4293);
nor U17139 (N_17139,N_5275,N_1273);
and U17140 (N_17140,N_7654,N_4361);
and U17141 (N_17141,N_2569,N_9229);
nor U17142 (N_17142,N_4596,N_8925);
and U17143 (N_17143,N_4453,N_9362);
nand U17144 (N_17144,N_3400,N_5114);
nand U17145 (N_17145,N_2665,N_220);
nand U17146 (N_17146,N_2788,N_4148);
or U17147 (N_17147,N_6990,N_8149);
or U17148 (N_17148,N_5874,N_5209);
or U17149 (N_17149,N_4949,N_320);
or U17150 (N_17150,N_3901,N_7538);
xor U17151 (N_17151,N_8562,N_9915);
or U17152 (N_17152,N_4904,N_1700);
nand U17153 (N_17153,N_8275,N_5900);
xor U17154 (N_17154,N_7594,N_3369);
nor U17155 (N_17155,N_2623,N_7077);
and U17156 (N_17156,N_1029,N_3979);
and U17157 (N_17157,N_3190,N_719);
and U17158 (N_17158,N_9601,N_562);
xnor U17159 (N_17159,N_5061,N_9570);
and U17160 (N_17160,N_3373,N_6874);
and U17161 (N_17161,N_9531,N_8231);
nor U17162 (N_17162,N_4234,N_2399);
nor U17163 (N_17163,N_1084,N_3658);
nand U17164 (N_17164,N_8796,N_6393);
or U17165 (N_17165,N_8081,N_9446);
nor U17166 (N_17166,N_3647,N_930);
nor U17167 (N_17167,N_6695,N_2348);
or U17168 (N_17168,N_3740,N_7069);
or U17169 (N_17169,N_2398,N_8716);
and U17170 (N_17170,N_8498,N_3415);
and U17171 (N_17171,N_1366,N_4942);
nor U17172 (N_17172,N_6815,N_7652);
xnor U17173 (N_17173,N_9196,N_3489);
or U17174 (N_17174,N_1778,N_8348);
nor U17175 (N_17175,N_5018,N_8999);
and U17176 (N_17176,N_3072,N_3791);
nand U17177 (N_17177,N_5264,N_5163);
nor U17178 (N_17178,N_1919,N_1857);
nor U17179 (N_17179,N_5971,N_5823);
nand U17180 (N_17180,N_8030,N_6048);
nand U17181 (N_17181,N_9469,N_4617);
xnor U17182 (N_17182,N_9373,N_8266);
and U17183 (N_17183,N_8525,N_6737);
and U17184 (N_17184,N_2113,N_6961);
nand U17185 (N_17185,N_858,N_3462);
or U17186 (N_17186,N_876,N_7344);
and U17187 (N_17187,N_3232,N_9822);
and U17188 (N_17188,N_5336,N_5110);
or U17189 (N_17189,N_88,N_1292);
nor U17190 (N_17190,N_6225,N_5817);
and U17191 (N_17191,N_4748,N_4325);
nand U17192 (N_17192,N_7948,N_7925);
and U17193 (N_17193,N_7308,N_5147);
and U17194 (N_17194,N_1197,N_247);
or U17195 (N_17195,N_2630,N_6563);
nand U17196 (N_17196,N_2700,N_1314);
or U17197 (N_17197,N_4633,N_5789);
xor U17198 (N_17198,N_46,N_5360);
nor U17199 (N_17199,N_4333,N_2778);
and U17200 (N_17200,N_7080,N_5695);
or U17201 (N_17201,N_4757,N_5115);
and U17202 (N_17202,N_9210,N_4287);
or U17203 (N_17203,N_5548,N_8294);
nand U17204 (N_17204,N_120,N_457);
nand U17205 (N_17205,N_3478,N_6441);
nand U17206 (N_17206,N_393,N_3000);
or U17207 (N_17207,N_52,N_4985);
and U17208 (N_17208,N_657,N_1595);
or U17209 (N_17209,N_4986,N_3019);
or U17210 (N_17210,N_2442,N_8361);
nand U17211 (N_17211,N_5274,N_6636);
nor U17212 (N_17212,N_7387,N_6316);
nor U17213 (N_17213,N_5445,N_6291);
and U17214 (N_17214,N_353,N_3375);
and U17215 (N_17215,N_661,N_2160);
nor U17216 (N_17216,N_3925,N_4191);
or U17217 (N_17217,N_8081,N_6662);
or U17218 (N_17218,N_8801,N_2275);
or U17219 (N_17219,N_4537,N_1876);
nand U17220 (N_17220,N_8929,N_9382);
or U17221 (N_17221,N_3497,N_8493);
nand U17222 (N_17222,N_6421,N_5859);
or U17223 (N_17223,N_558,N_4482);
xnor U17224 (N_17224,N_8310,N_8722);
xor U17225 (N_17225,N_9359,N_5643);
and U17226 (N_17226,N_6887,N_9685);
and U17227 (N_17227,N_7070,N_3664);
nand U17228 (N_17228,N_2112,N_4151);
xor U17229 (N_17229,N_3654,N_7889);
nand U17230 (N_17230,N_1123,N_1429);
nor U17231 (N_17231,N_72,N_4969);
and U17232 (N_17232,N_5710,N_2573);
nor U17233 (N_17233,N_3361,N_599);
nand U17234 (N_17234,N_5895,N_1539);
nand U17235 (N_17235,N_5298,N_5662);
or U17236 (N_17236,N_6429,N_4940);
nor U17237 (N_17237,N_9922,N_4551);
and U17238 (N_17238,N_4638,N_7093);
nor U17239 (N_17239,N_5913,N_5709);
and U17240 (N_17240,N_5262,N_9835);
xnor U17241 (N_17241,N_736,N_3835);
nor U17242 (N_17242,N_5083,N_4291);
and U17243 (N_17243,N_7820,N_3254);
or U17244 (N_17244,N_1607,N_951);
or U17245 (N_17245,N_7427,N_380);
and U17246 (N_17246,N_9510,N_1907);
nand U17247 (N_17247,N_7818,N_1846);
nor U17248 (N_17248,N_7393,N_6616);
and U17249 (N_17249,N_2753,N_5911);
nor U17250 (N_17250,N_3235,N_1927);
and U17251 (N_17251,N_286,N_2517);
nand U17252 (N_17252,N_7680,N_7828);
or U17253 (N_17253,N_9591,N_2918);
nand U17254 (N_17254,N_9100,N_2972);
or U17255 (N_17255,N_5646,N_9054);
xor U17256 (N_17256,N_6308,N_1558);
and U17257 (N_17257,N_5359,N_5422);
nor U17258 (N_17258,N_5380,N_2337);
xnor U17259 (N_17259,N_687,N_3604);
nor U17260 (N_17260,N_8049,N_9715);
nor U17261 (N_17261,N_7252,N_3426);
nand U17262 (N_17262,N_7022,N_2903);
or U17263 (N_17263,N_482,N_857);
nand U17264 (N_17264,N_2693,N_1744);
nand U17265 (N_17265,N_8466,N_4558);
nor U17266 (N_17266,N_7929,N_7345);
and U17267 (N_17267,N_9458,N_1947);
and U17268 (N_17268,N_6767,N_2844);
nor U17269 (N_17269,N_1452,N_5797);
nor U17270 (N_17270,N_4337,N_9048);
xor U17271 (N_17271,N_5969,N_1200);
nand U17272 (N_17272,N_7586,N_7222);
nand U17273 (N_17273,N_6095,N_254);
or U17274 (N_17274,N_7976,N_367);
nand U17275 (N_17275,N_7274,N_2140);
or U17276 (N_17276,N_1192,N_6549);
nor U17277 (N_17277,N_7405,N_9434);
nand U17278 (N_17278,N_3533,N_377);
nand U17279 (N_17279,N_3129,N_2678);
nand U17280 (N_17280,N_1963,N_665);
and U17281 (N_17281,N_9601,N_8717);
and U17282 (N_17282,N_4545,N_8084);
nor U17283 (N_17283,N_124,N_6123);
nor U17284 (N_17284,N_2988,N_4207);
or U17285 (N_17285,N_5706,N_851);
and U17286 (N_17286,N_9900,N_3058);
or U17287 (N_17287,N_9816,N_434);
nor U17288 (N_17288,N_5391,N_388);
and U17289 (N_17289,N_353,N_7483);
nor U17290 (N_17290,N_9922,N_4685);
nand U17291 (N_17291,N_3316,N_218);
nand U17292 (N_17292,N_1247,N_8992);
or U17293 (N_17293,N_6212,N_1882);
and U17294 (N_17294,N_5464,N_2755);
or U17295 (N_17295,N_7480,N_9404);
or U17296 (N_17296,N_3046,N_6098);
or U17297 (N_17297,N_8748,N_8863);
nand U17298 (N_17298,N_8944,N_5712);
nor U17299 (N_17299,N_8319,N_5699);
or U17300 (N_17300,N_3742,N_8687);
xor U17301 (N_17301,N_4324,N_95);
or U17302 (N_17302,N_8380,N_6868);
or U17303 (N_17303,N_5983,N_2539);
nand U17304 (N_17304,N_2075,N_6032);
and U17305 (N_17305,N_8407,N_6814);
or U17306 (N_17306,N_3869,N_9868);
and U17307 (N_17307,N_8352,N_1861);
or U17308 (N_17308,N_7855,N_5727);
nand U17309 (N_17309,N_1989,N_6945);
and U17310 (N_17310,N_7458,N_631);
or U17311 (N_17311,N_8543,N_350);
and U17312 (N_17312,N_5914,N_4400);
and U17313 (N_17313,N_8416,N_8689);
or U17314 (N_17314,N_7020,N_1024);
and U17315 (N_17315,N_3628,N_6711);
or U17316 (N_17316,N_5543,N_5695);
or U17317 (N_17317,N_4635,N_9251);
nand U17318 (N_17318,N_4474,N_8683);
nand U17319 (N_17319,N_7998,N_5859);
nor U17320 (N_17320,N_1968,N_9630);
nand U17321 (N_17321,N_3054,N_7715);
nand U17322 (N_17322,N_6272,N_6079);
or U17323 (N_17323,N_5335,N_224);
nor U17324 (N_17324,N_8239,N_9398);
and U17325 (N_17325,N_4029,N_6982);
nor U17326 (N_17326,N_3580,N_953);
xor U17327 (N_17327,N_3192,N_6729);
and U17328 (N_17328,N_4848,N_7100);
nand U17329 (N_17329,N_8686,N_3927);
or U17330 (N_17330,N_5458,N_4598);
nor U17331 (N_17331,N_3374,N_9565);
or U17332 (N_17332,N_1750,N_7082);
or U17333 (N_17333,N_3295,N_2030);
nand U17334 (N_17334,N_3,N_3954);
nand U17335 (N_17335,N_5570,N_8984);
nand U17336 (N_17336,N_2272,N_7294);
nand U17337 (N_17337,N_7848,N_1270);
or U17338 (N_17338,N_2913,N_9243);
nand U17339 (N_17339,N_6533,N_9211);
or U17340 (N_17340,N_1328,N_3344);
and U17341 (N_17341,N_7070,N_9582);
or U17342 (N_17342,N_4078,N_5846);
and U17343 (N_17343,N_8998,N_8988);
and U17344 (N_17344,N_4788,N_3778);
nand U17345 (N_17345,N_2997,N_7246);
xnor U17346 (N_17346,N_6559,N_7065);
nand U17347 (N_17347,N_1389,N_5959);
and U17348 (N_17348,N_9360,N_4100);
nor U17349 (N_17349,N_2177,N_7194);
and U17350 (N_17350,N_1714,N_8682);
nand U17351 (N_17351,N_6963,N_4962);
and U17352 (N_17352,N_5832,N_7571);
or U17353 (N_17353,N_6579,N_8522);
or U17354 (N_17354,N_7987,N_4321);
and U17355 (N_17355,N_7027,N_1288);
and U17356 (N_17356,N_6837,N_7977);
nor U17357 (N_17357,N_2917,N_8823);
and U17358 (N_17358,N_7141,N_1022);
or U17359 (N_17359,N_4475,N_5626);
or U17360 (N_17360,N_2551,N_880);
nand U17361 (N_17361,N_6560,N_4644);
and U17362 (N_17362,N_3338,N_3515);
or U17363 (N_17363,N_8081,N_7620);
nand U17364 (N_17364,N_3314,N_8185);
xnor U17365 (N_17365,N_8555,N_2812);
and U17366 (N_17366,N_2890,N_6349);
nand U17367 (N_17367,N_2729,N_4057);
nor U17368 (N_17368,N_916,N_4388);
or U17369 (N_17369,N_4297,N_2513);
or U17370 (N_17370,N_1476,N_4508);
nand U17371 (N_17371,N_6580,N_6819);
nor U17372 (N_17372,N_2648,N_5608);
nand U17373 (N_17373,N_1670,N_3494);
or U17374 (N_17374,N_1295,N_8647);
nor U17375 (N_17375,N_5677,N_5785);
or U17376 (N_17376,N_9923,N_1458);
or U17377 (N_17377,N_9626,N_3564);
nand U17378 (N_17378,N_7779,N_6742);
or U17379 (N_17379,N_8447,N_9445);
nor U17380 (N_17380,N_557,N_6706);
nand U17381 (N_17381,N_5765,N_6194);
nor U17382 (N_17382,N_4482,N_3765);
nand U17383 (N_17383,N_5594,N_1563);
nor U17384 (N_17384,N_8077,N_33);
or U17385 (N_17385,N_5404,N_806);
or U17386 (N_17386,N_9782,N_9251);
nor U17387 (N_17387,N_7342,N_8401);
and U17388 (N_17388,N_951,N_683);
and U17389 (N_17389,N_6472,N_168);
nor U17390 (N_17390,N_3885,N_8936);
or U17391 (N_17391,N_169,N_6890);
xnor U17392 (N_17392,N_2195,N_3010);
xor U17393 (N_17393,N_1199,N_9956);
and U17394 (N_17394,N_8822,N_4413);
nor U17395 (N_17395,N_3139,N_8450);
or U17396 (N_17396,N_6608,N_9247);
and U17397 (N_17397,N_589,N_1806);
and U17398 (N_17398,N_3148,N_8588);
xnor U17399 (N_17399,N_1605,N_7824);
nand U17400 (N_17400,N_9653,N_8873);
nor U17401 (N_17401,N_634,N_4144);
nor U17402 (N_17402,N_2159,N_221);
xnor U17403 (N_17403,N_4477,N_1073);
nand U17404 (N_17404,N_880,N_6958);
or U17405 (N_17405,N_6892,N_5088);
or U17406 (N_17406,N_9165,N_4232);
and U17407 (N_17407,N_6904,N_8201);
and U17408 (N_17408,N_934,N_3261);
or U17409 (N_17409,N_6850,N_3097);
and U17410 (N_17410,N_9156,N_1652);
and U17411 (N_17411,N_4729,N_6186);
nand U17412 (N_17412,N_7849,N_6451);
and U17413 (N_17413,N_6508,N_5166);
and U17414 (N_17414,N_219,N_6000);
nand U17415 (N_17415,N_6317,N_7399);
nor U17416 (N_17416,N_3942,N_9651);
xor U17417 (N_17417,N_9676,N_3134);
or U17418 (N_17418,N_610,N_4685);
nor U17419 (N_17419,N_1880,N_1472);
and U17420 (N_17420,N_7030,N_9981);
or U17421 (N_17421,N_6511,N_5121);
nand U17422 (N_17422,N_4905,N_8674);
or U17423 (N_17423,N_3405,N_3434);
nor U17424 (N_17424,N_1359,N_1307);
nor U17425 (N_17425,N_1443,N_1110);
nor U17426 (N_17426,N_9941,N_2140);
nor U17427 (N_17427,N_5763,N_5468);
or U17428 (N_17428,N_8562,N_9771);
xor U17429 (N_17429,N_9313,N_5069);
or U17430 (N_17430,N_9973,N_77);
or U17431 (N_17431,N_1027,N_2065);
nor U17432 (N_17432,N_730,N_3632);
and U17433 (N_17433,N_3086,N_6777);
nand U17434 (N_17434,N_8501,N_7434);
xor U17435 (N_17435,N_8102,N_1241);
nor U17436 (N_17436,N_2451,N_4084);
nor U17437 (N_17437,N_110,N_5136);
nand U17438 (N_17438,N_356,N_5604);
nand U17439 (N_17439,N_3151,N_8988);
and U17440 (N_17440,N_3472,N_8697);
nand U17441 (N_17441,N_6606,N_5583);
or U17442 (N_17442,N_6954,N_6777);
nor U17443 (N_17443,N_4527,N_8953);
nand U17444 (N_17444,N_3961,N_2012);
nor U17445 (N_17445,N_3778,N_8156);
or U17446 (N_17446,N_1448,N_4166);
nand U17447 (N_17447,N_8489,N_8947);
nor U17448 (N_17448,N_4122,N_7633);
nand U17449 (N_17449,N_8860,N_6703);
or U17450 (N_17450,N_4485,N_2492);
nand U17451 (N_17451,N_4323,N_8598);
nand U17452 (N_17452,N_8316,N_935);
and U17453 (N_17453,N_9135,N_7112);
nor U17454 (N_17454,N_9183,N_3825);
nor U17455 (N_17455,N_6858,N_9765);
or U17456 (N_17456,N_4416,N_5572);
nor U17457 (N_17457,N_2393,N_9477);
nand U17458 (N_17458,N_2463,N_6316);
or U17459 (N_17459,N_3325,N_8606);
and U17460 (N_17460,N_2441,N_5979);
nand U17461 (N_17461,N_7386,N_30);
and U17462 (N_17462,N_1509,N_4563);
and U17463 (N_17463,N_9374,N_8872);
or U17464 (N_17464,N_9759,N_9148);
nor U17465 (N_17465,N_7491,N_6283);
nand U17466 (N_17466,N_7788,N_6336);
nand U17467 (N_17467,N_1383,N_5714);
nor U17468 (N_17468,N_1120,N_8680);
and U17469 (N_17469,N_8664,N_7060);
and U17470 (N_17470,N_2997,N_7320);
and U17471 (N_17471,N_2703,N_9229);
nand U17472 (N_17472,N_7957,N_2658);
nand U17473 (N_17473,N_1581,N_6880);
and U17474 (N_17474,N_5832,N_5528);
nand U17475 (N_17475,N_3818,N_1209);
nand U17476 (N_17476,N_6797,N_3048);
nor U17477 (N_17477,N_9223,N_1877);
nand U17478 (N_17478,N_447,N_162);
and U17479 (N_17479,N_8059,N_4594);
nor U17480 (N_17480,N_1837,N_6047);
and U17481 (N_17481,N_8698,N_5557);
or U17482 (N_17482,N_2949,N_5960);
or U17483 (N_17483,N_1557,N_4012);
and U17484 (N_17484,N_2178,N_1206);
nand U17485 (N_17485,N_3573,N_8164);
nor U17486 (N_17486,N_3752,N_5027);
and U17487 (N_17487,N_5916,N_9325);
and U17488 (N_17488,N_7356,N_5193);
nand U17489 (N_17489,N_3613,N_9939);
nor U17490 (N_17490,N_2332,N_3593);
nand U17491 (N_17491,N_3517,N_4426);
or U17492 (N_17492,N_7976,N_8800);
and U17493 (N_17493,N_2107,N_1393);
or U17494 (N_17494,N_8310,N_9166);
nand U17495 (N_17495,N_9574,N_7918);
nor U17496 (N_17496,N_7188,N_2150);
and U17497 (N_17497,N_7218,N_6267);
and U17498 (N_17498,N_114,N_2840);
and U17499 (N_17499,N_5366,N_2736);
or U17500 (N_17500,N_3602,N_9252);
nor U17501 (N_17501,N_1394,N_7996);
nand U17502 (N_17502,N_8526,N_4194);
nor U17503 (N_17503,N_9523,N_4825);
or U17504 (N_17504,N_8656,N_7751);
or U17505 (N_17505,N_1024,N_6243);
or U17506 (N_17506,N_9382,N_2372);
xnor U17507 (N_17507,N_9377,N_5971);
or U17508 (N_17508,N_2761,N_8024);
and U17509 (N_17509,N_7148,N_1163);
nand U17510 (N_17510,N_5289,N_2360);
or U17511 (N_17511,N_3205,N_835);
or U17512 (N_17512,N_3580,N_6951);
nor U17513 (N_17513,N_4224,N_858);
or U17514 (N_17514,N_9538,N_8192);
nand U17515 (N_17515,N_6620,N_5511);
nor U17516 (N_17516,N_6265,N_9503);
nand U17517 (N_17517,N_4825,N_2957);
nor U17518 (N_17518,N_4818,N_1999);
nand U17519 (N_17519,N_1680,N_4012);
nand U17520 (N_17520,N_377,N_6806);
nor U17521 (N_17521,N_4069,N_2971);
nor U17522 (N_17522,N_3582,N_9047);
or U17523 (N_17523,N_1998,N_3305);
and U17524 (N_17524,N_8504,N_8108);
xnor U17525 (N_17525,N_3749,N_4679);
nor U17526 (N_17526,N_3295,N_833);
nand U17527 (N_17527,N_5306,N_600);
nor U17528 (N_17528,N_6188,N_5963);
and U17529 (N_17529,N_9211,N_5375);
or U17530 (N_17530,N_2627,N_1890);
nand U17531 (N_17531,N_2126,N_1197);
and U17532 (N_17532,N_1140,N_8775);
nand U17533 (N_17533,N_4565,N_2333);
and U17534 (N_17534,N_9288,N_2247);
nor U17535 (N_17535,N_2986,N_5879);
and U17536 (N_17536,N_1886,N_6567);
xnor U17537 (N_17537,N_2678,N_4427);
nor U17538 (N_17538,N_5095,N_743);
nor U17539 (N_17539,N_8918,N_5952);
nor U17540 (N_17540,N_3963,N_1825);
nor U17541 (N_17541,N_9272,N_5631);
nor U17542 (N_17542,N_3936,N_7020);
and U17543 (N_17543,N_1429,N_7652);
or U17544 (N_17544,N_8692,N_9062);
nor U17545 (N_17545,N_2849,N_2122);
xnor U17546 (N_17546,N_6451,N_573);
and U17547 (N_17547,N_6983,N_1269);
nor U17548 (N_17548,N_3967,N_1106);
or U17549 (N_17549,N_7565,N_1327);
xor U17550 (N_17550,N_4409,N_4050);
nor U17551 (N_17551,N_2419,N_5823);
nand U17552 (N_17552,N_5546,N_7544);
or U17553 (N_17553,N_5009,N_6550);
or U17554 (N_17554,N_153,N_4827);
or U17555 (N_17555,N_1912,N_5233);
nand U17556 (N_17556,N_6220,N_8420);
nand U17557 (N_17557,N_8860,N_1061);
nand U17558 (N_17558,N_9077,N_8037);
and U17559 (N_17559,N_5312,N_181);
or U17560 (N_17560,N_3932,N_5172);
nor U17561 (N_17561,N_1677,N_5373);
or U17562 (N_17562,N_9526,N_7772);
or U17563 (N_17563,N_8214,N_3343);
or U17564 (N_17564,N_838,N_5288);
nor U17565 (N_17565,N_693,N_3288);
nand U17566 (N_17566,N_4650,N_8911);
xnor U17567 (N_17567,N_6185,N_4288);
and U17568 (N_17568,N_8522,N_8389);
nor U17569 (N_17569,N_7974,N_6396);
nor U17570 (N_17570,N_1170,N_5725);
nor U17571 (N_17571,N_9935,N_9846);
and U17572 (N_17572,N_8835,N_6084);
and U17573 (N_17573,N_322,N_4889);
and U17574 (N_17574,N_4561,N_5739);
or U17575 (N_17575,N_8286,N_9494);
nor U17576 (N_17576,N_5191,N_1756);
or U17577 (N_17577,N_2922,N_3849);
nor U17578 (N_17578,N_2762,N_7164);
nor U17579 (N_17579,N_4963,N_9405);
nor U17580 (N_17580,N_7399,N_7751);
nor U17581 (N_17581,N_7382,N_2636);
nand U17582 (N_17582,N_7776,N_4047);
or U17583 (N_17583,N_1102,N_6464);
and U17584 (N_17584,N_6219,N_2133);
xor U17585 (N_17585,N_983,N_3886);
xor U17586 (N_17586,N_5531,N_6768);
nor U17587 (N_17587,N_3609,N_8318);
nor U17588 (N_17588,N_2977,N_4254);
nor U17589 (N_17589,N_8604,N_9575);
or U17590 (N_17590,N_6192,N_8479);
and U17591 (N_17591,N_982,N_3387);
or U17592 (N_17592,N_8012,N_8367);
and U17593 (N_17593,N_5503,N_4858);
xor U17594 (N_17594,N_1191,N_3191);
or U17595 (N_17595,N_5789,N_4274);
nor U17596 (N_17596,N_2660,N_5380);
or U17597 (N_17597,N_5363,N_3097);
nor U17598 (N_17598,N_7301,N_5134);
and U17599 (N_17599,N_5211,N_6824);
and U17600 (N_17600,N_4511,N_7703);
or U17601 (N_17601,N_6132,N_2204);
and U17602 (N_17602,N_9673,N_9467);
nand U17603 (N_17603,N_6271,N_719);
or U17604 (N_17604,N_9829,N_9525);
and U17605 (N_17605,N_7132,N_7880);
and U17606 (N_17606,N_7556,N_4034);
nand U17607 (N_17607,N_3867,N_5617);
xor U17608 (N_17608,N_4001,N_4703);
or U17609 (N_17609,N_5307,N_713);
and U17610 (N_17610,N_2603,N_27);
and U17611 (N_17611,N_3940,N_6408);
and U17612 (N_17612,N_6732,N_9516);
and U17613 (N_17613,N_7091,N_6785);
nand U17614 (N_17614,N_8245,N_5965);
or U17615 (N_17615,N_3450,N_4257);
and U17616 (N_17616,N_4304,N_1528);
nor U17617 (N_17617,N_6416,N_6652);
nor U17618 (N_17618,N_4116,N_8898);
and U17619 (N_17619,N_9422,N_7662);
nor U17620 (N_17620,N_933,N_7079);
nor U17621 (N_17621,N_4645,N_7639);
nor U17622 (N_17622,N_7039,N_1451);
and U17623 (N_17623,N_6872,N_5831);
or U17624 (N_17624,N_859,N_6749);
or U17625 (N_17625,N_3151,N_2788);
nand U17626 (N_17626,N_2915,N_2186);
nor U17627 (N_17627,N_4822,N_632);
and U17628 (N_17628,N_2463,N_7985);
nand U17629 (N_17629,N_5062,N_5092);
nand U17630 (N_17630,N_6053,N_838);
nand U17631 (N_17631,N_5458,N_9943);
and U17632 (N_17632,N_1179,N_4607);
and U17633 (N_17633,N_9451,N_6745);
or U17634 (N_17634,N_2369,N_4583);
xor U17635 (N_17635,N_5075,N_2740);
nor U17636 (N_17636,N_7253,N_9362);
and U17637 (N_17637,N_8004,N_6087);
nor U17638 (N_17638,N_5161,N_89);
nor U17639 (N_17639,N_4263,N_2127);
xnor U17640 (N_17640,N_9373,N_3880);
nor U17641 (N_17641,N_319,N_5470);
nor U17642 (N_17642,N_3738,N_4095);
nand U17643 (N_17643,N_7368,N_6225);
or U17644 (N_17644,N_5267,N_4082);
nor U17645 (N_17645,N_2561,N_5666);
or U17646 (N_17646,N_9142,N_8512);
or U17647 (N_17647,N_3813,N_8559);
or U17648 (N_17648,N_1707,N_2190);
and U17649 (N_17649,N_6074,N_6181);
nor U17650 (N_17650,N_7269,N_2615);
or U17651 (N_17651,N_384,N_769);
nor U17652 (N_17652,N_4198,N_8126);
nor U17653 (N_17653,N_417,N_3214);
xor U17654 (N_17654,N_6717,N_7877);
and U17655 (N_17655,N_5072,N_8866);
nor U17656 (N_17656,N_7677,N_9438);
and U17657 (N_17657,N_5601,N_8461);
xnor U17658 (N_17658,N_8178,N_5576);
nor U17659 (N_17659,N_3091,N_9268);
and U17660 (N_17660,N_5758,N_9326);
nand U17661 (N_17661,N_3478,N_8989);
or U17662 (N_17662,N_2622,N_499);
nand U17663 (N_17663,N_5555,N_8839);
nor U17664 (N_17664,N_5557,N_4144);
or U17665 (N_17665,N_6114,N_8711);
nand U17666 (N_17666,N_3575,N_4433);
nand U17667 (N_17667,N_9468,N_2261);
nand U17668 (N_17668,N_6554,N_1911);
nor U17669 (N_17669,N_9730,N_5602);
nand U17670 (N_17670,N_2121,N_2056);
nor U17671 (N_17671,N_9756,N_1468);
and U17672 (N_17672,N_9588,N_6624);
nor U17673 (N_17673,N_8948,N_3305);
nand U17674 (N_17674,N_5511,N_919);
and U17675 (N_17675,N_3288,N_5125);
nor U17676 (N_17676,N_4694,N_4276);
xnor U17677 (N_17677,N_3477,N_3574);
and U17678 (N_17678,N_4160,N_678);
xor U17679 (N_17679,N_5903,N_610);
and U17680 (N_17680,N_246,N_3207);
or U17681 (N_17681,N_1207,N_2086);
nor U17682 (N_17682,N_1142,N_9915);
nand U17683 (N_17683,N_8122,N_6290);
nand U17684 (N_17684,N_6061,N_4511);
or U17685 (N_17685,N_3130,N_6652);
nand U17686 (N_17686,N_9156,N_3539);
or U17687 (N_17687,N_8062,N_2964);
nor U17688 (N_17688,N_3198,N_7093);
and U17689 (N_17689,N_1008,N_6431);
and U17690 (N_17690,N_2566,N_4718);
or U17691 (N_17691,N_7616,N_310);
and U17692 (N_17692,N_1162,N_2840);
or U17693 (N_17693,N_9654,N_1388);
and U17694 (N_17694,N_3913,N_4975);
and U17695 (N_17695,N_5720,N_4652);
or U17696 (N_17696,N_14,N_6581);
nor U17697 (N_17697,N_8326,N_5129);
or U17698 (N_17698,N_1107,N_2196);
nor U17699 (N_17699,N_3450,N_8572);
xor U17700 (N_17700,N_5198,N_6244);
nand U17701 (N_17701,N_2513,N_9641);
nand U17702 (N_17702,N_2719,N_6833);
nor U17703 (N_17703,N_6819,N_8123);
nor U17704 (N_17704,N_7358,N_4272);
or U17705 (N_17705,N_9369,N_8216);
and U17706 (N_17706,N_1039,N_2050);
xnor U17707 (N_17707,N_5463,N_6990);
and U17708 (N_17708,N_5315,N_716);
and U17709 (N_17709,N_6412,N_6748);
and U17710 (N_17710,N_1214,N_428);
nor U17711 (N_17711,N_6871,N_9741);
or U17712 (N_17712,N_1274,N_7318);
or U17713 (N_17713,N_4657,N_8636);
xor U17714 (N_17714,N_8978,N_9246);
and U17715 (N_17715,N_4864,N_6737);
nand U17716 (N_17716,N_5251,N_3796);
nand U17717 (N_17717,N_855,N_5998);
and U17718 (N_17718,N_9400,N_7125);
or U17719 (N_17719,N_1579,N_3456);
nor U17720 (N_17720,N_5984,N_9053);
nand U17721 (N_17721,N_6734,N_6500);
xnor U17722 (N_17722,N_753,N_1412);
and U17723 (N_17723,N_5964,N_413);
nand U17724 (N_17724,N_8863,N_5626);
nor U17725 (N_17725,N_6416,N_4802);
or U17726 (N_17726,N_3256,N_7941);
nand U17727 (N_17727,N_9064,N_1569);
or U17728 (N_17728,N_9055,N_7252);
nand U17729 (N_17729,N_9817,N_5550);
xor U17730 (N_17730,N_7078,N_6064);
and U17731 (N_17731,N_8455,N_6571);
and U17732 (N_17732,N_3640,N_5026);
nor U17733 (N_17733,N_8276,N_4278);
xor U17734 (N_17734,N_1020,N_5288);
nand U17735 (N_17735,N_9308,N_6994);
and U17736 (N_17736,N_3415,N_3326);
xnor U17737 (N_17737,N_4649,N_647);
nor U17738 (N_17738,N_1324,N_2938);
nand U17739 (N_17739,N_8806,N_9870);
nand U17740 (N_17740,N_3858,N_5313);
or U17741 (N_17741,N_5621,N_5719);
nand U17742 (N_17742,N_4756,N_8986);
and U17743 (N_17743,N_6300,N_3114);
nand U17744 (N_17744,N_4489,N_156);
or U17745 (N_17745,N_4901,N_2912);
xor U17746 (N_17746,N_2260,N_1006);
or U17747 (N_17747,N_9944,N_4739);
xnor U17748 (N_17748,N_761,N_4103);
nand U17749 (N_17749,N_6864,N_2700);
nor U17750 (N_17750,N_577,N_9456);
nor U17751 (N_17751,N_2272,N_2583);
nor U17752 (N_17752,N_9152,N_9015);
xnor U17753 (N_17753,N_5968,N_7373);
and U17754 (N_17754,N_6737,N_8553);
nor U17755 (N_17755,N_3016,N_258);
or U17756 (N_17756,N_5537,N_5757);
and U17757 (N_17757,N_8935,N_1446);
and U17758 (N_17758,N_221,N_6042);
nor U17759 (N_17759,N_9131,N_7991);
and U17760 (N_17760,N_2641,N_1810);
nor U17761 (N_17761,N_8759,N_4579);
nand U17762 (N_17762,N_4616,N_3456);
or U17763 (N_17763,N_7333,N_4391);
xor U17764 (N_17764,N_4361,N_3629);
and U17765 (N_17765,N_5128,N_1720);
and U17766 (N_17766,N_2437,N_8033);
nand U17767 (N_17767,N_2595,N_4477);
nand U17768 (N_17768,N_7177,N_2066);
xnor U17769 (N_17769,N_6238,N_3246);
or U17770 (N_17770,N_3863,N_1913);
or U17771 (N_17771,N_956,N_1443);
or U17772 (N_17772,N_100,N_1775);
or U17773 (N_17773,N_7600,N_5779);
xnor U17774 (N_17774,N_320,N_6914);
nor U17775 (N_17775,N_2910,N_3634);
and U17776 (N_17776,N_2419,N_7842);
nand U17777 (N_17777,N_9074,N_6459);
and U17778 (N_17778,N_3727,N_7716);
nor U17779 (N_17779,N_7246,N_1459);
and U17780 (N_17780,N_5779,N_4507);
nor U17781 (N_17781,N_4232,N_4739);
and U17782 (N_17782,N_5979,N_8464);
or U17783 (N_17783,N_2855,N_3654);
and U17784 (N_17784,N_6470,N_9789);
and U17785 (N_17785,N_1372,N_697);
or U17786 (N_17786,N_7951,N_7981);
and U17787 (N_17787,N_1313,N_4150);
nor U17788 (N_17788,N_6451,N_9406);
xnor U17789 (N_17789,N_9610,N_3333);
nor U17790 (N_17790,N_6106,N_9533);
nor U17791 (N_17791,N_88,N_5157);
or U17792 (N_17792,N_6606,N_2129);
or U17793 (N_17793,N_6630,N_5090);
and U17794 (N_17794,N_9190,N_1101);
or U17795 (N_17795,N_9687,N_4640);
and U17796 (N_17796,N_6669,N_7038);
or U17797 (N_17797,N_8359,N_9119);
nand U17798 (N_17798,N_7548,N_6635);
or U17799 (N_17799,N_9527,N_7991);
nand U17800 (N_17800,N_5481,N_6865);
or U17801 (N_17801,N_8189,N_2255);
nand U17802 (N_17802,N_2660,N_6382);
and U17803 (N_17803,N_8308,N_7801);
and U17804 (N_17804,N_6132,N_2224);
nand U17805 (N_17805,N_8725,N_7576);
and U17806 (N_17806,N_3540,N_1730);
nor U17807 (N_17807,N_9759,N_9235);
xnor U17808 (N_17808,N_4569,N_1296);
nand U17809 (N_17809,N_9184,N_455);
or U17810 (N_17810,N_5566,N_8036);
nand U17811 (N_17811,N_2723,N_7736);
or U17812 (N_17812,N_6887,N_2699);
and U17813 (N_17813,N_3474,N_9962);
nor U17814 (N_17814,N_8555,N_6616);
nor U17815 (N_17815,N_7065,N_6926);
nand U17816 (N_17816,N_5751,N_4999);
or U17817 (N_17817,N_4504,N_1400);
or U17818 (N_17818,N_2258,N_33);
nor U17819 (N_17819,N_6774,N_5742);
and U17820 (N_17820,N_6931,N_7103);
and U17821 (N_17821,N_3256,N_6945);
nand U17822 (N_17822,N_8892,N_9005);
nand U17823 (N_17823,N_8392,N_3276);
nor U17824 (N_17824,N_6650,N_2164);
nor U17825 (N_17825,N_4523,N_7795);
nor U17826 (N_17826,N_7599,N_5325);
xor U17827 (N_17827,N_9270,N_7090);
nor U17828 (N_17828,N_7630,N_2405);
nor U17829 (N_17829,N_5187,N_4670);
and U17830 (N_17830,N_5059,N_4312);
nor U17831 (N_17831,N_2158,N_9911);
nor U17832 (N_17832,N_4835,N_6051);
and U17833 (N_17833,N_7264,N_8921);
nor U17834 (N_17834,N_9504,N_3229);
or U17835 (N_17835,N_7489,N_545);
or U17836 (N_17836,N_2407,N_9633);
and U17837 (N_17837,N_8329,N_2750);
or U17838 (N_17838,N_3248,N_4542);
or U17839 (N_17839,N_3961,N_6747);
nor U17840 (N_17840,N_3400,N_2028);
and U17841 (N_17841,N_9866,N_8958);
xor U17842 (N_17842,N_8485,N_484);
xor U17843 (N_17843,N_6035,N_6942);
or U17844 (N_17844,N_3666,N_3964);
or U17845 (N_17845,N_1787,N_1242);
nand U17846 (N_17846,N_3416,N_9484);
or U17847 (N_17847,N_9166,N_3583);
or U17848 (N_17848,N_3639,N_1061);
or U17849 (N_17849,N_9050,N_1882);
or U17850 (N_17850,N_5295,N_6918);
xor U17851 (N_17851,N_445,N_2773);
and U17852 (N_17852,N_544,N_7651);
and U17853 (N_17853,N_3300,N_6685);
or U17854 (N_17854,N_9435,N_1809);
nor U17855 (N_17855,N_5279,N_1242);
xor U17856 (N_17856,N_3168,N_2564);
and U17857 (N_17857,N_6413,N_1638);
and U17858 (N_17858,N_4596,N_6104);
or U17859 (N_17859,N_2548,N_567);
nor U17860 (N_17860,N_3580,N_9251);
or U17861 (N_17861,N_9258,N_1076);
nand U17862 (N_17862,N_9759,N_426);
or U17863 (N_17863,N_8961,N_6409);
nor U17864 (N_17864,N_2039,N_9742);
xnor U17865 (N_17865,N_2480,N_2211);
and U17866 (N_17866,N_9791,N_3140);
and U17867 (N_17867,N_7394,N_4679);
and U17868 (N_17868,N_6610,N_6691);
nor U17869 (N_17869,N_1725,N_6141);
or U17870 (N_17870,N_9847,N_1711);
or U17871 (N_17871,N_3749,N_2160);
nand U17872 (N_17872,N_3474,N_9925);
or U17873 (N_17873,N_4749,N_9203);
and U17874 (N_17874,N_335,N_7737);
nor U17875 (N_17875,N_3909,N_3265);
or U17876 (N_17876,N_2706,N_8950);
nand U17877 (N_17877,N_9449,N_9242);
xnor U17878 (N_17878,N_3484,N_6760);
xnor U17879 (N_17879,N_1674,N_9442);
nor U17880 (N_17880,N_9756,N_5944);
nor U17881 (N_17881,N_4404,N_612);
or U17882 (N_17882,N_2564,N_1551);
nor U17883 (N_17883,N_2643,N_7218);
xor U17884 (N_17884,N_8511,N_4221);
and U17885 (N_17885,N_7421,N_8175);
nor U17886 (N_17886,N_9552,N_7365);
and U17887 (N_17887,N_2585,N_4100);
or U17888 (N_17888,N_6583,N_3899);
and U17889 (N_17889,N_1364,N_6881);
xnor U17890 (N_17890,N_8610,N_5507);
and U17891 (N_17891,N_4755,N_6023);
and U17892 (N_17892,N_704,N_8229);
nand U17893 (N_17893,N_9894,N_5480);
and U17894 (N_17894,N_5901,N_4231);
nor U17895 (N_17895,N_9504,N_1954);
and U17896 (N_17896,N_8535,N_8360);
nor U17897 (N_17897,N_4754,N_6285);
and U17898 (N_17898,N_4462,N_9749);
or U17899 (N_17899,N_5539,N_4085);
nand U17900 (N_17900,N_3412,N_6998);
xnor U17901 (N_17901,N_1471,N_5331);
or U17902 (N_17902,N_3214,N_8479);
or U17903 (N_17903,N_2281,N_6848);
nand U17904 (N_17904,N_296,N_9478);
nor U17905 (N_17905,N_499,N_1684);
xnor U17906 (N_17906,N_7366,N_4044);
xor U17907 (N_17907,N_822,N_3201);
or U17908 (N_17908,N_9700,N_4728);
and U17909 (N_17909,N_6393,N_8066);
or U17910 (N_17910,N_3827,N_8273);
xnor U17911 (N_17911,N_3128,N_3125);
nor U17912 (N_17912,N_747,N_1791);
or U17913 (N_17913,N_2354,N_415);
nor U17914 (N_17914,N_250,N_2580);
nor U17915 (N_17915,N_1402,N_9070);
or U17916 (N_17916,N_1962,N_8917);
or U17917 (N_17917,N_9244,N_6009);
nor U17918 (N_17918,N_3658,N_5839);
nor U17919 (N_17919,N_4811,N_2386);
or U17920 (N_17920,N_7849,N_955);
or U17921 (N_17921,N_2994,N_5145);
and U17922 (N_17922,N_1099,N_1414);
and U17923 (N_17923,N_7918,N_2610);
or U17924 (N_17924,N_8225,N_4778);
nor U17925 (N_17925,N_3012,N_8880);
nor U17926 (N_17926,N_4293,N_8907);
and U17927 (N_17927,N_3554,N_728);
and U17928 (N_17928,N_6574,N_5668);
nor U17929 (N_17929,N_4255,N_8103);
or U17930 (N_17930,N_4952,N_5862);
nor U17931 (N_17931,N_7822,N_1767);
or U17932 (N_17932,N_8456,N_2820);
xor U17933 (N_17933,N_6081,N_2735);
nand U17934 (N_17934,N_6960,N_2258);
and U17935 (N_17935,N_9368,N_2229);
xnor U17936 (N_17936,N_3677,N_9069);
or U17937 (N_17937,N_1185,N_9422);
xnor U17938 (N_17938,N_2064,N_3535);
nand U17939 (N_17939,N_1598,N_862);
nor U17940 (N_17940,N_122,N_4179);
nand U17941 (N_17941,N_5034,N_4402);
or U17942 (N_17942,N_9775,N_3844);
nand U17943 (N_17943,N_7878,N_4468);
nor U17944 (N_17944,N_2149,N_4513);
nor U17945 (N_17945,N_6911,N_812);
or U17946 (N_17946,N_3651,N_3862);
nand U17947 (N_17947,N_9399,N_7061);
and U17948 (N_17948,N_1055,N_314);
and U17949 (N_17949,N_3748,N_8354);
nor U17950 (N_17950,N_4758,N_1117);
or U17951 (N_17951,N_9432,N_6153);
nand U17952 (N_17952,N_5402,N_2308);
and U17953 (N_17953,N_9429,N_7463);
xor U17954 (N_17954,N_2228,N_6011);
or U17955 (N_17955,N_4781,N_4169);
nand U17956 (N_17956,N_2564,N_5059);
nand U17957 (N_17957,N_386,N_9111);
or U17958 (N_17958,N_9084,N_4970);
xor U17959 (N_17959,N_1,N_6958);
nor U17960 (N_17960,N_7334,N_9747);
nand U17961 (N_17961,N_1450,N_5236);
and U17962 (N_17962,N_238,N_1711);
or U17963 (N_17963,N_6816,N_8590);
nor U17964 (N_17964,N_912,N_4704);
and U17965 (N_17965,N_3943,N_6776);
or U17966 (N_17966,N_9087,N_8382);
nor U17967 (N_17967,N_7380,N_1417);
nand U17968 (N_17968,N_8753,N_9281);
xor U17969 (N_17969,N_4967,N_1260);
xor U17970 (N_17970,N_9047,N_2980);
nor U17971 (N_17971,N_3127,N_3839);
and U17972 (N_17972,N_5241,N_4460);
nand U17973 (N_17973,N_2179,N_9224);
nand U17974 (N_17974,N_8051,N_5460);
nand U17975 (N_17975,N_8460,N_1269);
or U17976 (N_17976,N_2760,N_4363);
or U17977 (N_17977,N_1302,N_2423);
and U17978 (N_17978,N_2947,N_143);
and U17979 (N_17979,N_842,N_1525);
or U17980 (N_17980,N_4018,N_6233);
nor U17981 (N_17981,N_2488,N_2907);
or U17982 (N_17982,N_6451,N_5398);
nand U17983 (N_17983,N_1879,N_8815);
nand U17984 (N_17984,N_8823,N_3003);
and U17985 (N_17985,N_8462,N_8970);
nor U17986 (N_17986,N_2923,N_1554);
nor U17987 (N_17987,N_483,N_5622);
or U17988 (N_17988,N_7474,N_576);
or U17989 (N_17989,N_7940,N_1774);
xor U17990 (N_17990,N_6441,N_9754);
and U17991 (N_17991,N_1501,N_5190);
xor U17992 (N_17992,N_6820,N_5618);
and U17993 (N_17993,N_9692,N_4761);
or U17994 (N_17994,N_7765,N_5753);
nor U17995 (N_17995,N_7588,N_9930);
or U17996 (N_17996,N_680,N_9310);
nor U17997 (N_17997,N_7834,N_5792);
nand U17998 (N_17998,N_1885,N_195);
nand U17999 (N_17999,N_3916,N_7139);
nand U18000 (N_18000,N_9921,N_7308);
nand U18001 (N_18001,N_6409,N_6327);
nand U18002 (N_18002,N_4679,N_2942);
or U18003 (N_18003,N_4527,N_844);
and U18004 (N_18004,N_4866,N_8762);
and U18005 (N_18005,N_9128,N_490);
and U18006 (N_18006,N_8574,N_1865);
and U18007 (N_18007,N_4861,N_7645);
or U18008 (N_18008,N_7083,N_3206);
and U18009 (N_18009,N_5099,N_1883);
nor U18010 (N_18010,N_751,N_473);
xnor U18011 (N_18011,N_8834,N_6847);
and U18012 (N_18012,N_1620,N_6816);
nand U18013 (N_18013,N_2166,N_8635);
and U18014 (N_18014,N_4013,N_4428);
xnor U18015 (N_18015,N_249,N_3711);
and U18016 (N_18016,N_2287,N_1295);
or U18017 (N_18017,N_183,N_9249);
nand U18018 (N_18018,N_519,N_1032);
nand U18019 (N_18019,N_9442,N_4043);
and U18020 (N_18020,N_1451,N_3425);
and U18021 (N_18021,N_6,N_5875);
nor U18022 (N_18022,N_7285,N_1975);
or U18023 (N_18023,N_6315,N_2609);
nand U18024 (N_18024,N_1788,N_9831);
and U18025 (N_18025,N_6240,N_1573);
nor U18026 (N_18026,N_8807,N_9349);
nand U18027 (N_18027,N_5718,N_4015);
nor U18028 (N_18028,N_9851,N_8980);
or U18029 (N_18029,N_9994,N_9556);
and U18030 (N_18030,N_5291,N_1451);
nand U18031 (N_18031,N_6416,N_2053);
nor U18032 (N_18032,N_3400,N_8011);
nor U18033 (N_18033,N_1312,N_594);
nor U18034 (N_18034,N_1574,N_3421);
nand U18035 (N_18035,N_7005,N_7129);
and U18036 (N_18036,N_3401,N_3594);
or U18037 (N_18037,N_3833,N_367);
or U18038 (N_18038,N_3666,N_9179);
nor U18039 (N_18039,N_8779,N_2255);
nand U18040 (N_18040,N_9428,N_1065);
nand U18041 (N_18041,N_322,N_4426);
nand U18042 (N_18042,N_4288,N_3313);
nor U18043 (N_18043,N_2921,N_4972);
xnor U18044 (N_18044,N_8129,N_4540);
xnor U18045 (N_18045,N_9712,N_4760);
or U18046 (N_18046,N_7259,N_5621);
nand U18047 (N_18047,N_3386,N_6515);
nand U18048 (N_18048,N_4513,N_3078);
nand U18049 (N_18049,N_1285,N_187);
nor U18050 (N_18050,N_4535,N_552);
nor U18051 (N_18051,N_1510,N_1250);
and U18052 (N_18052,N_9712,N_3299);
or U18053 (N_18053,N_7941,N_8239);
nand U18054 (N_18054,N_9603,N_5543);
and U18055 (N_18055,N_2194,N_4036);
xor U18056 (N_18056,N_6270,N_7005);
nor U18057 (N_18057,N_356,N_8056);
xor U18058 (N_18058,N_7425,N_9183);
and U18059 (N_18059,N_1227,N_7525);
and U18060 (N_18060,N_5912,N_8266);
nand U18061 (N_18061,N_6863,N_844);
nor U18062 (N_18062,N_547,N_9941);
and U18063 (N_18063,N_3889,N_4136);
or U18064 (N_18064,N_6222,N_7915);
and U18065 (N_18065,N_9134,N_8418);
and U18066 (N_18066,N_7531,N_9369);
xor U18067 (N_18067,N_7974,N_9550);
or U18068 (N_18068,N_6847,N_6964);
nand U18069 (N_18069,N_3590,N_2750);
nand U18070 (N_18070,N_368,N_1441);
and U18071 (N_18071,N_5883,N_8614);
nor U18072 (N_18072,N_1797,N_7552);
nand U18073 (N_18073,N_3634,N_2671);
nor U18074 (N_18074,N_2165,N_1602);
nand U18075 (N_18075,N_2626,N_2268);
and U18076 (N_18076,N_6369,N_8802);
nand U18077 (N_18077,N_1600,N_2879);
or U18078 (N_18078,N_6007,N_7118);
or U18079 (N_18079,N_1734,N_207);
xnor U18080 (N_18080,N_8273,N_8684);
and U18081 (N_18081,N_8273,N_2947);
nand U18082 (N_18082,N_8265,N_6173);
xnor U18083 (N_18083,N_2074,N_1344);
and U18084 (N_18084,N_3094,N_7748);
nand U18085 (N_18085,N_8180,N_6953);
or U18086 (N_18086,N_9172,N_599);
nor U18087 (N_18087,N_1462,N_6196);
nor U18088 (N_18088,N_8619,N_7887);
or U18089 (N_18089,N_27,N_2070);
nor U18090 (N_18090,N_5142,N_2506);
nand U18091 (N_18091,N_4198,N_9198);
xor U18092 (N_18092,N_8727,N_6525);
or U18093 (N_18093,N_3202,N_3068);
nand U18094 (N_18094,N_201,N_7622);
xnor U18095 (N_18095,N_4873,N_7975);
and U18096 (N_18096,N_9520,N_393);
nand U18097 (N_18097,N_7446,N_4108);
or U18098 (N_18098,N_2186,N_2173);
nor U18099 (N_18099,N_4199,N_9627);
nand U18100 (N_18100,N_7514,N_6680);
nor U18101 (N_18101,N_2167,N_9672);
nor U18102 (N_18102,N_9203,N_6603);
or U18103 (N_18103,N_3097,N_3285);
and U18104 (N_18104,N_1583,N_5906);
and U18105 (N_18105,N_5655,N_1616);
or U18106 (N_18106,N_2943,N_8870);
nor U18107 (N_18107,N_8124,N_3846);
or U18108 (N_18108,N_6608,N_1929);
or U18109 (N_18109,N_1483,N_4745);
or U18110 (N_18110,N_3407,N_7438);
nand U18111 (N_18111,N_684,N_7017);
and U18112 (N_18112,N_2812,N_7628);
and U18113 (N_18113,N_6842,N_2209);
or U18114 (N_18114,N_2966,N_9017);
or U18115 (N_18115,N_7762,N_2784);
xor U18116 (N_18116,N_5843,N_1387);
or U18117 (N_18117,N_2799,N_463);
nor U18118 (N_18118,N_7919,N_6339);
and U18119 (N_18119,N_807,N_9968);
or U18120 (N_18120,N_1843,N_1531);
nand U18121 (N_18121,N_7659,N_4594);
nor U18122 (N_18122,N_921,N_4870);
and U18123 (N_18123,N_96,N_7834);
xnor U18124 (N_18124,N_4425,N_1116);
nor U18125 (N_18125,N_4391,N_7957);
or U18126 (N_18126,N_6639,N_7411);
nand U18127 (N_18127,N_6500,N_8938);
nand U18128 (N_18128,N_5059,N_4757);
or U18129 (N_18129,N_7849,N_5380);
or U18130 (N_18130,N_2178,N_3452);
or U18131 (N_18131,N_4755,N_6736);
and U18132 (N_18132,N_850,N_7853);
and U18133 (N_18133,N_5789,N_1709);
nand U18134 (N_18134,N_6562,N_2051);
or U18135 (N_18135,N_1416,N_4193);
and U18136 (N_18136,N_1811,N_6094);
nor U18137 (N_18137,N_8548,N_6704);
nor U18138 (N_18138,N_570,N_5634);
or U18139 (N_18139,N_2006,N_4758);
nand U18140 (N_18140,N_8250,N_5551);
nor U18141 (N_18141,N_8382,N_3795);
or U18142 (N_18142,N_4980,N_4087);
and U18143 (N_18143,N_633,N_8937);
or U18144 (N_18144,N_6794,N_9397);
and U18145 (N_18145,N_7204,N_7812);
and U18146 (N_18146,N_3219,N_1766);
nand U18147 (N_18147,N_2788,N_2531);
or U18148 (N_18148,N_3582,N_131);
xnor U18149 (N_18149,N_7578,N_8121);
and U18150 (N_18150,N_7632,N_8792);
nor U18151 (N_18151,N_3906,N_3031);
and U18152 (N_18152,N_6856,N_4821);
nand U18153 (N_18153,N_9751,N_1267);
xor U18154 (N_18154,N_1975,N_1155);
or U18155 (N_18155,N_4500,N_9957);
nor U18156 (N_18156,N_3228,N_4094);
or U18157 (N_18157,N_2083,N_4137);
xor U18158 (N_18158,N_8449,N_1590);
nor U18159 (N_18159,N_7839,N_9565);
or U18160 (N_18160,N_3473,N_2540);
nor U18161 (N_18161,N_5953,N_36);
nor U18162 (N_18162,N_7051,N_1330);
or U18163 (N_18163,N_226,N_9342);
and U18164 (N_18164,N_242,N_959);
and U18165 (N_18165,N_3143,N_8044);
nand U18166 (N_18166,N_9150,N_2640);
or U18167 (N_18167,N_6523,N_5017);
or U18168 (N_18168,N_1981,N_4373);
nand U18169 (N_18169,N_8499,N_9922);
and U18170 (N_18170,N_7001,N_9827);
and U18171 (N_18171,N_7707,N_3203);
or U18172 (N_18172,N_5692,N_4978);
nor U18173 (N_18173,N_9134,N_984);
nor U18174 (N_18174,N_1167,N_8629);
or U18175 (N_18175,N_9223,N_4345);
and U18176 (N_18176,N_6736,N_7542);
nand U18177 (N_18177,N_9788,N_545);
nor U18178 (N_18178,N_6836,N_5151);
xor U18179 (N_18179,N_224,N_5873);
and U18180 (N_18180,N_1769,N_8994);
or U18181 (N_18181,N_6841,N_7239);
nor U18182 (N_18182,N_2649,N_897);
xor U18183 (N_18183,N_5464,N_9755);
nand U18184 (N_18184,N_9986,N_4954);
and U18185 (N_18185,N_7808,N_8594);
and U18186 (N_18186,N_4781,N_6319);
nor U18187 (N_18187,N_3486,N_8772);
nor U18188 (N_18188,N_2322,N_6682);
xor U18189 (N_18189,N_9078,N_9661);
and U18190 (N_18190,N_9212,N_5441);
xor U18191 (N_18191,N_4422,N_4449);
nor U18192 (N_18192,N_697,N_2071);
and U18193 (N_18193,N_4464,N_496);
nand U18194 (N_18194,N_305,N_7070);
or U18195 (N_18195,N_6513,N_6434);
nor U18196 (N_18196,N_4335,N_3287);
and U18197 (N_18197,N_6677,N_3614);
xnor U18198 (N_18198,N_2380,N_5732);
nand U18199 (N_18199,N_5727,N_2258);
and U18200 (N_18200,N_2050,N_1629);
nand U18201 (N_18201,N_8952,N_6181);
nor U18202 (N_18202,N_154,N_1020);
or U18203 (N_18203,N_7353,N_3495);
nand U18204 (N_18204,N_2894,N_9801);
nor U18205 (N_18205,N_9901,N_4689);
nor U18206 (N_18206,N_9790,N_670);
and U18207 (N_18207,N_7411,N_9334);
nor U18208 (N_18208,N_1959,N_2860);
nor U18209 (N_18209,N_4104,N_9620);
nand U18210 (N_18210,N_9180,N_9238);
or U18211 (N_18211,N_2374,N_9472);
xnor U18212 (N_18212,N_6066,N_2568);
nor U18213 (N_18213,N_4807,N_3895);
and U18214 (N_18214,N_8560,N_6008);
xor U18215 (N_18215,N_9712,N_9764);
nand U18216 (N_18216,N_5422,N_5902);
and U18217 (N_18217,N_405,N_8926);
and U18218 (N_18218,N_1974,N_2487);
nand U18219 (N_18219,N_6822,N_1376);
and U18220 (N_18220,N_9280,N_3042);
and U18221 (N_18221,N_6425,N_7952);
nand U18222 (N_18222,N_461,N_6847);
nor U18223 (N_18223,N_9153,N_7217);
and U18224 (N_18224,N_5366,N_7067);
or U18225 (N_18225,N_9866,N_6040);
nor U18226 (N_18226,N_5619,N_4924);
nor U18227 (N_18227,N_7697,N_3500);
nor U18228 (N_18228,N_6116,N_5060);
or U18229 (N_18229,N_2225,N_4357);
nor U18230 (N_18230,N_5226,N_7768);
or U18231 (N_18231,N_4853,N_9724);
and U18232 (N_18232,N_9685,N_5865);
or U18233 (N_18233,N_3070,N_355);
nand U18234 (N_18234,N_1451,N_687);
or U18235 (N_18235,N_489,N_8851);
nand U18236 (N_18236,N_6443,N_4094);
or U18237 (N_18237,N_9471,N_5382);
and U18238 (N_18238,N_5568,N_7779);
and U18239 (N_18239,N_1106,N_367);
nand U18240 (N_18240,N_2052,N_4712);
or U18241 (N_18241,N_9865,N_2625);
or U18242 (N_18242,N_6237,N_2775);
and U18243 (N_18243,N_6292,N_2109);
nor U18244 (N_18244,N_9908,N_7712);
and U18245 (N_18245,N_3312,N_6075);
nand U18246 (N_18246,N_1920,N_4959);
nand U18247 (N_18247,N_9164,N_692);
or U18248 (N_18248,N_8009,N_8180);
nand U18249 (N_18249,N_2040,N_843);
nand U18250 (N_18250,N_2233,N_562);
and U18251 (N_18251,N_615,N_1242);
xnor U18252 (N_18252,N_2249,N_9197);
nor U18253 (N_18253,N_8114,N_4473);
or U18254 (N_18254,N_9652,N_9229);
or U18255 (N_18255,N_8698,N_5375);
nand U18256 (N_18256,N_7910,N_4353);
and U18257 (N_18257,N_6668,N_1830);
xor U18258 (N_18258,N_3146,N_7029);
nand U18259 (N_18259,N_4586,N_7844);
and U18260 (N_18260,N_3243,N_8714);
nor U18261 (N_18261,N_796,N_2756);
nand U18262 (N_18262,N_9699,N_1502);
nand U18263 (N_18263,N_702,N_8557);
nor U18264 (N_18264,N_1838,N_3649);
and U18265 (N_18265,N_3121,N_3214);
or U18266 (N_18266,N_28,N_8078);
nor U18267 (N_18267,N_9133,N_6564);
nor U18268 (N_18268,N_2599,N_4533);
nor U18269 (N_18269,N_9405,N_4675);
and U18270 (N_18270,N_6706,N_9437);
and U18271 (N_18271,N_3494,N_7823);
nand U18272 (N_18272,N_9860,N_1216);
or U18273 (N_18273,N_4764,N_715);
nor U18274 (N_18274,N_2546,N_8379);
and U18275 (N_18275,N_2236,N_1844);
nand U18276 (N_18276,N_3555,N_488);
nor U18277 (N_18277,N_6117,N_89);
nor U18278 (N_18278,N_7700,N_6771);
and U18279 (N_18279,N_6763,N_7842);
and U18280 (N_18280,N_4993,N_1204);
nand U18281 (N_18281,N_1504,N_6170);
or U18282 (N_18282,N_5564,N_2825);
or U18283 (N_18283,N_4400,N_3899);
nor U18284 (N_18284,N_258,N_2230);
nor U18285 (N_18285,N_1681,N_2433);
and U18286 (N_18286,N_3970,N_2924);
and U18287 (N_18287,N_3992,N_9846);
and U18288 (N_18288,N_1885,N_911);
and U18289 (N_18289,N_6493,N_2775);
and U18290 (N_18290,N_9907,N_4158);
nand U18291 (N_18291,N_8102,N_5836);
or U18292 (N_18292,N_3082,N_250);
xor U18293 (N_18293,N_3462,N_1703);
nor U18294 (N_18294,N_8380,N_8847);
nor U18295 (N_18295,N_774,N_9024);
nor U18296 (N_18296,N_3177,N_8520);
and U18297 (N_18297,N_3885,N_7882);
nor U18298 (N_18298,N_6889,N_2803);
or U18299 (N_18299,N_5612,N_7259);
or U18300 (N_18300,N_1147,N_2124);
or U18301 (N_18301,N_3247,N_7802);
nor U18302 (N_18302,N_8347,N_9852);
nand U18303 (N_18303,N_6061,N_5912);
nor U18304 (N_18304,N_9456,N_4679);
nor U18305 (N_18305,N_4190,N_8590);
nand U18306 (N_18306,N_0,N_566);
or U18307 (N_18307,N_1666,N_8241);
or U18308 (N_18308,N_7212,N_4486);
or U18309 (N_18309,N_2782,N_5607);
nor U18310 (N_18310,N_9823,N_596);
nor U18311 (N_18311,N_8843,N_2413);
or U18312 (N_18312,N_761,N_2808);
and U18313 (N_18313,N_6873,N_1586);
and U18314 (N_18314,N_4353,N_197);
and U18315 (N_18315,N_1316,N_4218);
nand U18316 (N_18316,N_4641,N_4279);
or U18317 (N_18317,N_4875,N_5054);
or U18318 (N_18318,N_5683,N_3397);
xnor U18319 (N_18319,N_9800,N_9852);
and U18320 (N_18320,N_3719,N_3849);
xor U18321 (N_18321,N_3186,N_7570);
nand U18322 (N_18322,N_5763,N_8245);
nor U18323 (N_18323,N_5296,N_4009);
or U18324 (N_18324,N_1411,N_5395);
nor U18325 (N_18325,N_1497,N_6244);
and U18326 (N_18326,N_4836,N_2990);
nand U18327 (N_18327,N_2398,N_5099);
and U18328 (N_18328,N_3904,N_4909);
and U18329 (N_18329,N_8168,N_3113);
or U18330 (N_18330,N_5273,N_4431);
nor U18331 (N_18331,N_4514,N_7121);
and U18332 (N_18332,N_7455,N_7473);
or U18333 (N_18333,N_5446,N_2423);
nor U18334 (N_18334,N_673,N_4094);
and U18335 (N_18335,N_5354,N_9721);
nor U18336 (N_18336,N_3583,N_6260);
nand U18337 (N_18337,N_9735,N_5422);
nor U18338 (N_18338,N_2337,N_9448);
and U18339 (N_18339,N_5904,N_677);
nand U18340 (N_18340,N_4548,N_6550);
nor U18341 (N_18341,N_2060,N_9984);
and U18342 (N_18342,N_9137,N_7624);
xor U18343 (N_18343,N_5434,N_501);
nand U18344 (N_18344,N_3057,N_609);
nor U18345 (N_18345,N_6585,N_3988);
nand U18346 (N_18346,N_2211,N_1162);
nand U18347 (N_18347,N_6109,N_1455);
or U18348 (N_18348,N_1942,N_7944);
and U18349 (N_18349,N_6546,N_784);
nand U18350 (N_18350,N_1486,N_4115);
xnor U18351 (N_18351,N_3955,N_9895);
or U18352 (N_18352,N_6280,N_9034);
and U18353 (N_18353,N_1510,N_4142);
xnor U18354 (N_18354,N_5149,N_8303);
or U18355 (N_18355,N_9019,N_3231);
and U18356 (N_18356,N_897,N_5265);
and U18357 (N_18357,N_5357,N_9585);
and U18358 (N_18358,N_9647,N_2706);
or U18359 (N_18359,N_9730,N_7029);
and U18360 (N_18360,N_409,N_405);
or U18361 (N_18361,N_3530,N_2386);
xor U18362 (N_18362,N_5690,N_7071);
nand U18363 (N_18363,N_8908,N_6728);
xor U18364 (N_18364,N_1782,N_5258);
or U18365 (N_18365,N_3921,N_1877);
and U18366 (N_18366,N_1533,N_1183);
nand U18367 (N_18367,N_2814,N_73);
or U18368 (N_18368,N_4793,N_38);
and U18369 (N_18369,N_9295,N_7772);
or U18370 (N_18370,N_3298,N_5743);
nand U18371 (N_18371,N_6864,N_2333);
and U18372 (N_18372,N_4853,N_5591);
nand U18373 (N_18373,N_4334,N_669);
nand U18374 (N_18374,N_6851,N_1755);
nand U18375 (N_18375,N_3843,N_8663);
and U18376 (N_18376,N_4757,N_1687);
and U18377 (N_18377,N_9444,N_4606);
and U18378 (N_18378,N_4085,N_676);
nand U18379 (N_18379,N_2605,N_7834);
or U18380 (N_18380,N_9757,N_4057);
nor U18381 (N_18381,N_5291,N_7996);
nand U18382 (N_18382,N_9106,N_3095);
nor U18383 (N_18383,N_3682,N_6081);
nand U18384 (N_18384,N_2197,N_4900);
xor U18385 (N_18385,N_653,N_5905);
and U18386 (N_18386,N_2224,N_734);
nor U18387 (N_18387,N_5378,N_3470);
nand U18388 (N_18388,N_1552,N_4321);
nand U18389 (N_18389,N_1949,N_3412);
or U18390 (N_18390,N_351,N_2658);
nand U18391 (N_18391,N_9691,N_4100);
or U18392 (N_18392,N_2002,N_6154);
nor U18393 (N_18393,N_8575,N_6304);
nor U18394 (N_18394,N_6750,N_3870);
or U18395 (N_18395,N_322,N_8119);
nand U18396 (N_18396,N_9479,N_956);
or U18397 (N_18397,N_1290,N_1495);
nand U18398 (N_18398,N_2824,N_7953);
xnor U18399 (N_18399,N_3698,N_8336);
xor U18400 (N_18400,N_3476,N_5927);
nor U18401 (N_18401,N_4998,N_3655);
and U18402 (N_18402,N_4219,N_2658);
and U18403 (N_18403,N_997,N_8949);
or U18404 (N_18404,N_4181,N_237);
nor U18405 (N_18405,N_5618,N_387);
or U18406 (N_18406,N_6407,N_9404);
and U18407 (N_18407,N_4099,N_2503);
and U18408 (N_18408,N_644,N_3818);
and U18409 (N_18409,N_5749,N_3237);
nand U18410 (N_18410,N_9580,N_3350);
and U18411 (N_18411,N_5142,N_5818);
nor U18412 (N_18412,N_2897,N_355);
and U18413 (N_18413,N_5809,N_3383);
nand U18414 (N_18414,N_3526,N_9941);
and U18415 (N_18415,N_2490,N_1082);
and U18416 (N_18416,N_250,N_4540);
nand U18417 (N_18417,N_1601,N_6026);
nor U18418 (N_18418,N_5615,N_8487);
or U18419 (N_18419,N_8679,N_1680);
nor U18420 (N_18420,N_5407,N_4979);
nor U18421 (N_18421,N_5771,N_4825);
and U18422 (N_18422,N_7686,N_6316);
or U18423 (N_18423,N_9847,N_7410);
nand U18424 (N_18424,N_9914,N_5266);
or U18425 (N_18425,N_5045,N_7408);
nand U18426 (N_18426,N_1257,N_2511);
nor U18427 (N_18427,N_6338,N_7273);
nand U18428 (N_18428,N_9208,N_1842);
and U18429 (N_18429,N_7608,N_3722);
or U18430 (N_18430,N_771,N_1747);
xor U18431 (N_18431,N_5917,N_3692);
nor U18432 (N_18432,N_5205,N_961);
nand U18433 (N_18433,N_921,N_6565);
nor U18434 (N_18434,N_8453,N_1021);
and U18435 (N_18435,N_2604,N_8657);
nor U18436 (N_18436,N_2724,N_8465);
nand U18437 (N_18437,N_5630,N_2787);
and U18438 (N_18438,N_1391,N_8366);
nand U18439 (N_18439,N_4957,N_2919);
nand U18440 (N_18440,N_1600,N_5218);
and U18441 (N_18441,N_3903,N_6464);
nand U18442 (N_18442,N_4347,N_7691);
nand U18443 (N_18443,N_6899,N_7393);
or U18444 (N_18444,N_8432,N_2911);
or U18445 (N_18445,N_3848,N_3333);
nand U18446 (N_18446,N_3923,N_278);
nor U18447 (N_18447,N_7854,N_7690);
or U18448 (N_18448,N_7216,N_2220);
nand U18449 (N_18449,N_8213,N_5069);
nor U18450 (N_18450,N_2711,N_5474);
nand U18451 (N_18451,N_8076,N_8451);
and U18452 (N_18452,N_2076,N_2822);
or U18453 (N_18453,N_6127,N_2629);
nand U18454 (N_18454,N_5258,N_4534);
nand U18455 (N_18455,N_5721,N_5409);
or U18456 (N_18456,N_6088,N_5749);
and U18457 (N_18457,N_3932,N_4756);
or U18458 (N_18458,N_1763,N_8198);
nand U18459 (N_18459,N_8473,N_4764);
nor U18460 (N_18460,N_6792,N_4427);
or U18461 (N_18461,N_2721,N_6760);
nor U18462 (N_18462,N_9284,N_923);
nor U18463 (N_18463,N_7892,N_7334);
or U18464 (N_18464,N_4352,N_8207);
nor U18465 (N_18465,N_1739,N_441);
and U18466 (N_18466,N_2820,N_8053);
and U18467 (N_18467,N_6142,N_1733);
nor U18468 (N_18468,N_8495,N_6118);
nor U18469 (N_18469,N_7328,N_446);
or U18470 (N_18470,N_8527,N_7477);
nor U18471 (N_18471,N_2523,N_3139);
and U18472 (N_18472,N_1845,N_5350);
and U18473 (N_18473,N_8163,N_1086);
and U18474 (N_18474,N_7778,N_4312);
nor U18475 (N_18475,N_6527,N_9939);
and U18476 (N_18476,N_3927,N_2798);
and U18477 (N_18477,N_7099,N_5355);
nor U18478 (N_18478,N_3688,N_6098);
nor U18479 (N_18479,N_6464,N_6413);
or U18480 (N_18480,N_6185,N_2491);
or U18481 (N_18481,N_3052,N_4040);
nand U18482 (N_18482,N_2516,N_3341);
nor U18483 (N_18483,N_8206,N_1458);
nor U18484 (N_18484,N_4064,N_7378);
or U18485 (N_18485,N_8872,N_861);
or U18486 (N_18486,N_7477,N_450);
xor U18487 (N_18487,N_5607,N_8519);
or U18488 (N_18488,N_3018,N_6611);
nor U18489 (N_18489,N_8033,N_6279);
nor U18490 (N_18490,N_6299,N_5438);
nand U18491 (N_18491,N_5,N_6439);
nand U18492 (N_18492,N_3150,N_4978);
nand U18493 (N_18493,N_2979,N_8550);
nor U18494 (N_18494,N_6905,N_5248);
and U18495 (N_18495,N_2446,N_8777);
xnor U18496 (N_18496,N_3246,N_8811);
nor U18497 (N_18497,N_9843,N_9611);
xor U18498 (N_18498,N_9693,N_897);
and U18499 (N_18499,N_3625,N_3652);
and U18500 (N_18500,N_4078,N_7998);
and U18501 (N_18501,N_5322,N_9997);
and U18502 (N_18502,N_1898,N_9244);
nand U18503 (N_18503,N_4527,N_5919);
nand U18504 (N_18504,N_1746,N_7600);
and U18505 (N_18505,N_2579,N_8000);
and U18506 (N_18506,N_5236,N_8166);
xor U18507 (N_18507,N_6355,N_5222);
nand U18508 (N_18508,N_500,N_3951);
nor U18509 (N_18509,N_9217,N_1345);
or U18510 (N_18510,N_4401,N_5928);
xnor U18511 (N_18511,N_4367,N_795);
nor U18512 (N_18512,N_4746,N_5114);
or U18513 (N_18513,N_9621,N_1596);
xor U18514 (N_18514,N_4643,N_3463);
nor U18515 (N_18515,N_1969,N_5169);
xor U18516 (N_18516,N_5783,N_4216);
xnor U18517 (N_18517,N_7923,N_6122);
nand U18518 (N_18518,N_5070,N_7751);
and U18519 (N_18519,N_954,N_4903);
nand U18520 (N_18520,N_2090,N_4883);
or U18521 (N_18521,N_7076,N_3382);
nand U18522 (N_18522,N_7398,N_9639);
and U18523 (N_18523,N_9771,N_3159);
or U18524 (N_18524,N_7381,N_9132);
nand U18525 (N_18525,N_4079,N_770);
and U18526 (N_18526,N_984,N_9038);
nand U18527 (N_18527,N_7324,N_9177);
nor U18528 (N_18528,N_6600,N_3072);
and U18529 (N_18529,N_8778,N_5790);
xor U18530 (N_18530,N_2245,N_5302);
and U18531 (N_18531,N_975,N_6831);
or U18532 (N_18532,N_3862,N_9801);
and U18533 (N_18533,N_6007,N_7651);
nor U18534 (N_18534,N_8754,N_2791);
xnor U18535 (N_18535,N_6446,N_8931);
and U18536 (N_18536,N_462,N_7910);
nor U18537 (N_18537,N_1591,N_145);
and U18538 (N_18538,N_3258,N_6384);
nor U18539 (N_18539,N_4151,N_455);
and U18540 (N_18540,N_8776,N_7005);
or U18541 (N_18541,N_8815,N_1891);
nor U18542 (N_18542,N_1926,N_3687);
nor U18543 (N_18543,N_3863,N_2176);
and U18544 (N_18544,N_5373,N_6608);
nand U18545 (N_18545,N_6893,N_3363);
nor U18546 (N_18546,N_6246,N_6679);
and U18547 (N_18547,N_6282,N_2804);
and U18548 (N_18548,N_825,N_4082);
and U18549 (N_18549,N_7837,N_5224);
and U18550 (N_18550,N_5941,N_5074);
or U18551 (N_18551,N_4657,N_3493);
nor U18552 (N_18552,N_6003,N_8805);
xnor U18553 (N_18553,N_1075,N_29);
nand U18554 (N_18554,N_232,N_4108);
xor U18555 (N_18555,N_1788,N_8312);
nor U18556 (N_18556,N_7500,N_3822);
or U18557 (N_18557,N_2858,N_3262);
and U18558 (N_18558,N_3572,N_5548);
nor U18559 (N_18559,N_5300,N_8813);
nor U18560 (N_18560,N_3277,N_4371);
nand U18561 (N_18561,N_5926,N_2368);
xnor U18562 (N_18562,N_4915,N_8918);
nand U18563 (N_18563,N_920,N_6724);
nor U18564 (N_18564,N_434,N_3734);
xnor U18565 (N_18565,N_1557,N_1371);
or U18566 (N_18566,N_3182,N_4600);
or U18567 (N_18567,N_2100,N_7285);
nand U18568 (N_18568,N_2599,N_4001);
and U18569 (N_18569,N_8271,N_3059);
nor U18570 (N_18570,N_5603,N_5247);
nand U18571 (N_18571,N_4548,N_2964);
or U18572 (N_18572,N_6718,N_4069);
nand U18573 (N_18573,N_9936,N_9625);
nor U18574 (N_18574,N_4473,N_7900);
nor U18575 (N_18575,N_6638,N_9901);
xor U18576 (N_18576,N_6703,N_8447);
or U18577 (N_18577,N_3520,N_178);
nor U18578 (N_18578,N_764,N_3926);
nor U18579 (N_18579,N_2734,N_7839);
or U18580 (N_18580,N_2637,N_1588);
xor U18581 (N_18581,N_1914,N_2024);
nor U18582 (N_18582,N_5172,N_7027);
xnor U18583 (N_18583,N_7862,N_9054);
nand U18584 (N_18584,N_8987,N_1116);
nand U18585 (N_18585,N_4689,N_5698);
and U18586 (N_18586,N_5225,N_4808);
nor U18587 (N_18587,N_9649,N_1377);
nor U18588 (N_18588,N_3673,N_9199);
or U18589 (N_18589,N_5217,N_8577);
nor U18590 (N_18590,N_7404,N_3201);
or U18591 (N_18591,N_3840,N_8490);
xor U18592 (N_18592,N_809,N_9095);
nor U18593 (N_18593,N_5581,N_2101);
and U18594 (N_18594,N_838,N_5654);
or U18595 (N_18595,N_3961,N_3441);
nor U18596 (N_18596,N_5396,N_4886);
or U18597 (N_18597,N_3771,N_1354);
nor U18598 (N_18598,N_4485,N_834);
nor U18599 (N_18599,N_1175,N_5050);
nor U18600 (N_18600,N_3217,N_9125);
or U18601 (N_18601,N_7663,N_525);
xnor U18602 (N_18602,N_7535,N_1579);
nor U18603 (N_18603,N_7933,N_1126);
nor U18604 (N_18604,N_5604,N_9780);
nand U18605 (N_18605,N_8136,N_2707);
or U18606 (N_18606,N_2025,N_7644);
or U18607 (N_18607,N_8815,N_7110);
nor U18608 (N_18608,N_8945,N_453);
nor U18609 (N_18609,N_6632,N_4700);
and U18610 (N_18610,N_7902,N_4817);
nor U18611 (N_18611,N_1472,N_7756);
and U18612 (N_18612,N_1880,N_5287);
nand U18613 (N_18613,N_7552,N_2988);
and U18614 (N_18614,N_5298,N_7704);
xor U18615 (N_18615,N_196,N_360);
and U18616 (N_18616,N_5964,N_4972);
and U18617 (N_18617,N_2173,N_6615);
nand U18618 (N_18618,N_1503,N_2358);
nor U18619 (N_18619,N_6732,N_1861);
nor U18620 (N_18620,N_5893,N_6316);
and U18621 (N_18621,N_9922,N_8016);
or U18622 (N_18622,N_5984,N_3782);
nor U18623 (N_18623,N_2502,N_580);
or U18624 (N_18624,N_4994,N_1294);
or U18625 (N_18625,N_9743,N_9400);
nor U18626 (N_18626,N_5950,N_4786);
or U18627 (N_18627,N_2418,N_6679);
and U18628 (N_18628,N_9807,N_7335);
nand U18629 (N_18629,N_7228,N_2887);
nor U18630 (N_18630,N_289,N_8545);
or U18631 (N_18631,N_5213,N_7370);
nor U18632 (N_18632,N_6122,N_8666);
nor U18633 (N_18633,N_8392,N_3893);
or U18634 (N_18634,N_5775,N_5665);
or U18635 (N_18635,N_719,N_1155);
and U18636 (N_18636,N_9310,N_5339);
nor U18637 (N_18637,N_5719,N_7956);
or U18638 (N_18638,N_2508,N_3473);
nand U18639 (N_18639,N_8735,N_9919);
nor U18640 (N_18640,N_3086,N_41);
nand U18641 (N_18641,N_6069,N_8951);
and U18642 (N_18642,N_2323,N_9319);
or U18643 (N_18643,N_7234,N_6337);
nor U18644 (N_18644,N_1784,N_7835);
nand U18645 (N_18645,N_6606,N_7871);
nand U18646 (N_18646,N_245,N_2863);
nor U18647 (N_18647,N_2042,N_9220);
xnor U18648 (N_18648,N_1895,N_1001);
nor U18649 (N_18649,N_1335,N_696);
or U18650 (N_18650,N_5956,N_6);
xnor U18651 (N_18651,N_468,N_5251);
nand U18652 (N_18652,N_6074,N_8440);
nor U18653 (N_18653,N_8567,N_2417);
or U18654 (N_18654,N_7399,N_8825);
and U18655 (N_18655,N_3500,N_3982);
nor U18656 (N_18656,N_3166,N_1836);
nor U18657 (N_18657,N_6935,N_8022);
nand U18658 (N_18658,N_5232,N_5936);
xnor U18659 (N_18659,N_8966,N_2564);
or U18660 (N_18660,N_2363,N_1323);
or U18661 (N_18661,N_1097,N_3667);
or U18662 (N_18662,N_5688,N_1529);
or U18663 (N_18663,N_4218,N_4072);
nand U18664 (N_18664,N_4132,N_1615);
nor U18665 (N_18665,N_6797,N_9036);
or U18666 (N_18666,N_1585,N_1447);
nor U18667 (N_18667,N_7235,N_8904);
xor U18668 (N_18668,N_8954,N_7541);
nor U18669 (N_18669,N_7911,N_9277);
nand U18670 (N_18670,N_7796,N_1566);
nand U18671 (N_18671,N_4112,N_5541);
nor U18672 (N_18672,N_9682,N_1453);
or U18673 (N_18673,N_7471,N_2312);
and U18674 (N_18674,N_7924,N_2268);
and U18675 (N_18675,N_6520,N_3638);
nand U18676 (N_18676,N_5571,N_8807);
and U18677 (N_18677,N_4232,N_523);
and U18678 (N_18678,N_442,N_9199);
nor U18679 (N_18679,N_9111,N_5408);
or U18680 (N_18680,N_7206,N_5429);
nand U18681 (N_18681,N_3803,N_5810);
and U18682 (N_18682,N_7942,N_8030);
or U18683 (N_18683,N_2683,N_1641);
or U18684 (N_18684,N_2974,N_2488);
nor U18685 (N_18685,N_3496,N_2752);
xor U18686 (N_18686,N_9168,N_6531);
or U18687 (N_18687,N_3135,N_1335);
nor U18688 (N_18688,N_6282,N_9797);
nand U18689 (N_18689,N_8407,N_3802);
and U18690 (N_18690,N_5823,N_7198);
xnor U18691 (N_18691,N_7970,N_9034);
and U18692 (N_18692,N_5952,N_659);
or U18693 (N_18693,N_4444,N_5347);
nor U18694 (N_18694,N_2678,N_536);
and U18695 (N_18695,N_1197,N_280);
nand U18696 (N_18696,N_1626,N_1970);
or U18697 (N_18697,N_8024,N_3306);
xor U18698 (N_18698,N_492,N_8934);
and U18699 (N_18699,N_8244,N_6710);
and U18700 (N_18700,N_3289,N_3972);
or U18701 (N_18701,N_8049,N_1724);
nand U18702 (N_18702,N_3777,N_1975);
and U18703 (N_18703,N_6458,N_9217);
nor U18704 (N_18704,N_7447,N_6155);
nor U18705 (N_18705,N_9432,N_2317);
or U18706 (N_18706,N_4643,N_2635);
nor U18707 (N_18707,N_4309,N_5366);
and U18708 (N_18708,N_1305,N_8176);
or U18709 (N_18709,N_5632,N_1100);
nor U18710 (N_18710,N_9058,N_3699);
nor U18711 (N_18711,N_1228,N_8332);
or U18712 (N_18712,N_9147,N_519);
or U18713 (N_18713,N_3680,N_7441);
nand U18714 (N_18714,N_2589,N_3935);
and U18715 (N_18715,N_7131,N_8196);
nor U18716 (N_18716,N_4743,N_5414);
nand U18717 (N_18717,N_1609,N_8473);
nand U18718 (N_18718,N_504,N_948);
xor U18719 (N_18719,N_1891,N_6802);
nor U18720 (N_18720,N_8868,N_5815);
and U18721 (N_18721,N_7042,N_4363);
nand U18722 (N_18722,N_2425,N_921);
or U18723 (N_18723,N_6854,N_2387);
nand U18724 (N_18724,N_4223,N_740);
xor U18725 (N_18725,N_2944,N_7386);
or U18726 (N_18726,N_2962,N_6286);
nor U18727 (N_18727,N_1374,N_7754);
nor U18728 (N_18728,N_945,N_582);
nor U18729 (N_18729,N_5288,N_3376);
nand U18730 (N_18730,N_6952,N_7677);
nand U18731 (N_18731,N_4961,N_2102);
nor U18732 (N_18732,N_3930,N_5254);
or U18733 (N_18733,N_5757,N_2746);
nor U18734 (N_18734,N_5235,N_9891);
nand U18735 (N_18735,N_7970,N_1970);
nor U18736 (N_18736,N_9509,N_1806);
or U18737 (N_18737,N_2349,N_1152);
or U18738 (N_18738,N_6101,N_3560);
nand U18739 (N_18739,N_7462,N_7649);
nand U18740 (N_18740,N_7734,N_2152);
nand U18741 (N_18741,N_4474,N_4993);
nor U18742 (N_18742,N_16,N_9366);
or U18743 (N_18743,N_2192,N_7997);
nand U18744 (N_18744,N_3482,N_6371);
nand U18745 (N_18745,N_7231,N_2494);
and U18746 (N_18746,N_1244,N_3977);
nor U18747 (N_18747,N_5315,N_7742);
nand U18748 (N_18748,N_428,N_8665);
xnor U18749 (N_18749,N_7409,N_1685);
and U18750 (N_18750,N_690,N_7035);
and U18751 (N_18751,N_9379,N_7840);
or U18752 (N_18752,N_5672,N_2884);
or U18753 (N_18753,N_8262,N_4941);
and U18754 (N_18754,N_8287,N_6386);
and U18755 (N_18755,N_3998,N_3337);
and U18756 (N_18756,N_8145,N_9544);
and U18757 (N_18757,N_6686,N_6123);
xor U18758 (N_18758,N_6746,N_9013);
nor U18759 (N_18759,N_3821,N_7993);
nand U18760 (N_18760,N_2938,N_9335);
nand U18761 (N_18761,N_3678,N_7642);
nor U18762 (N_18762,N_6894,N_8906);
and U18763 (N_18763,N_8073,N_6371);
nand U18764 (N_18764,N_2390,N_8299);
and U18765 (N_18765,N_8836,N_6164);
nor U18766 (N_18766,N_9941,N_9953);
nor U18767 (N_18767,N_5485,N_1740);
or U18768 (N_18768,N_9831,N_7321);
and U18769 (N_18769,N_366,N_8291);
and U18770 (N_18770,N_9500,N_8381);
or U18771 (N_18771,N_1155,N_6200);
nor U18772 (N_18772,N_2326,N_5928);
nor U18773 (N_18773,N_6040,N_9394);
and U18774 (N_18774,N_2914,N_8577);
and U18775 (N_18775,N_6974,N_7752);
nor U18776 (N_18776,N_5171,N_4509);
nor U18777 (N_18777,N_6862,N_1478);
and U18778 (N_18778,N_7111,N_6036);
or U18779 (N_18779,N_7662,N_8921);
nor U18780 (N_18780,N_6137,N_8412);
xnor U18781 (N_18781,N_8762,N_8973);
and U18782 (N_18782,N_9716,N_2383);
nand U18783 (N_18783,N_5663,N_9585);
and U18784 (N_18784,N_2426,N_2083);
or U18785 (N_18785,N_4080,N_3028);
nand U18786 (N_18786,N_8719,N_4936);
nand U18787 (N_18787,N_9966,N_1089);
nor U18788 (N_18788,N_7656,N_8957);
or U18789 (N_18789,N_1468,N_8012);
or U18790 (N_18790,N_7365,N_1823);
nor U18791 (N_18791,N_1638,N_6733);
and U18792 (N_18792,N_6911,N_9786);
xnor U18793 (N_18793,N_8000,N_3695);
and U18794 (N_18794,N_512,N_871);
or U18795 (N_18795,N_2497,N_1356);
or U18796 (N_18796,N_5067,N_7342);
nor U18797 (N_18797,N_1220,N_2986);
nor U18798 (N_18798,N_9674,N_6375);
or U18799 (N_18799,N_4713,N_1181);
nor U18800 (N_18800,N_2028,N_6548);
and U18801 (N_18801,N_4896,N_2889);
and U18802 (N_18802,N_773,N_5291);
nand U18803 (N_18803,N_1251,N_6711);
nand U18804 (N_18804,N_1726,N_2422);
nand U18805 (N_18805,N_6323,N_1156);
and U18806 (N_18806,N_6810,N_3615);
nor U18807 (N_18807,N_8243,N_7920);
or U18808 (N_18808,N_3416,N_6791);
or U18809 (N_18809,N_9353,N_6757);
and U18810 (N_18810,N_27,N_1398);
nand U18811 (N_18811,N_1924,N_2591);
or U18812 (N_18812,N_692,N_4924);
nor U18813 (N_18813,N_1863,N_2260);
nor U18814 (N_18814,N_1392,N_9563);
or U18815 (N_18815,N_3314,N_9940);
xor U18816 (N_18816,N_53,N_8372);
and U18817 (N_18817,N_1875,N_8919);
and U18818 (N_18818,N_4150,N_7308);
and U18819 (N_18819,N_7676,N_7678);
and U18820 (N_18820,N_8808,N_3871);
or U18821 (N_18821,N_2673,N_3358);
or U18822 (N_18822,N_6325,N_1644);
and U18823 (N_18823,N_1842,N_6395);
or U18824 (N_18824,N_6175,N_3662);
and U18825 (N_18825,N_8113,N_9125);
or U18826 (N_18826,N_6245,N_3019);
and U18827 (N_18827,N_2750,N_3164);
nor U18828 (N_18828,N_2596,N_3599);
and U18829 (N_18829,N_7925,N_390);
xor U18830 (N_18830,N_1325,N_2707);
nand U18831 (N_18831,N_8419,N_1843);
and U18832 (N_18832,N_4095,N_1870);
and U18833 (N_18833,N_9913,N_4782);
or U18834 (N_18834,N_3732,N_9437);
and U18835 (N_18835,N_6929,N_3812);
and U18836 (N_18836,N_4842,N_6660);
xor U18837 (N_18837,N_8487,N_1072);
and U18838 (N_18838,N_93,N_2711);
and U18839 (N_18839,N_5139,N_566);
and U18840 (N_18840,N_8685,N_2851);
or U18841 (N_18841,N_5825,N_4933);
nand U18842 (N_18842,N_3338,N_5994);
nor U18843 (N_18843,N_4176,N_6359);
xnor U18844 (N_18844,N_9180,N_1197);
or U18845 (N_18845,N_2068,N_6818);
xor U18846 (N_18846,N_2642,N_1318);
and U18847 (N_18847,N_2879,N_5661);
nand U18848 (N_18848,N_2574,N_3263);
nor U18849 (N_18849,N_5410,N_7791);
or U18850 (N_18850,N_3677,N_4309);
or U18851 (N_18851,N_7497,N_7384);
or U18852 (N_18852,N_9787,N_9246);
nor U18853 (N_18853,N_3303,N_7436);
and U18854 (N_18854,N_5436,N_672);
nand U18855 (N_18855,N_1902,N_4257);
and U18856 (N_18856,N_7224,N_8016);
and U18857 (N_18857,N_4173,N_3547);
xnor U18858 (N_18858,N_4872,N_1818);
nand U18859 (N_18859,N_6954,N_5424);
nor U18860 (N_18860,N_9296,N_1044);
xor U18861 (N_18861,N_1010,N_40);
and U18862 (N_18862,N_8185,N_7813);
and U18863 (N_18863,N_4472,N_5064);
or U18864 (N_18864,N_2008,N_7126);
nand U18865 (N_18865,N_29,N_7885);
and U18866 (N_18866,N_3449,N_4733);
xor U18867 (N_18867,N_8049,N_5283);
nor U18868 (N_18868,N_5700,N_6636);
nor U18869 (N_18869,N_7220,N_4414);
and U18870 (N_18870,N_6967,N_2189);
or U18871 (N_18871,N_6771,N_9702);
nand U18872 (N_18872,N_7106,N_7182);
nor U18873 (N_18873,N_269,N_5416);
and U18874 (N_18874,N_6555,N_2153);
and U18875 (N_18875,N_1921,N_1120);
nor U18876 (N_18876,N_9369,N_3427);
nand U18877 (N_18877,N_9435,N_6145);
nor U18878 (N_18878,N_4997,N_9009);
nand U18879 (N_18879,N_4890,N_1862);
and U18880 (N_18880,N_2673,N_5958);
nand U18881 (N_18881,N_5547,N_8127);
or U18882 (N_18882,N_9820,N_2935);
or U18883 (N_18883,N_2216,N_9715);
or U18884 (N_18884,N_5692,N_4328);
nor U18885 (N_18885,N_3753,N_5963);
and U18886 (N_18886,N_417,N_1170);
nor U18887 (N_18887,N_2561,N_2368);
nand U18888 (N_18888,N_511,N_6663);
or U18889 (N_18889,N_1153,N_8533);
xnor U18890 (N_18890,N_4877,N_7339);
or U18891 (N_18891,N_2271,N_830);
xnor U18892 (N_18892,N_1973,N_6777);
nor U18893 (N_18893,N_9083,N_2705);
and U18894 (N_18894,N_4980,N_1555);
nor U18895 (N_18895,N_7007,N_6525);
or U18896 (N_18896,N_4760,N_4531);
nor U18897 (N_18897,N_7968,N_3361);
nor U18898 (N_18898,N_4930,N_2931);
nand U18899 (N_18899,N_9216,N_5984);
nor U18900 (N_18900,N_4520,N_136);
or U18901 (N_18901,N_9806,N_7852);
xor U18902 (N_18902,N_2461,N_1737);
nand U18903 (N_18903,N_3510,N_8925);
nand U18904 (N_18904,N_244,N_3130);
and U18905 (N_18905,N_4147,N_3720);
nor U18906 (N_18906,N_9540,N_6214);
or U18907 (N_18907,N_8161,N_480);
nor U18908 (N_18908,N_1786,N_9521);
nor U18909 (N_18909,N_423,N_8549);
nor U18910 (N_18910,N_1014,N_5864);
nor U18911 (N_18911,N_6,N_4979);
or U18912 (N_18912,N_7174,N_5385);
nand U18913 (N_18913,N_1220,N_5167);
nand U18914 (N_18914,N_5917,N_4725);
or U18915 (N_18915,N_5055,N_3825);
and U18916 (N_18916,N_7790,N_6251);
nor U18917 (N_18917,N_3105,N_8034);
nor U18918 (N_18918,N_5266,N_6671);
nand U18919 (N_18919,N_4282,N_2001);
nor U18920 (N_18920,N_3939,N_2035);
or U18921 (N_18921,N_6164,N_8648);
nor U18922 (N_18922,N_6652,N_1793);
nor U18923 (N_18923,N_3897,N_5593);
or U18924 (N_18924,N_3292,N_6610);
or U18925 (N_18925,N_2383,N_517);
nand U18926 (N_18926,N_9380,N_7498);
and U18927 (N_18927,N_1692,N_6549);
nor U18928 (N_18928,N_2055,N_3065);
and U18929 (N_18929,N_460,N_6014);
nor U18930 (N_18930,N_8945,N_2286);
nor U18931 (N_18931,N_4683,N_3422);
or U18932 (N_18932,N_1264,N_6917);
and U18933 (N_18933,N_897,N_3064);
and U18934 (N_18934,N_9015,N_1332);
nor U18935 (N_18935,N_6474,N_2671);
xnor U18936 (N_18936,N_6179,N_4114);
nand U18937 (N_18937,N_5039,N_593);
nand U18938 (N_18938,N_2579,N_2123);
xor U18939 (N_18939,N_4132,N_7033);
nand U18940 (N_18940,N_6402,N_7138);
and U18941 (N_18941,N_4832,N_5907);
nor U18942 (N_18942,N_3338,N_9733);
or U18943 (N_18943,N_8286,N_6594);
and U18944 (N_18944,N_5885,N_975);
nand U18945 (N_18945,N_7900,N_684);
nand U18946 (N_18946,N_3668,N_9238);
or U18947 (N_18947,N_6733,N_1909);
nand U18948 (N_18948,N_529,N_894);
nand U18949 (N_18949,N_6808,N_3882);
nor U18950 (N_18950,N_7654,N_5581);
nand U18951 (N_18951,N_1424,N_6431);
or U18952 (N_18952,N_4473,N_3058);
nor U18953 (N_18953,N_7091,N_2334);
nand U18954 (N_18954,N_7373,N_3);
nor U18955 (N_18955,N_2850,N_8654);
or U18956 (N_18956,N_5128,N_6613);
nor U18957 (N_18957,N_2411,N_9031);
and U18958 (N_18958,N_9543,N_9783);
xor U18959 (N_18959,N_9542,N_6799);
and U18960 (N_18960,N_8600,N_4707);
nand U18961 (N_18961,N_2875,N_6092);
or U18962 (N_18962,N_8771,N_6789);
nand U18963 (N_18963,N_6608,N_4713);
and U18964 (N_18964,N_8684,N_5014);
or U18965 (N_18965,N_9868,N_6542);
and U18966 (N_18966,N_4824,N_1344);
xor U18967 (N_18967,N_2017,N_4933);
and U18968 (N_18968,N_5641,N_3456);
nor U18969 (N_18969,N_6525,N_8828);
nand U18970 (N_18970,N_9391,N_7263);
nor U18971 (N_18971,N_6827,N_7041);
nand U18972 (N_18972,N_8189,N_4354);
nand U18973 (N_18973,N_3315,N_118);
nand U18974 (N_18974,N_9248,N_9945);
nor U18975 (N_18975,N_7742,N_1789);
nand U18976 (N_18976,N_4079,N_7443);
and U18977 (N_18977,N_8982,N_4456);
or U18978 (N_18978,N_8301,N_4239);
and U18979 (N_18979,N_9344,N_3001);
and U18980 (N_18980,N_6952,N_8257);
xor U18981 (N_18981,N_4756,N_1526);
nand U18982 (N_18982,N_8728,N_363);
nor U18983 (N_18983,N_84,N_4169);
or U18984 (N_18984,N_2836,N_1832);
and U18985 (N_18985,N_5844,N_1596);
or U18986 (N_18986,N_1554,N_5141);
nand U18987 (N_18987,N_7812,N_8742);
xor U18988 (N_18988,N_5899,N_5123);
nor U18989 (N_18989,N_7619,N_8838);
and U18990 (N_18990,N_8038,N_827);
or U18991 (N_18991,N_7855,N_6700);
nor U18992 (N_18992,N_3979,N_5572);
and U18993 (N_18993,N_9850,N_9704);
nor U18994 (N_18994,N_2665,N_1616);
and U18995 (N_18995,N_4730,N_6345);
and U18996 (N_18996,N_8733,N_7224);
nor U18997 (N_18997,N_4128,N_340);
and U18998 (N_18998,N_8484,N_7291);
nor U18999 (N_18999,N_6495,N_3915);
nor U19000 (N_19000,N_2975,N_6981);
or U19001 (N_19001,N_6934,N_8123);
xnor U19002 (N_19002,N_5004,N_6171);
nand U19003 (N_19003,N_5431,N_4644);
nand U19004 (N_19004,N_5479,N_9743);
xor U19005 (N_19005,N_9816,N_8088);
nor U19006 (N_19006,N_2674,N_333);
nand U19007 (N_19007,N_7851,N_4584);
nor U19008 (N_19008,N_1722,N_3724);
xor U19009 (N_19009,N_795,N_8042);
nand U19010 (N_19010,N_3402,N_5153);
nand U19011 (N_19011,N_3928,N_6431);
nor U19012 (N_19012,N_3291,N_2539);
nor U19013 (N_19013,N_4752,N_1795);
nor U19014 (N_19014,N_6875,N_5802);
nor U19015 (N_19015,N_6391,N_9025);
and U19016 (N_19016,N_6156,N_735);
and U19017 (N_19017,N_4453,N_2658);
xnor U19018 (N_19018,N_8208,N_9527);
nor U19019 (N_19019,N_5743,N_9299);
nand U19020 (N_19020,N_83,N_3084);
nand U19021 (N_19021,N_6602,N_1635);
nor U19022 (N_19022,N_2924,N_3709);
and U19023 (N_19023,N_1900,N_4298);
nor U19024 (N_19024,N_9616,N_2125);
nand U19025 (N_19025,N_4194,N_5370);
or U19026 (N_19026,N_2632,N_1887);
nand U19027 (N_19027,N_4355,N_610);
xnor U19028 (N_19028,N_462,N_2886);
nand U19029 (N_19029,N_6775,N_5260);
and U19030 (N_19030,N_8642,N_1408);
and U19031 (N_19031,N_9206,N_689);
or U19032 (N_19032,N_3826,N_1180);
nor U19033 (N_19033,N_5610,N_2885);
nor U19034 (N_19034,N_7393,N_1603);
and U19035 (N_19035,N_3150,N_9973);
nand U19036 (N_19036,N_431,N_9206);
and U19037 (N_19037,N_869,N_5502);
or U19038 (N_19038,N_1118,N_6727);
or U19039 (N_19039,N_9452,N_8398);
and U19040 (N_19040,N_3995,N_1702);
and U19041 (N_19041,N_1043,N_3284);
xor U19042 (N_19042,N_9586,N_8281);
or U19043 (N_19043,N_2280,N_6921);
xnor U19044 (N_19044,N_3918,N_5417);
or U19045 (N_19045,N_650,N_2467);
nand U19046 (N_19046,N_487,N_5183);
and U19047 (N_19047,N_3215,N_4032);
or U19048 (N_19048,N_7353,N_5613);
and U19049 (N_19049,N_5070,N_5323);
or U19050 (N_19050,N_2099,N_1220);
or U19051 (N_19051,N_293,N_3408);
nand U19052 (N_19052,N_9115,N_6210);
nand U19053 (N_19053,N_8672,N_9404);
nor U19054 (N_19054,N_2725,N_4961);
or U19055 (N_19055,N_9243,N_1759);
nand U19056 (N_19056,N_2254,N_6521);
nand U19057 (N_19057,N_8196,N_950);
and U19058 (N_19058,N_3344,N_5342);
nor U19059 (N_19059,N_7357,N_7645);
nand U19060 (N_19060,N_677,N_2274);
and U19061 (N_19061,N_8,N_963);
nand U19062 (N_19062,N_1847,N_8649);
and U19063 (N_19063,N_6963,N_549);
nand U19064 (N_19064,N_5173,N_577);
or U19065 (N_19065,N_5517,N_6896);
or U19066 (N_19066,N_8320,N_1568);
nand U19067 (N_19067,N_4845,N_3697);
or U19068 (N_19068,N_1495,N_5051);
nor U19069 (N_19069,N_9113,N_5524);
nand U19070 (N_19070,N_5450,N_7558);
or U19071 (N_19071,N_2456,N_6793);
and U19072 (N_19072,N_1331,N_9065);
and U19073 (N_19073,N_7292,N_7594);
and U19074 (N_19074,N_3070,N_2560);
nand U19075 (N_19075,N_5677,N_2661);
and U19076 (N_19076,N_7083,N_5185);
and U19077 (N_19077,N_1332,N_7423);
nand U19078 (N_19078,N_8441,N_8384);
and U19079 (N_19079,N_502,N_2318);
or U19080 (N_19080,N_7975,N_8238);
or U19081 (N_19081,N_4722,N_7458);
nor U19082 (N_19082,N_191,N_5046);
nand U19083 (N_19083,N_8144,N_3313);
or U19084 (N_19084,N_6779,N_808);
nor U19085 (N_19085,N_5898,N_3154);
nand U19086 (N_19086,N_4531,N_5286);
xor U19087 (N_19087,N_4862,N_3644);
nand U19088 (N_19088,N_9889,N_4974);
nor U19089 (N_19089,N_3486,N_9185);
nor U19090 (N_19090,N_7697,N_9342);
or U19091 (N_19091,N_806,N_1785);
nor U19092 (N_19092,N_7378,N_527);
xor U19093 (N_19093,N_5012,N_6800);
or U19094 (N_19094,N_8609,N_5493);
nand U19095 (N_19095,N_1210,N_2856);
and U19096 (N_19096,N_9552,N_3880);
and U19097 (N_19097,N_3125,N_9330);
or U19098 (N_19098,N_114,N_2264);
and U19099 (N_19099,N_2145,N_3734);
and U19100 (N_19100,N_3219,N_5073);
nand U19101 (N_19101,N_5601,N_72);
xnor U19102 (N_19102,N_8722,N_7863);
and U19103 (N_19103,N_3183,N_2545);
nand U19104 (N_19104,N_6408,N_4624);
nand U19105 (N_19105,N_2886,N_5284);
xnor U19106 (N_19106,N_4761,N_1799);
nand U19107 (N_19107,N_7927,N_8808);
nand U19108 (N_19108,N_9345,N_2289);
or U19109 (N_19109,N_1242,N_8801);
or U19110 (N_19110,N_7827,N_3885);
nand U19111 (N_19111,N_6431,N_1101);
nand U19112 (N_19112,N_4345,N_1574);
nand U19113 (N_19113,N_3603,N_7030);
and U19114 (N_19114,N_6507,N_1662);
nand U19115 (N_19115,N_3453,N_5039);
nand U19116 (N_19116,N_3971,N_3592);
nand U19117 (N_19117,N_9213,N_9930);
xor U19118 (N_19118,N_4882,N_5080);
or U19119 (N_19119,N_6687,N_925);
nor U19120 (N_19120,N_4619,N_1922);
nand U19121 (N_19121,N_2666,N_8980);
nor U19122 (N_19122,N_7646,N_2356);
or U19123 (N_19123,N_5529,N_189);
or U19124 (N_19124,N_4913,N_5477);
nor U19125 (N_19125,N_5578,N_7781);
and U19126 (N_19126,N_5041,N_3792);
nor U19127 (N_19127,N_361,N_0);
or U19128 (N_19128,N_1146,N_4564);
nand U19129 (N_19129,N_9191,N_8595);
nand U19130 (N_19130,N_4740,N_781);
xnor U19131 (N_19131,N_5740,N_9021);
or U19132 (N_19132,N_9036,N_6388);
nor U19133 (N_19133,N_2687,N_3667);
nor U19134 (N_19134,N_4558,N_4814);
nor U19135 (N_19135,N_8790,N_8330);
and U19136 (N_19136,N_4984,N_452);
and U19137 (N_19137,N_3179,N_2778);
nand U19138 (N_19138,N_143,N_1508);
or U19139 (N_19139,N_3877,N_7667);
and U19140 (N_19140,N_3822,N_3535);
nor U19141 (N_19141,N_7318,N_3924);
nand U19142 (N_19142,N_6546,N_99);
nor U19143 (N_19143,N_7252,N_6552);
or U19144 (N_19144,N_3915,N_3580);
nor U19145 (N_19145,N_3841,N_1598);
nand U19146 (N_19146,N_4383,N_8683);
nand U19147 (N_19147,N_410,N_6674);
xor U19148 (N_19148,N_7526,N_5034);
and U19149 (N_19149,N_1260,N_8232);
nand U19150 (N_19150,N_8346,N_3571);
or U19151 (N_19151,N_5767,N_8313);
and U19152 (N_19152,N_6524,N_4268);
nor U19153 (N_19153,N_4055,N_1210);
xnor U19154 (N_19154,N_7829,N_8895);
nor U19155 (N_19155,N_2672,N_5314);
and U19156 (N_19156,N_9145,N_3150);
nor U19157 (N_19157,N_2885,N_5691);
nand U19158 (N_19158,N_3806,N_1489);
and U19159 (N_19159,N_7025,N_1601);
and U19160 (N_19160,N_4549,N_5282);
or U19161 (N_19161,N_639,N_2854);
nor U19162 (N_19162,N_1942,N_4452);
nand U19163 (N_19163,N_2672,N_6242);
nand U19164 (N_19164,N_3237,N_7065);
and U19165 (N_19165,N_125,N_9929);
nand U19166 (N_19166,N_8410,N_3031);
nand U19167 (N_19167,N_4573,N_6517);
nor U19168 (N_19168,N_3836,N_4395);
nand U19169 (N_19169,N_9554,N_3453);
nand U19170 (N_19170,N_6446,N_3947);
nor U19171 (N_19171,N_7749,N_3105);
or U19172 (N_19172,N_7994,N_2372);
or U19173 (N_19173,N_5958,N_1787);
nand U19174 (N_19174,N_3005,N_45);
and U19175 (N_19175,N_1262,N_2165);
xor U19176 (N_19176,N_1718,N_6925);
nand U19177 (N_19177,N_8057,N_7295);
or U19178 (N_19178,N_891,N_5125);
nor U19179 (N_19179,N_1411,N_2377);
or U19180 (N_19180,N_4399,N_300);
and U19181 (N_19181,N_806,N_686);
nor U19182 (N_19182,N_636,N_3289);
or U19183 (N_19183,N_6485,N_3292);
or U19184 (N_19184,N_9372,N_7547);
and U19185 (N_19185,N_3786,N_3242);
and U19186 (N_19186,N_3584,N_1009);
nand U19187 (N_19187,N_4979,N_1464);
or U19188 (N_19188,N_7574,N_2592);
and U19189 (N_19189,N_7438,N_866);
and U19190 (N_19190,N_8463,N_2686);
xnor U19191 (N_19191,N_128,N_6388);
and U19192 (N_19192,N_6804,N_7788);
or U19193 (N_19193,N_5461,N_4345);
nand U19194 (N_19194,N_2159,N_73);
nor U19195 (N_19195,N_5345,N_801);
and U19196 (N_19196,N_953,N_8585);
nor U19197 (N_19197,N_8210,N_5872);
nand U19198 (N_19198,N_6439,N_9930);
nor U19199 (N_19199,N_1240,N_8892);
nand U19200 (N_19200,N_9369,N_3189);
or U19201 (N_19201,N_1022,N_2510);
and U19202 (N_19202,N_5135,N_3387);
or U19203 (N_19203,N_2595,N_6562);
or U19204 (N_19204,N_3475,N_4239);
nor U19205 (N_19205,N_6687,N_3356);
and U19206 (N_19206,N_5885,N_2184);
nor U19207 (N_19207,N_692,N_6999);
nand U19208 (N_19208,N_4605,N_4463);
nor U19209 (N_19209,N_8947,N_8128);
and U19210 (N_19210,N_3925,N_6380);
and U19211 (N_19211,N_4994,N_4165);
xnor U19212 (N_19212,N_4329,N_8147);
nor U19213 (N_19213,N_2159,N_7185);
xor U19214 (N_19214,N_8875,N_6236);
nand U19215 (N_19215,N_1585,N_6532);
nand U19216 (N_19216,N_9639,N_4257);
or U19217 (N_19217,N_7021,N_1281);
and U19218 (N_19218,N_5181,N_9971);
or U19219 (N_19219,N_5625,N_6059);
nand U19220 (N_19220,N_198,N_9240);
nand U19221 (N_19221,N_9831,N_8125);
nor U19222 (N_19222,N_1165,N_1794);
and U19223 (N_19223,N_1590,N_161);
or U19224 (N_19224,N_1965,N_9814);
nand U19225 (N_19225,N_4573,N_3810);
nand U19226 (N_19226,N_4934,N_6573);
and U19227 (N_19227,N_6992,N_4413);
and U19228 (N_19228,N_4086,N_8138);
and U19229 (N_19229,N_3951,N_9910);
or U19230 (N_19230,N_6443,N_4888);
or U19231 (N_19231,N_5557,N_5863);
xor U19232 (N_19232,N_1182,N_7671);
nand U19233 (N_19233,N_96,N_4514);
nand U19234 (N_19234,N_1525,N_4646);
xnor U19235 (N_19235,N_3494,N_4371);
nand U19236 (N_19236,N_1561,N_6364);
nand U19237 (N_19237,N_567,N_6649);
xor U19238 (N_19238,N_764,N_3587);
nor U19239 (N_19239,N_236,N_8930);
nand U19240 (N_19240,N_3034,N_5450);
nand U19241 (N_19241,N_3537,N_4351);
and U19242 (N_19242,N_1451,N_1616);
nand U19243 (N_19243,N_6277,N_8821);
or U19244 (N_19244,N_3677,N_302);
xnor U19245 (N_19245,N_2247,N_8612);
nand U19246 (N_19246,N_3057,N_1578);
or U19247 (N_19247,N_9068,N_2253);
nor U19248 (N_19248,N_9708,N_3843);
nor U19249 (N_19249,N_5360,N_4375);
nand U19250 (N_19250,N_1074,N_6799);
or U19251 (N_19251,N_7375,N_9617);
xnor U19252 (N_19252,N_9847,N_9780);
or U19253 (N_19253,N_3485,N_2495);
nor U19254 (N_19254,N_7083,N_1825);
xnor U19255 (N_19255,N_5020,N_4387);
nand U19256 (N_19256,N_659,N_7518);
nand U19257 (N_19257,N_878,N_3879);
nand U19258 (N_19258,N_6905,N_6663);
or U19259 (N_19259,N_4044,N_1955);
nand U19260 (N_19260,N_5100,N_4852);
or U19261 (N_19261,N_465,N_6799);
or U19262 (N_19262,N_34,N_1852);
nand U19263 (N_19263,N_4716,N_3623);
nand U19264 (N_19264,N_1095,N_4540);
nand U19265 (N_19265,N_5035,N_5378);
nor U19266 (N_19266,N_5962,N_8835);
nand U19267 (N_19267,N_1165,N_1417);
or U19268 (N_19268,N_5956,N_3983);
nor U19269 (N_19269,N_8669,N_9284);
nand U19270 (N_19270,N_3763,N_6622);
nor U19271 (N_19271,N_8040,N_4878);
nor U19272 (N_19272,N_5596,N_8381);
nand U19273 (N_19273,N_3455,N_654);
and U19274 (N_19274,N_7526,N_7326);
nand U19275 (N_19275,N_6987,N_7384);
nor U19276 (N_19276,N_2867,N_3512);
or U19277 (N_19277,N_6228,N_2743);
nor U19278 (N_19278,N_7664,N_3937);
nand U19279 (N_19279,N_7014,N_3571);
nor U19280 (N_19280,N_486,N_866);
and U19281 (N_19281,N_580,N_8276);
or U19282 (N_19282,N_957,N_3345);
xnor U19283 (N_19283,N_4203,N_7914);
and U19284 (N_19284,N_8684,N_8868);
and U19285 (N_19285,N_5787,N_640);
and U19286 (N_19286,N_6861,N_402);
nand U19287 (N_19287,N_8356,N_7282);
and U19288 (N_19288,N_7070,N_5555);
nor U19289 (N_19289,N_6883,N_1738);
nor U19290 (N_19290,N_169,N_4144);
nand U19291 (N_19291,N_2927,N_8154);
and U19292 (N_19292,N_5971,N_7902);
nand U19293 (N_19293,N_6017,N_2638);
nor U19294 (N_19294,N_9876,N_7711);
and U19295 (N_19295,N_1233,N_8669);
nor U19296 (N_19296,N_2250,N_2435);
nand U19297 (N_19297,N_6946,N_9942);
nand U19298 (N_19298,N_3531,N_2389);
or U19299 (N_19299,N_9630,N_9272);
nand U19300 (N_19300,N_4024,N_3036);
nand U19301 (N_19301,N_7371,N_3444);
nor U19302 (N_19302,N_9739,N_1360);
nand U19303 (N_19303,N_396,N_1214);
nor U19304 (N_19304,N_2937,N_4);
and U19305 (N_19305,N_3758,N_5634);
and U19306 (N_19306,N_8759,N_75);
or U19307 (N_19307,N_5642,N_7445);
nor U19308 (N_19308,N_464,N_6488);
and U19309 (N_19309,N_5046,N_8439);
or U19310 (N_19310,N_5389,N_58);
or U19311 (N_19311,N_326,N_1981);
and U19312 (N_19312,N_199,N_5158);
or U19313 (N_19313,N_2396,N_1701);
and U19314 (N_19314,N_5236,N_3527);
nor U19315 (N_19315,N_3890,N_5460);
nand U19316 (N_19316,N_5195,N_6285);
nand U19317 (N_19317,N_602,N_8552);
nor U19318 (N_19318,N_1681,N_3656);
nor U19319 (N_19319,N_764,N_504);
nor U19320 (N_19320,N_3562,N_7811);
or U19321 (N_19321,N_3720,N_2629);
nand U19322 (N_19322,N_6348,N_9983);
xnor U19323 (N_19323,N_7119,N_5086);
nand U19324 (N_19324,N_858,N_5145);
nor U19325 (N_19325,N_1058,N_4068);
and U19326 (N_19326,N_4186,N_358);
or U19327 (N_19327,N_2327,N_5653);
xor U19328 (N_19328,N_6892,N_6483);
and U19329 (N_19329,N_4549,N_3872);
nand U19330 (N_19330,N_4205,N_855);
nand U19331 (N_19331,N_5316,N_8568);
nand U19332 (N_19332,N_2881,N_5853);
nor U19333 (N_19333,N_8368,N_7719);
or U19334 (N_19334,N_3505,N_908);
and U19335 (N_19335,N_5046,N_9398);
and U19336 (N_19336,N_3583,N_6753);
xnor U19337 (N_19337,N_2929,N_9308);
and U19338 (N_19338,N_5770,N_9993);
nor U19339 (N_19339,N_7826,N_4247);
nor U19340 (N_19340,N_676,N_6347);
xnor U19341 (N_19341,N_1709,N_2283);
or U19342 (N_19342,N_8976,N_6684);
or U19343 (N_19343,N_3937,N_8852);
nor U19344 (N_19344,N_9486,N_7828);
and U19345 (N_19345,N_804,N_3229);
or U19346 (N_19346,N_8821,N_606);
nor U19347 (N_19347,N_762,N_9465);
xor U19348 (N_19348,N_2292,N_4133);
xor U19349 (N_19349,N_3013,N_6192);
and U19350 (N_19350,N_3983,N_7429);
nor U19351 (N_19351,N_5767,N_4391);
nand U19352 (N_19352,N_5237,N_6958);
nor U19353 (N_19353,N_8494,N_1848);
nor U19354 (N_19354,N_4186,N_1263);
nand U19355 (N_19355,N_9440,N_3885);
nand U19356 (N_19356,N_2120,N_7143);
and U19357 (N_19357,N_8862,N_4894);
and U19358 (N_19358,N_8478,N_1424);
or U19359 (N_19359,N_9554,N_4629);
nand U19360 (N_19360,N_3643,N_8683);
nand U19361 (N_19361,N_38,N_496);
xnor U19362 (N_19362,N_1416,N_6233);
and U19363 (N_19363,N_6171,N_2653);
or U19364 (N_19364,N_6227,N_7110);
nand U19365 (N_19365,N_8330,N_1249);
or U19366 (N_19366,N_2784,N_9805);
or U19367 (N_19367,N_6683,N_8007);
or U19368 (N_19368,N_277,N_744);
or U19369 (N_19369,N_1070,N_961);
nor U19370 (N_19370,N_3188,N_448);
and U19371 (N_19371,N_7624,N_8765);
and U19372 (N_19372,N_814,N_929);
or U19373 (N_19373,N_6597,N_4280);
and U19374 (N_19374,N_8582,N_2668);
and U19375 (N_19375,N_5820,N_1185);
xor U19376 (N_19376,N_6193,N_6664);
and U19377 (N_19377,N_1584,N_8357);
and U19378 (N_19378,N_3568,N_8545);
or U19379 (N_19379,N_8476,N_2139);
nor U19380 (N_19380,N_9407,N_8251);
nand U19381 (N_19381,N_5728,N_11);
nand U19382 (N_19382,N_3817,N_5962);
nand U19383 (N_19383,N_8743,N_3864);
nor U19384 (N_19384,N_2017,N_1374);
and U19385 (N_19385,N_2305,N_4972);
nand U19386 (N_19386,N_6167,N_8631);
or U19387 (N_19387,N_1015,N_5658);
nand U19388 (N_19388,N_4246,N_8582);
or U19389 (N_19389,N_8185,N_5573);
or U19390 (N_19390,N_2529,N_9163);
nor U19391 (N_19391,N_7754,N_6206);
nor U19392 (N_19392,N_3784,N_4690);
and U19393 (N_19393,N_4680,N_2706);
nand U19394 (N_19394,N_2453,N_9400);
nand U19395 (N_19395,N_2663,N_7956);
and U19396 (N_19396,N_9197,N_9906);
nand U19397 (N_19397,N_4245,N_2489);
nor U19398 (N_19398,N_9739,N_1371);
nand U19399 (N_19399,N_3567,N_8886);
nand U19400 (N_19400,N_9880,N_6209);
nand U19401 (N_19401,N_5764,N_6801);
nor U19402 (N_19402,N_3334,N_3207);
nor U19403 (N_19403,N_3238,N_4306);
nand U19404 (N_19404,N_9507,N_4516);
nand U19405 (N_19405,N_2821,N_7492);
or U19406 (N_19406,N_9651,N_3274);
or U19407 (N_19407,N_8429,N_3502);
nor U19408 (N_19408,N_4746,N_3946);
and U19409 (N_19409,N_8034,N_1407);
and U19410 (N_19410,N_1774,N_8481);
and U19411 (N_19411,N_9146,N_4302);
nor U19412 (N_19412,N_9608,N_2173);
or U19413 (N_19413,N_9366,N_574);
nor U19414 (N_19414,N_626,N_2919);
or U19415 (N_19415,N_1698,N_2160);
or U19416 (N_19416,N_5608,N_1729);
nor U19417 (N_19417,N_9897,N_2993);
nor U19418 (N_19418,N_5685,N_7393);
or U19419 (N_19419,N_867,N_2754);
xnor U19420 (N_19420,N_6655,N_9795);
or U19421 (N_19421,N_6414,N_7104);
nand U19422 (N_19422,N_3056,N_6724);
nor U19423 (N_19423,N_6701,N_7580);
nor U19424 (N_19424,N_2350,N_9836);
nand U19425 (N_19425,N_4945,N_6422);
nand U19426 (N_19426,N_9157,N_6086);
nor U19427 (N_19427,N_5630,N_7866);
xor U19428 (N_19428,N_2536,N_729);
and U19429 (N_19429,N_1849,N_2162);
and U19430 (N_19430,N_6286,N_4339);
nor U19431 (N_19431,N_680,N_5220);
xor U19432 (N_19432,N_4068,N_9899);
or U19433 (N_19433,N_2470,N_5954);
nor U19434 (N_19434,N_3936,N_9749);
or U19435 (N_19435,N_7962,N_1608);
and U19436 (N_19436,N_9507,N_7735);
or U19437 (N_19437,N_343,N_3774);
and U19438 (N_19438,N_5859,N_423);
and U19439 (N_19439,N_3057,N_1758);
and U19440 (N_19440,N_546,N_8920);
xnor U19441 (N_19441,N_2423,N_5905);
xor U19442 (N_19442,N_1846,N_4641);
nor U19443 (N_19443,N_9801,N_2023);
nand U19444 (N_19444,N_7161,N_7284);
nand U19445 (N_19445,N_2130,N_8199);
nor U19446 (N_19446,N_1275,N_495);
nand U19447 (N_19447,N_7064,N_9592);
nor U19448 (N_19448,N_5822,N_6090);
nand U19449 (N_19449,N_6926,N_1648);
nand U19450 (N_19450,N_2070,N_5509);
or U19451 (N_19451,N_4713,N_7534);
xnor U19452 (N_19452,N_4299,N_1694);
nand U19453 (N_19453,N_9796,N_9005);
or U19454 (N_19454,N_6282,N_8233);
xnor U19455 (N_19455,N_9162,N_2044);
nor U19456 (N_19456,N_8034,N_145);
nor U19457 (N_19457,N_6236,N_6914);
nor U19458 (N_19458,N_9588,N_3826);
or U19459 (N_19459,N_1100,N_943);
nor U19460 (N_19460,N_9486,N_2277);
or U19461 (N_19461,N_7253,N_4257);
and U19462 (N_19462,N_1629,N_7634);
nor U19463 (N_19463,N_1263,N_2057);
nand U19464 (N_19464,N_4137,N_7558);
or U19465 (N_19465,N_8429,N_9084);
nor U19466 (N_19466,N_7343,N_7692);
and U19467 (N_19467,N_7958,N_7406);
and U19468 (N_19468,N_2733,N_1535);
nand U19469 (N_19469,N_8357,N_823);
or U19470 (N_19470,N_8617,N_57);
nand U19471 (N_19471,N_4193,N_9533);
nand U19472 (N_19472,N_4057,N_8913);
nand U19473 (N_19473,N_5788,N_674);
nor U19474 (N_19474,N_9992,N_2572);
nand U19475 (N_19475,N_1643,N_192);
nor U19476 (N_19476,N_1774,N_6068);
xnor U19477 (N_19477,N_4732,N_1598);
and U19478 (N_19478,N_3559,N_9312);
nand U19479 (N_19479,N_1138,N_7590);
nand U19480 (N_19480,N_6029,N_6085);
nor U19481 (N_19481,N_3394,N_9638);
nor U19482 (N_19482,N_7087,N_2703);
nor U19483 (N_19483,N_8719,N_5489);
and U19484 (N_19484,N_9084,N_292);
and U19485 (N_19485,N_6967,N_3584);
or U19486 (N_19486,N_7337,N_3025);
or U19487 (N_19487,N_1887,N_2409);
xnor U19488 (N_19488,N_9495,N_2744);
nand U19489 (N_19489,N_9544,N_2616);
or U19490 (N_19490,N_3897,N_5306);
and U19491 (N_19491,N_7725,N_6258);
xnor U19492 (N_19492,N_9238,N_9312);
nand U19493 (N_19493,N_1120,N_8344);
or U19494 (N_19494,N_5843,N_7688);
and U19495 (N_19495,N_5699,N_9975);
xnor U19496 (N_19496,N_8279,N_8202);
nand U19497 (N_19497,N_2588,N_2041);
or U19498 (N_19498,N_9347,N_6251);
or U19499 (N_19499,N_9419,N_1603);
or U19500 (N_19500,N_5114,N_5134);
and U19501 (N_19501,N_7561,N_8720);
nor U19502 (N_19502,N_1388,N_7145);
nor U19503 (N_19503,N_2263,N_605);
or U19504 (N_19504,N_1604,N_8632);
and U19505 (N_19505,N_212,N_8202);
and U19506 (N_19506,N_2550,N_8271);
xnor U19507 (N_19507,N_8795,N_8370);
nor U19508 (N_19508,N_3456,N_7923);
nand U19509 (N_19509,N_8114,N_9574);
xor U19510 (N_19510,N_5857,N_2191);
nor U19511 (N_19511,N_1878,N_5736);
or U19512 (N_19512,N_7232,N_8894);
and U19513 (N_19513,N_8291,N_8176);
and U19514 (N_19514,N_3130,N_5236);
nand U19515 (N_19515,N_5861,N_5417);
and U19516 (N_19516,N_8631,N_5328);
or U19517 (N_19517,N_2632,N_8704);
xnor U19518 (N_19518,N_733,N_6023);
or U19519 (N_19519,N_690,N_5880);
xnor U19520 (N_19520,N_7846,N_7176);
nand U19521 (N_19521,N_9838,N_6854);
nor U19522 (N_19522,N_5828,N_5355);
or U19523 (N_19523,N_6110,N_7484);
nor U19524 (N_19524,N_703,N_3606);
and U19525 (N_19525,N_7681,N_4154);
and U19526 (N_19526,N_2178,N_2904);
and U19527 (N_19527,N_4933,N_3624);
nor U19528 (N_19528,N_788,N_5638);
or U19529 (N_19529,N_8849,N_1077);
and U19530 (N_19530,N_5041,N_8316);
nand U19531 (N_19531,N_1528,N_4348);
nor U19532 (N_19532,N_7444,N_3843);
nor U19533 (N_19533,N_7918,N_1223);
nand U19534 (N_19534,N_1771,N_1062);
or U19535 (N_19535,N_5008,N_9587);
nor U19536 (N_19536,N_5181,N_9256);
and U19537 (N_19537,N_1751,N_2971);
and U19538 (N_19538,N_1045,N_8846);
xor U19539 (N_19539,N_6675,N_5385);
or U19540 (N_19540,N_4522,N_4815);
xor U19541 (N_19541,N_6979,N_7765);
xor U19542 (N_19542,N_687,N_8804);
xnor U19543 (N_19543,N_519,N_6209);
or U19544 (N_19544,N_6151,N_2095);
xor U19545 (N_19545,N_4623,N_4090);
nor U19546 (N_19546,N_409,N_6780);
nor U19547 (N_19547,N_7596,N_3668);
xor U19548 (N_19548,N_3977,N_4066);
xor U19549 (N_19549,N_5373,N_2991);
or U19550 (N_19550,N_6305,N_5611);
xnor U19551 (N_19551,N_565,N_5976);
nor U19552 (N_19552,N_9716,N_5878);
or U19553 (N_19553,N_9482,N_8977);
nor U19554 (N_19554,N_7844,N_4696);
nor U19555 (N_19555,N_7567,N_4602);
nand U19556 (N_19556,N_5993,N_7435);
or U19557 (N_19557,N_7313,N_5906);
and U19558 (N_19558,N_7340,N_7890);
and U19559 (N_19559,N_6918,N_7503);
or U19560 (N_19560,N_8171,N_2538);
or U19561 (N_19561,N_703,N_3451);
and U19562 (N_19562,N_8708,N_7205);
or U19563 (N_19563,N_2310,N_8285);
and U19564 (N_19564,N_8892,N_3034);
nand U19565 (N_19565,N_6457,N_2989);
nor U19566 (N_19566,N_5974,N_3492);
nand U19567 (N_19567,N_1384,N_1933);
xnor U19568 (N_19568,N_3854,N_5829);
xnor U19569 (N_19569,N_2695,N_3500);
nand U19570 (N_19570,N_7351,N_9430);
and U19571 (N_19571,N_5023,N_4932);
nor U19572 (N_19572,N_561,N_8954);
nor U19573 (N_19573,N_3276,N_2518);
nand U19574 (N_19574,N_7454,N_8797);
xnor U19575 (N_19575,N_6200,N_4396);
nor U19576 (N_19576,N_7676,N_7518);
nand U19577 (N_19577,N_1369,N_2993);
nor U19578 (N_19578,N_1571,N_1452);
and U19579 (N_19579,N_7416,N_790);
and U19580 (N_19580,N_3332,N_4090);
xnor U19581 (N_19581,N_7960,N_1722);
nor U19582 (N_19582,N_8328,N_2709);
and U19583 (N_19583,N_443,N_6752);
or U19584 (N_19584,N_382,N_5512);
and U19585 (N_19585,N_6209,N_6676);
or U19586 (N_19586,N_589,N_8294);
or U19587 (N_19587,N_1375,N_5146);
nor U19588 (N_19588,N_6264,N_5133);
nor U19589 (N_19589,N_3892,N_4272);
and U19590 (N_19590,N_4976,N_4498);
or U19591 (N_19591,N_3425,N_991);
or U19592 (N_19592,N_1503,N_5931);
xor U19593 (N_19593,N_9356,N_1110);
or U19594 (N_19594,N_5780,N_538);
xor U19595 (N_19595,N_7623,N_6202);
or U19596 (N_19596,N_2376,N_6840);
xnor U19597 (N_19597,N_1394,N_9921);
nand U19598 (N_19598,N_9050,N_92);
nand U19599 (N_19599,N_6625,N_9613);
or U19600 (N_19600,N_3141,N_1348);
or U19601 (N_19601,N_7116,N_5939);
nand U19602 (N_19602,N_470,N_2394);
and U19603 (N_19603,N_58,N_6819);
nor U19604 (N_19604,N_4017,N_966);
or U19605 (N_19605,N_2592,N_5612);
nor U19606 (N_19606,N_5543,N_5895);
nor U19607 (N_19607,N_9598,N_4009);
or U19608 (N_19608,N_2170,N_7679);
or U19609 (N_19609,N_1617,N_4800);
nor U19610 (N_19610,N_8887,N_8152);
or U19611 (N_19611,N_573,N_3755);
and U19612 (N_19612,N_6638,N_6252);
and U19613 (N_19613,N_7487,N_4392);
and U19614 (N_19614,N_8286,N_7270);
nor U19615 (N_19615,N_1868,N_9199);
and U19616 (N_19616,N_206,N_4219);
nand U19617 (N_19617,N_1495,N_1535);
and U19618 (N_19618,N_6286,N_9048);
nor U19619 (N_19619,N_9081,N_5888);
nand U19620 (N_19620,N_104,N_4941);
nand U19621 (N_19621,N_5524,N_7356);
or U19622 (N_19622,N_2712,N_9841);
and U19623 (N_19623,N_1176,N_2811);
xor U19624 (N_19624,N_6586,N_950);
nand U19625 (N_19625,N_1708,N_7232);
or U19626 (N_19626,N_7341,N_7776);
and U19627 (N_19627,N_5792,N_2997);
nand U19628 (N_19628,N_3537,N_1679);
nor U19629 (N_19629,N_6879,N_9456);
nor U19630 (N_19630,N_8556,N_2646);
nand U19631 (N_19631,N_9424,N_5010);
and U19632 (N_19632,N_7856,N_1475);
nor U19633 (N_19633,N_4139,N_4815);
nand U19634 (N_19634,N_8774,N_6959);
and U19635 (N_19635,N_8040,N_5702);
nor U19636 (N_19636,N_3371,N_8860);
nand U19637 (N_19637,N_5751,N_8560);
and U19638 (N_19638,N_7028,N_2679);
nand U19639 (N_19639,N_6476,N_6201);
nor U19640 (N_19640,N_9692,N_3952);
nand U19641 (N_19641,N_7145,N_8041);
xor U19642 (N_19642,N_3173,N_8651);
and U19643 (N_19643,N_4794,N_1244);
nand U19644 (N_19644,N_1441,N_3702);
nand U19645 (N_19645,N_8366,N_4808);
nand U19646 (N_19646,N_9086,N_6260);
or U19647 (N_19647,N_6640,N_5112);
or U19648 (N_19648,N_8377,N_5532);
nor U19649 (N_19649,N_3386,N_3937);
and U19650 (N_19650,N_2802,N_7991);
nand U19651 (N_19651,N_632,N_2227);
and U19652 (N_19652,N_4541,N_4255);
nand U19653 (N_19653,N_7290,N_2180);
and U19654 (N_19654,N_7254,N_8210);
or U19655 (N_19655,N_5455,N_3302);
nand U19656 (N_19656,N_8867,N_3482);
nand U19657 (N_19657,N_5264,N_7575);
and U19658 (N_19658,N_5359,N_3686);
and U19659 (N_19659,N_7286,N_2631);
nand U19660 (N_19660,N_2813,N_7767);
nand U19661 (N_19661,N_6283,N_520);
or U19662 (N_19662,N_1666,N_6678);
xor U19663 (N_19663,N_6226,N_6008);
xnor U19664 (N_19664,N_7178,N_3950);
or U19665 (N_19665,N_2481,N_3594);
nand U19666 (N_19666,N_6801,N_668);
nor U19667 (N_19667,N_8184,N_5532);
and U19668 (N_19668,N_2286,N_4978);
nand U19669 (N_19669,N_8155,N_5755);
or U19670 (N_19670,N_4215,N_7389);
or U19671 (N_19671,N_7866,N_9800);
and U19672 (N_19672,N_6764,N_9002);
xor U19673 (N_19673,N_1758,N_8149);
and U19674 (N_19674,N_2650,N_3199);
nand U19675 (N_19675,N_6663,N_4066);
and U19676 (N_19676,N_7985,N_368);
or U19677 (N_19677,N_6345,N_3189);
nor U19678 (N_19678,N_1506,N_1160);
and U19679 (N_19679,N_1832,N_122);
nand U19680 (N_19680,N_3610,N_4723);
nor U19681 (N_19681,N_1429,N_389);
or U19682 (N_19682,N_9421,N_8680);
nor U19683 (N_19683,N_8797,N_7570);
or U19684 (N_19684,N_9788,N_3271);
nand U19685 (N_19685,N_4600,N_2429);
and U19686 (N_19686,N_707,N_4331);
or U19687 (N_19687,N_7683,N_8385);
or U19688 (N_19688,N_3440,N_5842);
and U19689 (N_19689,N_2774,N_5157);
nor U19690 (N_19690,N_9023,N_390);
xor U19691 (N_19691,N_6190,N_3570);
or U19692 (N_19692,N_1115,N_6500);
nor U19693 (N_19693,N_144,N_2942);
and U19694 (N_19694,N_6136,N_6011);
and U19695 (N_19695,N_3172,N_9910);
nor U19696 (N_19696,N_8699,N_6240);
nand U19697 (N_19697,N_6953,N_3629);
nand U19698 (N_19698,N_9929,N_1635);
or U19699 (N_19699,N_4022,N_5319);
nor U19700 (N_19700,N_5082,N_6163);
nand U19701 (N_19701,N_5797,N_2413);
and U19702 (N_19702,N_7629,N_2671);
and U19703 (N_19703,N_962,N_8292);
or U19704 (N_19704,N_7541,N_3346);
nand U19705 (N_19705,N_2564,N_7154);
and U19706 (N_19706,N_2900,N_8885);
nand U19707 (N_19707,N_7531,N_6214);
or U19708 (N_19708,N_5025,N_6861);
nand U19709 (N_19709,N_1500,N_4175);
and U19710 (N_19710,N_7379,N_4486);
nor U19711 (N_19711,N_1207,N_7100);
nand U19712 (N_19712,N_1893,N_618);
nor U19713 (N_19713,N_1877,N_1495);
or U19714 (N_19714,N_6285,N_7071);
or U19715 (N_19715,N_370,N_2205);
xor U19716 (N_19716,N_3017,N_7151);
and U19717 (N_19717,N_2389,N_8461);
or U19718 (N_19718,N_879,N_7403);
or U19719 (N_19719,N_9111,N_5999);
nor U19720 (N_19720,N_2625,N_5150);
and U19721 (N_19721,N_4977,N_3255);
or U19722 (N_19722,N_6060,N_2725);
nor U19723 (N_19723,N_792,N_9627);
nand U19724 (N_19724,N_3780,N_5786);
or U19725 (N_19725,N_5438,N_5329);
nand U19726 (N_19726,N_7186,N_5579);
nor U19727 (N_19727,N_7637,N_6357);
nand U19728 (N_19728,N_7366,N_3865);
nand U19729 (N_19729,N_6589,N_3539);
nand U19730 (N_19730,N_3374,N_7564);
xnor U19731 (N_19731,N_4165,N_4006);
nand U19732 (N_19732,N_2476,N_130);
or U19733 (N_19733,N_1272,N_5904);
and U19734 (N_19734,N_146,N_4981);
nand U19735 (N_19735,N_3036,N_1677);
nand U19736 (N_19736,N_3362,N_5611);
xnor U19737 (N_19737,N_8760,N_3396);
nor U19738 (N_19738,N_4223,N_634);
xor U19739 (N_19739,N_2025,N_9660);
xnor U19740 (N_19740,N_3304,N_1341);
or U19741 (N_19741,N_8205,N_2968);
nor U19742 (N_19742,N_8003,N_2553);
or U19743 (N_19743,N_9089,N_845);
xnor U19744 (N_19744,N_2044,N_5213);
or U19745 (N_19745,N_9847,N_3875);
and U19746 (N_19746,N_2776,N_4178);
and U19747 (N_19747,N_1053,N_7137);
nor U19748 (N_19748,N_4993,N_3247);
or U19749 (N_19749,N_4320,N_9980);
and U19750 (N_19750,N_5586,N_151);
nor U19751 (N_19751,N_7293,N_3451);
nor U19752 (N_19752,N_4531,N_3746);
nand U19753 (N_19753,N_2819,N_8739);
and U19754 (N_19754,N_7621,N_3792);
nand U19755 (N_19755,N_8042,N_9338);
nand U19756 (N_19756,N_8121,N_3300);
nor U19757 (N_19757,N_7922,N_6371);
nor U19758 (N_19758,N_4686,N_7571);
nor U19759 (N_19759,N_2446,N_7159);
nand U19760 (N_19760,N_2534,N_1819);
xnor U19761 (N_19761,N_5780,N_5695);
xnor U19762 (N_19762,N_4554,N_8314);
nor U19763 (N_19763,N_2159,N_3386);
nand U19764 (N_19764,N_4287,N_1193);
and U19765 (N_19765,N_5649,N_7044);
and U19766 (N_19766,N_9023,N_7294);
xor U19767 (N_19767,N_6161,N_3159);
nand U19768 (N_19768,N_7956,N_5178);
nor U19769 (N_19769,N_1652,N_5967);
and U19770 (N_19770,N_9435,N_5350);
and U19771 (N_19771,N_9535,N_4947);
or U19772 (N_19772,N_3302,N_9900);
nor U19773 (N_19773,N_2643,N_4734);
or U19774 (N_19774,N_1675,N_5918);
or U19775 (N_19775,N_3106,N_331);
nor U19776 (N_19776,N_6663,N_4529);
nand U19777 (N_19777,N_4786,N_1661);
or U19778 (N_19778,N_9523,N_8048);
or U19779 (N_19779,N_6949,N_4353);
nor U19780 (N_19780,N_7937,N_1320);
or U19781 (N_19781,N_4873,N_6907);
or U19782 (N_19782,N_1184,N_9849);
nand U19783 (N_19783,N_402,N_8582);
xor U19784 (N_19784,N_2749,N_1485);
nand U19785 (N_19785,N_953,N_9373);
nand U19786 (N_19786,N_8717,N_7759);
or U19787 (N_19787,N_1925,N_8863);
nor U19788 (N_19788,N_8685,N_3855);
or U19789 (N_19789,N_4403,N_1439);
nor U19790 (N_19790,N_1577,N_4304);
nor U19791 (N_19791,N_1655,N_5107);
nor U19792 (N_19792,N_2191,N_1041);
or U19793 (N_19793,N_5744,N_4758);
and U19794 (N_19794,N_9152,N_3412);
nand U19795 (N_19795,N_3500,N_5880);
and U19796 (N_19796,N_910,N_6596);
or U19797 (N_19797,N_9670,N_5273);
or U19798 (N_19798,N_9227,N_4142);
nor U19799 (N_19799,N_7513,N_9168);
or U19800 (N_19800,N_4533,N_4685);
or U19801 (N_19801,N_3805,N_9355);
or U19802 (N_19802,N_9388,N_3514);
and U19803 (N_19803,N_1253,N_1929);
and U19804 (N_19804,N_2669,N_6983);
or U19805 (N_19805,N_3817,N_844);
and U19806 (N_19806,N_5030,N_3343);
or U19807 (N_19807,N_3349,N_8500);
or U19808 (N_19808,N_9264,N_7766);
and U19809 (N_19809,N_8488,N_5311);
or U19810 (N_19810,N_9424,N_661);
or U19811 (N_19811,N_6579,N_1043);
or U19812 (N_19812,N_4305,N_902);
or U19813 (N_19813,N_7187,N_6364);
nor U19814 (N_19814,N_8917,N_9972);
or U19815 (N_19815,N_5527,N_6604);
and U19816 (N_19816,N_5482,N_488);
nor U19817 (N_19817,N_4754,N_8275);
or U19818 (N_19818,N_1150,N_6065);
nor U19819 (N_19819,N_4246,N_3403);
nor U19820 (N_19820,N_4897,N_3794);
xor U19821 (N_19821,N_9854,N_8469);
nand U19822 (N_19822,N_6834,N_3900);
and U19823 (N_19823,N_5081,N_4547);
nor U19824 (N_19824,N_7730,N_6578);
and U19825 (N_19825,N_4508,N_9795);
or U19826 (N_19826,N_8771,N_1265);
xnor U19827 (N_19827,N_8408,N_8564);
or U19828 (N_19828,N_1141,N_2740);
or U19829 (N_19829,N_6781,N_9305);
and U19830 (N_19830,N_8078,N_381);
and U19831 (N_19831,N_8017,N_3635);
or U19832 (N_19832,N_1534,N_8580);
or U19833 (N_19833,N_1870,N_3836);
nand U19834 (N_19834,N_7767,N_9574);
nand U19835 (N_19835,N_1335,N_8526);
and U19836 (N_19836,N_5210,N_8749);
or U19837 (N_19837,N_7947,N_581);
xor U19838 (N_19838,N_9773,N_6745);
or U19839 (N_19839,N_2913,N_377);
nor U19840 (N_19840,N_3715,N_2906);
nand U19841 (N_19841,N_2726,N_811);
and U19842 (N_19842,N_5455,N_1031);
nor U19843 (N_19843,N_2921,N_1027);
nand U19844 (N_19844,N_9559,N_6577);
and U19845 (N_19845,N_7653,N_3124);
and U19846 (N_19846,N_1813,N_1719);
and U19847 (N_19847,N_732,N_9234);
xnor U19848 (N_19848,N_9724,N_4135);
nand U19849 (N_19849,N_9362,N_8254);
nand U19850 (N_19850,N_2874,N_3357);
or U19851 (N_19851,N_7857,N_6159);
nand U19852 (N_19852,N_5328,N_6910);
nor U19853 (N_19853,N_3113,N_997);
or U19854 (N_19854,N_4609,N_4728);
nor U19855 (N_19855,N_3084,N_9272);
and U19856 (N_19856,N_2516,N_1432);
and U19857 (N_19857,N_4909,N_799);
or U19858 (N_19858,N_5826,N_8267);
nand U19859 (N_19859,N_4288,N_7031);
nor U19860 (N_19860,N_8305,N_7312);
or U19861 (N_19861,N_5862,N_1390);
and U19862 (N_19862,N_2165,N_2549);
nand U19863 (N_19863,N_3715,N_3898);
or U19864 (N_19864,N_6671,N_9785);
nand U19865 (N_19865,N_4052,N_9720);
or U19866 (N_19866,N_7628,N_7248);
nand U19867 (N_19867,N_9481,N_7315);
nor U19868 (N_19868,N_946,N_4665);
or U19869 (N_19869,N_3233,N_7129);
and U19870 (N_19870,N_1093,N_5272);
nor U19871 (N_19871,N_7790,N_2448);
nand U19872 (N_19872,N_7532,N_8797);
nand U19873 (N_19873,N_6983,N_5585);
and U19874 (N_19874,N_1579,N_9035);
nand U19875 (N_19875,N_1742,N_7337);
nand U19876 (N_19876,N_4006,N_1444);
and U19877 (N_19877,N_6294,N_6760);
nand U19878 (N_19878,N_5743,N_5139);
and U19879 (N_19879,N_1620,N_4457);
or U19880 (N_19880,N_6077,N_6595);
nor U19881 (N_19881,N_3095,N_5088);
nor U19882 (N_19882,N_1293,N_2523);
or U19883 (N_19883,N_7554,N_1033);
nor U19884 (N_19884,N_7358,N_2180);
or U19885 (N_19885,N_8496,N_4023);
nor U19886 (N_19886,N_6779,N_7075);
or U19887 (N_19887,N_3845,N_6738);
nand U19888 (N_19888,N_9905,N_4373);
nand U19889 (N_19889,N_8867,N_834);
nand U19890 (N_19890,N_7479,N_3596);
and U19891 (N_19891,N_6391,N_8751);
and U19892 (N_19892,N_1229,N_7138);
nor U19893 (N_19893,N_9570,N_8451);
and U19894 (N_19894,N_3080,N_8581);
or U19895 (N_19895,N_5609,N_7365);
or U19896 (N_19896,N_4583,N_5895);
xnor U19897 (N_19897,N_691,N_1209);
or U19898 (N_19898,N_7482,N_3647);
nand U19899 (N_19899,N_8491,N_7705);
nand U19900 (N_19900,N_4605,N_5343);
and U19901 (N_19901,N_6258,N_9098);
xnor U19902 (N_19902,N_9900,N_3875);
nor U19903 (N_19903,N_1498,N_2379);
or U19904 (N_19904,N_4312,N_9844);
nor U19905 (N_19905,N_8479,N_4232);
nor U19906 (N_19906,N_2001,N_9312);
or U19907 (N_19907,N_4208,N_1397);
nand U19908 (N_19908,N_9488,N_1660);
or U19909 (N_19909,N_1013,N_8702);
xnor U19910 (N_19910,N_5443,N_7065);
nor U19911 (N_19911,N_4335,N_1234);
or U19912 (N_19912,N_6344,N_6);
nor U19913 (N_19913,N_6575,N_8098);
nand U19914 (N_19914,N_9511,N_3154);
nand U19915 (N_19915,N_6446,N_7046);
nor U19916 (N_19916,N_3863,N_804);
and U19917 (N_19917,N_1830,N_3068);
or U19918 (N_19918,N_4522,N_7870);
xnor U19919 (N_19919,N_4007,N_3004);
nor U19920 (N_19920,N_2300,N_8394);
nor U19921 (N_19921,N_9859,N_6701);
and U19922 (N_19922,N_4573,N_1108);
nand U19923 (N_19923,N_477,N_5982);
nand U19924 (N_19924,N_5341,N_4361);
nor U19925 (N_19925,N_395,N_7932);
nand U19926 (N_19926,N_1325,N_3054);
or U19927 (N_19927,N_1733,N_8523);
and U19928 (N_19928,N_5289,N_2322);
or U19929 (N_19929,N_6124,N_1536);
xor U19930 (N_19930,N_9625,N_4563);
or U19931 (N_19931,N_8502,N_1265);
or U19932 (N_19932,N_6692,N_9368);
xor U19933 (N_19933,N_183,N_8574);
nand U19934 (N_19934,N_450,N_2649);
and U19935 (N_19935,N_2092,N_4088);
or U19936 (N_19936,N_4303,N_9270);
nand U19937 (N_19937,N_344,N_8634);
nand U19938 (N_19938,N_8672,N_5466);
and U19939 (N_19939,N_1714,N_230);
nor U19940 (N_19940,N_2970,N_9157);
nand U19941 (N_19941,N_6277,N_7803);
nor U19942 (N_19942,N_1940,N_222);
nor U19943 (N_19943,N_6998,N_8000);
nor U19944 (N_19944,N_7453,N_3216);
or U19945 (N_19945,N_3556,N_2175);
nor U19946 (N_19946,N_2734,N_6473);
and U19947 (N_19947,N_4333,N_5057);
and U19948 (N_19948,N_40,N_3601);
nor U19949 (N_19949,N_2004,N_2806);
nor U19950 (N_19950,N_5216,N_363);
nor U19951 (N_19951,N_5342,N_1865);
or U19952 (N_19952,N_2141,N_5558);
nor U19953 (N_19953,N_1225,N_1919);
nand U19954 (N_19954,N_671,N_1440);
or U19955 (N_19955,N_604,N_6451);
nand U19956 (N_19956,N_8284,N_3914);
nor U19957 (N_19957,N_1585,N_4091);
and U19958 (N_19958,N_3709,N_9090);
nand U19959 (N_19959,N_7066,N_6592);
or U19960 (N_19960,N_1191,N_717);
and U19961 (N_19961,N_2914,N_3794);
nor U19962 (N_19962,N_9802,N_1386);
nor U19963 (N_19963,N_8456,N_7979);
nor U19964 (N_19964,N_6509,N_5645);
or U19965 (N_19965,N_4970,N_4018);
or U19966 (N_19966,N_2662,N_1054);
or U19967 (N_19967,N_338,N_7025);
nor U19968 (N_19968,N_3584,N_2749);
xor U19969 (N_19969,N_2151,N_5600);
and U19970 (N_19970,N_3194,N_2210);
or U19971 (N_19971,N_2335,N_3198);
and U19972 (N_19972,N_5865,N_6028);
nand U19973 (N_19973,N_8994,N_8080);
and U19974 (N_19974,N_7038,N_5548);
xor U19975 (N_19975,N_5459,N_1582);
xnor U19976 (N_19976,N_2476,N_6685);
and U19977 (N_19977,N_5540,N_846);
nor U19978 (N_19978,N_7567,N_1838);
and U19979 (N_19979,N_3661,N_3856);
nand U19980 (N_19980,N_2210,N_6767);
or U19981 (N_19981,N_2833,N_5033);
nand U19982 (N_19982,N_8144,N_3960);
or U19983 (N_19983,N_5009,N_5928);
nand U19984 (N_19984,N_7865,N_7280);
xnor U19985 (N_19985,N_5440,N_5376);
nor U19986 (N_19986,N_4879,N_6457);
and U19987 (N_19987,N_1994,N_9873);
nor U19988 (N_19988,N_5079,N_2829);
nand U19989 (N_19989,N_6382,N_1480);
nand U19990 (N_19990,N_3381,N_7853);
nor U19991 (N_19991,N_5131,N_6247);
or U19992 (N_19992,N_6249,N_3411);
nand U19993 (N_19993,N_5621,N_214);
and U19994 (N_19994,N_9748,N_2517);
or U19995 (N_19995,N_4271,N_7885);
and U19996 (N_19996,N_9327,N_9437);
or U19997 (N_19997,N_7542,N_8566);
or U19998 (N_19998,N_7879,N_9618);
nand U19999 (N_19999,N_1424,N_6517);
and U20000 (N_20000,N_16145,N_15798);
nor U20001 (N_20001,N_10843,N_15609);
nor U20002 (N_20002,N_12622,N_16782);
nand U20003 (N_20003,N_15163,N_12069);
nor U20004 (N_20004,N_17952,N_14313);
and U20005 (N_20005,N_19933,N_19378);
or U20006 (N_20006,N_18378,N_17385);
and U20007 (N_20007,N_18429,N_12771);
and U20008 (N_20008,N_19942,N_18802);
or U20009 (N_20009,N_10550,N_16913);
and U20010 (N_20010,N_19062,N_18336);
and U20011 (N_20011,N_19253,N_10886);
nor U20012 (N_20012,N_13720,N_12170);
nand U20013 (N_20013,N_18966,N_10385);
and U20014 (N_20014,N_18829,N_18386);
and U20015 (N_20015,N_10303,N_17799);
xor U20016 (N_20016,N_19588,N_18854);
or U20017 (N_20017,N_13792,N_12264);
nand U20018 (N_20018,N_18831,N_19424);
nand U20019 (N_20019,N_11529,N_19739);
and U20020 (N_20020,N_17395,N_19830);
nor U20021 (N_20021,N_16176,N_12661);
or U20022 (N_20022,N_16970,N_17364);
nor U20023 (N_20023,N_18865,N_18475);
or U20024 (N_20024,N_16151,N_15262);
or U20025 (N_20025,N_15119,N_10906);
or U20026 (N_20026,N_15156,N_15277);
nand U20027 (N_20027,N_15837,N_17989);
nor U20028 (N_20028,N_19510,N_11234);
and U20029 (N_20029,N_19391,N_18684);
nor U20030 (N_20030,N_19372,N_14979);
nor U20031 (N_20031,N_18081,N_19072);
nor U20032 (N_20032,N_14527,N_18894);
nand U20033 (N_20033,N_13717,N_14236);
or U20034 (N_20034,N_13713,N_14326);
xnor U20035 (N_20035,N_11103,N_10893);
and U20036 (N_20036,N_12626,N_11134);
and U20037 (N_20037,N_18295,N_19808);
nor U20038 (N_20038,N_14186,N_17782);
or U20039 (N_20039,N_14916,N_17037);
nor U20040 (N_20040,N_16191,N_12013);
nand U20041 (N_20041,N_15496,N_15605);
or U20042 (N_20042,N_10549,N_10800);
nor U20043 (N_20043,N_16420,N_17715);
and U20044 (N_20044,N_18626,N_12516);
nor U20045 (N_20045,N_18342,N_15195);
and U20046 (N_20046,N_11487,N_15634);
and U20047 (N_20047,N_11098,N_15726);
nor U20048 (N_20048,N_19406,N_13835);
nor U20049 (N_20049,N_16582,N_17387);
or U20050 (N_20050,N_14135,N_17948);
nor U20051 (N_20051,N_15376,N_17704);
xnor U20052 (N_20052,N_15225,N_14548);
nand U20053 (N_20053,N_18754,N_10947);
and U20054 (N_20054,N_14910,N_11442);
or U20055 (N_20055,N_15470,N_15695);
nand U20056 (N_20056,N_18725,N_16687);
nand U20057 (N_20057,N_14219,N_13970);
nand U20058 (N_20058,N_10747,N_16999);
or U20059 (N_20059,N_18983,N_11105);
and U20060 (N_20060,N_16006,N_12790);
nand U20061 (N_20061,N_18516,N_19914);
nor U20062 (N_20062,N_15189,N_13111);
and U20063 (N_20063,N_18168,N_16923);
nor U20064 (N_20064,N_17055,N_18108);
nor U20065 (N_20065,N_10287,N_11754);
nand U20066 (N_20066,N_15118,N_18703);
nand U20067 (N_20067,N_16067,N_16453);
and U20068 (N_20068,N_10838,N_16048);
nand U20069 (N_20069,N_19023,N_12322);
nand U20070 (N_20070,N_13594,N_15629);
and U20071 (N_20071,N_10235,N_18412);
or U20072 (N_20072,N_18551,N_12256);
nor U20073 (N_20073,N_10286,N_14486);
and U20074 (N_20074,N_10433,N_13569);
nand U20075 (N_20075,N_11657,N_16032);
nand U20076 (N_20076,N_19851,N_10655);
nand U20077 (N_20077,N_14700,N_16513);
and U20078 (N_20078,N_19737,N_15797);
xor U20079 (N_20079,N_12357,N_18066);
nand U20080 (N_20080,N_18897,N_14083);
nand U20081 (N_20081,N_11341,N_16182);
and U20082 (N_20082,N_13666,N_13909);
and U20083 (N_20083,N_13616,N_10976);
nand U20084 (N_20084,N_19943,N_11252);
and U20085 (N_20085,N_12396,N_17409);
nor U20086 (N_20086,N_14944,N_12894);
xnor U20087 (N_20087,N_18032,N_17103);
nand U20088 (N_20088,N_15024,N_11015);
nand U20089 (N_20089,N_15446,N_16316);
nor U20090 (N_20090,N_15744,N_18648);
nor U20091 (N_20091,N_15557,N_12783);
or U20092 (N_20092,N_18491,N_10950);
nor U20093 (N_20093,N_16165,N_12455);
nand U20094 (N_20094,N_14908,N_19094);
xnor U20095 (N_20095,N_15848,N_11834);
and U20096 (N_20096,N_14407,N_10003);
or U20097 (N_20097,N_14725,N_17116);
nor U20098 (N_20098,N_13967,N_14786);
nor U20099 (N_20099,N_12282,N_15380);
nor U20100 (N_20100,N_14775,N_11711);
nand U20101 (N_20101,N_10635,N_15468);
and U20102 (N_20102,N_12454,N_16174);
and U20103 (N_20103,N_18227,N_13622);
xnor U20104 (N_20104,N_17611,N_19069);
or U20105 (N_20105,N_13833,N_19055);
xnor U20106 (N_20106,N_13269,N_14662);
nor U20107 (N_20107,N_11839,N_17299);
and U20108 (N_20108,N_15092,N_15227);
xor U20109 (N_20109,N_16585,N_11799);
nor U20110 (N_20110,N_11750,N_11936);
and U20111 (N_20111,N_11063,N_16347);
xnor U20112 (N_20112,N_16510,N_15103);
nor U20113 (N_20113,N_11583,N_18490);
and U20114 (N_20114,N_18415,N_13268);
and U20115 (N_20115,N_16371,N_16426);
and U20116 (N_20116,N_16500,N_17755);
nand U20117 (N_20117,N_18945,N_10474);
or U20118 (N_20118,N_13810,N_11037);
or U20119 (N_20119,N_11517,N_14035);
nand U20120 (N_20120,N_16203,N_18577);
and U20121 (N_20121,N_19027,N_11635);
xor U20122 (N_20122,N_19869,N_10046);
nand U20123 (N_20123,N_11587,N_16543);
or U20124 (N_20124,N_11380,N_10511);
nor U20125 (N_20125,N_18467,N_14619);
or U20126 (N_20126,N_18206,N_16801);
nor U20127 (N_20127,N_14715,N_19707);
or U20128 (N_20128,N_12685,N_19931);
nand U20129 (N_20129,N_19936,N_15234);
or U20130 (N_20130,N_19007,N_10837);
nand U20131 (N_20131,N_12280,N_10570);
nor U20132 (N_20132,N_18561,N_19556);
and U20133 (N_20133,N_15702,N_14465);
nor U20134 (N_20134,N_17711,N_13132);
and U20135 (N_20135,N_13438,N_15300);
nor U20136 (N_20136,N_19895,N_18417);
and U20137 (N_20137,N_16236,N_10610);
nor U20138 (N_20138,N_12506,N_14671);
xnor U20139 (N_20139,N_10817,N_19671);
and U20140 (N_20140,N_14383,N_19093);
or U20141 (N_20141,N_19147,N_10401);
nand U20142 (N_20142,N_17886,N_17283);
nand U20143 (N_20143,N_18827,N_18483);
nand U20144 (N_20144,N_15898,N_17644);
or U20145 (N_20145,N_13261,N_12347);
nand U20146 (N_20146,N_14508,N_18468);
and U20147 (N_20147,N_18004,N_15715);
nor U20148 (N_20148,N_19196,N_10486);
nor U20149 (N_20149,N_10249,N_18184);
nand U20150 (N_20150,N_17958,N_19102);
nor U20151 (N_20151,N_16608,N_15155);
or U20152 (N_20152,N_14626,N_18679);
and U20153 (N_20153,N_14966,N_16377);
and U20154 (N_20154,N_19300,N_13094);
or U20155 (N_20155,N_15378,N_10853);
nor U20156 (N_20156,N_19364,N_14356);
nor U20157 (N_20157,N_14951,N_12141);
or U20158 (N_20158,N_19243,N_13695);
and U20159 (N_20159,N_10971,N_13347);
nand U20160 (N_20160,N_12832,N_13276);
nand U20161 (N_20161,N_15064,N_17767);
nand U20162 (N_20162,N_19440,N_16264);
nand U20163 (N_20163,N_14180,N_15266);
nand U20164 (N_20164,N_16947,N_14649);
xnor U20165 (N_20165,N_19469,N_10146);
or U20166 (N_20166,N_15154,N_12067);
and U20167 (N_20167,N_12024,N_15908);
nand U20168 (N_20168,N_18987,N_19322);
nand U20169 (N_20169,N_11574,N_18165);
nand U20170 (N_20170,N_16992,N_13873);
or U20171 (N_20171,N_18989,N_15691);
and U20172 (N_20172,N_13487,N_10760);
nor U20173 (N_20173,N_13066,N_14831);
and U20174 (N_20174,N_19742,N_12393);
nand U20175 (N_20175,N_16899,N_18678);
and U20176 (N_20176,N_14431,N_12418);
nor U20177 (N_20177,N_16778,N_13669);
nor U20178 (N_20178,N_19946,N_13500);
nand U20179 (N_20179,N_16987,N_13034);
and U20180 (N_20180,N_11299,N_15739);
nor U20181 (N_20181,N_17049,N_19115);
and U20182 (N_20182,N_11162,N_16647);
nand U20183 (N_20183,N_17874,N_17238);
nand U20184 (N_20184,N_17041,N_12018);
nor U20185 (N_20185,N_18400,N_19838);
nand U20186 (N_20186,N_16574,N_10456);
nand U20187 (N_20187,N_18597,N_12496);
nand U20188 (N_20188,N_10767,N_16486);
nand U20189 (N_20189,N_14697,N_13402);
or U20190 (N_20190,N_13121,N_17268);
nand U20191 (N_20191,N_10031,N_14770);
nand U20192 (N_20192,N_14880,N_19290);
or U20193 (N_20193,N_17553,N_17211);
or U20194 (N_20194,N_13981,N_10794);
or U20195 (N_20195,N_10108,N_18898);
or U20196 (N_20196,N_10823,N_13912);
nor U20197 (N_20197,N_18602,N_17454);
nor U20198 (N_20198,N_15508,N_15895);
xnor U20199 (N_20199,N_16271,N_11766);
nor U20200 (N_20200,N_11680,N_18572);
and U20201 (N_20201,N_17453,N_18702);
or U20202 (N_20202,N_13295,N_14339);
nand U20203 (N_20203,N_12411,N_16502);
nor U20204 (N_20204,N_13257,N_14772);
nand U20205 (N_20205,N_18875,N_13263);
xor U20206 (N_20206,N_15777,N_19345);
xor U20207 (N_20207,N_15563,N_18789);
or U20208 (N_20208,N_14375,N_12546);
and U20209 (N_20209,N_15230,N_18394);
xnor U20210 (N_20210,N_15348,N_18076);
nand U20211 (N_20211,N_16818,N_13950);
nor U20212 (N_20212,N_12964,N_15520);
nor U20213 (N_20213,N_10464,N_15045);
nor U20214 (N_20214,N_11402,N_12556);
xnor U20215 (N_20215,N_14917,N_13396);
nand U20216 (N_20216,N_13504,N_11664);
nand U20217 (N_20217,N_19765,N_14126);
nand U20218 (N_20218,N_18884,N_16884);
nor U20219 (N_20219,N_19220,N_12521);
or U20220 (N_20220,N_13529,N_17583);
and U20221 (N_20221,N_19729,N_13310);
and U20222 (N_20222,N_18607,N_19884);
or U20223 (N_20223,N_17460,N_19398);
nor U20224 (N_20224,N_17209,N_19494);
and U20225 (N_20225,N_17178,N_11374);
nand U20226 (N_20226,N_11119,N_18482);
nor U20227 (N_20227,N_10231,N_19122);
and U20228 (N_20228,N_15580,N_16861);
nor U20229 (N_20229,N_13158,N_11684);
nand U20230 (N_20230,N_14437,N_11699);
nand U20231 (N_20231,N_15682,N_10214);
or U20232 (N_20232,N_13378,N_10058);
and U20233 (N_20233,N_10815,N_17911);
nand U20234 (N_20234,N_18244,N_19698);
nand U20235 (N_20235,N_18877,N_12284);
and U20236 (N_20236,N_17607,N_14381);
and U20237 (N_20237,N_17359,N_10674);
or U20238 (N_20238,N_16830,N_13341);
xor U20239 (N_20239,N_11740,N_13308);
nor U20240 (N_20240,N_15211,N_14468);
nor U20241 (N_20241,N_19258,N_18039);
nor U20242 (N_20242,N_10264,N_15914);
or U20243 (N_20243,N_13100,N_16382);
or U20244 (N_20244,N_14747,N_18781);
nand U20245 (N_20245,N_11367,N_10894);
or U20246 (N_20246,N_16017,N_18264);
and U20247 (N_20247,N_16731,N_10224);
nand U20248 (N_20248,N_13030,N_13324);
and U20249 (N_20249,N_12497,N_13973);
and U20250 (N_20250,N_16883,N_13822);
nand U20251 (N_20251,N_14791,N_18233);
and U20252 (N_20252,N_19908,N_12165);
or U20253 (N_20253,N_19218,N_12842);
nand U20254 (N_20254,N_13612,N_18376);
nor U20255 (N_20255,N_17648,N_19539);
nor U20256 (N_20256,N_10453,N_12490);
nand U20257 (N_20257,N_12400,N_13319);
or U20258 (N_20258,N_10504,N_12997);
and U20259 (N_20259,N_19558,N_18649);
nand U20260 (N_20260,N_12344,N_11040);
and U20261 (N_20261,N_16832,N_12057);
and U20262 (N_20262,N_19294,N_12804);
xor U20263 (N_20263,N_11533,N_15392);
or U20264 (N_20264,N_14382,N_11117);
nor U20265 (N_20265,N_13627,N_14585);
nor U20266 (N_20266,N_15000,N_14078);
nand U20267 (N_20267,N_15866,N_18586);
nor U20268 (N_20268,N_17568,N_16653);
and U20269 (N_20269,N_11530,N_18513);
nand U20270 (N_20270,N_15410,N_13510);
and U20271 (N_20271,N_19767,N_14530);
nand U20272 (N_20272,N_18056,N_15107);
nand U20273 (N_20273,N_11602,N_10186);
and U20274 (N_20274,N_16196,N_12920);
nand U20275 (N_20275,N_11389,N_13591);
nor U20276 (N_20276,N_12718,N_17516);
or U20277 (N_20277,N_11439,N_10983);
nand U20278 (N_20278,N_16454,N_10603);
or U20279 (N_20279,N_15342,N_13808);
or U20280 (N_20280,N_15864,N_17507);
xnor U20281 (N_20281,N_12656,N_13953);
nand U20282 (N_20282,N_15492,N_19392);
or U20283 (N_20283,N_13174,N_14643);
or U20284 (N_20284,N_18177,N_13856);
nor U20285 (N_20285,N_15823,N_18292);
xor U20286 (N_20286,N_17245,N_17430);
nor U20287 (N_20287,N_14852,N_11798);
nor U20288 (N_20288,N_10062,N_11783);
nand U20289 (N_20289,N_17270,N_11434);
or U20290 (N_20290,N_12243,N_13566);
nand U20291 (N_20291,N_10079,N_16589);
or U20292 (N_20292,N_16945,N_13831);
nand U20293 (N_20293,N_15919,N_10707);
or U20294 (N_20294,N_18954,N_19959);
and U20295 (N_20295,N_12432,N_15149);
or U20296 (N_20296,N_17484,N_17408);
nand U20297 (N_20297,N_14361,N_10721);
nand U20298 (N_20298,N_14600,N_18795);
or U20299 (N_20299,N_14642,N_12011);
nor U20300 (N_20300,N_13462,N_12873);
nand U20301 (N_20301,N_15199,N_19413);
and U20302 (N_20302,N_12876,N_13692);
or U20303 (N_20303,N_19816,N_18105);
nand U20304 (N_20304,N_19474,N_14255);
and U20305 (N_20305,N_16355,N_18212);
nand U20306 (N_20306,N_16240,N_16729);
nand U20307 (N_20307,N_18101,N_16706);
nor U20308 (N_20308,N_15180,N_14307);
nand U20309 (N_20309,N_14553,N_10898);
nand U20310 (N_20310,N_12985,N_18576);
and U20311 (N_20311,N_16673,N_12975);
nor U20312 (N_20312,N_10432,N_12169);
nand U20313 (N_20313,N_19041,N_11851);
nand U20314 (N_20314,N_19214,N_14137);
nand U20315 (N_20315,N_15491,N_10080);
nor U20316 (N_20316,N_18353,N_14647);
xnor U20317 (N_20317,N_12047,N_16696);
xor U20318 (N_20318,N_19454,N_18084);
xor U20319 (N_20319,N_12316,N_16385);
nor U20320 (N_20320,N_13760,N_17649);
nor U20321 (N_20321,N_19414,N_14761);
nor U20322 (N_20322,N_15831,N_17341);
nor U20323 (N_20323,N_10148,N_13334);
and U20324 (N_20324,N_19075,N_17119);
or U20325 (N_20325,N_10035,N_16774);
or U20326 (N_20326,N_12200,N_17301);
nand U20327 (N_20327,N_13196,N_17258);
and U20328 (N_20328,N_16935,N_18852);
nand U20329 (N_20329,N_14146,N_13367);
xor U20330 (N_20330,N_13489,N_17397);
and U20331 (N_20331,N_12222,N_18747);
and U20332 (N_20332,N_17700,N_11941);
and U20333 (N_20333,N_19501,N_13073);
nor U20334 (N_20334,N_18769,N_15521);
nand U20335 (N_20335,N_16550,N_17318);
xor U20336 (N_20336,N_19691,N_19705);
and U20337 (N_20337,N_11112,N_13383);
nand U20338 (N_20338,N_19160,N_18616);
nor U20339 (N_20339,N_15100,N_12690);
and U20340 (N_20340,N_18711,N_15417);
nor U20341 (N_20341,N_16091,N_19119);
or U20342 (N_20342,N_18362,N_19436);
or U20343 (N_20343,N_14018,N_10125);
nand U20344 (N_20344,N_19939,N_11360);
and U20345 (N_20345,N_13989,N_13182);
or U20346 (N_20346,N_18167,N_14388);
nor U20347 (N_20347,N_12734,N_15819);
nand U20348 (N_20348,N_18760,N_11942);
and U20349 (N_20349,N_18872,N_13446);
nor U20350 (N_20350,N_11713,N_13918);
or U20351 (N_20351,N_15556,N_19216);
nand U20352 (N_20352,N_13744,N_14445);
and U20353 (N_20353,N_12472,N_10615);
and U20354 (N_20354,N_14542,N_19423);
nor U20355 (N_20355,N_17146,N_18188);
and U20356 (N_20356,N_16120,N_10200);
and U20357 (N_20357,N_12445,N_18634);
nand U20358 (N_20358,N_10775,N_15612);
or U20359 (N_20359,N_15430,N_15809);
nor U20360 (N_20360,N_10447,N_19648);
nor U20361 (N_20361,N_19898,N_14765);
or U20362 (N_20362,N_11629,N_11430);
nand U20363 (N_20363,N_18030,N_13032);
nor U20364 (N_20364,N_19308,N_13765);
and U20365 (N_20365,N_16425,N_10923);
nor U20366 (N_20366,N_14670,N_14947);
and U20367 (N_20367,N_18220,N_14797);
nand U20368 (N_20368,N_13598,N_10710);
and U20369 (N_20369,N_10663,N_17087);
or U20370 (N_20370,N_16139,N_11106);
and U20371 (N_20371,N_13645,N_11688);
nand U20372 (N_20372,N_18202,N_19295);
nor U20373 (N_20373,N_17861,N_14351);
nand U20374 (N_20374,N_17127,N_16705);
xnor U20375 (N_20375,N_12305,N_17466);
nand U20376 (N_20376,N_17424,N_11893);
nand U20377 (N_20377,N_12801,N_18473);
nor U20378 (N_20378,N_16819,N_11366);
or U20379 (N_20379,N_18973,N_15686);
nor U20380 (N_20380,N_16522,N_18425);
xor U20381 (N_20381,N_11515,N_18826);
nor U20382 (N_20382,N_10203,N_13702);
nand U20383 (N_20383,N_10283,N_10400);
or U20384 (N_20384,N_15684,N_17512);
and U20385 (N_20385,N_17601,N_15037);
and U20386 (N_20386,N_12713,N_19383);
nor U20387 (N_20387,N_18825,N_11096);
or U20388 (N_20388,N_14172,N_16545);
nand U20389 (N_20389,N_16914,N_19449);
xnor U20390 (N_20390,N_10170,N_12738);
nor U20391 (N_20391,N_16432,N_14191);
nor U20392 (N_20392,N_11945,N_16759);
nand U20393 (N_20393,N_19944,N_14892);
xnor U20394 (N_20394,N_15731,N_16736);
nor U20395 (N_20395,N_18284,N_12761);
nor U20396 (N_20396,N_18990,N_19177);
and U20397 (N_20397,N_13718,N_10359);
xor U20398 (N_20398,N_18221,N_11612);
and U20399 (N_20399,N_15899,N_16666);
xnor U20400 (N_20400,N_18050,N_10904);
and U20401 (N_20401,N_12770,N_12823);
nor U20402 (N_20402,N_19042,N_14107);
and U20403 (N_20403,N_15801,N_12388);
nand U20404 (N_20404,N_14568,N_18409);
nor U20405 (N_20405,N_12935,N_13404);
or U20406 (N_20406,N_15409,N_15800);
nand U20407 (N_20407,N_17216,N_18563);
nor U20408 (N_20408,N_14130,N_13600);
and U20409 (N_20409,N_18106,N_18591);
nor U20410 (N_20410,N_11048,N_15012);
or U20411 (N_20411,N_17994,N_11128);
and U20412 (N_20412,N_14036,N_15770);
and U20413 (N_20413,N_14278,N_19883);
nor U20414 (N_20414,N_12740,N_18505);
and U20415 (N_20415,N_10226,N_11013);
xnor U20416 (N_20416,N_19754,N_19254);
nand U20417 (N_20417,N_10706,N_17647);
or U20418 (N_20418,N_14833,N_16202);
and U20419 (N_20419,N_13248,N_17795);
or U20420 (N_20420,N_13513,N_13919);
and U20421 (N_20421,N_19467,N_14332);
or U20422 (N_20422,N_11308,N_13472);
nand U20423 (N_20423,N_14194,N_16132);
or U20424 (N_20424,N_10051,N_10419);
and U20425 (N_20425,N_18932,N_17990);
or U20426 (N_20426,N_16364,N_13388);
nand U20427 (N_20427,N_19048,N_11372);
and U20428 (N_20428,N_14701,N_10605);
or U20429 (N_20429,N_15948,N_18833);
and U20430 (N_20430,N_14764,N_15534);
xnor U20431 (N_20431,N_19636,N_18621);
nor U20432 (N_20432,N_16835,N_11722);
and U20433 (N_20433,N_13551,N_12232);
or U20434 (N_20434,N_11057,N_10441);
nand U20435 (N_20435,N_19906,N_13398);
or U20436 (N_20436,N_18488,N_13162);
nor U20437 (N_20437,N_11120,N_13900);
nand U20438 (N_20438,N_14014,N_17546);
nand U20439 (N_20439,N_18959,N_14080);
and U20440 (N_20440,N_10854,N_14319);
or U20441 (N_20441,N_16243,N_17319);
nand U20442 (N_20442,N_13773,N_12444);
and U20443 (N_20443,N_10417,N_13145);
nand U20444 (N_20444,N_18904,N_14788);
xor U20445 (N_20445,N_13210,N_14462);
or U20446 (N_20446,N_17683,N_18097);
xor U20447 (N_20447,N_15734,N_11455);
and U20448 (N_20448,N_12541,N_15383);
and U20449 (N_20449,N_12756,N_19080);
nor U20450 (N_20450,N_12511,N_19609);
or U20451 (N_20451,N_15991,N_10420);
or U20452 (N_20452,N_16026,N_14011);
and U20453 (N_20453,N_18133,N_10418);
and U20454 (N_20454,N_10580,N_16002);
and U20455 (N_20455,N_19841,N_18532);
nor U20456 (N_20456,N_10814,N_14519);
or U20457 (N_20457,N_18015,N_15411);
xor U20458 (N_20458,N_11697,N_11328);
xnor U20459 (N_20459,N_19086,N_11695);
nand U20460 (N_20460,N_12270,N_10221);
and U20461 (N_20461,N_16200,N_17848);
or U20462 (N_20462,N_14438,N_12074);
nor U20463 (N_20463,N_13571,N_17112);
nand U20464 (N_20464,N_15650,N_11449);
or U20465 (N_20465,N_13401,N_18594);
nor U20466 (N_20466,N_12125,N_15335);
nand U20467 (N_20467,N_14592,N_16721);
and U20468 (N_20468,N_13239,N_14022);
or U20469 (N_20469,N_15829,N_12566);
nand U20470 (N_20470,N_17016,N_19833);
nand U20471 (N_20471,N_17936,N_10495);
nand U20472 (N_20472,N_13786,N_19357);
nand U20473 (N_20473,N_15670,N_13540);
or U20474 (N_20474,N_15497,N_16526);
or U20475 (N_20475,N_12466,N_14760);
nor U20476 (N_20476,N_18028,N_14932);
and U20477 (N_20477,N_19486,N_11866);
nand U20478 (N_20478,N_14962,N_17377);
xnor U20479 (N_20479,N_10295,N_17001);
and U20480 (N_20480,N_19514,N_10074);
nor U20481 (N_20481,N_19587,N_17698);
nand U20482 (N_20482,N_15029,N_16788);
nand U20483 (N_20483,N_10805,N_13603);
or U20484 (N_20484,N_16609,N_16224);
nand U20485 (N_20485,N_10064,N_13457);
nand U20486 (N_20486,N_17339,N_15501);
and U20487 (N_20487,N_17889,N_19778);
nand U20488 (N_20488,N_14805,N_12360);
nor U20489 (N_20489,N_13002,N_18873);
nand U20490 (N_20490,N_16905,N_17233);
nor U20491 (N_20491,N_18855,N_14494);
or U20492 (N_20492,N_14961,N_18350);
nor U20493 (N_20493,N_10779,N_18224);
xor U20494 (N_20494,N_13924,N_15441);
nand U20495 (N_20495,N_19517,N_12769);
and U20496 (N_20496,N_19015,N_11445);
nand U20497 (N_20497,N_17515,N_18250);
nor U20498 (N_20498,N_17605,N_15913);
nand U20499 (N_20499,N_19134,N_16979);
nand U20500 (N_20500,N_18900,N_13920);
and U20501 (N_20501,N_10571,N_13763);
and U20502 (N_20502,N_12422,N_19704);
or U20503 (N_20503,N_12932,N_10658);
or U20504 (N_20504,N_14893,N_13508);
nor U20505 (N_20505,N_19969,N_17951);
and U20506 (N_20506,N_14090,N_16433);
nand U20507 (N_20507,N_16577,N_10618);
nand U20508 (N_20508,N_18985,N_18200);
nor U20509 (N_20509,N_12374,N_18263);
and U20510 (N_20510,N_14869,N_19269);
or U20511 (N_20511,N_11431,N_19475);
or U20512 (N_20512,N_19664,N_10820);
or U20513 (N_20513,N_16124,N_12505);
and U20514 (N_20514,N_19133,N_11420);
and U20515 (N_20515,N_12574,N_15964);
and U20516 (N_20516,N_13387,N_17901);
or U20517 (N_20517,N_16015,N_15827);
nor U20518 (N_20518,N_19770,N_16390);
or U20519 (N_20519,N_12077,N_15165);
and U20520 (N_20520,N_13783,N_18557);
and U20521 (N_20521,N_16564,N_12272);
and U20522 (N_20522,N_12318,N_17326);
nor U20523 (N_20523,N_10672,N_17243);
or U20524 (N_20524,N_12750,N_10006);
nand U20525 (N_20525,N_10201,N_12321);
nand U20526 (N_20526,N_14546,N_18969);
nor U20527 (N_20527,N_17346,N_17248);
nor U20528 (N_20528,N_10182,N_16904);
nand U20529 (N_20529,N_13068,N_13678);
or U20530 (N_20530,N_16926,N_15934);
or U20531 (N_20531,N_16590,N_10827);
nand U20532 (N_20532,N_15836,N_13202);
xnor U20533 (N_20533,N_13582,N_10253);
and U20534 (N_20534,N_14976,N_19994);
or U20535 (N_20535,N_10860,N_19082);
xnor U20536 (N_20536,N_14963,N_11330);
nor U20537 (N_20537,N_19232,N_15388);
nand U20538 (N_20538,N_18778,N_10387);
and U20539 (N_20539,N_10951,N_13284);
or U20540 (N_20540,N_10689,N_17150);
and U20541 (N_20541,N_15402,N_18289);
and U20542 (N_20542,N_17493,N_16291);
or U20543 (N_20543,N_11543,N_19495);
nand U20544 (N_20544,N_10491,N_18564);
and U20545 (N_20545,N_18753,N_18587);
and U20546 (N_20546,N_14132,N_15939);
and U20547 (N_20547,N_10268,N_16210);
nand U20548 (N_20548,N_18145,N_17297);
nor U20549 (N_20549,N_15906,N_16537);
nor U20550 (N_20550,N_12250,N_14795);
and U20551 (N_20551,N_19791,N_12767);
nand U20552 (N_20552,N_11816,N_17059);
or U20553 (N_20553,N_15428,N_15785);
nand U20554 (N_20554,N_15636,N_19256);
and U20555 (N_20555,N_13085,N_14677);
or U20556 (N_20556,N_12676,N_17187);
or U20557 (N_20557,N_14338,N_13381);
nand U20558 (N_20558,N_19755,N_14498);
or U20559 (N_20559,N_11710,N_18837);
or U20560 (N_20560,N_11157,N_13816);
nor U20561 (N_20561,N_12308,N_11746);
xnor U20562 (N_20562,N_11237,N_17392);
nand U20563 (N_20563,N_19342,N_13966);
and U20564 (N_20564,N_13634,N_10336);
nand U20565 (N_20565,N_17955,N_19162);
nor U20566 (N_20566,N_19565,N_12206);
and U20567 (N_20567,N_15998,N_16702);
and U20568 (N_20568,N_18044,N_11671);
xnor U20569 (N_20569,N_10771,N_11762);
and U20570 (N_20570,N_12604,N_14998);
and U20571 (N_20571,N_10668,N_15067);
nor U20572 (N_20572,N_18078,N_13335);
and U20573 (N_20573,N_18629,N_12555);
and U20574 (N_20574,N_13371,N_10131);
and U20575 (N_20575,N_10684,N_15741);
or U20576 (N_20576,N_18928,N_14844);
nand U20577 (N_20577,N_18123,N_11407);
or U20578 (N_20578,N_16780,N_15135);
and U20579 (N_20579,N_17943,N_11604);
nand U20580 (N_20580,N_15796,N_11287);
and U20581 (N_20581,N_16791,N_18309);
or U20582 (N_20582,N_19650,N_15054);
nor U20583 (N_20583,N_10828,N_17157);
and U20584 (N_20584,N_15989,N_16627);
nor U20585 (N_20585,N_19912,N_11167);
and U20586 (N_20586,N_14259,N_12923);
and U20587 (N_20587,N_12635,N_14913);
and U20588 (N_20588,N_10124,N_17020);
nor U20589 (N_20589,N_17391,N_16299);
xor U20590 (N_20590,N_10786,N_16255);
and U20591 (N_20591,N_10157,N_19780);
or U20592 (N_20592,N_12345,N_12902);
or U20593 (N_20593,N_12515,N_19998);
nor U20594 (N_20594,N_13927,N_11319);
xor U20595 (N_20595,N_15483,N_12926);
nor U20596 (N_20596,N_17776,N_17923);
nand U20597 (N_20597,N_14628,N_19934);
nand U20598 (N_20598,N_11582,N_19081);
xnor U20599 (N_20599,N_17739,N_14825);
or U20600 (N_20600,N_11944,N_13313);
or U20601 (N_20601,N_14767,N_14418);
or U20602 (N_20602,N_18484,N_14896);
nor U20603 (N_20603,N_15585,N_10716);
or U20604 (N_20604,N_15389,N_11613);
nor U20605 (N_20605,N_13222,N_15477);
nand U20606 (N_20606,N_19288,N_12868);
and U20607 (N_20607,N_11853,N_17534);
or U20608 (N_20608,N_19555,N_18502);
xnor U20609 (N_20609,N_10502,N_10025);
or U20610 (N_20610,N_12226,N_13008);
or U20611 (N_20611,N_11058,N_18571);
or U20612 (N_20612,N_11884,N_15905);
and U20613 (N_20613,N_14837,N_12230);
xnor U20614 (N_20614,N_14613,N_13775);
and U20615 (N_20615,N_14826,N_18096);
or U20616 (N_20616,N_16903,N_10220);
nor U20617 (N_20617,N_18298,N_17149);
or U20618 (N_20618,N_13821,N_17860);
nor U20619 (N_20619,N_16665,N_14596);
and U20620 (N_20620,N_11969,N_14425);
and U20621 (N_20621,N_14127,N_18950);
nor U20622 (N_20622,N_12957,N_18688);
nand U20623 (N_20623,N_13680,N_12408);
or U20624 (N_20624,N_13844,N_12911);
or U20625 (N_20625,N_11669,N_13573);
nor U20626 (N_20626,N_12379,N_18034);
or U20627 (N_20627,N_13498,N_14806);
and U20628 (N_20628,N_13350,N_11871);
and U20629 (N_20629,N_10442,N_11401);
and U20630 (N_20630,N_19500,N_17986);
and U20631 (N_20631,N_14807,N_15060);
nor U20632 (N_20632,N_13080,N_10755);
and U20633 (N_20633,N_11879,N_10749);
or U20634 (N_20634,N_17887,N_16667);
nor U20635 (N_20635,N_11548,N_13558);
nor U20636 (N_20636,N_10119,N_10555);
nand U20637 (N_20637,N_19624,N_19489);
nand U20638 (N_20638,N_10228,N_11404);
nand U20639 (N_20639,N_19916,N_16285);
nor U20640 (N_20640,N_15122,N_14652);
nand U20641 (N_20641,N_11682,N_12727);
nor U20642 (N_20642,N_18099,N_19402);
nand U20643 (N_20643,N_17810,N_18146);
and U20644 (N_20644,N_17508,N_17148);
or U20645 (N_20645,N_16836,N_13863);
nor U20646 (N_20646,N_10503,N_13562);
nand U20647 (N_20647,N_19656,N_15968);
nand U20648 (N_20648,N_14506,N_18141);
nor U20649 (N_20649,N_10241,N_12399);
nand U20650 (N_20650,N_19649,N_10151);
or U20651 (N_20651,N_16248,N_17394);
and U20652 (N_20652,N_10057,N_15552);
nor U20653 (N_20653,N_12395,N_15644);
nor U20654 (N_20654,N_16761,N_19123);
or U20655 (N_20655,N_15860,N_17764);
or U20656 (N_20656,N_10880,N_10413);
or U20657 (N_20657,N_18210,N_14502);
nor U20658 (N_20658,N_18439,N_18065);
and U20659 (N_20659,N_13887,N_13436);
nor U20660 (N_20660,N_18686,N_14380);
and U20661 (N_20661,N_17521,N_12421);
or U20662 (N_20662,N_14975,N_11450);
and U20663 (N_20663,N_15865,N_14363);
xor U20664 (N_20664,N_15010,N_10634);
or U20665 (N_20665,N_10473,N_13320);
and U20666 (N_20666,N_10890,N_13014);
nor U20667 (N_20667,N_11763,N_10351);
and U20668 (N_20668,N_15641,N_15938);
nor U20669 (N_20669,N_13391,N_15361);
nand U20670 (N_20670,N_12708,N_19409);
or U20671 (N_20671,N_18531,N_19144);
or U20672 (N_20672,N_11080,N_17573);
and U20673 (N_20673,N_10242,N_10691);
nand U20674 (N_20674,N_16869,N_14450);
nor U20675 (N_20675,N_14340,N_11557);
nand U20676 (N_20676,N_17646,N_15778);
or U20677 (N_20677,N_19330,N_16393);
or U20678 (N_20678,N_16456,N_13007);
nand U20679 (N_20679,N_15790,N_14496);
nor U20680 (N_20680,N_15545,N_18981);
nor U20681 (N_20681,N_10540,N_10300);
nor U20682 (N_20682,N_18726,N_12413);
or U20683 (N_20683,N_17817,N_18625);
nand U20684 (N_20684,N_13703,N_16876);
nor U20685 (N_20685,N_17048,N_10412);
nand U20686 (N_20686,N_17545,N_19642);
xor U20687 (N_20687,N_14741,N_14302);
nand U20688 (N_20688,N_12262,N_16223);
and U20689 (N_20689,N_12737,N_14633);
or U20690 (N_20690,N_16854,N_11812);
nand U20691 (N_20691,N_17634,N_18555);
or U20692 (N_20692,N_16887,N_14115);
xnor U20693 (N_20693,N_19150,N_19832);
and U20694 (N_20694,N_10979,N_15298);
nand U20695 (N_20695,N_18411,N_15197);
nor U20696 (N_20696,N_11737,N_12747);
nor U20697 (N_20697,N_12475,N_11661);
and U20698 (N_20698,N_13670,N_12487);
or U20699 (N_20699,N_17797,N_10554);
nand U20700 (N_20700,N_13312,N_19516);
nor U20701 (N_20701,N_15274,N_16871);
xnor U20702 (N_20702,N_10531,N_12136);
and U20703 (N_20703,N_10492,N_12438);
and U20704 (N_20704,N_16828,N_16515);
nand U20705 (N_20705,N_19678,N_16900);
nor U20706 (N_20706,N_14708,N_10252);
xor U20707 (N_20707,N_15314,N_16917);
nand U20708 (N_20708,N_18528,N_18414);
or U20709 (N_20709,N_15033,N_17458);
or U20710 (N_20710,N_12211,N_17063);
xnor U20711 (N_20711,N_14742,N_19405);
and U20712 (N_20712,N_16029,N_11745);
and U20713 (N_20713,N_12443,N_13771);
or U20714 (N_20714,N_11731,N_15594);
xnor U20715 (N_20715,N_14784,N_17821);
and U20716 (N_20716,N_13711,N_12274);
nor U20717 (N_20717,N_16288,N_12150);
xnor U20718 (N_20718,N_19272,N_14776);
nand U20719 (N_20719,N_14283,N_15498);
nor U20720 (N_20720,N_17575,N_11008);
or U20721 (N_20721,N_19411,N_19868);
and U20722 (N_20722,N_17082,N_14160);
xnor U20723 (N_20723,N_15952,N_17025);
xor U20724 (N_20724,N_12450,N_13701);
nor U20725 (N_20725,N_15728,N_14271);
nand U20726 (N_20726,N_10259,N_18256);
nand U20727 (N_20727,N_10468,N_11828);
and U20728 (N_20728,N_12287,N_16910);
and U20729 (N_20729,N_18714,N_13021);
nand U20730 (N_20730,N_15773,N_17447);
nor U20731 (N_20731,N_10704,N_18804);
or U20732 (N_20732,N_10928,N_11491);
and U20733 (N_20733,N_17040,N_18705);
nor U20734 (N_20734,N_12053,N_17617);
nand U20735 (N_20735,N_11971,N_12323);
and U20736 (N_20736,N_19084,N_10440);
and U20737 (N_20737,N_17350,N_12174);
nand U20738 (N_20738,N_14549,N_19697);
nor U20739 (N_20739,N_13445,N_19738);
xnor U20740 (N_20740,N_12480,N_12020);
or U20741 (N_20741,N_10012,N_11030);
or U20742 (N_20742,N_14387,N_16039);
or U20743 (N_20743,N_11980,N_17723);
nor U20744 (N_20744,N_18961,N_11470);
nor U20745 (N_20745,N_16314,N_19477);
nor U20746 (N_20746,N_14885,N_10307);
and U20747 (N_20747,N_19151,N_12215);
nor U20748 (N_20748,N_12075,N_12087);
nand U20749 (N_20749,N_16056,N_11647);
nand U20750 (N_20750,N_14591,N_18025);
and U20751 (N_20751,N_11031,N_11553);
nor U20752 (N_20752,N_17287,N_14056);
and U20753 (N_20753,N_11474,N_17363);
nor U20754 (N_20754,N_12609,N_18019);
nor U20755 (N_20755,N_10518,N_13455);
nor U20756 (N_20756,N_17244,N_15071);
xnor U20757 (N_20757,N_10757,N_14930);
nor U20758 (N_20758,N_19618,N_11344);
and U20759 (N_20759,N_12089,N_10713);
or U20760 (N_20760,N_17381,N_17626);
nor U20761 (N_20761,N_14617,N_13448);
or U20762 (N_20762,N_11068,N_14605);
nand U20763 (N_20763,N_16310,N_17618);
or U20764 (N_20764,N_12491,N_10097);
nor U20765 (N_20765,N_18290,N_19181);
nor U20766 (N_20766,N_18234,N_16599);
nor U20767 (N_20767,N_11077,N_17778);
or U20768 (N_20768,N_11735,N_15538);
or U20769 (N_20769,N_19061,N_10092);
nor U20770 (N_20770,N_10551,N_15957);
nor U20771 (N_20771,N_14290,N_16695);
nand U20772 (N_20772,N_16231,N_15216);
or U20773 (N_20773,N_19843,N_18740);
nand U20774 (N_20774,N_10437,N_14804);
xnor U20775 (N_20775,N_16095,N_15742);
xor U20776 (N_20776,N_18020,N_12818);
xnor U20777 (N_20777,N_15282,N_19465);
nor U20778 (N_20778,N_12901,N_13672);
nand U20779 (N_20779,N_18535,N_11904);
nand U20780 (N_20780,N_15111,N_19658);
and U20781 (N_20781,N_17478,N_17892);
nand U20782 (N_20782,N_14364,N_12372);
or U20783 (N_20783,N_19067,N_15662);
nor U20784 (N_20784,N_18344,N_10248);
or U20785 (N_20785,N_14785,N_11133);
or U20786 (N_20786,N_17740,N_11922);
nand U20787 (N_20787,N_15170,N_11300);
and U20788 (N_20788,N_16356,N_16156);
nor U20789 (N_20789,N_18435,N_17905);
nor U20790 (N_20790,N_15942,N_11107);
nor U20791 (N_20791,N_12633,N_15231);
xor U20792 (N_20792,N_19370,N_18335);
or U20793 (N_20793,N_12822,N_16096);
or U20794 (N_20794,N_16554,N_14419);
nand U20795 (N_20795,N_11188,N_13377);
nor U20796 (N_20796,N_13651,N_15705);
nor U20797 (N_20797,N_12110,N_15370);
and U20798 (N_20798,N_12513,N_16329);
or U20799 (N_20799,N_12430,N_19878);
nor U20800 (N_20800,N_12135,N_11622);
nor U20801 (N_20801,N_11046,N_17499);
nor U20802 (N_20802,N_17088,N_14231);
or U20803 (N_20803,N_17973,N_18451);
xor U20804 (N_20804,N_12692,N_14451);
nor U20805 (N_20805,N_12986,N_11819);
nor U20806 (N_20806,N_13845,N_14734);
or U20807 (N_20807,N_11920,N_13605);
and U20808 (N_20808,N_11747,N_15222);
or U20809 (N_20809,N_14595,N_19471);
nand U20810 (N_20810,N_17084,N_11415);
nor U20811 (N_20811,N_14969,N_15725);
nand U20812 (N_20812,N_11393,N_17434);
and U20813 (N_20813,N_13192,N_19749);
nor U20814 (N_20814,N_11829,N_14249);
and U20815 (N_20815,N_15013,N_14594);
and U20816 (N_20816,N_19515,N_19677);
or U20817 (N_20817,N_12971,N_16055);
or U20818 (N_20818,N_11859,N_19619);
nor U20819 (N_20819,N_15805,N_16009);
or U20820 (N_20820,N_17981,N_17783);
nor U20821 (N_20821,N_14886,N_12792);
nor U20822 (N_20822,N_12291,N_19240);
nor U20823 (N_20823,N_10011,N_13664);
xor U20824 (N_20824,N_16948,N_19992);
xnor U20825 (N_20825,N_17047,N_18142);
and U20826 (N_20826,N_14724,N_13755);
or U20827 (N_20827,N_11454,N_10831);
nor U20828 (N_20828,N_13351,N_18757);
or U20829 (N_20829,N_17304,N_11124);
or U20830 (N_20830,N_16752,N_15787);
nand U20831 (N_20831,N_11545,N_15788);
or U20832 (N_20832,N_15614,N_17004);
nor U20833 (N_20833,N_18860,N_11110);
and U20834 (N_20834,N_19132,N_10692);
or U20835 (N_20835,N_18474,N_11625);
and U20836 (N_20836,N_12904,N_17678);
nor U20837 (N_20837,N_13223,N_10350);
and U20838 (N_20838,N_14094,N_16807);
nor U20839 (N_20839,N_15365,N_11914);
nor U20840 (N_20840,N_17717,N_10389);
nor U20841 (N_20841,N_14493,N_12937);
nand U20842 (N_20842,N_12046,N_16684);
nor U20843 (N_20843,N_17188,N_19487);
nor U20844 (N_20844,N_14346,N_13240);
and U20845 (N_20845,N_14817,N_11443);
xor U20846 (N_20846,N_15622,N_11966);
or U20847 (N_20847,N_11976,N_12637);
nand U20848 (N_20848,N_14012,N_12889);
xor U20849 (N_20849,N_14678,N_19993);
nor U20850 (N_20850,N_19314,N_18632);
nor U20851 (N_20851,N_15871,N_12908);
xor U20852 (N_20852,N_12554,N_11787);
nand U20853 (N_20853,N_14650,N_19688);
or U20854 (N_20854,N_16568,N_14082);
or U20855 (N_20855,N_16654,N_15730);
and U20856 (N_20856,N_14543,N_14396);
nor U20857 (N_20857,N_13877,N_10280);
or U20858 (N_20858,N_14748,N_16942);
or U20859 (N_20859,N_19473,N_12577);
nand U20860 (N_20860,N_16457,N_12848);
or U20861 (N_20861,N_14328,N_19098);
nand U20862 (N_20862,N_14739,N_11220);
or U20863 (N_20863,N_17608,N_17998);
xnor U20864 (N_20864,N_14489,N_12309);
or U20865 (N_20865,N_15332,N_17472);
and U20866 (N_20866,N_19603,N_19178);
nor U20867 (N_20867,N_10136,N_13155);
nand U20868 (N_20868,N_18160,N_12351);
nor U20869 (N_20869,N_19175,N_11703);
or U20870 (N_20870,N_15995,N_17807);
and U20871 (N_20871,N_17875,N_13724);
and U20872 (N_20872,N_17633,N_10363);
and U20873 (N_20873,N_11091,N_16166);
nand U20874 (N_20874,N_10366,N_15813);
nand U20875 (N_20875,N_13675,N_10731);
or U20876 (N_20876,N_15117,N_13386);
nor U20877 (N_20877,N_17570,N_13168);
nor U20878 (N_20878,N_17449,N_19375);
and U20879 (N_20879,N_15279,N_16540);
or U20880 (N_20880,N_14349,N_11095);
nand U20881 (N_20881,N_14663,N_14689);
nand U20882 (N_20882,N_14226,N_13083);
or U20883 (N_20883,N_14156,N_19675);
or U20884 (N_20884,N_11067,N_10187);
or U20885 (N_20885,N_19815,N_18751);
or U20886 (N_20886,N_11973,N_10380);
nand U20887 (N_20887,N_19255,N_18500);
nand U20888 (N_20888,N_13235,N_19444);
or U20889 (N_20889,N_15717,N_16881);
nand U20890 (N_20890,N_10609,N_17069);
or U20891 (N_20891,N_17292,N_16941);
nor U20892 (N_20892,N_17859,N_14882);
nor U20893 (N_20893,N_13317,N_11693);
nand U20894 (N_20894,N_11298,N_12489);
xor U20895 (N_20895,N_16571,N_11744);
nor U20896 (N_20896,N_15127,N_19238);
nand U20897 (N_20897,N_12041,N_13247);
nand U20898 (N_20898,N_18863,N_18548);
nor U20899 (N_20899,N_10619,N_12531);
or U20900 (N_20900,N_11297,N_16785);
and U20901 (N_20901,N_11278,N_16770);
nand U20902 (N_20902,N_12797,N_17221);
or U20903 (N_20903,N_17619,N_11927);
nand U20904 (N_20904,N_11466,N_16756);
xnor U20905 (N_20905,N_10402,N_17729);
nor U20906 (N_20906,N_13801,N_10493);
nor U20907 (N_20907,N_18283,N_13957);
or U20908 (N_20908,N_16476,N_10465);
nor U20909 (N_20909,N_17984,N_14836);
nor U20910 (N_20910,N_11805,N_10260);
nand U20911 (N_20911,N_10878,N_14622);
or U20912 (N_20912,N_13751,N_13348);
nor U20913 (N_20913,N_13668,N_15595);
nor U20914 (N_20914,N_17086,N_16890);
xor U20915 (N_20915,N_12884,N_16130);
or U20916 (N_20916,N_12257,N_15138);
nand U20917 (N_20917,N_10245,N_16193);
nand U20918 (N_20918,N_13805,N_16459);
xnor U20919 (N_20919,N_15587,N_14420);
nor U20920 (N_20920,N_10472,N_18619);
and U20921 (N_20921,N_11377,N_15359);
or U20922 (N_20922,N_19553,N_18257);
nor U20923 (N_20923,N_18403,N_15607);
nor U20924 (N_20924,N_14184,N_14353);
nand U20925 (N_20925,N_13004,N_17770);
or U20926 (N_20926,N_15651,N_16792);
nand U20927 (N_20927,N_18169,N_19719);
nor U20928 (N_20928,N_13169,N_11223);
and U20929 (N_20929,N_18080,N_13704);
xor U20930 (N_20930,N_16268,N_13642);
xor U20931 (N_20931,N_19230,N_10274);
and U20932 (N_20932,N_18410,N_17410);
and U20933 (N_20933,N_15746,N_14469);
nor U20934 (N_20934,N_16350,N_15986);
and U20935 (N_20935,N_15269,N_12778);
nor U20936 (N_20936,N_15646,N_11329);
or U20937 (N_20937,N_12325,N_13277);
or U20938 (N_20938,N_14994,N_17895);
and U20939 (N_20939,N_18090,N_19760);
nand U20940 (N_20940,N_10397,N_18903);
xnor U20941 (N_20941,N_14832,N_19149);
nor U20942 (N_20942,N_16082,N_12482);
nor U20943 (N_20943,N_12187,N_15701);
or U20944 (N_20944,N_13188,N_13241);
nor U20945 (N_20945,N_14737,N_19652);
nand U20946 (N_20946,N_19348,N_14798);
or U20947 (N_20947,N_14329,N_18673);
and U20948 (N_20948,N_11155,N_16634);
nand U20949 (N_20949,N_13012,N_16762);
nor U20950 (N_20950,N_10071,N_12867);
nand U20951 (N_20951,N_12817,N_13654);
nand U20952 (N_20952,N_14171,N_11650);
nand U20953 (N_20953,N_14850,N_11172);
nor U20954 (N_20954,N_10873,N_13964);
or U20955 (N_20955,N_12665,N_12117);
nor U20956 (N_20956,N_16373,N_11753);
or U20957 (N_20957,N_14125,N_19478);
or U20958 (N_20958,N_17597,N_11649);
nand U20959 (N_20959,N_19853,N_12246);
nand U20960 (N_20960,N_11705,N_14923);
xnor U20961 (N_20961,N_12424,N_16059);
xnor U20962 (N_20962,N_16583,N_12026);
nor U20963 (N_20963,N_11121,N_14333);
nand U20964 (N_20964,N_19720,N_14783);
and U20965 (N_20965,N_19990,N_13520);
nor U20966 (N_20966,N_15371,N_10036);
or U20967 (N_20967,N_14105,N_10147);
or U20968 (N_20968,N_14293,N_15966);
and U20969 (N_20969,N_16078,N_13843);
or U20970 (N_20970,N_18286,N_14141);
or U20971 (N_20971,N_11483,N_14441);
or U20972 (N_20972,N_17111,N_16391);
and U20973 (N_20973,N_17712,N_17504);
xor U20974 (N_20974,N_16633,N_10723);
nand U20975 (N_20975,N_14109,N_12009);
or U20976 (N_20976,N_17379,N_12561);
or U20977 (N_20977,N_18523,N_19722);
nand U20978 (N_20978,N_15206,N_12373);
nor U20979 (N_20979,N_13303,N_15185);
nor U20980 (N_20980,N_11522,N_15542);
or U20981 (N_20981,N_16467,N_13940);
nor U20982 (N_20982,N_11748,N_11949);
xnor U20983 (N_20983,N_13866,N_13060);
nor U20984 (N_20984,N_16208,N_17541);
xnor U20985 (N_20985,N_18114,N_19286);
or U20986 (N_20986,N_19246,N_10111);
or U20987 (N_20987,N_19207,N_17374);
xnor U20988 (N_20988,N_18957,N_14167);
nor U20989 (N_20989,N_15176,N_19750);
or U20990 (N_20990,N_10556,N_16129);
nor U20991 (N_20991,N_12145,N_10341);
nor U20992 (N_20992,N_14607,N_11608);
and U20993 (N_20993,N_12807,N_14945);
and U20994 (N_20994,N_13832,N_18956);
and U20995 (N_20995,N_18946,N_14086);
or U20996 (N_20996,N_14002,N_18450);
nand U20997 (N_20997,N_11371,N_18338);
nand U20998 (N_20998,N_14583,N_15272);
xnor U20999 (N_20999,N_18371,N_12623);
and U21000 (N_21000,N_17230,N_12019);
and U21001 (N_21001,N_11887,N_18544);
nor U21002 (N_21002,N_12514,N_10195);
nand U21003 (N_21003,N_12582,N_14043);
nand U21004 (N_21004,N_19277,N_17839);
or U21005 (N_21005,N_16831,N_16386);
nand U21006 (N_21006,N_12225,N_10858);
xor U21007 (N_21007,N_12071,N_14906);
nand U21008 (N_21008,N_16043,N_13161);
nor U21009 (N_21009,N_15824,N_10095);
nor U21010 (N_21010,N_13005,N_17196);
nor U21011 (N_21011,N_14878,N_13857);
nor U21012 (N_21012,N_13607,N_16838);
and U21013 (N_21013,N_14134,N_13293);
and U21014 (N_21014,N_17897,N_19285);
nand U21015 (N_21015,N_18530,N_16747);
and U21016 (N_21016,N_10103,N_11508);
xnor U21017 (N_21017,N_11959,N_17524);
nor U21018 (N_21018,N_15970,N_18808);
and U21019 (N_21019,N_11492,N_12732);
nor U21020 (N_21020,N_17303,N_12231);
and U21021 (N_21021,N_18436,N_14296);
nand U21022 (N_21022,N_18846,N_16990);
nand U21023 (N_21023,N_18077,N_18433);
xnor U21024 (N_21024,N_16548,N_17124);
nand U21025 (N_21025,N_19584,N_17147);
or U21026 (N_21026,N_12789,N_10592);
and U21027 (N_21027,N_14731,N_15600);
nand U21028 (N_21028,N_19842,N_19902);
nand U21029 (N_21029,N_10501,N_10616);
xnor U21030 (N_21030,N_10457,N_14193);
xor U21031 (N_21031,N_12478,N_13302);
nand U21032 (N_21032,N_16640,N_16119);
nand U21033 (N_21033,N_19035,N_19879);
xor U21034 (N_21034,N_16446,N_18399);
xnor U21035 (N_21035,N_16122,N_15878);
nand U21036 (N_21036,N_16084,N_15727);
nor U21037 (N_21037,N_17768,N_16636);
or U21038 (N_21038,N_12319,N_11668);
nand U21039 (N_21039,N_16441,N_10202);
xor U21040 (N_21040,N_17490,N_13840);
and U21041 (N_21041,N_10935,N_16116);
or U21042 (N_21042,N_13803,N_17599);
nor U21043 (N_21043,N_18185,N_19551);
xnor U21044 (N_21044,N_14183,N_12657);
nand U21045 (N_21045,N_10190,N_10314);
nand U21046 (N_21046,N_18331,N_17321);
xnor U21047 (N_21047,N_10348,N_19235);
and U21048 (N_21048,N_18395,N_11426);
nand U21049 (N_21049,N_14696,N_10100);
or U21050 (N_21050,N_18496,N_19625);
and U21051 (N_21051,N_17275,N_14030);
and U21052 (N_21052,N_19038,N_17935);
or U21053 (N_21053,N_14229,N_14060);
and U21054 (N_21054,N_17547,N_13630);
nor U21055 (N_21055,N_14021,N_13727);
nand U21056 (N_21056,N_17893,N_19684);
nand U21057 (N_21057,N_18938,N_12733);
xnor U21058 (N_21058,N_18193,N_14031);
and U21059 (N_21059,N_11208,N_16001);
nand U21060 (N_21060,N_16225,N_13409);
nor U21061 (N_21061,N_18905,N_12639);
nand U21062 (N_21062,N_19638,N_11245);
xnor U21063 (N_21063,N_13854,N_10138);
or U21064 (N_21064,N_18023,N_16298);
nor U21065 (N_21065,N_11701,N_19544);
xnor U21066 (N_21066,N_11233,N_16272);
or U21067 (N_21067,N_17266,N_12385);
xor U21068 (N_21068,N_16858,N_19401);
and U21069 (N_21069,N_12082,N_13283);
nor U21070 (N_21070,N_13352,N_14661);
nand U21071 (N_21071,N_14702,N_18604);
nor U21072 (N_21072,N_16283,N_16841);
nand U21073 (N_21073,N_10334,N_17500);
or U21074 (N_21074,N_10485,N_17885);
nor U21075 (N_21075,N_17670,N_11578);
or U21076 (N_21076,N_15453,N_15901);
and U21077 (N_21077,N_16376,N_15588);
nand U21078 (N_21078,N_13706,N_13874);
nand U21079 (N_21079,N_18982,N_13237);
nand U21080 (N_21080,N_10982,N_11303);
nor U21081 (N_21081,N_11947,N_14248);
xnor U21082 (N_21082,N_18637,N_18247);
nor U21083 (N_21083,N_19747,N_19745);
nand U21084 (N_21084,N_19326,N_15438);
nor U21085 (N_21085,N_11632,N_17226);
nand U21086 (N_21086,N_14102,N_12979);
nand U21087 (N_21087,N_19617,N_13787);
or U21088 (N_21088,N_14207,N_15867);
xor U21089 (N_21089,N_16644,N_10547);
or U21090 (N_21090,N_10431,N_11148);
and U21091 (N_21091,N_18359,N_12389);
or U21092 (N_21092,N_14439,N_17963);
nor U21093 (N_21093,N_11743,N_17792);
nor U21094 (N_21094,N_13534,N_12175);
nand U21095 (N_21095,N_12320,N_14474);
xor U21096 (N_21096,N_11406,N_11915);
nor U21097 (N_21097,N_13238,N_15363);
xnor U21098 (N_21098,N_16558,N_19050);
nand U21099 (N_21099,N_10497,N_14576);
and U21100 (N_21100,N_10291,N_14555);
xnor U21101 (N_21101,N_14013,N_11028);
nand U21102 (N_21102,N_19920,N_14796);
or U21103 (N_21103,N_15018,N_19831);
nor U21104 (N_21104,N_19446,N_17100);
nand U21105 (N_21105,N_13536,N_17549);
and U21106 (N_21106,N_14273,N_15252);
nand U21107 (N_21107,N_16786,N_14378);
or U21108 (N_21108,N_10104,N_18912);
or U21109 (N_21109,N_16491,N_14263);
and U21110 (N_21110,N_13260,N_14925);
and U21111 (N_21111,N_14635,N_12483);
or U21112 (N_21112,N_11484,N_12434);
xor U21113 (N_21113,N_15023,N_12470);
or U21114 (N_21114,N_11379,N_16247);
and U21115 (N_21115,N_17066,N_14884);
nand U21116 (N_21116,N_15843,N_13730);
nor U21117 (N_21117,N_18205,N_13870);
or U21118 (N_21118,N_18672,N_12922);
or U21119 (N_21119,N_12998,N_19877);
nor U21120 (N_21120,N_17295,N_11217);
or U21121 (N_21121,N_18495,N_16530);
xor U21122 (N_21122,N_16098,N_18055);
or U21123 (N_21123,N_17688,N_12641);
and U21124 (N_21124,N_17259,N_18355);
and U21125 (N_21125,N_11258,N_16259);
xnor U21126 (N_21126,N_16149,N_18219);
and U21127 (N_21127,N_13527,N_10098);
nand U21128 (N_21128,N_19338,N_11822);
xnor U21129 (N_21129,N_13983,N_14456);
and U21130 (N_21130,N_18297,N_14999);
and U21131 (N_21131,N_18878,N_16260);
xnor U21132 (N_21132,N_17853,N_17002);
nand U21133 (N_21133,N_12085,N_19152);
nand U21134 (N_21134,N_17136,N_17085);
or U21135 (N_21135,N_19574,N_16187);
or U21136 (N_21136,N_17322,N_11796);
and U21137 (N_21137,N_16911,N_11071);
and U21138 (N_21138,N_18953,N_19986);
nand U21139 (N_21139,N_12334,N_15762);
nand U21140 (N_21140,N_14718,N_11097);
and U21141 (N_21141,N_11797,N_16354);
nor U21142 (N_21142,N_10734,N_16511);
nor U21143 (N_21143,N_15751,N_14841);
nand U21144 (N_21144,N_18770,N_14954);
and U21145 (N_21145,N_11218,N_14454);
nor U21146 (N_21146,N_12144,N_10029);
or U21147 (N_21147,N_10980,N_18651);
nand U21148 (N_21148,N_19211,N_16366);
or U21149 (N_21149,N_19455,N_14174);
nand U21150 (N_21150,N_14004,N_11269);
nor U21151 (N_21151,N_17581,N_14076);
or U21152 (N_21152,N_10194,N_11186);
xor U21153 (N_21153,N_18272,N_13140);
xor U21154 (N_21154,N_11198,N_19226);
and U21155 (N_21155,N_16183,N_13673);
or U21156 (N_21156,N_18471,N_17932);
or U21157 (N_21157,N_14049,N_14901);
and U21158 (N_21158,N_12650,N_19693);
and U21159 (N_21159,N_17557,N_14648);
nor U21160 (N_21160,N_16889,N_10967);
nor U21161 (N_21161,N_10576,N_14655);
nand U21162 (N_21162,N_18558,N_15980);
and U21163 (N_21163,N_11723,N_18180);
nor U21164 (N_21164,N_16440,N_10562);
nor U21165 (N_21165,N_15435,N_12918);
nor U21166 (N_21166,N_11720,N_15589);
nor U21167 (N_21167,N_18388,N_19427);
or U21168 (N_21168,N_16848,N_10613);
and U21169 (N_21169,N_11070,N_17896);
xnor U21170 (N_21170,N_11419,N_13049);
nand U21171 (N_21171,N_17343,N_19829);
or U21172 (N_21172,N_14294,N_17137);
and U21173 (N_21173,N_14552,N_18807);
xor U21174 (N_21174,N_15113,N_10667);
nor U21175 (N_21175,N_13734,N_13271);
nand U21176 (N_21176,N_15973,N_19955);
and U21177 (N_21177,N_14537,N_15756);
nand U21178 (N_21178,N_17529,N_11194);
nand U21179 (N_21179,N_13907,N_19757);
or U21180 (N_21180,N_14603,N_13657);
and U21181 (N_21181,N_12620,N_16997);
or U21182 (N_21182,N_14265,N_16931);
or U21183 (N_21183,N_16117,N_15284);
and U21184 (N_21184,N_11963,N_19021);
and U21185 (N_21185,N_11144,N_18914);
xnor U21186 (N_21186,N_15425,N_12462);
nor U21187 (N_21187,N_12042,N_12409);
or U21188 (N_21188,N_16381,N_10807);
or U21189 (N_21189,N_18494,N_11677);
nor U21190 (N_21190,N_12228,N_12104);
nand U21191 (N_21191,N_17420,N_17140);
or U21192 (N_21192,N_13061,N_12942);
and U21193 (N_21193,N_12961,N_12522);
or U21194 (N_21194,N_12520,N_16408);
and U21195 (N_21195,N_17734,N_16177);
or U21196 (N_21196,N_10265,N_10659);
and U21197 (N_21197,N_14429,N_14683);
nand U21198 (N_21198,N_15395,N_19626);
or U21199 (N_21199,N_15172,N_10423);
or U21200 (N_21200,N_10797,N_17985);
and U21201 (N_21201,N_15601,N_10753);
nand U21202 (N_21202,N_18173,N_19360);
nor U21203 (N_21203,N_14280,N_14447);
or U21204 (N_21204,N_17907,N_14266);
nand U21205 (N_21205,N_19748,N_19358);
nor U21206 (N_21206,N_14403,N_15712);
or U21207 (N_21207,N_18977,N_11885);
nand U21208 (N_21208,N_16204,N_14510);
and U21209 (N_21209,N_10399,N_16487);
nor U21210 (N_21210,N_16037,N_18815);
nor U21211 (N_21211,N_13897,N_12914);
or U21212 (N_21212,N_16228,N_12921);
xor U21213 (N_21213,N_16595,N_17422);
nor U21214 (N_21214,N_18427,N_13679);
xnor U21215 (N_21215,N_16005,N_11781);
xor U21216 (N_21216,N_12972,N_14522);
or U21217 (N_21217,N_14970,N_19457);
or U21218 (N_21218,N_12965,N_18269);
nand U21219 (N_21219,N_13360,N_13812);
nor U21220 (N_21220,N_10583,N_10766);
or U21221 (N_21221,N_19913,N_18910);
xor U21222 (N_21222,N_14532,N_12766);
xor U21223 (N_21223,N_13588,N_14414);
or U21224 (N_21224,N_16822,N_10569);
or U21225 (N_21225,N_19340,N_11339);
nor U21226 (N_21226,N_10567,N_19972);
xor U21227 (N_21227,N_16065,N_10430);
xnor U21228 (N_21228,N_14240,N_12584);
and U21229 (N_21229,N_10516,N_11570);
nand U21230 (N_21230,N_18948,N_14287);
nor U21231 (N_21231,N_10778,N_10239);
nor U21232 (N_21232,N_19090,N_19208);
or U21233 (N_21233,N_15096,N_15687);
and U21234 (N_21234,N_14871,N_13615);
and U21235 (N_21235,N_16205,N_16019);
or U21236 (N_21236,N_12502,N_14038);
and U21237 (N_21237,N_19802,N_17922);
or U21238 (N_21238,N_15879,N_18773);
nand U21239 (N_21239,N_11512,N_17718);
or U21240 (N_21240,N_10992,N_13499);
nor U21241 (N_21241,N_11346,N_18009);
nand U21242 (N_21242,N_17992,N_11654);
nand U21243 (N_21243,N_18104,N_11857);
and U21244 (N_21244,N_12051,N_19417);
nor U21245 (N_21245,N_15432,N_11810);
xnor U21246 (N_21246,N_19560,N_14922);
and U21247 (N_21247,N_12342,N_14598);
or U21248 (N_21248,N_16638,N_10596);
and U21249 (N_21249,N_10386,N_10988);
xnor U21250 (N_21250,N_17699,N_19562);
nand U21251 (N_21251,N_11092,N_17909);
and U21252 (N_21252,N_14840,N_14392);
and U21253 (N_21253,N_11176,N_13357);
nor U21254 (N_21254,N_15674,N_18006);
nor U21255 (N_21255,N_12252,N_15079);
nand U21256 (N_21256,N_15140,N_16505);
and U21257 (N_21257,N_11532,N_16600);
or U21258 (N_21258,N_15115,N_18787);
xor U21259 (N_21259,N_13855,N_19397);
or U21260 (N_21260,N_18707,N_16344);
and U21261 (N_21261,N_12146,N_17345);
or U21262 (N_21262,N_18379,N_18951);
and U21263 (N_21263,N_15063,N_19973);
and U21264 (N_21264,N_10899,N_15659);
xor U21265 (N_21265,N_13126,N_15559);
nor U21266 (N_21266,N_16184,N_14570);
and U21267 (N_21267,N_10022,N_16070);
and U21268 (N_21268,N_11702,N_19511);
nor U21269 (N_21269,N_14460,N_10310);
or U21270 (N_21270,N_16951,N_12364);
or U21271 (N_21271,N_12869,N_12862);
nor U21272 (N_21272,N_19267,N_10483);
and U21273 (N_21273,N_18402,N_12005);
nor U21274 (N_21274,N_14045,N_18143);
nand U21275 (N_21275,N_19124,N_12209);
or U21276 (N_21276,N_12467,N_17416);
nor U21277 (N_21277,N_10541,N_13568);
nor U21278 (N_21278,N_12100,N_19527);
nor U21279 (N_21279,N_12636,N_14624);
and U21280 (N_21280,N_10677,N_14895);
xor U21281 (N_21281,N_14919,N_14492);
and U21282 (N_21282,N_13988,N_12133);
and U21283 (N_21283,N_16328,N_15338);
nand U21284 (N_21284,N_13102,N_15811);
nand U21285 (N_21285,N_19583,N_15479);
nand U21286 (N_21286,N_17182,N_13757);
and U21287 (N_21287,N_10574,N_15205);
nor U21288 (N_21288,N_11061,N_17035);
nand U21289 (N_21289,N_10137,N_17155);
nor U21290 (N_21290,N_10534,N_15125);
nand U21291 (N_21291,N_17369,N_12575);
or U21292 (N_21292,N_18130,N_16569);
and U21293 (N_21293,N_18593,N_18656);
nor U21294 (N_21294,N_11540,N_11556);
nand U21295 (N_21295,N_16125,N_10462);
nand U21296 (N_21296,N_16383,N_18851);
nor U21297 (N_21297,N_19399,N_12435);
and U21298 (N_21298,N_12288,N_16755);
or U21299 (N_21299,N_15457,N_14927);
nor U21300 (N_21300,N_15775,N_12608);
and U21301 (N_21301,N_12384,N_10670);
or U21302 (N_21302,N_16879,N_10818);
or U21303 (N_21303,N_17959,N_11416);
or U21304 (N_21304,N_10564,N_16419);
and U21305 (N_21305,N_16290,N_14679);
nand U21306 (N_21306,N_18086,N_17033);
or U21307 (N_21307,N_10455,N_11513);
xor U21308 (N_21308,N_18430,N_11313);
and U21309 (N_21309,N_14164,N_13264);
nand U21310 (N_21310,N_11581,N_19775);
and U21311 (N_21311,N_12236,N_10288);
nand U21312 (N_21312,N_19529,N_17707);
and U21313 (N_21313,N_11023,N_13246);
or U21314 (N_21314,N_14268,N_10027);
xnor U21315 (N_21315,N_11064,N_11673);
nand U21316 (N_21316,N_16164,N_10471);
and U21317 (N_21317,N_15993,N_16662);
and U21318 (N_21318,N_17229,N_11383);
and U21319 (N_21319,N_10752,N_16995);
nor U21320 (N_21320,N_14693,N_11656);
or U21321 (N_21321,N_11357,N_11974);
nor U21322 (N_21322,N_11029,N_15035);
nor U21323 (N_21323,N_12180,N_10135);
nor U21324 (N_21324,N_17445,N_18947);
nand U21325 (N_21325,N_18001,N_16254);
and U21326 (N_21326,N_14272,N_13814);
and U21327 (N_21327,N_19561,N_12535);
xnor U21328 (N_21328,N_16169,N_10263);
and U21329 (N_21329,N_12557,N_16570);
nor U21330 (N_21330,N_19498,N_14627);
and U21331 (N_21331,N_11638,N_13686);
nor U21332 (N_21332,N_15930,N_11784);
nor U21333 (N_21333,N_15517,N_15513);
nand U21334 (N_21334,N_12983,N_17944);
or U21335 (N_21335,N_12401,N_10703);
or U21336 (N_21336,N_18788,N_12905);
nor U21337 (N_21337,N_10016,N_16418);
and U21338 (N_21338,N_16281,N_15910);
or U21339 (N_21339,N_19903,N_18708);
or U21340 (N_21340,N_10697,N_13502);
nor U21341 (N_21341,N_14376,N_13328);
nand U21342 (N_21342,N_19173,N_13969);
nor U21343 (N_21343,N_18479,N_10927);
and U21344 (N_21344,N_17495,N_11523);
and U21345 (N_21345,N_12368,N_12545);
nand U21346 (N_21346,N_16214,N_14039);
or U21347 (N_21347,N_19012,N_13322);
nor U21348 (N_21348,N_18230,N_16085);
nand U21349 (N_21349,N_10144,N_13199);
or U21350 (N_21350,N_13839,N_13003);
and U21351 (N_21351,N_19785,N_15217);
nor U21352 (N_21352,N_17654,N_13806);
and U21353 (N_21353,N_14205,N_10278);
nor U21354 (N_21354,N_12021,N_16332);
or U21355 (N_21355,N_14843,N_10780);
nand U21356 (N_21356,N_11083,N_12916);
nor U21357 (N_21357,N_11764,N_16277);
and U21358 (N_21358,N_15752,N_13728);
or U21359 (N_21359,N_18398,N_15904);
nand U21360 (N_21360,N_19145,N_14066);
nand U21361 (N_21361,N_16292,N_16430);
or U21362 (N_21362,N_12129,N_10743);
nor U21363 (N_21363,N_18870,N_16642);
or U21364 (N_21364,N_14315,N_10445);
nand U21365 (N_21365,N_11630,N_11210);
nor U21366 (N_21366,N_17327,N_17533);
nand U21367 (N_21367,N_12826,N_17809);
nor U21368 (N_21368,N_13103,N_13086);
and U21369 (N_21369,N_19051,N_15765);
or U21370 (N_21370,N_14397,N_14544);
or U21371 (N_21371,N_18907,N_13779);
and U21372 (N_21372,N_15982,N_11820);
nand U21373 (N_21373,N_15621,N_19818);
xor U21374 (N_21374,N_16359,N_10094);
nor U21375 (N_21375,N_17544,N_15384);
nand U21376 (N_21376,N_17286,N_19323);
or U21377 (N_21377,N_16319,N_13511);
or U21378 (N_21378,N_16894,N_16768);
or U21379 (N_21379,N_15539,N_11627);
nand U21380 (N_21380,N_11875,N_19863);
nor U21381 (N_21381,N_14814,N_11051);
nor U21382 (N_21382,N_11765,N_18437);
xor U21383 (N_21383,N_11542,N_10782);
or U21384 (N_21384,N_11149,N_11480);
or U21385 (N_21385,N_13883,N_14835);
xnor U21386 (N_21386,N_10175,N_10088);
or U21387 (N_21387,N_16760,N_18848);
nor U21388 (N_21388,N_17190,N_11852);
and U21389 (N_21389,N_12632,N_18974);
and U21390 (N_21390,N_19044,N_16167);
and U21391 (N_21391,N_16798,N_11355);
and U21392 (N_21392,N_17769,N_16966);
and U21393 (N_21393,N_14993,N_13022);
or U21394 (N_21394,N_16625,N_13807);
or U21395 (N_21395,N_19388,N_15141);
nor U21396 (N_21396,N_17660,N_14295);
nand U21397 (N_21397,N_11511,N_19166);
nand U21398 (N_21398,N_12213,N_12006);
and U21399 (N_21399,N_17823,N_19708);
nor U21400 (N_21400,N_12458,N_12453);
xnor U21401 (N_21401,N_11052,N_11979);
nand U21402 (N_21402,N_17121,N_13435);
or U21403 (N_21403,N_19187,N_10394);
nand U21404 (N_21404,N_11085,N_11498);
and U21405 (N_21405,N_15146,N_10206);
or U21406 (N_21406,N_16834,N_11580);
or U21407 (N_21407,N_19205,N_13986);
nand U21408 (N_21408,N_12173,N_19957);
or U21409 (N_21409,N_19657,N_19096);
or U21410 (N_21410,N_14587,N_12996);
nand U21411 (N_21411,N_15445,N_10177);
or U21412 (N_21412,N_11094,N_13901);
or U21413 (N_21413,N_14239,N_10601);
nor U21414 (N_21414,N_14881,N_11691);
or U21415 (N_21415,N_11759,N_15194);
and U21416 (N_21416,N_17005,N_16748);
nand U21417 (N_21417,N_12123,N_10127);
and U21418 (N_21418,N_11728,N_12107);
or U21419 (N_21419,N_16020,N_18213);
or U21420 (N_21420,N_14222,N_10318);
and U21421 (N_21421,N_12105,N_12227);
nor U21422 (N_21422,N_16488,N_12079);
xnor U21423 (N_21423,N_16955,N_18800);
nor U21424 (N_21424,N_14815,N_18801);
and U21425 (N_21425,N_15826,N_15058);
nand U21426 (N_21426,N_19662,N_19932);
nor U21427 (N_21427,N_19282,N_10237);
xnor U21428 (N_21428,N_16784,N_18170);
or U21429 (N_21429,N_15414,N_11992);
nand U21430 (N_21430,N_16294,N_17808);
and U21431 (N_21431,N_16697,N_16025);
nand U21432 (N_21432,N_13624,N_15130);
nor U21433 (N_21433,N_12102,N_16977);
nand U21434 (N_21434,N_19481,N_13620);
and U21435 (N_21435,N_12518,N_14978);
nor U21436 (N_21436,N_13794,N_15337);
or U21437 (N_21437,N_13010,N_17062);
and U21438 (N_21438,N_18658,N_11192);
nor U21439 (N_21439,N_18749,N_13011);
or U21440 (N_21440,N_15123,N_16991);
and U21441 (N_21441,N_16793,N_19857);
nor U21442 (N_21442,N_15570,N_10892);
and U21443 (N_21443,N_15540,N_16159);
or U21444 (N_21444,N_14398,N_13867);
or U21445 (N_21445,N_19823,N_10694);
and U21446 (N_21446,N_12397,N_11054);
nand U21447 (N_21447,N_14865,N_16507);
nor U21448 (N_21448,N_12940,N_13092);
nand U21449 (N_21449,N_10154,N_18199);
and U21450 (N_21450,N_16560,N_16323);
xnor U21451 (N_21451,N_19088,N_10724);
nand U21452 (N_21452,N_12758,N_19312);
nand U21453 (N_21453,N_12880,N_16980);
and U21454 (N_21454,N_10806,N_17215);
and U21455 (N_21455,N_19968,N_13207);
and U21456 (N_21456,N_19744,N_10343);
nand U21457 (N_21457,N_15036,N_17122);
nand U21458 (N_21458,N_14929,N_16146);
xnor U21459 (N_21459,N_11876,N_13343);
nor U21460 (N_21460,N_19792,N_19001);
and U21461 (N_21461,N_16763,N_11793);
and U21462 (N_21462,N_17000,N_19441);
and U21463 (N_21463,N_10322,N_12066);
nor U21464 (N_21464,N_12781,N_15810);
or U21465 (N_21465,N_11259,N_19890);
nand U21466 (N_21466,N_14698,N_12312);
and U21467 (N_21467,N_13629,N_17272);
or U21468 (N_21468,N_17580,N_12293);
xnor U21469 (N_21469,N_17991,N_11665);
nand U21470 (N_21470,N_19484,N_14238);
or U21471 (N_21471,N_17043,N_10589);
nand U21472 (N_21472,N_16631,N_15568);
or U21473 (N_21473,N_10538,N_17203);
or U21474 (N_21474,N_11824,N_13893);
and U21475 (N_21475,N_11932,N_12970);
nor U21476 (N_21476,N_13716,N_16308);
nor U21477 (N_21477,N_15655,N_12547);
nand U21478 (N_21478,N_10109,N_14909);
or U21479 (N_21479,N_10939,N_19390);
nor U21480 (N_21480,N_12550,N_10711);
or U21481 (N_21481,N_11078,N_14097);
xnor U21482 (N_21482,N_16309,N_16937);
nor U21483 (N_21483,N_13518,N_16021);
nand U21484 (N_21484,N_10159,N_11813);
or U21485 (N_21485,N_17191,N_11689);
nor U21486 (N_21486,N_16924,N_11860);
xor U21487 (N_21487,N_11955,N_11087);
and U21488 (N_21488,N_14738,N_11199);
or U21489 (N_21489,N_14244,N_15642);
nor U21490 (N_21490,N_12383,N_17089);
and U21491 (N_21491,N_16908,N_14562);
and U21492 (N_21492,N_15729,N_17091);
xnor U21493 (N_21493,N_16352,N_13535);
nand U21494 (N_21494,N_12993,N_17497);
and U21495 (N_21495,N_13374,N_10514);
xor U21496 (N_21496,N_14177,N_14625);
and U21497 (N_21497,N_17017,N_15784);
and U21498 (N_21498,N_15382,N_19204);
and U21499 (N_21499,N_12000,N_15179);
xor U21500 (N_21500,N_12070,N_12893);
xnor U21501 (N_21501,N_11905,N_11072);
xor U21502 (N_21502,N_13146,N_18174);
xnor U21503 (N_21503,N_13099,N_11179);
and U21504 (N_21504,N_13219,N_11539);
or U21505 (N_21505,N_15114,N_12078);
or U21506 (N_21506,N_15548,N_15947);
nand U21507 (N_21507,N_18861,N_15555);
and U21508 (N_21508,N_16539,N_11601);
nor U21509 (N_21509,N_11169,N_19806);
nand U21510 (N_21510,N_16688,N_18349);
nor U21511 (N_21511,N_14830,N_13028);
or U21512 (N_21512,N_15937,N_13300);
nor U21513 (N_21513,N_16796,N_12666);
nor U21514 (N_21514,N_15412,N_13138);
and U21515 (N_21515,N_17110,N_18510);
and U21516 (N_21516,N_15722,N_15672);
nor U21517 (N_21517,N_17185,N_15868);
nor U21518 (N_21518,N_18775,N_16958);
nand U21519 (N_21519,N_15833,N_17176);
nor U21520 (N_21520,N_14495,N_15052);
nand U21521 (N_21521,N_15015,N_13613);
xnor U21522 (N_21522,N_16544,N_11653);
and U21523 (N_21523,N_15597,N_10812);
xnor U21524 (N_21524,N_14072,N_10007);
nor U21525 (N_21525,N_17818,N_17904);
nand U21526 (N_21526,N_11146,N_17329);
nor U21527 (N_21527,N_11843,N_15858);
nor U21528 (N_21528,N_17925,N_16449);
nand U21529 (N_21529,N_12764,N_14934);
nand U21530 (N_21530,N_14204,N_15265);
nand U21531 (N_21531,N_17181,N_10174);
nor U21532 (N_21532,N_19777,N_17872);
or U21533 (N_21533,N_18715,N_13262);
nor U21534 (N_21534,N_16405,N_18514);
nor U21535 (N_21535,N_17727,N_15200);
or U21536 (N_21536,N_19803,N_11832);
nand U21537 (N_21537,N_17917,N_16671);
nand U21538 (N_21538,N_14984,N_16353);
nor U21539 (N_21539,N_15367,N_13563);
or U21540 (N_21540,N_14443,N_14075);
and U21541 (N_21541,N_11934,N_10000);
nor U21542 (N_21542,N_13496,N_12261);
and U21543 (N_21543,N_17596,N_16394);
nand U21544 (N_21544,N_11953,N_10466);
nand U21545 (N_21545,N_14247,N_15573);
or U21546 (N_21546,N_10142,N_13042);
or U21547 (N_21547,N_13886,N_13039);
nor U21548 (N_21548,N_13190,N_14971);
or U21549 (N_21549,N_10395,N_11164);
or U21550 (N_21550,N_11001,N_12586);
and U21551 (N_21551,N_19466,N_13423);
nor U21552 (N_21552,N_15537,N_11348);
nor U21553 (N_21553,N_17771,N_13490);
or U21554 (N_21554,N_18911,N_17962);
and U21555 (N_21555,N_18830,N_19174);
nand U21556 (N_21556,N_15444,N_18443);
nor U21557 (N_21557,N_13602,N_13567);
and U21558 (N_21558,N_15313,N_16180);
xor U21559 (N_21559,N_16076,N_10304);
and U21560 (N_21560,N_18151,N_14150);
nor U21561 (N_21561,N_13084,N_14942);
nor U21562 (N_21562,N_10859,N_10910);
xor U21563 (N_21563,N_18756,N_14754);
nor U21564 (N_21564,N_10415,N_10626);
nand U21565 (N_21565,N_14155,N_15461);
and U21566 (N_21566,N_15721,N_17179);
and U21567 (N_21567,N_13586,N_17078);
nor U21568 (N_21568,N_18931,N_14572);
nor U21569 (N_21569,N_15354,N_13063);
and U21570 (N_21570,N_11154,N_10297);
nor U21571 (N_21571,N_15070,N_12219);
nand U21572 (N_21572,N_18158,N_14334);
and U21573 (N_21573,N_13149,N_12492);
or U21574 (N_21574,N_19680,N_10120);
nor U21575 (N_21575,N_12785,N_18606);
xnor U21576 (N_21576,N_18275,N_11026);
xor U21577 (N_21577,N_13197,N_13830);
or U21578 (N_21578,N_11002,N_15567);
or U21579 (N_21579,N_16197,N_19066);
nor U21580 (N_21580,N_13315,N_15635);
and U21581 (N_21581,N_10643,N_19714);
or U21582 (N_21582,N_19103,N_19683);
nor U21583 (N_21583,N_15677,N_13889);
nand U21584 (N_21584,N_12929,N_14845);
or U21585 (N_21585,N_14235,N_10727);
or U21586 (N_21586,N_15330,N_14640);
xor U21587 (N_21587,N_12015,N_10591);
nand U21588 (N_21588,N_11716,N_11687);
and U21589 (N_21589,N_12304,N_12634);
nor U21590 (N_21590,N_12212,N_11135);
or U21591 (N_21591,N_13243,N_18327);
or U21592 (N_21592,N_11562,N_15907);
or U21593 (N_21593,N_16969,N_11895);
nand U21594 (N_21594,N_16274,N_12702);
nand U21595 (N_21595,N_15420,N_17746);
nand U21596 (N_21596,N_13181,N_17520);
xnor U21597 (N_21597,N_18195,N_14849);
nor U21598 (N_21598,N_18611,N_19071);
nor U21599 (N_21599,N_16939,N_18970);
or U21600 (N_21600,N_19213,N_10799);
xor U21601 (N_21601,N_14890,N_11282);
nand U21602 (N_21602,N_13906,N_12235);
nand U21603 (N_21603,N_16250,N_16712);
or U21604 (N_21604,N_19087,N_17762);
or U21605 (N_21605,N_16303,N_15229);
or U21606 (N_21606,N_17759,N_15977);
or U21607 (N_21607,N_14564,N_11079);
or U21608 (N_21608,N_11411,N_15974);
and U21609 (N_21609,N_19380,N_18925);
or U21610 (N_21610,N_16618,N_14959);
xnor U21611 (N_21611,N_13405,N_14991);
or U21612 (N_21612,N_15802,N_13976);
or U21613 (N_21613,N_14520,N_14539);
or U21614 (N_21614,N_19605,N_18455);
or U21615 (N_21615,N_17602,N_15897);
nor U21616 (N_21616,N_18098,N_17631);
and U21617 (N_21617,N_14608,N_14616);
and U21618 (N_21618,N_18704,N_16567);
and U21619 (N_21619,N_11472,N_11641);
nand U21620 (N_21620,N_17940,N_14654);
nor U21621 (N_21621,N_13449,N_14921);
nor U21622 (N_21622,N_17250,N_13231);
nand U21623 (N_21623,N_18463,N_18018);
or U21624 (N_21624,N_15933,N_14203);
nor U21625 (N_21625,N_12239,N_17979);
nor U21626 (N_21626,N_18967,N_17983);
nand U21627 (N_21627,N_14048,N_12035);
nand U21628 (N_21628,N_13318,N_12565);
or U21629 (N_21629,N_16964,N_17019);
and U21630 (N_21630,N_17010,N_15527);
or U21631 (N_21631,N_16862,N_19476);
or U21632 (N_21632,N_14285,N_11326);
or U21633 (N_21633,N_17532,N_18838);
and U21634 (N_21634,N_14829,N_11435);
nand U21635 (N_21635,N_12354,N_17919);
and U21636 (N_21636,N_18822,N_18109);
nand U21637 (N_21637,N_15451,N_16270);
and U21638 (N_21638,N_15192,N_14846);
nand U21639 (N_21639,N_16994,N_14224);
nand U21640 (N_21640,N_16635,N_10745);
nand U21641 (N_21641,N_11044,N_11273);
nand U21642 (N_21642,N_11831,N_10122);
nor U21643 (N_21643,N_16934,N_16704);
or U21644 (N_21644,N_14712,N_14778);
nand U21645 (N_21645,N_10298,N_16817);
nand U21646 (N_21646,N_10920,N_17357);
nand U21647 (N_21647,N_17642,N_14253);
and U21648 (N_21648,N_10052,N_17130);
and U21649 (N_21649,N_18421,N_10978);
nand U21650 (N_21650,N_16045,N_17125);
or U21651 (N_21651,N_10666,N_11528);
or U21652 (N_21652,N_11724,N_19249);
or U21653 (N_21653,N_19353,N_19278);
and U21654 (N_21654,N_18241,N_17200);
nor U21655 (N_21655,N_14623,N_11440);
nor U21656 (N_21656,N_16246,N_13777);
xor U21657 (N_21657,N_11946,N_19265);
or U21658 (N_21658,N_16616,N_16902);
nand U21659 (N_21659,N_16103,N_16375);
nor U21660 (N_21660,N_10577,N_13929);
nor U21661 (N_21661,N_13023,N_15434);
nand U21662 (N_21662,N_19938,N_10744);
nor U21663 (N_21663,N_19502,N_19492);
nor U21664 (N_21664,N_17396,N_12245);
xor U21665 (N_21665,N_12031,N_11552);
and U21666 (N_21666,N_17910,N_17957);
nor U21667 (N_21667,N_11977,N_14320);
nor U21668 (N_21668,N_10509,N_12775);
nor U21669 (N_21669,N_15386,N_12154);
nor U21670 (N_21670,N_18461,N_11605);
nand U21671 (N_21671,N_12457,N_11158);
nor U21672 (N_21672,N_17842,N_19999);
xnor U21673 (N_21673,N_17501,N_14377);
nor U21674 (N_21674,N_12717,N_14515);
nor U21675 (N_21675,N_17673,N_15385);
xnor U21676 (N_21676,N_19753,N_19164);
or U21677 (N_21677,N_14634,N_11968);
or U21678 (N_21678,N_18457,N_10040);
nor U21679 (N_21679,N_18072,N_19589);
nand U21680 (N_21680,N_13397,N_11166);
and U21681 (N_21681,N_18472,N_19995);
or U21682 (N_21682,N_15048,N_18226);
nor U21683 (N_21683,N_14464,N_13733);
nor U21684 (N_21684,N_11985,N_10301);
and U21685 (N_21685,N_10623,N_14875);
nor U21686 (N_21686,N_11423,N_11521);
and U21687 (N_21687,N_12276,N_16395);
and U21688 (N_21688,N_17131,N_12697);
nor U21689 (N_21689,N_17811,N_11490);
or U21690 (N_21690,N_11320,N_11168);
and U21691 (N_21691,N_17609,N_18235);
nand U21692 (N_21692,N_12617,N_13784);
or U21693 (N_21693,N_15714,N_17480);
or U21694 (N_21694,N_12594,N_13521);
nor U21695 (N_21695,N_12210,N_12856);
or U21696 (N_21696,N_14408,N_18780);
nor U21697 (N_21697,N_18325,N_17253);
xnor U21698 (N_21698,N_12166,N_14187);
or U21699 (N_21699,N_19382,N_17060);
xor U21700 (N_21700,N_13815,N_19179);
nor U21701 (N_21701,N_15495,N_14368);
nor U21702 (N_21702,N_18083,N_16421);
nand U21703 (N_21703,N_10459,N_17972);
nand U21704 (N_21704,N_15120,N_14675);
and U21705 (N_21705,N_11846,N_15139);
and U21706 (N_21706,N_16555,N_19817);
or U21707 (N_21707,N_14241,N_14216);
nand U21708 (N_21708,N_11361,N_18999);
or U21709 (N_21709,N_16998,N_17384);
nand U21710 (N_21710,N_13707,N_16185);
or U21711 (N_21711,N_10740,N_13166);
and U21712 (N_21712,N_16639,N_11600);
nor U21713 (N_21713,N_12777,N_11643);
nor U21714 (N_21714,N_17623,N_18282);
or U21715 (N_21715,N_16741,N_18129);
or U21716 (N_21716,N_10411,N_13097);
and U21717 (N_21717,N_17735,N_14973);
and U21718 (N_21718,N_11049,N_15697);
or U21719 (N_21719,N_12779,N_12196);
and U21720 (N_21720,N_11125,N_19590);
xor U21721 (N_21721,N_17659,N_13537);
xor U21722 (N_21722,N_19293,N_14990);
and U21723 (N_21723,N_10931,N_18519);
nand U21724 (N_21724,N_13663,N_12910);
and U21725 (N_21725,N_12439,N_18646);
nand U21726 (N_21726,N_10372,N_14143);
nor U21727 (N_21727,N_12329,N_11815);
nor U21728 (N_21728,N_17794,N_14250);
nand U21729 (N_21729,N_10991,N_12471);
nand U21730 (N_21730,N_11205,N_17606);
or U21731 (N_21731,N_18809,N_10317);
or U21732 (N_21732,N_14824,N_12028);
nand U21733 (N_21733,N_15912,N_16128);
nand U21734 (N_21734,N_14058,N_15157);
nor U21735 (N_21735,N_10638,N_16708);
nor U21736 (N_21736,N_18420,N_18137);
and U21737 (N_21737,N_10795,N_14641);
nor U21738 (N_21738,N_17667,N_14116);
nor U21739 (N_21739,N_15042,N_17015);
nand U21740 (N_21740,N_10008,N_17293);
nor U21741 (N_21741,N_14327,N_16163);
nor U21742 (N_21742,N_16337,N_17279);
nand U21743 (N_21743,N_16717,N_12086);
and U21744 (N_21744,N_10082,N_10841);
nor U21745 (N_21745,N_14117,N_11414);
and U21746 (N_21746,N_19192,N_18314);
and U21747 (N_21747,N_17918,N_16844);
or U21748 (N_21748,N_15647,N_15669);
nand U21749 (N_21749,N_13163,N_14119);
nor U21750 (N_21750,N_12726,N_10728);
nor U21751 (N_21751,N_15090,N_17790);
and U21752 (N_21752,N_11667,N_13998);
or U21753 (N_21753,N_15803,N_14331);
nand U21754 (N_21754,N_11441,N_13054);
and U21755 (N_21755,N_12587,N_17982);
and U21756 (N_21756,N_19548,N_13349);
or U21757 (N_21757,N_18923,N_13337);
and U21758 (N_21758,N_10087,N_11623);
nand U21759 (N_21759,N_15059,N_19582);
and U21760 (N_21760,N_15637,N_14481);
nand U21761 (N_21761,N_19610,N_15535);
nand U21762 (N_21762,N_11337,N_19333);
and U21763 (N_21763,N_10361,N_16320);
nand U21764 (N_21764,N_19977,N_11572);
nor U21765 (N_21765,N_19404,N_10233);
nor U21766 (N_21766,N_19315,N_18718);
nor U21767 (N_21767,N_15196,N_19958);
nand U21768 (N_21768,N_12528,N_13211);
nand U21769 (N_21769,N_16013,N_12244);
nor U21770 (N_21770,N_12654,N_13325);
nand U21771 (N_21771,N_19577,N_19710);
nor U21772 (N_21772,N_11721,N_10702);
and U21773 (N_21773,N_14308,N_10362);
nor U21774 (N_21774,N_17115,N_10872);
and U21775 (N_21775,N_16730,N_16651);
nand U21776 (N_21776,N_14463,N_18163);
and U21777 (N_21777,N_19060,N_10118);
xor U21778 (N_21778,N_14274,N_16244);
nor U21779 (N_21779,N_10463,N_11730);
nor U21780 (N_21780,N_17961,N_18204);
and U21781 (N_21781,N_17540,N_13696);
and U21782 (N_21782,N_16921,N_14703);
or U21783 (N_21783,N_16289,N_19524);
nor U21784 (N_21784,N_13674,N_13858);
and U21785 (N_21785,N_15131,N_10597);
nor U21786 (N_21786,N_10360,N_17878);
or U21787 (N_21787,N_10266,N_11153);
and U21788 (N_21788,N_15129,N_19758);
and U21789 (N_21789,N_14753,N_13228);
nor U21790 (N_21790,N_19141,N_18058);
or U21791 (N_21791,N_11670,N_16226);
nand U21792 (N_21792,N_19947,N_16893);
nor U21793 (N_21793,N_14027,N_12300);
or U21794 (N_21794,N_18755,N_18949);
and U21795 (N_21795,N_11069,N_11325);
and U21796 (N_21796,N_14299,N_17620);
and U21797 (N_21797,N_12992,N_15001);
nor U21798 (N_21798,N_11510,N_16847);
or U21799 (N_21799,N_19268,N_13425);
xnor U21800 (N_21800,N_15818,N_12119);
or U21801 (N_21801,N_18074,N_16296);
and U21802 (N_21802,N_10527,N_10256);
xor U21803 (N_21803,N_16547,N_19229);
nor U21804 (N_21804,N_15876,N_15839);
and U21805 (N_21805,N_10262,N_13923);
or U21806 (N_21806,N_14726,N_18192);
nand U21807 (N_21807,N_16049,N_19266);
nand U21808 (N_21808,N_13171,N_11331);
xor U21809 (N_21809,N_13817,N_14485);
nand U21810 (N_21810,N_12630,N_17567);
nor U21811 (N_21811,N_11790,N_11368);
and U21812 (N_21812,N_15519,N_17600);
or U21813 (N_21813,N_16023,N_15267);
or U21814 (N_21814,N_15515,N_13935);
and U21815 (N_21815,N_16079,N_15485);
nor U21816 (N_21816,N_14952,N_18828);
nor U21817 (N_21817,N_13275,N_10030);
nand U21818 (N_21818,N_19718,N_18573);
or U21819 (N_21819,N_17709,N_15516);
nand U21820 (N_21820,N_17774,N_19824);
and U21821 (N_21821,N_10517,N_15564);
nor U21822 (N_21822,N_18538,N_16617);
or U21823 (N_21823,N_18660,N_19359);
nand U21824 (N_21824,N_15055,N_14762);
nand U21825 (N_21825,N_16135,N_11566);
and U21826 (N_21826,N_15880,N_18031);
nand U21827 (N_21827,N_15711,N_16677);
nand U21828 (N_21828,N_15352,N_11173);
and U21829 (N_21829,N_16802,N_16588);
nor U21830 (N_21830,N_11970,N_10836);
and U21831 (N_21831,N_14000,N_12377);
nand U21832 (N_21832,N_11777,N_18268);
and U21833 (N_21833,N_10328,N_15221);
or U21834 (N_21834,N_13229,N_14926);
and U21835 (N_21835,N_17798,N_19271);
nor U21836 (N_21836,N_16621,N_11514);
nand U21837 (N_21837,N_18211,N_19176);
and U21838 (N_21838,N_16956,N_14209);
xnor U21839 (N_21839,N_13338,N_14015);
or U21840 (N_21840,N_19431,N_15116);
nor U21841 (N_21841,N_15460,N_11242);
xor U21842 (N_21842,N_15245,N_13385);
xor U21843 (N_21843,N_16988,N_19788);
nand U21844 (N_21844,N_13421,N_18209);
or U21845 (N_21845,N_19011,N_13025);
or U21846 (N_21846,N_10258,N_11886);
nor U21847 (N_21847,N_11384,N_14803);
nor U21848 (N_21848,N_15419,N_14477);
or U21849 (N_21849,N_16190,N_19646);
nor U21850 (N_21850,N_14864,N_17868);
or U21851 (N_21851,N_18322,N_14823);
or U21852 (N_21852,N_14629,N_19033);
nor U21853 (N_21853,N_18426,N_13065);
nand U21854 (N_21854,N_14288,N_10379);
nor U21855 (N_21855,N_19126,N_16275);
nand U21856 (N_21856,N_15678,N_14799);
or U21857 (N_21857,N_13486,N_12969);
or U21858 (N_21858,N_10234,N_13129);
nand U21859 (N_21859,N_16849,N_10632);
or U21860 (N_21860,N_11585,N_11525);
and U21861 (N_21861,N_17183,N_12980);
nor U21862 (N_21862,N_19941,N_11101);
nand U21863 (N_21863,N_11883,N_10001);
nand U21864 (N_21864,N_11499,N_14430);
nor U21865 (N_21865,N_14140,N_12548);
xor U21866 (N_21866,N_11088,N_10897);
and U21867 (N_21867,N_13292,N_18719);
nor U21868 (N_21868,N_18354,N_12569);
and U21869 (N_21869,N_11226,N_18111);
or U21870 (N_21870,N_18779,N_12529);
or U21871 (N_21871,N_10942,N_13691);
and U21872 (N_21872,N_16918,N_15184);
and U21873 (N_21873,N_17058,N_12301);
nor U21874 (N_21874,N_18644,N_13434);
nor U21875 (N_21875,N_18734,N_17126);
nor U21876 (N_21876,N_17404,N_10277);
or U21877 (N_21877,N_11446,N_19125);
nor U21878 (N_21878,N_16219,N_16957);
nand U21879 (N_21879,N_13996,N_11151);
xnor U21880 (N_21880,N_18061,N_11209);
nand U21881 (N_21881,N_17308,N_10510);
and U21882 (N_21882,N_16141,N_12290);
nor U21883 (N_21883,N_19746,N_17595);
nand U21884 (N_21884,N_11006,N_18155);
xor U21885 (N_21885,N_16485,N_13987);
xor U21886 (N_21886,N_12674,N_15073);
nor U21887 (N_21887,N_13577,N_11354);
nor U21888 (N_21888,N_16815,N_11972);
nor U21889 (N_21889,N_15173,N_11161);
nand U21890 (N_21890,N_13150,N_11369);
nor U21891 (N_21891,N_18569,N_15944);
nand U21892 (N_21892,N_15923,N_11500);
nor U21893 (N_21893,N_10049,N_10622);
and U21894 (N_21894,N_12437,N_12647);
or U21895 (N_21895,N_18449,N_11997);
xor U21896 (N_21896,N_16267,N_16378);
or U21897 (N_21897,N_12081,N_15608);
or U21898 (N_21898,N_12669,N_14538);
nand U21899 (N_21899,N_11850,N_15768);
and U21900 (N_21900,N_17720,N_19318);
or U21901 (N_21901,N_17686,N_19368);
and U21902 (N_21902,N_18893,N_10522);
and U21903 (N_21903,N_17486,N_16607);
and U21904 (N_21904,N_11898,N_19919);
xor U21905 (N_21905,N_15518,N_16414);
and U21906 (N_21906,N_11356,N_19367);
nor U21907 (N_21907,N_11284,N_14504);
or U21908 (N_21908,N_19331,N_11555);
nand U21909 (N_21909,N_19135,N_15243);
or U21910 (N_21910,N_12860,N_16241);
and U21911 (N_21911,N_19573,N_12780);
and U21912 (N_21912,N_17438,N_10705);
nand U21913 (N_21913,N_19575,N_18590);
nand U21914 (N_21914,N_10349,N_10368);
and U21915 (N_21915,N_17578,N_13865);
nor U21916 (N_21916,N_12101,N_16797);
xor U21917 (N_21917,N_12465,N_17144);
and U21918 (N_21918,N_15760,N_15575);
or U21919 (N_21919,N_12618,N_19980);
nor U21920 (N_21920,N_11929,N_11011);
nor U21921 (N_21921,N_10306,N_10593);
or U21922 (N_21922,N_12182,N_13553);
or U21923 (N_21923,N_17517,N_14561);
and U21924 (N_21924,N_15368,N_12890);
nor U21925 (N_21925,N_16984,N_11911);
xor U21926 (N_21926,N_12503,N_16650);
nand U21927 (N_21927,N_18027,N_11503);
or U21928 (N_21928,N_16579,N_11425);
nand U21929 (N_21929,N_12132,N_10785);
or U21930 (N_21930,N_10039,N_19104);
nand U21931 (N_21931,N_15815,N_19660);
and U21932 (N_21932,N_10765,N_11891);
nand U21933 (N_21933,N_11142,N_19740);
xor U21934 (N_21934,N_15318,N_14114);
nor U21935 (N_21935,N_13738,N_15072);
xor U21936 (N_21936,N_11840,N_18060);
nor U21937 (N_21937,N_16895,N_17457);
nand U21938 (N_21938,N_14071,N_19389);
nor U21939 (N_21939,N_14176,N_17535);
nor U21940 (N_21940,N_16468,N_12456);
and U21941 (N_21941,N_18820,N_12423);
nand U21942 (N_21942,N_13159,N_15758);
or U21943 (N_21943,N_10735,N_18351);
nor U21944 (N_21944,N_10646,N_17247);
nor U21945 (N_21945,N_18570,N_10520);
and U21946 (N_21946,N_12605,N_15979);
or U21947 (N_21947,N_15259,N_17257);
and U21948 (N_21948,N_17423,N_16745);
and U21949 (N_21949,N_14727,N_18347);
nor U21950 (N_21950,N_10896,N_15835);
and U21951 (N_21951,N_17622,N_10068);
or U21952 (N_21952,N_13932,N_16875);
nor U21953 (N_21953,N_18584,N_11801);
nor U21954 (N_21954,N_12885,N_15124);
and U21955 (N_21955,N_11873,N_13758);
and U21956 (N_21956,N_10640,N_19142);
or U21957 (N_21957,N_16035,N_16397);
nor U21958 (N_21958,N_15779,N_10944);
or U21959 (N_21959,N_16443,N_16689);
nor U21960 (N_21960,N_18630,N_16431);
or U21961 (N_21961,N_17640,N_10041);
or U21962 (N_21962,N_19613,N_11536);
nor U21963 (N_21963,N_11845,N_10403);
xor U21964 (N_21964,N_19762,N_11956);
or U21965 (N_21965,N_18812,N_15224);
nand U21966 (N_21966,N_16901,N_13095);
or U21967 (N_21967,N_15772,N_15465);
nand U21968 (N_21968,N_13249,N_18818);
xnor U21969 (N_21969,N_14230,N_17632);
and U21970 (N_21970,N_16012,N_13768);
nand U21971 (N_21971,N_10585,N_13990);
nand U21972 (N_21972,N_19611,N_17796);
nor U21973 (N_21973,N_17924,N_11899);
or U21974 (N_21974,N_18929,N_17280);
or U21975 (N_21975,N_17539,N_15214);
or U21976 (N_21976,N_18313,N_11413);
and U21977 (N_21977,N_14466,N_12590);
nor U21978 (N_21978,N_19242,N_10066);
xor U21979 (N_21979,N_12927,N_12137);
and U21980 (N_21980,N_11584,N_15084);
nor U21981 (N_21981,N_10067,N_15002);
or U21982 (N_21982,N_19221,N_18382);
nand U21983 (N_21983,N_13494,N_16531);
or U21984 (N_21984,N_10914,N_18240);
nor U21985 (N_21985,N_17378,N_17439);
xnor U21986 (N_21986,N_15679,N_16936);
nor U21987 (N_21987,N_17843,N_19377);
nor U21988 (N_21988,N_13978,N_13641);
and U21989 (N_21989,N_13266,N_16750);
xnor U21990 (N_21990,N_16341,N_11204);
nand U21991 (N_21991,N_17315,N_19915);
nor U21992 (N_21992,N_12951,N_19673);
and U21993 (N_21993,N_11708,N_16435);
nand U21994 (N_21994,N_14672,N_12092);
and U21995 (N_21995,N_18207,N_11219);
or U21996 (N_21996,N_17219,N_13299);
and U21997 (N_21997,N_13467,N_15296);
nand U21998 (N_21998,N_11990,N_15766);
or U21999 (N_21999,N_16557,N_17710);
nand U22000 (N_22000,N_18466,N_18310);
and U22001 (N_22001,N_11310,N_16886);
nor U22002 (N_22002,N_10089,N_15295);
or U22003 (N_22003,N_18509,N_12333);
nor U22004 (N_22004,N_10185,N_12579);
or U22005 (N_22005,N_17011,N_16853);
nand U22006 (N_22006,N_11715,N_18255);
nor U22007 (N_22007,N_12501,N_19361);
nor U22008 (N_22008,N_13137,N_17558);
nor U22009 (N_22009,N_11334,N_10671);
nor U22010 (N_22010,N_15786,N_11854);
nor U22011 (N_22011,N_12427,N_19470);
nand U22012 (N_22012,N_12607,N_13752);
nand U22013 (N_22013,N_14008,N_11644);
xnor U22014 (N_22014,N_10851,N_14879);
nand U22015 (N_22015,N_15577,N_14309);
xor U22016 (N_22016,N_10117,N_17325);
and U22017 (N_22017,N_10404,N_14195);
and U22018 (N_22018,N_15065,N_12896);
or U22019 (N_22019,N_17680,N_12192);
nor U22020 (N_22020,N_19867,N_16816);
and U22021 (N_22021,N_14768,N_15560);
nand U22022 (N_22022,N_13913,N_14153);
and U22023 (N_22023,N_11170,N_19420);
and U22024 (N_22024,N_17692,N_17926);
nor U22025 (N_22025,N_16606,N_17206);
xnor U22026 (N_22026,N_18922,N_13862);
nor U22027 (N_22027,N_18103,N_17763);
or U22028 (N_22028,N_18068,N_12111);
and U22029 (N_22029,N_13369,N_15972);
or U22030 (N_22030,N_10840,N_12143);
and U22031 (N_22031,N_10198,N_11791);
nand U22032 (N_22032,N_18222,N_12772);
and U22033 (N_22033,N_13156,N_19332);
nor U22034 (N_22034,N_10537,N_18618);
xor U22035 (N_22035,N_18881,N_17376);
or U22036 (N_22036,N_14800,N_15703);
nor U22037 (N_22037,N_12723,N_11586);
or U22038 (N_22038,N_11814,N_18042);
nand U22039 (N_22039,N_19601,N_11718);
and U22040 (N_22040,N_12055,N_18432);
or U22041 (N_22041,N_16071,N_17903);
or U22042 (N_22042,N_11655,N_17432);
xor U22043 (N_22043,N_15396,N_14182);
or U22044 (N_22044,N_18786,N_11662);
or U22045 (N_22045,N_10496,N_10093);
or U22046 (N_22046,N_19279,N_11417);
and U22047 (N_22047,N_16573,N_15108);
or U22048 (N_22048,N_14874,N_11055);
and U22049 (N_22049,N_10536,N_11676);
xnor U22050 (N_22050,N_16794,N_19576);
xor U22051 (N_22051,N_14578,N_15894);
or U22052 (N_22052,N_11453,N_11255);
xnor U22053 (N_22053,N_11281,N_11998);
nand U22054 (N_22054,N_15603,N_11564);
nand U22055 (N_22055,N_13802,N_17865);
nor U22056 (N_22056,N_12913,N_18913);
nor U22057 (N_22057,N_13272,N_12204);
xnor U22058 (N_22058,N_15631,N_15017);
and U22059 (N_22059,N_19483,N_11569);
nor U22060 (N_22060,N_19728,N_19328);
nor U22061 (N_22061,N_13662,N_18722);
nor U22062 (N_22062,N_12837,N_15749);
nand U22063 (N_22063,N_13045,N_12593);
and U22064 (N_22064,N_19480,N_13549);
nand U22065 (N_22065,N_14792,N_19676);
and U22066 (N_22066,N_18434,N_14059);
nor U22067 (N_22067,N_18635,N_12925);
or U22068 (N_22068,N_13165,N_11312);
nand U22069 (N_22069,N_11590,N_10690);
and U22070 (N_22070,N_13316,N_19252);
nor U22071 (N_22071,N_12164,N_18859);
nor U22072 (N_22072,N_16160,N_17801);
and U22073 (N_22073,N_16701,N_13345);
and U22074 (N_22074,N_12390,N_16508);
nor U22075 (N_22075,N_19416,N_16044);
or U22076 (N_22076,N_11686,N_18696);
and U22077 (N_22077,N_11524,N_18002);
and U22078 (N_22078,N_18729,N_14876);
and U22079 (N_22079,N_14432,N_14393);
or U22080 (N_22080,N_17916,N_10742);
and U22081 (N_22081,N_10957,N_14136);
nor U22082 (N_22082,N_12648,N_13440);
nor U22083 (N_22083,N_19275,N_16192);
xor U22084 (N_22084,N_16158,N_18201);
xor U22085 (N_22085,N_13606,N_11527);
nor U22086 (N_22086,N_17006,N_15250);
nand U22087 (N_22087,N_13708,N_13288);
or U22088 (N_22088,N_13618,N_15278);
nor U22089 (N_22089,N_16534,N_15366);
and U22090 (N_22090,N_14421,N_12892);
xor U22091 (N_22091,N_16472,N_13429);
or U22092 (N_22092,N_14559,N_10529);
nor U22093 (N_22093,N_12681,N_18343);
and U22094 (N_22094,N_17311,N_15442);
and U22095 (N_22095,N_11903,N_12436);
and U22096 (N_22096,N_15305,N_18805);
nor U22097 (N_22097,N_11285,N_19871);
and U22098 (N_22098,N_17419,N_15091);
xnor U22099 (N_22099,N_11039,N_14740);
or U22100 (N_22100,N_19546,N_17668);
nor U22101 (N_22101,N_19349,N_17751);
and U22102 (N_22102,N_13029,N_11531);
and U22103 (N_22103,N_14085,N_10302);
and U22104 (N_22104,N_13059,N_19910);
and U22105 (N_22105,N_18784,N_10661);
or U22106 (N_22106,N_13225,N_11769);
nor U22107 (N_22107,N_13619,N_10998);
xnor U22108 (N_22108,N_16276,N_10015);
xnor U22109 (N_22109,N_12742,N_16445);
nand U22110 (N_22110,N_11302,N_18908);
or U22111 (N_22111,N_13356,N_15736);
nor U22112 (N_22112,N_15482,N_17785);
nand U22113 (N_22113,N_17820,N_11129);
nand U22114 (N_22114,N_19419,N_11335);
nor U22115 (N_22115,N_17775,N_18237);
and U22116 (N_22116,N_16336,N_13280);
or U22117 (N_22117,N_10409,N_18867);
nand U22118 (N_22118,N_14898,N_13117);
nor U22119 (N_22119,N_11719,N_13186);
and U22120 (N_22120,N_12099,N_17336);
xnor U22121 (N_22121,N_11005,N_15658);
and U22122 (N_22122,N_18605,N_16437);
nand U22123 (N_22123,N_13485,N_17862);
nor U22124 (N_22124,N_13236,N_16518);
and U22125 (N_22125,N_11235,N_14165);
nor U22126 (N_22126,N_19888,N_15870);
and U22127 (N_22127,N_19227,N_12485);
or U22128 (N_22128,N_14811,N_17027);
and U22129 (N_22129,N_13491,N_19006);
or U22130 (N_22130,N_14936,N_12952);
or U22131 (N_22131,N_13390,N_13926);
nand U22132 (N_22132,N_16656,N_16492);
or U22133 (N_22133,N_12158,N_18416);
nand U22134 (N_22134,N_11074,N_16080);
and U22135 (N_22135,N_17856,N_10217);
and U22136 (N_22136,N_12711,N_19025);
nor U22137 (N_22137,N_13938,N_13437);
nor U22138 (N_22138,N_19580,N_13647);
nor U22139 (N_22139,N_17721,N_13172);
nand U22140 (N_22140,N_10188,N_17222);
xnor U22141 (N_22141,N_17527,N_15323);
nand U22142 (N_22142,N_13648,N_15248);
or U22143 (N_22143,N_19384,N_15877);
xnor U22144 (N_22144,N_19063,N_11045);
and U22145 (N_22145,N_17053,N_15057);
and U22146 (N_22146,N_10581,N_15808);
nand U22147 (N_22147,N_18370,N_14005);
nand U22148 (N_22148,N_12967,N_13124);
nor U22149 (N_22149,N_19924,N_16983);
and U22150 (N_22150,N_18891,N_19655);
xnor U22151 (N_22151,N_13200,N_12331);
or U22152 (N_22152,N_15041,N_18062);
and U22153 (N_22153,N_14722,N_18832);
and U22154 (N_22154,N_16962,N_12468);
nor U22155 (N_22155,N_18664,N_19118);
or U22156 (N_22156,N_10917,N_13078);
nor U22157 (N_22157,N_17353,N_16436);
and U22158 (N_22158,N_15401,N_13947);
xnor U22159 (N_22159,N_14213,N_16929);
and U22160 (N_22160,N_10181,N_17672);
nand U22161 (N_22161,N_15403,N_12403);
or U22162 (N_22162,N_15882,N_11433);
and U22163 (N_22163,N_13353,N_14540);
and U22164 (N_22164,N_15638,N_11617);
nand U22165 (N_22165,N_11138,N_15604);
or U22166 (N_22166,N_11855,N_16198);
nand U22167 (N_22167,N_13596,N_14088);
and U22168 (N_22168,N_11786,N_17165);
nand U22169 (N_22169,N_18010,N_11640);
and U22170 (N_22170,N_19350,N_11014);
and U22171 (N_22171,N_10999,N_14318);
or U22172 (N_22172,N_10688,N_18853);
xnor U22173 (N_22173,N_18423,N_11274);
nand U22174 (N_22174,N_12394,N_11706);
or U22175 (N_22175,N_19442,N_13346);
and U22176 (N_22176,N_19695,N_10396);
and U22177 (N_22177,N_16641,N_13327);
and U22178 (N_22178,N_18127,N_16062);
or U22179 (N_22179,N_15167,N_14550);
nand U22180 (N_22180,N_19003,N_13736);
nor U22181 (N_22181,N_19316,N_18652);
xnor U22182 (N_22182,N_11376,N_19429);
nor U22183 (N_22183,N_17559,N_16880);
xnor U22184 (N_22184,N_19482,N_13650);
and U22185 (N_22185,N_14751,N_14159);
nor U22186 (N_22186,N_15449,N_14590);
nor U22187 (N_22187,N_16718,N_13847);
nand U22188 (N_22188,N_17427,N_10255);
or U22189 (N_22189,N_16351,N_15524);
and U22190 (N_22190,N_16411,N_13898);
nor U22191 (N_22191,N_13309,N_17496);
or U22192 (N_22192,N_14560,N_18582);
and U22193 (N_22193,N_15804,N_11340);
and U22194 (N_22194,N_12853,N_18357);
nand U22195 (N_22195,N_13290,N_17800);
xnor U22196 (N_22196,N_10922,N_15128);
or U22197 (N_22197,N_17906,N_13062);
nand U22198 (N_22198,N_18986,N_16669);
nor U22199 (N_22199,N_12744,N_11756);
nand U22200 (N_22200,N_10126,N_13408);
nand U22201 (N_22201,N_13997,N_18005);
nand U22202 (N_22202,N_18175,N_13051);
nand U22203 (N_22203,N_17641,N_13456);
and U22204 (N_22204,N_10625,N_18144);
or U22205 (N_22205,N_17372,N_17032);
or U22206 (N_22206,N_11456,N_19320);
and U22207 (N_22207,N_17163,N_15549);
nand U22208 (N_22208,N_11576,N_10081);
xnor U22209 (N_22209,N_14860,N_18847);
nor U22210 (N_22210,N_10421,N_11311);
and U22211 (N_22211,N_18203,N_11294);
or U22212 (N_22212,N_13631,N_11837);
nand U22213 (N_22213,N_16766,N_12836);
or U22214 (N_22214,N_15421,N_11546);
nand U22215 (N_22215,N_17579,N_13937);
nand U22216 (N_22216,N_13753,N_19121);
nor U22217 (N_22217,N_15329,N_14054);
nor U22218 (N_22218,N_19865,N_18138);
nand U22219 (N_22219,N_16083,N_13431);
or U22220 (N_22220,N_13804,N_14602);
or U22221 (N_22221,N_11960,N_14717);
xnor U22222 (N_22222,N_10169,N_10844);
and U22223 (N_22223,N_14360,N_16872);
xor U22224 (N_22224,N_13105,N_17205);
or U22225 (N_22225,N_19633,N_10949);
or U22226 (N_22226,N_19073,N_12589);
nand U22227 (N_22227,N_11591,N_17722);
nand U22228 (N_22228,N_18730,N_15924);
nand U22229 (N_22229,N_12958,N_18391);
nand U22230 (N_22230,N_13689,N_16870);
nand U22231 (N_22231,N_12714,N_15683);
nand U22232 (N_22232,N_19930,N_12879);
xor U22233 (N_22233,N_17645,N_14842);
nor U22234 (N_22234,N_12122,N_19311);
and U22235 (N_22235,N_19846,N_18265);
or U22236 (N_22236,N_10382,N_13834);
nor U22237 (N_22237,N_15187,N_17870);
nor U22238 (N_22238,N_10193,N_12343);
and U22239 (N_22239,N_18208,N_13635);
or U22240 (N_22240,N_15925,N_19732);
nand U22241 (N_22241,N_11392,N_18601);
or U22242 (N_22242,N_10973,N_17193);
nor U22243 (N_22243,N_10560,N_14007);
nor U22244 (N_22244,N_12474,N_10229);
xor U22245 (N_22245,N_18668,N_10559);
nor U22246 (N_22246,N_10038,N_12710);
xnor U22247 (N_22247,N_17273,N_16691);
or U22248 (N_22248,N_15610,N_15309);
nor U22249 (N_22249,N_17949,N_17724);
nor U22250 (N_22250,N_19653,N_14185);
nor U22251 (N_22251,N_16321,N_14029);
xor U22252 (N_22252,N_10675,N_11633);
and U22253 (N_22253,N_16497,N_12956);
and U22254 (N_22254,N_17509,N_13682);
nor U22255 (N_22255,N_18858,N_18782);
and U22256 (N_22256,N_13825,N_12387);
or U22257 (N_22257,N_17510,N_19532);
nand U22258 (N_22258,N_11924,N_16461);
and U22259 (N_22259,N_16162,N_13314);
or U22260 (N_22260,N_17538,N_16041);
or U22261 (N_22261,N_16379,N_18441);
nand U22262 (N_22262,N_12613,N_16520);
xnor U22263 (N_22263,N_18431,N_18126);
nand U22264 (N_22264,N_14497,N_10313);
nor U22265 (N_22265,N_13963,N_14270);
nor U22266 (N_22266,N_14269,N_19909);
or U22267 (N_22267,N_13311,N_14704);
nand U22268 (N_22268,N_18968,N_10717);
nor U22269 (N_22269,N_19988,N_12134);
nor U22270 (N_22270,N_11930,N_18574);
nand U22271 (N_22271,N_18978,N_19703);
nand U22272 (N_22272,N_18790,N_16374);
or U22273 (N_22273,N_14514,N_11729);
nand U22274 (N_22274,N_15493,N_11165);
and U22275 (N_22275,N_14547,N_17401);
nand U22276 (N_22276,N_11502,N_19512);
xor U22277 (N_22277,N_10905,N_18294);
nor U22278 (N_22278,N_19801,N_13255);
and U22279 (N_22279,N_16670,N_11136);
nor U22280 (N_22280,N_14636,N_18926);
nor U22281 (N_22281,N_12481,N_10425);
or U22282 (N_22282,N_12191,N_17076);
nand U22283 (N_22283,N_12870,N_15394);
nand U22284 (N_22284,N_14245,N_18552);
or U22285 (N_22285,N_10210,N_13154);
nand U22286 (N_22286,N_12688,N_18497);
nor U22287 (N_22287,N_11295,N_18768);
xor U22288 (N_22288,N_13740,N_12601);
nor U22289 (N_22289,N_10042,N_18936);
and U22290 (N_22290,N_19784,N_19009);
nor U22291 (N_22291,N_13545,N_17467);
nor U22292 (N_22292,N_10665,N_11290);
and U22293 (N_22293,N_15820,N_10428);
or U22294 (N_22294,N_17018,N_18217);
nor U22295 (N_22295,N_18887,N_15169);
and U22296 (N_22296,N_10809,N_14020);
nand U22297 (N_22297,N_17390,N_16157);
or U22298 (N_22298,N_13861,N_15336);
or U22299 (N_22299,N_19741,N_13868);
or U22300 (N_22300,N_12716,N_17475);
nor U22301 (N_22301,N_13209,N_13851);
nand U22302 (N_22302,N_18636,N_10719);
nand U22303 (N_22303,N_17151,N_10650);
or U22304 (N_22304,N_16331,N_15792);
nor U22305 (N_22305,N_19099,N_16856);
or U22306 (N_22306,N_14524,N_10561);
nor U22307 (N_22307,N_15581,N_14122);
nand U22308 (N_22308,N_19209,N_18022);
or U22309 (N_22309,N_14112,N_16593);
nand U22310 (N_22310,N_13905,N_13447);
or U22311 (N_22311,N_17565,N_18930);
nor U22312 (N_22312,N_13403,N_16307);
or U22313 (N_22313,N_10162,N_11725);
xor U22314 (N_22314,N_11359,N_15475);
and U22315 (N_22315,N_15940,N_12595);
xnor U22316 (N_22316,N_10956,N_16234);
nor U22317 (N_22317,N_10512,N_15168);
nand U22318 (N_22318,N_17141,N_11180);
and U22319 (N_22319,N_18358,N_10121);
and U22320 (N_22320,N_10821,N_13452);
or U22321 (N_22321,N_17741,N_14051);
and U22322 (N_22322,N_14369,N_18407);
and U22323 (N_22323,N_17075,N_13052);
nand U22324 (N_22324,N_13460,N_17202);
nor U22325 (N_22325,N_10150,N_15484);
or U22326 (N_22326,N_12176,N_17708);
and U22327 (N_22327,N_18655,N_18915);
and U22328 (N_22328,N_14828,N_10149);
and U22329 (N_22329,N_12381,N_18281);
xnor U22330 (N_22330,N_17610,N_11364);
and U22331 (N_22331,N_14569,N_10981);
nand U22332 (N_22332,N_17135,N_18943);
nor U22333 (N_22333,N_10044,N_13979);
nand U22334 (N_22334,N_10636,N_19979);
nor U22335 (N_22335,N_15393,N_18975);
nor U22336 (N_22336,N_12283,N_19840);
and U22337 (N_22337,N_13015,N_13934);
and U22338 (N_22338,N_12417,N_14674);
or U22339 (N_22339,N_19199,N_13442);
and U22340 (N_22340,N_13410,N_12429);
and U22341 (N_22341,N_17161,N_10106);
or U22342 (N_22342,N_10572,N_16865);
xnor U22343 (N_22343,N_12147,N_19593);
and U22344 (N_22344,N_19571,N_11263);
nand U22345 (N_22345,N_10633,N_13212);
nor U22346 (N_22346,N_12917,N_15473);
and U22347 (N_22347,N_13742,N_12510);
xor U22348 (N_22348,N_18774,N_18764);
or U22349 (N_22349,N_10867,N_16615);
and U22350 (N_22350,N_17847,N_18993);
nor U22351 (N_22351,N_18368,N_18595);
nand U22352 (N_22352,N_15190,N_10374);
nand U22353 (N_22353,N_19864,N_11467);
or U22354 (N_22354,N_19773,N_12759);
nand U22355 (N_22355,N_16172,N_14609);
nand U22356 (N_22356,N_15422,N_10275);
and U22357 (N_22357,N_14645,N_16953);
and U22358 (N_22358,N_15237,N_16483);
nand U22359 (N_22359,N_17577,N_17109);
xor U22360 (N_22360,N_17966,N_17366);
nand U22361 (N_22361,N_11090,N_12537);
or U22362 (N_22362,N_18504,N_11771);
xor U22363 (N_22363,N_12691,N_14579);
nor U22364 (N_22364,N_12148,N_12037);
or U22365 (N_22365,N_10335,N_10869);
nand U22366 (N_22366,N_10783,N_13888);
nand U22367 (N_22367,N_19085,N_12114);
and U22368 (N_22368,N_19169,N_10460);
nor U22369 (N_22369,N_14192,N_10013);
or U22370 (N_22370,N_15743,N_11041);
or U22371 (N_22371,N_19725,N_12139);
xor U22372 (N_22372,N_10101,N_10435);
or U22373 (N_22373,N_15764,N_10847);
or U22374 (N_22374,N_10452,N_11009);
or U22375 (N_22375,N_15431,N_19602);
or U22376 (N_22376,N_19702,N_11838);
nor U22377 (N_22377,N_16154,N_19839);
nand U22378 (N_22378,N_18178,N_17177);
or U22379 (N_22379,N_19426,N_12179);
and U22380 (N_22380,N_15960,N_12719);
and U22381 (N_22381,N_17225,N_17748);
or U22382 (N_22382,N_14446,N_10480);
or U22383 (N_22383,N_17469,N_16709);
nand U22384 (N_22384,N_18720,N_11193);
nor U22385 (N_22385,N_18806,N_11448);
nand U22386 (N_22386,N_17815,N_17593);
nor U22387 (N_22387,N_14317,N_16280);
and U22388 (N_22388,N_18216,N_17854);
nand U22389 (N_22389,N_11065,N_10004);
or U22390 (N_22390,N_14111,N_12358);
or U22391 (N_22391,N_14467,N_18013);
xor U22392 (N_22392,N_13554,N_12285);
or U22393 (N_22393,N_14915,N_16406);
xor U22394 (N_22394,N_13850,N_12944);
and U22395 (N_22395,N_12649,N_17836);
and U22396 (N_22396,N_13941,N_14516);
nor U22397 (N_22397,N_13321,N_18792);
nand U22398 (N_22398,N_17077,N_12494);
or U22399 (N_22399,N_16127,N_14759);
or U22400 (N_22400,N_10273,N_17070);
xnor U22401 (N_22401,N_18320,N_11215);
xor U22402 (N_22402,N_15723,N_11506);
or U22403 (N_22403,N_12699,N_15807);
and U22404 (N_22404,N_17061,N_11526);
nand U22405 (N_22405,N_14914,N_11391);
nor U22406 (N_22406,N_13595,N_13046);
and U22407 (N_22407,N_14857,N_17242);
or U22408 (N_22408,N_16716,N_15249);
and U22409 (N_22409,N_10624,N_14101);
xor U22410 (N_22410,N_15183,N_17812);
nand U22411 (N_22411,N_16843,N_12845);
nor U22412 (N_22412,N_18117,N_14068);
nand U22413 (N_22413,N_13684,N_17464);
nor U22414 (N_22414,N_19726,N_11408);
nor U22415 (N_22415,N_17920,N_17305);
nor U22416 (N_22416,N_18845,N_11872);
nand U22417 (N_22417,N_12858,N_11102);
nor U22418 (N_22418,N_17264,N_11909);
xnor U22419 (N_22419,N_19430,N_11250);
xor U22420 (N_22420,N_13910,N_11261);
nor U22421 (N_22421,N_12126,N_12542);
nand U22422 (N_22422,N_12748,N_11230);
xnor U22423 (N_22423,N_16597,N_19543);
nand U22424 (N_22424,N_12029,N_14034);
or U22425 (N_22425,N_18000,N_16734);
or U22426 (N_22426,N_15978,N_19000);
xnor U22427 (N_22427,N_14877,N_19168);
xor U22428 (N_22428,N_16484,N_16737);
and U22429 (N_22429,N_19468,N_14374);
or U22430 (N_22430,N_10868,N_11471);
nand U22431 (N_22431,N_16075,N_15696);
nand U22432 (N_22432,N_16912,N_18499);
nand U22433 (N_22433,N_15988,N_15916);
xnor U22434 (N_22434,N_18918,N_19579);
xor U22435 (N_22435,N_19509,N_13916);
nor U22436 (N_22436,N_16152,N_15415);
and U22437 (N_22437,N_14728,N_11272);
nand U22438 (N_22438,N_12898,N_12348);
nor U22439 (N_22439,N_19109,N_14448);
nand U22440 (N_22440,N_18508,N_12588);
nand U22441 (N_22441,N_19825,N_10553);
nand U22442 (N_22442,N_12479,N_13406);
or U22443 (N_22443,N_11462,N_13903);
nand U22444 (N_22444,N_16054,N_18650);
or U22445 (N_22445,N_18333,N_10751);
nand U22446 (N_22446,N_15654,N_10152);
nand U22447 (N_22447,N_12036,N_14521);
or U22448 (N_22448,N_13628,N_13859);
or U22449 (N_22449,N_16804,N_14744);
nand U22450 (N_22450,N_19896,N_19796);
nor U22451 (N_22451,N_14168,N_15175);
or U22452 (N_22452,N_14065,N_16326);
nor U22453 (N_22453,N_11704,N_11306);
or U22454 (N_22454,N_19369,N_14138);
and U22455 (N_22455,N_16494,N_14736);
or U22456 (N_22456,N_16985,N_15003);
nor U22457 (N_22457,N_14001,N_16587);
or U22458 (N_22458,N_15583,N_13453);
and U22459 (N_22459,N_18933,N_16740);
or U22460 (N_22460,N_13767,N_17706);
or U22461 (N_22461,N_14676,N_15795);
and U22462 (N_22462,N_15161,N_12544);
nand U22463 (N_22463,N_18252,N_19197);
nand U22464 (N_22464,N_10565,N_15407);
or U22465 (N_22465,N_12162,N_16232);
nand U22466 (N_22466,N_13082,N_12793);
nor U22467 (N_22467,N_13481,N_18152);
nor U22468 (N_22468,N_10526,N_17425);
and U22469 (N_22469,N_17784,N_12571);
xor U22470 (N_22470,N_19927,N_12803);
nor U22471 (N_22471,N_16033,N_16338);
nand U22472 (N_22472,N_16212,N_11038);
xnor U22473 (N_22473,N_15755,N_14342);
or U22474 (N_22474,N_14053,N_19386);
nand U22475 (N_22475,N_17288,N_18935);
nand U22476 (N_22476,N_18549,N_13633);
nand U22477 (N_22477,N_19905,N_12625);
or U22478 (N_22478,N_11291,N_15565);
nor U22479 (N_22479,N_17677,N_11823);
nor U22480 (N_22480,N_17368,N_14243);
nand U22481 (N_22481,N_13096,N_18162);
and U22482 (N_22482,N_15832,N_15093);
and U22483 (N_22483,N_19004,N_15462);
nor U22484 (N_22484,N_10933,N_12157);
nand U22485 (N_22485,N_17468,N_12757);
or U22486 (N_22486,N_15198,N_16199);
nand U22487 (N_22487,N_11863,N_11494);
or U22488 (N_22488,N_16370,N_16771);
or U22489 (N_22489,N_17189,N_10578);
nor U22490 (N_22490,N_19303,N_12201);
xnor U22491 (N_22491,N_16842,N_18363);
or U22492 (N_22492,N_11868,N_13676);
or U22493 (N_22493,N_14256,N_12524);
or U22494 (N_22494,N_15050,N_11338);
nand U22495 (N_22495,N_16952,N_16286);
nor U22496 (N_22496,N_15885,N_17757);
nand U22497 (N_22497,N_19291,N_14173);
nor U22498 (N_22498,N_12527,N_17373);
nor U22499 (N_22499,N_12507,N_19996);
or U22500 (N_22500,N_15019,N_11910);
xnor U22501 (N_22501,N_10725,N_15362);
nand U22502 (N_22502,N_17701,N_17908);
nand U22503 (N_22503,N_14335,N_16646);
nand U22504 (N_22504,N_17098,N_17679);
and U22505 (N_22505,N_15203,N_13714);
nor U22506 (N_22506,N_11409,N_12361);
nor U22507 (N_22507,N_18553,N_19951);
and U22508 (N_22508,N_18592,N_13961);
nor U22509 (N_22509,N_19504,N_11679);
or U22510 (N_22510,N_11861,N_11611);
nor U22511 (N_22511,N_14017,N_12259);
nor U22512 (N_22512,N_19989,N_12677);
nor U22513 (N_22513,N_16053,N_12038);
xor U22514 (N_22514,N_18100,N_19731);
xor U22515 (N_22515,N_18842,N_12278);
and U22516 (N_22516,N_11352,N_11387);
nor U22517 (N_22517,N_17945,N_19018);
or U22518 (N_22518,N_11563,N_10086);
xor U22519 (N_22519,N_12559,N_15529);
or U22520 (N_22520,N_14221,N_19672);
xnor U22521 (N_22521,N_11848,N_19170);
and U22522 (N_22522,N_10687,N_19880);
nor U22523 (N_22523,N_16809,N_19183);
xnor U22524 (N_22524,N_18024,N_15660);
nor U22525 (N_22525,N_17186,N_16516);
nand U22526 (N_22526,N_16541,N_19687);
and U22527 (N_22527,N_12973,N_12197);
nand U22528 (N_22528,N_12658,N_15372);
nand U22529 (N_22529,N_11957,N_13667);
nor U22530 (N_22530,N_16643,N_18713);
and U22531 (N_22531,N_17204,N_18328);
and U22532 (N_22532,N_11082,N_13201);
xor U22533 (N_22533,N_12667,N_18739);
or U22534 (N_22534,N_15665,N_14551);
xor U22535 (N_22535,N_16220,N_16424);
xnor U22536 (N_22536,N_15028,N_10507);
xor U22537 (N_22537,N_15617,N_16150);
nand U22538 (N_22538,N_19017,N_17780);
nor U22539 (N_22539,N_13254,N_10290);
xor U22540 (N_22540,N_13164,N_12936);
or U22541 (N_22541,N_13726,N_16605);
and U22542 (N_22542,N_19953,N_18051);
or U22543 (N_22543,N_13593,N_14611);
or U22544 (N_22544,N_15109,N_19309);
xnor U22545 (N_22545,N_10930,N_16885);
nand U22546 (N_22546,N_15379,N_11336);
nand U22547 (N_22547,N_12452,N_11458);
or U22548 (N_22548,N_19225,N_18029);
xor U22549 (N_22549,N_15932,N_10855);
or U22550 (N_22550,N_10134,N_11752);
and U22551 (N_22551,N_19743,N_13842);
and U22552 (N_22552,N_14471,N_14424);
or U22553 (N_22553,N_14344,N_13340);
nand U22554 (N_22554,N_13643,N_11757);
nor U22555 (N_22555,N_18882,N_19925);
nand U22556 (N_22556,N_19668,N_18036);
nor U22557 (N_22557,N_13176,N_12459);
and U22558 (N_22558,N_10604,N_11385);
nand U22559 (N_22559,N_18239,N_12794);
or U22560 (N_22560,N_17830,N_10699);
nand U22561 (N_22561,N_10172,N_12281);
and U22562 (N_22562,N_14064,N_12025);
and U22563 (N_22563,N_13756,N_17277);
nor U22564 (N_22564,N_18813,N_14113);
nor U22565 (N_22565,N_10009,N_18296);
nor U22566 (N_22566,N_14157,N_14428);
nand U22567 (N_22567,N_10145,N_11658);
and U22568 (N_22568,N_14449,N_10311);
nor U22569 (N_22569,N_18567,N_18007);
and U22570 (N_22570,N_17274,N_16077);
and U22571 (N_22571,N_16427,N_17038);
or U22572 (N_22572,N_13896,N_17630);
xor U22573 (N_22573,N_11537,N_13112);
xor U22574 (N_22574,N_10533,N_15917);
nand U22575 (N_22575,N_12341,N_14660);
or U22576 (N_22576,N_11888,N_18492);
xnor U22577 (N_22577,N_12830,N_16295);
xnor U22578 (N_22578,N_17194,N_10712);
nand U22579 (N_22579,N_18465,N_19893);
xnor U22580 (N_22580,N_13995,N_19304);
nand U22581 (N_22581,N_13824,N_18670);
nor U22582 (N_22582,N_17813,N_10732);
or U22583 (N_22583,N_12168,N_10729);
nor U22584 (N_22584,N_11606,N_18816);
nor U22585 (N_22585,N_10986,N_16859);
nand U22586 (N_22586,N_14606,N_13774);
or U22587 (N_22587,N_13441,N_17101);
nor U22588 (N_22588,N_11634,N_14566);
xor U22589 (N_22589,N_12820,N_19858);
and U22590 (N_22590,N_15793,N_16528);
or U22591 (N_22591,N_18638,N_10017);
or U22592 (N_22592,N_13601,N_12984);
nand U22593 (N_22593,N_15151,N_19623);
and U22594 (N_22594,N_19900,N_13933);
nor U22595 (N_22595,N_19010,N_17506);
or U22596 (N_22596,N_19917,N_18136);
nand U22597 (N_22597,N_15503,N_16256);
and U22598 (N_22598,N_13688,N_13681);
nand U22599 (N_22599,N_10802,N_15143);
or U22600 (N_22600,N_18396,N_17123);
and U22601 (N_22601,N_15855,N_11734);
or U22602 (N_22602,N_17518,N_17589);
nor U22603 (N_22603,N_19191,N_17657);
or U22604 (N_22604,N_18736,N_12273);
or U22605 (N_22605,N_16265,N_18308);
and U22606 (N_22606,N_17884,N_17745);
and U22607 (N_22607,N_16950,N_15657);
or U22608 (N_22608,N_11827,N_10761);
nor U22609 (N_22609,N_15586,N_11275);
and U22610 (N_22610,N_10513,N_12184);
or U22611 (N_22611,N_13469,N_10033);
xor U22612 (N_22612,N_18186,N_19241);
nand U22613 (N_22613,N_12428,N_19503);
or U22614 (N_22614,N_18179,N_11189);
or U22615 (N_22615,N_11314,N_19964);
or U22616 (N_22616,N_15838,N_16330);
nor U22617 (N_22617,N_18776,N_10700);
nand U22618 (N_22618,N_11227,N_17429);
nor U22619 (N_22619,N_12498,N_12722);
nor U22620 (N_22620,N_12277,N_10499);
or U22621 (N_22621,N_10446,N_12532);
nand U22622 (N_22622,N_11109,N_19828);
nand U22623 (N_22623,N_17743,N_12460);
nor U22624 (N_22624,N_13599,N_10171);
nand U22625 (N_22625,N_16372,N_11104);
and U22626 (N_22626,N_19856,N_14389);
and U22627 (N_22627,N_10644,N_10856);
nand U22628 (N_22628,N_14199,N_17207);
xnor U22629 (N_22629,N_14499,N_18014);
or U22630 (N_22630,N_13144,N_17276);
or U22631 (N_22631,N_19283,N_13476);
nor U22632 (N_22632,N_10733,N_10128);
nor U22633 (N_22633,N_18120,N_17117);
or U22634 (N_22634,N_12703,N_19615);
or U22635 (N_22635,N_14687,N_19983);
nor U22636 (N_22636,N_19904,N_10614);
and U22637 (N_22637,N_11394,N_15021);
and U22638 (N_22638,N_10543,N_15718);
or U22639 (N_22639,N_16946,N_13731);
and U22640 (N_22640,N_16181,N_11965);
nand U22641 (N_22641,N_17282,N_16413);
nand U22642 (N_22642,N_17773,N_19872);
or U22643 (N_22643,N_10883,N_19537);
nor U22644 (N_22644,N_10211,N_13525);
xor U22645 (N_22645,N_15953,N_15085);
and U22646 (N_22646,N_19804,N_15842);
nor U22647 (N_22647,N_10438,N_19661);
or U22648 (N_22648,N_15360,N_19472);
and U22649 (N_22649,N_12795,N_18387);
nand U22650 (N_22650,N_18892,N_19922);
nor U22651 (N_22651,N_10450,N_19030);
nand U22652 (N_22652,N_13559,N_11017);
and U22653 (N_22653,N_12267,N_16478);
nor U22654 (N_22654,N_10964,N_15543);
nand U22655 (N_22655,N_11123,N_16074);
or U22656 (N_22656,N_12627,N_17738);
nand U22657 (N_22657,N_13047,N_15949);
nor U22658 (N_22658,N_16368,N_16024);
and U22659 (N_22659,N_14790,N_18980);
or U22660 (N_22660,N_13375,N_19764);
and U22661 (N_22661,N_14218,N_12567);
xor U22662 (N_22662,N_14305,N_13088);
or U22663 (N_22663,N_16361,N_12525);
nand U22664 (N_22664,N_15533,N_10434);
and U22665 (N_22665,N_11836,N_15466);
nor U22666 (N_22666,N_14304,N_15228);
nor U22667 (N_22667,N_12788,N_12002);
nor U22668 (N_22668,N_19887,N_12643);
or U22669 (N_22669,N_18458,N_11267);
or U22670 (N_22670,N_10238,N_16300);
and U22671 (N_22671,N_12404,N_19567);
or U22672 (N_22672,N_16610,N_13444);
and U22673 (N_22673,N_17371,N_11651);
nand U22674 (N_22674,N_10900,N_19479);
or U22675 (N_22675,N_18460,N_18743);
nor U22676 (N_22676,N_19950,N_12752);
nand U22677 (N_22677,N_19694,N_10261);
and U22678 (N_22678,N_19564,N_18536);
or U22679 (N_22679,N_18079,N_14630);
nor U22680 (N_22680,N_14041,N_15077);
xor U22681 (N_22681,N_14262,N_11024);
xnor U22682 (N_22682,N_14358,N_14554);
and U22683 (N_22683,N_18131,N_10874);
and U22684 (N_22684,N_17522,N_19889);
and U22685 (N_22685,N_14139,N_12671);
nor U22686 (N_22686,N_12493,N_14533);
nand U22687 (N_22687,N_15331,N_13992);
nand U22688 (N_22688,N_12461,N_16779);
and U22689 (N_22689,N_15649,N_16623);
nand U22690 (N_22690,N_18128,N_18522);
and U22691 (N_22691,N_10955,N_11181);
or U22692 (N_22692,N_18709,N_10600);
nor U22693 (N_22693,N_12008,N_15639);
nor U22694 (N_22694,N_10199,N_16470);
nor U22695 (N_22695,N_10825,N_18666);
or U22696 (N_22696,N_19376,N_16715);
xnor U22697 (N_22697,N_14487,N_13532);
nand U22698 (N_22698,N_14848,N_12949);
nand U22699 (N_22699,N_18139,N_11595);
nor U22700 (N_22700,N_10938,N_14571);
nand U22701 (N_22701,N_16874,N_14580);
or U22702 (N_22702,N_17437,N_18728);
xor U22703 (N_22703,N_16523,N_13013);
and U22704 (N_22704,N_13180,N_19569);
and U22705 (N_22705,N_14939,N_13115);
nor U22706 (N_22706,N_13071,N_16346);
nand U22707 (N_22707,N_13108,N_13053);
or U22708 (N_22708,N_18164,N_16230);
or U22709 (N_22709,N_16235,N_11257);
or U22710 (N_22710,N_12849,N_14169);
or U22711 (N_22711,N_11774,N_17142);
and U22712 (N_22712,N_11288,N_15355);
nand U22713 (N_22713,N_17281,N_13091);
or U22714 (N_22714,N_11324,N_15297);
nand U22715 (N_22715,N_11035,N_15874);
and U22716 (N_22716,N_13331,N_14891);
nor U22717 (N_22717,N_13339,N_19433);
nand U22718 (N_22718,N_19139,N_10165);
and U22719 (N_22719,N_13743,N_15571);
and U22720 (N_22720,N_17548,N_18667);
xor U22721 (N_22721,N_17208,N_18527);
nand U22722 (N_22722,N_12533,N_19645);
xnor U22723 (N_22723,N_11317,N_10340);
or U22724 (N_22724,N_15507,N_15884);
and U22725 (N_22725,N_18526,N_14802);
and U22726 (N_22726,N_14827,N_11229);
and U22727 (N_22727,N_18785,N_11573);
nor U22728 (N_22728,N_17481,N_16961);
xor U22729 (N_22729,N_10552,N_17844);
xnor U22730 (N_22730,N_15240,N_13407);
xor U22731 (N_22731,N_19076,N_19452);
nand U22732 (N_22732,N_13697,N_14861);
or U22733 (N_22733,N_10487,N_15439);
nor U22734 (N_22734,N_15663,N_14098);
nor U22735 (N_22735,N_11541,N_13653);
nand U22736 (N_22736,N_15693,N_13250);
nand U22737 (N_22737,N_16562,N_13640);
and U22738 (N_22738,N_13329,N_13153);
nand U22739 (N_22739,N_19260,N_19432);
or U22740 (N_22740,N_15456,N_12484);
or U22741 (N_22741,N_11113,N_14680);
and U22742 (N_22742,N_11696,N_15147);
or U22743 (N_22743,N_12440,N_18682);
xor U22744 (N_22744,N_14512,N_14756);
xnor U22745 (N_22745,N_14789,N_11350);
nor U22746 (N_22746,N_13943,N_11817);
nand U22747 (N_22747,N_16168,N_10060);
or U22748 (N_22748,N_19724,N_17787);
nor U22749 (N_22749,N_13827,N_10179);
nor U22750 (N_22750,N_12171,N_12402);
nor U22751 (N_22751,N_10611,N_11115);
nor U22752 (N_22752,N_14511,N_16495);
and U22753 (N_22753,N_17825,N_11926);
and U22754 (N_22754,N_16659,N_19604);
and U22755 (N_22755,N_14170,N_17271);
nand U22756 (N_22756,N_16201,N_12549);
and U22757 (N_22757,N_12854,N_15181);
and U22758 (N_22758,N_13798,N_17260);
or U22759 (N_22759,N_16959,N_18480);
nor U22760 (N_22760,N_14950,N_18008);
nand U22761 (N_22761,N_10176,N_18232);
or U22762 (N_22762,N_16178,N_14614);
nor U22763 (N_22763,N_15353,N_11878);
or U22764 (N_22764,N_14501,N_16266);
xnor U22765 (N_22765,N_17555,N_16906);
nor U22766 (N_22766,N_15854,N_11358);
or U22767 (N_22767,N_13433,N_19827);
or U22768 (N_22768,N_11709,N_17890);
and U22769 (N_22769,N_12040,N_15625);
nand U22770 (N_22770,N_13533,N_18190);
and U22771 (N_22771,N_14500,N_10077);
or U22772 (N_22772,N_13956,N_13458);
xnor U22773 (N_22773,N_12946,N_15340);
and U22774 (N_22774,N_14104,N_18242);
nor U22775 (N_22775,N_14210,N_13363);
nor U22776 (N_22776,N_11981,N_11559);
nand U22777 (N_22777,N_19651,N_10862);
xnor U22778 (N_22778,N_10436,N_18690);
nor U22779 (N_22779,N_17488,N_19507);
or U22780 (N_22780,N_18596,N_13364);
nand U22781 (N_22781,N_13959,N_17413);
and U22782 (N_22782,N_17604,N_13788);
nor U22783 (N_22783,N_18994,N_15494);
or U22784 (N_22784,N_13564,N_17349);
xnor U22785 (N_22785,N_19097,N_17697);
and U22786 (N_22786,N_13617,N_18122);
nand U22787 (N_22787,N_18107,N_17265);
or U22788 (N_22788,N_18440,N_11486);
nor U22789 (N_22789,N_13428,N_13853);
or U22790 (N_22790,N_19901,N_15757);
or U22791 (N_22791,N_12670,N_16744);
xor U22792 (N_22792,N_15780,N_11666);
and U22793 (N_22793,N_15740,N_10575);
nor U22794 (N_22794,N_10524,N_11203);
nor U22795 (N_22795,N_14646,N_14958);
or U22796 (N_22796,N_17152,N_11776);
nand U22797 (N_22797,N_14838,N_14905);
nor U22798 (N_22798,N_12476,N_17978);
nor U22799 (N_22799,N_16452,N_19163);
nand U22800 (N_22800,N_12255,N_11984);
nor U22801 (N_22801,N_10479,N_10299);
and U22802 (N_22802,N_12655,N_12030);
nor U22803 (N_22803,N_11844,N_12310);
or U22804 (N_22804,N_18059,N_19961);
and U22805 (N_22805,N_18356,N_12668);
nand U22806 (N_22806,N_17440,N_13167);
nor U22807 (N_22807,N_11727,N_17669);
and U22808 (N_22808,N_13516,N_10769);
nor U22809 (N_22809,N_16102,N_12642);
or U22810 (N_22810,N_15404,N_17614);
or U22811 (N_22811,N_15219,N_12058);
or U22812 (N_22812,N_19528,N_16790);
nand U22813 (N_22813,N_17310,N_13578);
nor U22814 (N_22814,N_16612,N_18477);
and U22815 (N_22815,N_16036,N_13694);
nor U22816 (N_22816,N_13818,N_14567);
or U22817 (N_22817,N_17079,N_15959);
or U22818 (N_22818,N_12930,N_14399);
xor U22819 (N_22819,N_12829,N_15399);
nor U22820 (N_22820,N_13074,N_17220);
and U22821 (N_22821,N_12686,N_19506);
xor U22822 (N_22822,N_12296,N_19559);
nand U22823 (N_22823,N_14964,N_19540);
or U22824 (N_22824,N_11056,N_16480);
and U22825 (N_22825,N_12712,N_18321);
xor U22826 (N_22826,N_11185,N_16175);
xnor U22827 (N_22827,N_14631,N_19393);
or U22828 (N_22828,N_16916,N_19821);
nand U22829 (N_22829,N_17802,N_10218);
or U22830 (N_22830,N_15929,N_14055);
xor U22831 (N_22831,N_14110,N_18306);
nand U22832 (N_22832,N_15275,N_11457);
nor U22833 (N_22833,N_18469,N_18901);
nand U22834 (N_22834,N_13273,N_17912);
or U22835 (N_22835,N_19193,N_10099);
nor U22836 (N_22836,N_12844,N_11749);
nand U22837 (N_22837,N_19421,N_13230);
or U22838 (N_22838,N_11254,N_14534);
or U22839 (N_22839,N_11010,N_17996);
nor U22840 (N_22840,N_15590,N_10881);
xnor U22841 (N_22841,N_19965,N_15391);
xnor U22842 (N_22842,N_11880,N_10451);
nor U22843 (N_22843,N_19031,N_10875);
nor U22844 (N_22844,N_14710,N_17629);
and U22845 (N_22845,N_13769,N_12839);
nand U22846 (N_22846,N_14763,N_12745);
nor U22847 (N_22847,N_11902,N_16532);
nor U22848 (N_22848,N_17355,N_13828);
nor U22849 (N_22849,N_16693,N_11127);
nand U22850 (N_22850,N_18254,N_16601);
nor U22851 (N_22851,N_14118,N_13592);
nor U22852 (N_22852,N_15288,N_16586);
nand U22853 (N_22853,N_19305,N_19374);
nand U22854 (N_22854,N_15075,N_11289);
nor U22855 (N_22855,N_19812,N_14133);
and U22856 (N_22856,N_16679,N_19526);
and U22857 (N_22857,N_10866,N_13116);
nor U22858 (N_22858,N_13994,N_10990);
and U22859 (N_22859,N_17050,N_12615);
nor U22860 (N_22860,N_17417,N_13064);
or U22861 (N_22861,N_11422,N_10996);
nor U22862 (N_22862,N_15909,N_16584);
nor U22863 (N_22863,N_10075,N_11588);
nor U22864 (N_22864,N_15310,N_16269);
nand U22865 (N_22865,N_15992,N_17456);
and U22866 (N_22866,N_18323,N_17551);
xor U22867 (N_22867,N_10695,N_18680);
and U22868 (N_22868,N_12335,N_13274);
nand U22869 (N_22869,N_10204,N_10736);
or U22870 (N_22870,N_13974,N_13395);
and U22871 (N_22871,N_12109,N_12012);
nor U22872 (N_22872,N_15841,N_13009);
nand U22873 (N_22873,N_12359,N_19158);
nand U22874 (N_22874,N_15290,N_13468);
or U22875 (N_22875,N_11775,N_13948);
nand U22876 (N_22876,N_10850,N_17566);
and U22877 (N_22877,N_17869,N_12289);
xor U22878 (N_22878,N_11733,N_12798);
or U22879 (N_22879,N_16348,N_15174);
and U22880 (N_22880,N_13305,N_11053);
and U22881 (N_22881,N_11788,N_10115);
xor U22882 (N_22882,N_10332,N_11928);
nor U22883 (N_22883,N_17252,N_13745);
nand U22884 (N_22884,N_17241,N_17051);
or U22885 (N_22885,N_14024,N_19876);
xnor U22886 (N_22886,N_14818,N_13041);
xor U22887 (N_22887,N_10143,N_18896);
or U22888 (N_22888,N_14586,N_10852);
and U22889 (N_22889,N_19231,N_13454);
nand U22890 (N_22890,N_16683,N_17479);
or U22891 (N_22891,N_17412,N_10315);
nand U22892 (N_22892,N_18876,N_18003);
nor U22893 (N_22893,N_13872,N_14200);
and U22894 (N_22894,N_14264,N_10682);
nand U22895 (N_22895,N_15097,N_17687);
nor U22896 (N_22896,N_19485,N_16933);
nor U22897 (N_22897,N_18609,N_17056);
nor U22898 (N_22898,N_17716,N_10388);
nand U22899 (N_22899,N_19274,N_10599);
nor U22900 (N_22900,N_11821,N_18685);
or U22901 (N_22901,N_13735,N_16469);
nand U22902 (N_22902,N_14821,N_16101);
or U22903 (N_22903,N_14750,N_14705);
and U22904 (N_22904,N_15926,N_19215);
xnor U22905 (N_22905,N_15619,N_17462);
nor U22906 (N_22906,N_15643,N_14928);
or U22907 (N_22907,N_12363,N_13766);
xor U22908 (N_22908,N_15632,N_16218);
xor U22909 (N_22909,N_13772,N_13737);
or U22910 (N_22910,N_15347,N_13217);
nand U22911 (N_22911,N_11620,N_10069);
nand U22912 (N_22912,N_17477,N_17344);
and U22913 (N_22913,N_14669,N_14801);
or U22914 (N_22914,N_13875,N_19807);
or U22915 (N_22915,N_17375,N_18181);
xnor U22916 (N_22916,N_10257,N_15945);
or U22917 (N_22917,N_14525,N_18424);
and U22918 (N_22918,N_16514,N_16580);
nor U22919 (N_22919,N_13090,N_10375);
nand U22920 (N_22920,N_15405,N_16140);
or U22921 (N_22921,N_16209,N_17160);
nor U22922 (N_22922,N_14459,N_19324);
nor U22923 (N_22923,N_11507,N_15892);
nand U22924 (N_22924,N_13826,N_17556);
nand U22925 (N_22925,N_14575,N_15821);
or U22926 (N_22926,N_16536,N_10325);
nor U22927 (N_22927,N_14144,N_16594);
nor U22928 (N_22928,N_16278,N_16503);
or U22929 (N_22929,N_14366,N_13125);
and U22930 (N_22930,N_15951,N_10498);
or U22931 (N_22931,N_18397,N_11497);
nand U22932 (N_22932,N_16460,N_16506);
nor U22933 (N_22933,N_12198,N_13543);
xor U22934 (N_22934,N_19064,N_18369);
or U22935 (N_22935,N_15502,N_19711);
or U22936 (N_22936,N_17857,N_13079);
nor U22937 (N_22937,N_11139,N_19783);
or U22938 (N_22938,N_14989,N_11833);
nand U22939 (N_22939,N_15936,N_12366);
nand U22940 (N_22940,N_10205,N_12419);
nand U22941 (N_22941,N_15806,N_10602);
and U22942 (N_22942,N_17065,N_14257);
and U22943 (N_22943,N_17388,N_16327);
or U22944 (N_22944,N_11327,N_10811);
and U22945 (N_22945,N_13376,N_13427);
and U22946 (N_22946,N_14121,N_17737);
or U22947 (N_22947,N_12328,N_18372);
nor U22948 (N_22948,N_19918,N_19794);
and U22949 (N_22949,N_15381,N_19299);
nand U22950 (N_22950,N_19450,N_19112);
xnor U22951 (N_22951,N_11610,N_11236);
and U22952 (N_22952,N_15523,N_16058);
and U22953 (N_22953,N_16322,N_10020);
nor U22954 (N_22954,N_16118,N_13157);
xnor U22955 (N_22955,N_16072,N_15522);
or U22956 (N_22956,N_16481,N_15301);
nand U22957 (N_22957,N_13006,N_19014);
nor U22958 (N_22958,N_15999,N_13069);
nand U22959 (N_22959,N_17612,N_19736);
nand U22960 (N_22960,N_19224,N_12819);
nand U22961 (N_22961,N_19422,N_13389);
and U22962 (N_22962,N_14491,N_16976);
or U22963 (N_22963,N_14933,N_16339);
or U22964 (N_22964,N_12730,N_12068);
xor U22965 (N_22965,N_13120,N_10762);
or U22966 (N_22966,N_12405,N_16698);
and U22967 (N_22967,N_19200,N_15984);
nor U22968 (N_22968,N_19696,N_11939);
and U22969 (N_22969,N_15616,N_10641);
and U22970 (N_22970,N_11432,N_11637);
and U22971 (N_22971,N_14442,N_15541);
and U22972 (N_22972,N_14416,N_13414);
or U22973 (N_22973,N_13253,N_13422);
xnor U22974 (N_22974,N_12784,N_18843);
nor U22975 (N_22975,N_14808,N_19045);
nor U22976 (N_22976,N_11382,N_19247);
and U22977 (N_22977,N_15186,N_11975);
or U22978 (N_22978,N_11084,N_12500);
xnor U22979 (N_22979,N_17036,N_18038);
nand U22980 (N_22980,N_16538,N_15783);
or U22981 (N_22981,N_15830,N_11130);
or U22982 (N_22982,N_10132,N_18377);
nor U22983 (N_22983,N_18135,N_13147);
or U22984 (N_22984,N_18902,N_11266);
nor U22985 (N_22985,N_18834,N_13882);
and U22986 (N_22986,N_14618,N_16965);
and U22987 (N_22987,N_18937,N_17765);
nand U22988 (N_22988,N_12866,N_13880);
nor U22989 (N_22989,N_12083,N_13637);
and U22990 (N_22990,N_13514,N_11468);
and U22991 (N_22991,N_12753,N_15698);
nor U22992 (N_22992,N_17744,N_10028);
xor U22993 (N_22993,N_19929,N_19549);
nand U22994 (N_22994,N_11050,N_10631);
nor U22995 (N_22995,N_16943,N_19987);
nor U22996 (N_22996,N_18517,N_13623);
and U22997 (N_22997,N_12741,N_11882);
nor U22998 (N_22998,N_11342,N_12564);
or U22999 (N_22999,N_15845,N_14282);
or U23000 (N_23000,N_19448,N_10932);
or U23001 (N_23001,N_17658,N_13878);
nor U23002 (N_23002,N_13552,N_11396);
nor U23003 (N_23003,N_16803,N_11547);
or U23004 (N_23004,N_19699,N_16846);
and U23005 (N_23005,N_17514,N_10968);
or U23006 (N_23006,N_16663,N_12800);
nand U23007 (N_23007,N_11114,N_19365);
nand U23008 (N_23008,N_17650,N_14345);
xnor U23009 (N_23009,N_17184,N_10153);
nand U23010 (N_23010,N_19161,N_17733);
and U23011 (N_23011,N_10139,N_14953);
or U23012 (N_23012,N_16207,N_12221);
and U23013 (N_23013,N_13965,N_10796);
nand U23014 (N_23014,N_19881,N_16681);
or U23015 (N_23015,N_18560,N_19400);
nand U23016 (N_23016,N_16591,N_12512);
nand U23017 (N_23017,N_15443,N_19425);
and U23018 (N_23018,N_15145,N_13881);
nor U23019 (N_23019,N_18401,N_17968);
or U23020 (N_23020,N_12652,N_19201);
nand U23021 (N_23021,N_13770,N_18869);
nor U23022 (N_23022,N_19395,N_12050);
nor U23023 (N_23023,N_10091,N_19855);
nor U23024 (N_23024,N_13837,N_15889);
and U23025 (N_23025,N_19437,N_14047);
xor U23026 (N_23026,N_14604,N_16360);
nor U23027 (N_23027,N_19568,N_13864);
and U23028 (N_23028,N_11190,N_15903);
or U23029 (N_23029,N_18043,N_16981);
nor U23030 (N_23030,N_18506,N_18693);
and U23031 (N_23031,N_16754,N_15038);
or U23032 (N_23032,N_12871,N_16474);
and U23033 (N_23033,N_19585,N_13216);
nand U23034 (N_23034,N_10929,N_12749);
xor U23035 (N_23035,N_19456,N_12763);
nand U23036 (N_23036,N_10476,N_19034);
and U23037 (N_23037,N_17995,N_13259);
and U23038 (N_23038,N_12217,N_13109);
nor U23039 (N_23039,N_19928,N_18444);
or U23040 (N_23040,N_10804,N_10083);
nand U23041 (N_23041,N_19036,N_12131);
and U23042 (N_23042,N_18481,N_15283);
xor U23043 (N_23043,N_10972,N_10243);
nand U23044 (N_23044,N_11579,N_14911);
or U23045 (N_23045,N_10679,N_17212);
nand U23046 (N_23046,N_19550,N_16442);
nand U23047 (N_23047,N_15319,N_18307);
nor U23048 (N_23048,N_19344,N_12223);
and U23049 (N_23049,N_18276,N_15328);
nand U23050 (N_23050,N_10919,N_18052);
nor U23051 (N_23051,N_19600,N_14582);
and U23052 (N_23052,N_11160,N_14003);
xor U23053 (N_23053,N_17950,N_17291);
nand U23054 (N_23054,N_10984,N_17129);
and U23055 (N_23055,N_17525,N_18110);
nand U23056 (N_23056,N_15158,N_16367);
nand U23057 (N_23057,N_11818,N_13528);
and U23058 (N_23058,N_16097,N_15544);
and U23059 (N_23059,N_17976,N_19190);
nor U23060 (N_23060,N_17228,N_18927);
nor U23061 (N_23061,N_11043,N_14639);
and U23062 (N_23062,N_17781,N_11881);
nand U23063 (N_23063,N_12852,N_18280);
xnor U23064 (N_23064,N_19127,N_16333);
or U23065 (N_23065,N_17023,N_12412);
nand U23066 (N_23066,N_16707,N_10223);
or U23067 (N_23067,N_17337,N_15299);
nor U23068 (N_23068,N_17324,N_17969);
nand U23069 (N_23069,N_19379,N_12523);
and U23070 (N_23070,N_10356,N_17705);
and U23071 (N_23071,N_12010,N_19325);
nor U23072 (N_23072,N_12415,N_10339);
nand U23073 (N_23073,N_12578,N_13416);
or U23074 (N_23074,N_18941,N_16692);
or U23075 (N_23075,N_15769,N_12576);
and U23076 (N_23076,N_16811,N_16724);
or U23077 (N_23077,N_18539,N_19488);
and U23078 (N_23078,N_13930,N_15426);
and U23079 (N_23079,N_13050,N_14757);
nor U23080 (N_23080,N_14426,N_17097);
nand U23081 (N_23081,N_16799,N_15888);
nand U23082 (N_23082,N_14223,N_19518);
and U23083 (N_23083,N_10903,N_12660);
xnor U23084 (N_23084,N_14069,N_15566);
and U23085 (N_23085,N_17894,N_18384);
or U23086 (N_23086,N_15315,N_10424);
nand U23087 (N_23087,N_19244,N_17846);
nand U23088 (N_23088,N_12611,N_14610);
xor U23089 (N_23089,N_13037,N_11538);
and U23090 (N_23090,N_15349,N_14941);
nor U23091 (N_23091,N_19862,N_17192);
nor U23092 (N_23092,N_17942,N_18246);
or U23093 (N_23093,N_12463,N_12063);
nand U23094 (N_23094,N_15624,N_18088);
and U23095 (N_23095,N_18823,N_12553);
or U23096 (N_23096,N_19596,N_10156);
nor U23097 (N_23097,N_12638,N_17804);
or U23098 (N_23098,N_11137,N_19143);
nor U23099 (N_23099,N_14275,N_15699);
or U23100 (N_23100,N_16592,N_12640);
and U23101 (N_23101,N_16028,N_10777);
xor U23102 (N_23102,N_13384,N_13611);
and U23103 (N_23103,N_11615,N_18543);
nor U23104 (N_23104,N_10378,N_10888);
nor U23105 (N_23105,N_13227,N_18172);
xnor U23106 (N_23106,N_13131,N_14422);
or U23107 (N_23107,N_14188,N_16227);
xor U23108 (N_23108,N_11631,N_18147);
or U23109 (N_23109,N_13067,N_10515);
and U23110 (N_23110,N_17414,N_11399);
and U23111 (N_23111,N_16233,N_16678);
xor U23112 (N_23112,N_10320,N_12181);
nand U23113 (N_23113,N_18958,N_19273);
nor U23114 (N_23114,N_16860,N_12982);
or U23115 (N_23115,N_16973,N_14212);
nand U23116 (N_23116,N_17473,N_19766);
xor U23117 (N_23117,N_17476,N_10053);
and U23118 (N_23118,N_18727,N_17888);
and U23119 (N_23119,N_16387,N_18035);
and U23120 (N_23120,N_13841,N_17719);
nor U23121 (N_23121,N_19186,N_11347);
and U23122 (N_23122,N_16365,N_14214);
and U23123 (N_23123,N_16529,N_16093);
and U23124 (N_23124,N_18639,N_13565);
and U23125 (N_23125,N_14032,N_10429);
nor U23126 (N_23126,N_16648,N_10061);
nand U23127 (N_23127,N_18796,N_17831);
nor U23128 (N_23128,N_19355,N_13610);
nand U23129 (N_23129,N_19310,N_10293);
nand U23130 (N_23130,N_13418,N_18732);
or U23131 (N_23131,N_12339,N_12931);
or U23132 (N_23132,N_13471,N_16810);
nand U23133 (N_23133,N_10236,N_17298);
or U23134 (N_23134,N_17590,N_19203);
nand U23135 (N_23135,N_14006,N_11410);
or U23136 (N_23136,N_19836,N_17956);
nor U23137 (N_23137,N_14794,N_18844);
and U23138 (N_23138,N_19189,N_16624);
xnor U23139 (N_23139,N_10741,N_14938);
and U23140 (N_23140,N_10055,N_18054);
or U23141 (N_23141,N_18575,N_19810);
or U23142 (N_23142,N_15226,N_18385);
and U23143 (N_23143,N_16975,N_19666);
or U23144 (N_23144,N_11386,N_17362);
nand U23145 (N_23145,N_12695,N_10244);
or U23146 (N_23146,N_13548,N_15260);
nor U23147 (N_23147,N_10369,N_13215);
nand U23148 (N_23148,N_10116,N_10587);
and U23149 (N_23149,N_19793,N_10648);
and U23150 (N_23150,N_13899,N_12195);
nor U23151 (N_23151,N_13152,N_14096);
or U23152 (N_23152,N_11624,N_18767);
and U23153 (N_23153,N_15450,N_11825);
and U23154 (N_23154,N_11228,N_17382);
nor U23155 (N_23155,N_17312,N_16813);
nand U23156 (N_23156,N_14103,N_10902);
or U23157 (N_23157,N_10709,N_13589);
nand U23158 (N_23158,N_15253,N_18681);
nand U23159 (N_23159,N_16622,N_18997);
nor U23160 (N_23160,N_11995,N_12127);
or U23161 (N_23161,N_16519,N_17866);
and U23162 (N_23162,N_17405,N_16974);
or U23163 (N_23163,N_17099,N_15286);
nand U23164 (N_23164,N_10342,N_12203);
xnor U23165 (N_23165,N_17451,N_11509);
and U23166 (N_23166,N_19366,N_16473);
or U23167 (N_23167,N_12248,N_17360);
nand U23168 (N_23168,N_16795,N_14472);
nor U23169 (N_23169,N_18285,N_11921);
or U23170 (N_23170,N_18885,N_11802);
nor U23171 (N_23171,N_10940,N_12477);
nor U23172 (N_23172,N_18600,N_11894);
nor U23173 (N_23173,N_19835,N_17073);
or U23174 (N_23174,N_12909,N_12084);
nor U23175 (N_23175,N_18520,N_18121);
and U23176 (N_23176,N_16099,N_12059);
or U23177 (N_23177,N_11978,N_19860);
nor U23178 (N_23178,N_19091,N_16821);
or U23179 (N_23179,N_19153,N_11388);
nor U23180 (N_23180,N_19387,N_15463);
xnor U23181 (N_23181,N_10161,N_12052);
nor U23182 (N_23182,N_13519,N_14201);
nor U23183 (N_23183,N_12693,N_13968);
nor U23184 (N_23184,N_19635,N_19092);
and U23185 (N_23185,N_15599,N_15872);
xor U23186 (N_23186,N_14099,N_10595);
xor U23187 (N_23187,N_18071,N_13658);
or U23188 (N_23188,N_17828,N_15688);
nor U23189 (N_23189,N_19701,N_15671);
nor U23190 (N_23190,N_16126,N_16450);
and U23191 (N_23191,N_14531,N_16864);
nand U23192 (N_23192,N_13018,N_19068);
and U23193 (N_23193,N_17643,N_14289);
and U23194 (N_23194,N_14573,N_11779);
nor U23195 (N_23195,N_12469,N_17442);
and U23196 (N_23196,N_19461,N_15427);
nor U23197 (N_23197,N_17693,N_18895);
or U23198 (N_23198,N_15293,N_14889);
xnor U23199 (N_23199,N_13860,N_10542);
and U23200 (N_23200,N_14063,N_15816);
nor U23201 (N_23201,N_15526,N_16155);
nor U23202 (N_23202,N_14372,N_17584);
nor U23203 (N_23203,N_12128,N_13114);
or U23204 (N_23204,N_18737,N_10686);
or U23205 (N_23205,N_10539,N_10490);
nand U23206 (N_23206,N_15306,N_13522);
nor U23207 (N_23207,N_10774,N_16743);
nor U23208 (N_23208,N_18952,N_12994);
or U23209 (N_23209,N_17435,N_13424);
xor U23210 (N_23210,N_17537,N_17094);
nand U23211 (N_23211,N_19016,N_19723);
nand U23212 (N_23212,N_17307,N_14362);
or U23213 (N_23213,N_16213,N_12861);
nand U23214 (N_23214,N_10078,N_12551);
and U23215 (N_23215,N_13113,N_19078);
or U23216 (N_23216,N_12762,N_14198);
nand U23217 (N_23217,N_13081,N_14062);
xor U23218 (N_23218,N_14084,N_15997);
or U23219 (N_23219,N_12540,N_15062);
nand U23220 (N_23220,N_14997,N_19713);
xor U23221 (N_23221,N_14526,N_16851);
nand U23222 (N_23222,N_14581,N_17827);
nor U23223 (N_23223,N_11436,N_17975);
nand U23224 (N_23224,N_19982,N_10864);
nor U23225 (N_23225,N_17591,N_16982);
or U23226 (N_23226,N_10945,N_15254);
nand U23227 (N_23227,N_14077,N_18647);
or U23228 (N_23228,N_16915,N_12570);
and U23229 (N_23229,N_17234,N_14972);
and U23230 (N_23230,N_17470,N_18542);
and U23231 (N_23231,N_13636,N_14206);
or U23232 (N_23232,N_18624,N_12045);
and U23233 (N_23233,N_19811,N_11238);
nor U23234 (N_23234,N_12159,N_11059);
nor U23235 (N_23235,N_10114,N_19566);
nand U23236 (N_23236,N_14866,N_19782);
xor U23237 (N_23237,N_14779,N_19415);
nor U23238 (N_23238,N_14016,N_10047);
or U23239 (N_23239,N_14325,N_10962);
and U23240 (N_23240,N_10155,N_16808);
nand U23241 (N_23241,N_13001,N_18183);
nand U23242 (N_23242,N_13871,N_14400);
nand U23243 (N_23243,N_13483,N_13333);
and U23244 (N_23244,N_17347,N_16061);
nor U23245 (N_23245,N_14478,N_19763);
and U23246 (N_23246,N_11316,N_16238);
nand U23247 (N_23247,N_12519,N_12167);
xor U23248 (N_23248,N_13574,N_16620);
or U23249 (N_23249,N_15846,N_14691);
nand U23250 (N_23250,N_10916,N_13480);
nand U23251 (N_23251,N_15834,N_14781);
or U23252 (N_23252,N_19343,N_13561);
nor U23253 (N_23253,N_17284,N_18871);
nor U23254 (N_23254,N_15648,N_18364);
nor U23255 (N_23255,N_14026,N_11075);
nor U23256 (N_23256,N_11800,N_17367);
or U23257 (N_23257,N_13183,N_10448);
nand U23258 (N_23258,N_19886,N_13148);
and U23259 (N_23259,N_10861,N_19117);
or U23260 (N_23260,N_17528,N_15289);
or U23261 (N_23261,N_18839,N_10076);
or U23262 (N_23262,N_15525,N_17386);
and U23263 (N_23263,N_17338,N_14822);
and U23264 (N_23264,N_18334,N_11938);
nor U23265 (N_23265,N_18332,N_18814);
nor U23266 (N_23266,N_17431,N_17034);
and U23267 (N_23267,N_11060,N_14793);
xnor U23268 (N_23268,N_19690,N_17806);
nor U23269 (N_23269,N_18249,N_16349);
xor U23270 (N_23270,N_11251,N_18124);
or U23271 (N_23271,N_15799,N_19289);
nor U23272 (N_23272,N_19262,N_12096);
nor U23273 (N_23273,N_11481,N_16863);
nor U23274 (N_23274,N_10819,N_11405);
nand U23275 (N_23275,N_10642,N_12064);
xor U23276 (N_23276,N_14907,N_16978);
nand U23277 (N_23277,N_19854,N_10925);
or U23278 (N_23278,N_15716,N_12098);
and U23279 (N_23279,N_12448,N_17937);
nor U23280 (N_23280,N_11363,N_16389);
and U23281 (N_23281,N_18654,N_15464);
nor U23282 (N_23282,N_10857,N_10810);
or U23283 (N_23283,N_14812,N_18392);
or U23284 (N_23284,N_18445,N_13952);
or U23285 (N_23285,N_12995,N_12306);
nor U23286 (N_23286,N_15754,N_12425);
nand U23287 (N_23287,N_19029,N_19351);
nand U23288 (N_23288,N_16824,N_10756);
nor U23289 (N_23289,N_18675,N_18324);
nand U23290 (N_23290,N_17603,N_14589);
nand U23291 (N_23291,N_17837,N_10410);
and U23292 (N_23292,N_14894,N_16521);
and U23293 (N_23293,N_12441,N_15668);
xnor U23294 (N_23294,N_16655,N_11496);
nor U23295 (N_23295,N_17482,N_16722);
xnor U23296 (N_23296,N_17093,N_18866);
nand U23297 (N_23297,N_17348,N_18366);
nor U23298 (N_23298,N_19620,N_13917);
and U23299 (N_23299,N_16313,N_14128);
and U23300 (N_23300,N_18633,N_10384);
nand U23301 (N_23301,N_12968,N_16253);
or U23302 (N_23302,N_12265,N_18070);
xor U23303 (N_23303,N_19522,N_12963);
nor U23304 (N_23304,N_13432,N_13057);
or U23305 (N_23305,N_11493,N_15424);
nand U23306 (N_23306,N_11283,N_17021);
and U23307 (N_23307,N_11286,N_17169);
or U23308 (N_23308,N_17365,N_10026);
nor U23309 (N_23309,N_11475,N_16112);
or U23310 (N_23310,N_11403,N_13373);
and U23311 (N_23311,N_14108,N_17938);
nor U23312 (N_23312,N_14365,N_15333);
nand U23313 (N_23313,N_16552,N_16057);
nand U23314 (N_23314,N_11996,N_17588);
nand U23315 (N_23315,N_18393,N_16422);
and U23316 (N_23316,N_18112,N_12619);
nor U23317 (N_23317,N_11309,N_11214);
or U23318 (N_23318,N_11378,N_10959);
and U23319 (N_23319,N_13344,N_10183);
nor U23320 (N_23320,N_19981,N_16711);
nand U23321 (N_23321,N_14638,N_11086);
and U23322 (N_23322,N_12229,N_17426);
xnor U23323 (N_23323,N_12809,N_10222);
and U23324 (N_23324,N_17052,N_18094);
nand U23325 (N_23325,N_18196,N_12039);
xor U23326 (N_23326,N_11830,N_16195);
nor U23327 (N_23327,N_10965,N_16614);
xnor U23328 (N_23328,N_18116,N_12049);
xnor U23329 (N_23329,N_12118,N_13710);
and U23330 (N_23330,N_19954,N_15789);
and U23331 (N_23331,N_16940,N_15553);
or U23332 (N_23332,N_14357,N_13547);
or U23333 (N_23333,N_19682,N_10481);
or U23334 (N_23334,N_19940,N_11305);
nor U23335 (N_23335,N_18723,N_19634);
xor U23336 (N_23336,N_17505,N_18762);
nor U23337 (N_23337,N_10895,N_11858);
or U23338 (N_23338,N_17993,N_11847);
nand U23339 (N_23339,N_19212,N_10737);
nor U23340 (N_23340,N_11916,N_15223);
nand U23341 (N_23341,N_15104,N_16242);
nand U23342 (N_23342,N_12707,N_15304);
and U23343 (N_23343,N_17316,N_18857);
nand U23344 (N_23344,N_13538,N_12032);
xnor U23345 (N_23345,N_16400,N_11568);
nor U23346 (N_23346,N_18701,N_17074);
nor U23347 (N_23347,N_14482,N_11594);
or U23348 (N_23348,N_18917,N_11683);
nor U23349 (N_23349,N_17840,N_12214);
or U23350 (N_23350,N_19870,N_19026);
nor U23351 (N_23351,N_10813,N_12811);
and U23352 (N_23352,N_10324,N_12612);
xor U23353 (N_23353,N_19911,N_14260);
and U23354 (N_23354,N_11520,N_10582);
nor U23355 (N_23355,N_18312,N_16919);
and U23356 (N_23356,N_14782,N_11232);
xor U23357 (N_23357,N_15162,N_15630);
and U23358 (N_23358,N_14394,N_10617);
nand U23359 (N_23359,N_19281,N_14455);
nand U23360 (N_23360,N_13419,N_15822);
nand U23361 (N_23361,N_14820,N_13705);
or U23362 (N_23362,N_12044,N_12447);
nor U23363 (N_23363,N_16345,N_18406);
or U23364 (N_23364,N_18890,N_16429);
nand U23365 (N_23365,N_17105,N_15006);
or U23366 (N_23366,N_19641,N_19771);
or U23367 (N_23367,N_18478,N_17246);
nor U23368 (N_23368,N_15825,N_17118);
or U23369 (N_23369,N_13739,N_15569);
xnor U23370 (N_23370,N_18810,N_13330);
and U23371 (N_23371,N_15532,N_18301);
and U23372 (N_23372,N_15397,N_15781);
nand U23373 (N_23373,N_12161,N_14920);
xor U23374 (N_23374,N_17902,N_17814);
and U23375 (N_23375,N_18404,N_16920);
and U23376 (N_23376,N_17402,N_17526);
nor U23377 (N_23377,N_17511,N_11246);
and U23378 (N_23378,N_11628,N_12315);
or U23379 (N_23379,N_19639,N_17441);
nor U23380 (N_23380,N_10954,N_17210);
and U23381 (N_23381,N_14123,N_12881);
nor U23382 (N_23382,N_19116,N_19730);
xnor U23383 (N_23383,N_16016,N_13306);
nor U23384 (N_23384,N_11000,N_15126);
nor U23385 (N_23385,N_15782,N_15316);
or U23386 (N_23386,N_18683,N_16664);
or U23387 (N_23387,N_19157,N_10594);
or U23388 (N_23388,N_12224,N_15596);
and U23389 (N_23389,N_15886,N_17236);
and U23390 (N_23390,N_11265,N_17822);
nor U23391 (N_23391,N_16412,N_13958);
nand U23392 (N_23392,N_11216,N_12295);
and U23393 (N_23393,N_15025,N_18311);
and U23394 (N_23394,N_14729,N_14162);
and U23395 (N_23395,N_13570,N_15080);
or U23396 (N_23396,N_19797,N_18545);
xor U23397 (N_23397,N_14758,N_13206);
xnor U23398 (N_23398,N_17871,N_16645);
nor U23399 (N_23399,N_14092,N_19385);
or U23400 (N_23400,N_10948,N_13055);
and U23401 (N_23401,N_15087,N_15134);
nand U23402 (N_23402,N_10037,N_12216);
and U23403 (N_23403,N_16812,N_15955);
or U23404 (N_23404,N_15454,N_11565);
xnor U23405 (N_23405,N_19991,N_11519);
and U23406 (N_23406,N_12054,N_17249);
nand U23407 (N_23407,N_19733,N_10835);
nand U23408 (N_23408,N_15034,N_11262);
nor U23409 (N_23409,N_12142,N_17407);
and U23410 (N_23410,N_16444,N_15144);
and U23411 (N_23411,N_11835,N_17513);
and U23412 (N_23412,N_16022,N_15418);
or U23413 (N_23413,N_15719,N_10269);
or U23414 (N_23414,N_10208,N_16553);
nor U23415 (N_23415,N_17636,N_17214);
nand U23416 (N_23416,N_12367,N_11958);
or U23417 (N_23417,N_18277,N_13451);
nand U23418 (N_23418,N_18390,N_13712);
nor U23419 (N_23419,N_18588,N_19976);
nor U23420 (N_23420,N_17653,N_11544);
nand U23421 (N_23421,N_14528,N_19882);
xor U23422 (N_23422,N_16396,N_17217);
or U23423 (N_23423,N_16273,N_18879);
nand U23424 (N_23424,N_11100,N_18819);
nand U23425 (N_23425,N_13951,N_10426);
nor U23426 (N_23426,N_12899,N_17114);
and U23427 (N_23427,N_17684,N_10449);
nand U23428 (N_23428,N_12787,N_14563);
and U23429 (N_23429,N_16287,N_12739);
nor U23430 (N_23430,N_11488,N_19108);
nor U23431 (N_23431,N_14145,N_13296);
nor U23432 (N_23432,N_11479,N_14129);
nand U23433 (N_23433,N_15881,N_16423);
nand U23434 (N_23434,N_15920,N_18447);
or U23435 (N_23435,N_16735,N_13278);
or U23436 (N_23436,N_11042,N_19182);
xnor U23437 (N_23437,N_16556,N_13746);
and U23438 (N_23438,N_17731,N_15582);
nor U23439 (N_23439,N_17702,N_13885);
nand U23440 (N_23440,N_13127,N_17929);
and U23441 (N_23441,N_15193,N_14311);
nor U23442 (N_23442,N_14900,N_15987);
and U23443 (N_23443,N_14079,N_15152);
nor U23444 (N_23444,N_15413,N_18303);
and U23445 (N_23445,N_10708,N_19554);
nand U23446 (N_23446,N_11698,N_15584);
or U23447 (N_23447,N_15455,N_15918);
xor U23448 (N_23448,N_19490,N_13493);
nor U23449 (N_23449,N_10354,N_10500);
and U23450 (N_23450,N_17530,N_10018);
nor U23451 (N_23451,N_11842,N_13506);
or U23452 (N_23452,N_15709,N_19892);
nor U23453 (N_23453,N_13252,N_15506);
xor U23454 (N_23454,N_13749,N_18367);
xnor U23455 (N_23455,N_12352,N_13729);
nor U23456 (N_23456,N_16399,N_17240);
and U23457 (N_23457,N_12120,N_19100);
nor U23458 (N_23458,N_11271,N_18082);
and U23459 (N_23459,N_14120,N_11782);
and U23460 (N_23460,N_12563,N_19371);
nor U23461 (N_23461,N_12398,N_11785);
and U23462 (N_23462,N_15656,N_13597);
nor U23463 (N_23463,N_11558,N_19937);
nand U23464 (N_23464,N_12562,N_13789);
nor U23465 (N_23465,N_19752,N_18889);
or U23466 (N_23466,N_16682,N_13747);
or U23467 (N_23467,N_13134,N_16251);
and U23468 (N_23468,N_17132,N_18777);
nor U23469 (N_23469,N_14050,N_13497);
nand U23470 (N_23470,N_14100,N_16855);
nand U23471 (N_23471,N_15510,N_14685);
nor U23472 (N_23472,N_16773,N_12017);
nor U23473 (N_23473,N_16357,N_12954);
xor U23474 (N_23474,N_16674,N_13781);
nor U23475 (N_23475,N_15713,N_14968);
or U23476 (N_23476,N_14246,N_17965);
and U23477 (N_23477,N_10494,N_19113);
or U23478 (N_23478,N_14087,N_15689);
nor U23479 (N_23479,N_16867,N_12140);
nor U23480 (N_23480,N_16402,N_10331);
or U23481 (N_23481,N_18613,N_10364);
nor U23482 (N_23482,N_12786,N_11027);
nand U23483 (N_23483,N_18772,N_11447);
nor U23484 (N_23484,N_12386,N_10129);
xor U23485 (N_23485,N_13488,N_19538);
or U23486 (N_23486,N_17029,N_11780);
or U23487 (N_23487,N_19608,N_12106);
nand U23488 (N_23488,N_11485,N_16302);
or U23489 (N_23489,N_13980,N_15472);
or U23490 (N_23490,N_10358,N_10482);
or U23491 (N_23491,N_19022,N_12365);
and U23492 (N_23492,N_11349,N_13232);
nor U23493 (N_23493,N_19545,N_16031);
or U23494 (N_23494,N_16465,N_19557);
and U23495 (N_23495,N_13587,N_10546);
nand U23496 (N_23496,N_10657,N_15941);
nor U23497 (N_23497,N_11174,N_14488);
and U23498 (N_23498,N_12895,N_16897);
xnor U23499 (N_23499,N_14412,N_14310);
nor U23500 (N_23500,N_14355,N_14713);
and U23501 (N_23501,N_14379,N_17703);
and U23502 (N_23502,N_11207,N_18315);
or U23503 (N_23503,N_17834,N_17380);
xnor U23504 (N_23504,N_10722,N_11212);
nor U23505 (N_23505,N_14774,N_11296);
nor U23506 (N_23506,N_12003,N_10808);
nand U23507 (N_23507,N_10467,N_14695);
nand U23508 (N_23508,N_13501,N_12831);
xor U23509 (N_23509,N_17997,N_15043);
nor U23510 (N_23510,N_10158,N_17934);
nor U23511 (N_23511,N_17582,N_19837);
or U23512 (N_23512,N_17356,N_13891);
and U23513 (N_23513,N_11619,N_13043);
nor U23514 (N_23514,N_19059,N_19899);
nand U23515 (N_23515,N_14529,N_14593);
nor U23516 (N_23516,N_11464,N_11429);
nand U23517 (N_23517,N_12048,N_16996);
and U23518 (N_23518,N_13495,N_18302);
xnor U23519 (N_23519,N_11890,N_10407);
or U23520 (N_23520,N_17550,N_19346);
nand U23521 (N_23521,N_13332,N_18251);
nand U23522 (N_23522,N_12178,N_13038);
nand U23523 (N_23523,N_17138,N_17452);
or U23524 (N_23524,N_12094,N_19248);
nand U23525 (N_23525,N_15976,N_11276);
or U23526 (N_23526,N_17448,N_19845);
nand U23527 (N_23527,N_12938,N_11609);
xor U23528 (N_23528,N_16837,N_19508);
nor U23529 (N_23529,N_19665,N_13759);
or U23530 (N_23530,N_17317,N_17953);
or U23531 (N_23531,N_10267,N_17946);
nor U23532 (N_23532,N_12773,N_11444);
or U23533 (N_23533,N_12882,N_19891);
nor U23534 (N_23534,N_14227,N_13382);
and U23535 (N_23535,N_13076,N_11482);
xnor U23536 (N_23536,N_12088,N_14370);
nand U23537 (N_23537,N_13846,N_10685);
and U23538 (N_23538,N_14769,N_19706);
nor U23539 (N_23539,N_19101,N_15602);
or U23540 (N_23540,N_18554,N_17418);
and U23541 (N_23541,N_19443,N_15264);
xnor U23542 (N_23542,N_15201,N_12720);
nand U23543 (N_23543,N_18874,N_10308);
or U23544 (N_23544,N_19148,N_12433);
or U23545 (N_23545,N_13590,N_13400);
nor U23546 (N_23546,N_18317,N_17855);
xnor U23547 (N_23547,N_17159,N_15350);
or U23548 (N_23548,N_18026,N_13542);
or U23549 (N_23549,N_13671,N_10096);
nand U23550 (N_23550,N_11222,N_12883);
xor U23551 (N_23551,N_17691,N_18064);
and U23552 (N_23552,N_18245,N_14912);
nor U23553 (N_23553,N_11240,N_16661);
nand U23554 (N_23554,N_18069,N_13583);
xnor U23555 (N_23555,N_12736,N_17172);
nor U23556 (N_23556,N_15710,N_18697);
and U23557 (N_23557,N_10772,N_13361);
or U23558 (N_23558,N_10338,N_17471);
and U23559 (N_23559,N_17914,N_17954);
nand U23560 (N_23560,N_16700,N_11592);
nor U23561 (N_23561,N_17941,N_18699);
nor U23562 (N_23562,N_10924,N_11200);
nand U23563 (N_23563,N_11025,N_19598);
nor U23564 (N_23564,N_12205,N_13179);
nor U23565 (N_23565,N_15488,N_19065);
nor U23566 (N_23566,N_19974,N_18750);
or U23567 (N_23567,N_12238,N_15074);
nor U23568 (N_23568,N_15312,N_12631);
nor U23569 (N_23569,N_14373,N_10523);
xor U23570 (N_23570,N_13914,N_14252);
nand U23571 (N_23571,N_13928,N_18171);
nor U23572 (N_23572,N_16967,N_13342);
and U23573 (N_23573,N_19926,N_17107);
and U23574 (N_23574,N_12591,N_16954);
or U23575 (N_23575,N_11397,N_12663);
or U23576 (N_23576,N_11642,N_15965);
nor U23577 (N_23577,N_11567,N_18150);
nand U23578 (N_23578,N_17411,N_17444);
nor U23579 (N_23579,N_19019,N_11047);
or U23580 (N_23580,N_15094,N_17845);
and U23581 (N_23581,N_12751,N_13101);
nand U23582 (N_23582,N_13797,N_17227);
or U23583 (N_23583,N_10987,N_15303);
nor U23584 (N_23584,N_18744,N_12706);
and U23585 (N_23585,N_15591,N_10276);
nand U23586 (N_23586,N_19525,N_16829);
or U23587 (N_23587,N_16727,N_11636);
and U23588 (N_23588,N_17014,N_16613);
and U23589 (N_23589,N_18657,N_13683);
nor U23590 (N_23590,N_15759,N_16046);
and U23591 (N_23591,N_19599,N_18261);
and U23592 (N_23592,N_11908,N_17485);
nor U23593 (N_23593,N_16170,N_14281);
xor U23594 (N_23594,N_19721,N_17398);
and U23595 (N_23595,N_19497,N_15896);
and U23596 (N_23596,N_11912,N_10720);
xor U23597 (N_23597,N_12989,N_12108);
or U23598 (N_23598,N_10918,N_10849);
nor U23599 (N_23599,N_12138,N_14977);
or U23600 (N_23600,N_15345,N_14558);
xor U23601 (N_23601,N_11004,N_11062);
or U23602 (N_23602,N_12933,N_19194);
nor U23603 (N_23603,N_11473,N_13991);
xnor U23604 (N_23604,N_17491,N_10296);
or U23605 (N_23605,N_11451,N_13778);
or U23606 (N_23606,N_12251,N_15078);
or U23607 (N_23607,N_11465,N_19438);
nor U23608 (N_23608,N_11690,N_13307);
nor U23609 (N_23609,N_16257,N_19859);
or U23610 (N_23610,N_13464,N_19513);
nor U23611 (N_23611,N_18916,N_13879);
and U23612 (N_23612,N_16369,N_19172);
and U23613 (N_23613,N_14402,N_15408);
nor U23614 (N_23614,N_15150,N_18546);
nand U23615 (N_23615,N_13813,N_10247);
nand U23616 (N_23616,N_17031,N_15005);
or U23617 (N_23617,N_15606,N_18706);
nor U23618 (N_23618,N_10133,N_11964);
or U23619 (N_23619,N_13399,N_12897);
or U23620 (N_23620,N_10824,N_15346);
nor U23621 (N_23621,N_19809,N_18645);
nand U23622 (N_23622,N_13982,N_12263);
and U23623 (N_23623,N_18166,N_14888);
or U23624 (N_23624,N_17489,N_16499);
and U23625 (N_23625,N_19533,N_15476);
nand U23626 (N_23626,N_17531,N_11260);
and U23627 (N_23627,N_12253,N_18187);
or U23628 (N_23628,N_15681,N_14452);
nand U23629 (N_23629,N_12271,N_12731);
nand U23630 (N_23630,N_12311,N_11241);
nand U23631 (N_23631,N_15733,N_13725);
and U23632 (N_23632,N_10912,N_10876);
xnor U23633 (N_23633,N_16725,N_19897);
nand U23634 (N_23634,N_14435,N_14343);
xnor U23635 (N_23635,N_14541,N_13474);
and U23636 (N_23636,N_15423,N_17977);
nor U23637 (N_23637,N_18340,N_14440);
and U23638 (N_23638,N_19654,N_12340);
xnor U23639 (N_23639,N_10787,N_10882);
or U23640 (N_23640,N_16050,N_14395);
nand U23641 (N_23641,N_17585,N_19616);
and U23642 (N_23642,N_14415,N_18803);
xnor U23643 (N_23643,N_19077,N_19967);
nand U23644 (N_23644,N_12153,N_11770);
and U23645 (N_23645,N_16827,N_18140);
nor U23646 (N_23646,N_16027,N_13626);
or U23647 (N_23647,N_13939,N_14859);
nor U23648 (N_23648,N_16989,N_19335);
nor U23649 (N_23649,N_15857,N_13721);
or U23650 (N_23650,N_17829,N_12802);
nor U23651 (N_23651,N_11145,N_15887);
or U23652 (N_23652,N_16758,N_18271);
and U23653 (N_23653,N_18944,N_11390);
or U23654 (N_23654,N_19850,N_19327);
and U23655 (N_23655,N_16882,N_18345);
and U23656 (N_23656,N_14242,N_19128);
nor U23657 (N_23657,N_10178,N_15776);
nor U23658 (N_23658,N_18057,N_12391);
xnor U23659 (N_23659,N_14904,N_16868);
or U23660 (N_23660,N_11551,N_12539);
or U23661 (N_23661,N_17713,N_17237);
nand U23662 (N_23662,N_11685,N_17054);
or U23663 (N_23663,N_18375,N_10995);
or U23664 (N_23664,N_13286,N_16757);
nand U23665 (N_23665,N_16007,N_12629);
nand U23666 (N_23666,N_18687,N_10191);
and U23667 (N_23667,N_15547,N_16723);
nand U23668 (N_23668,N_16878,N_10357);
or U23669 (N_23669,N_18048,N_15967);
nand U23670 (N_23670,N_10478,N_15068);
and U23671 (N_23671,N_12090,N_12662);
and U23672 (N_23672,N_14010,N_15369);
nand U23673 (N_23673,N_12673,N_10822);
or U23674 (N_23674,N_10637,N_12552);
and U23675 (N_23675,N_10414,N_10215);
xor U23676 (N_23676,N_18125,N_17351);
or U23677 (N_23677,N_12689,N_10353);
or U23678 (N_23678,N_17635,N_14924);
or U23679 (N_23679,N_16108,N_18456);
or U23680 (N_23680,N_10803,N_16839);
nand U23681 (N_23681,N_18793,N_17791);
and U23682 (N_23682,N_17560,N_17913);
and U23683 (N_23683,N_11351,N_14711);
or U23684 (N_23684,N_13118,N_13581);
xor U23685 (N_23685,N_17760,N_14809);
nor U23686 (N_23686,N_10282,N_16131);
or U23687 (N_23687,N_18712,N_13608);
nor U23688 (N_23688,N_11333,N_10292);
nor U23689 (N_23689,N_13089,N_10993);
nand U23690 (N_23690,N_16719,N_18620);
xnor U23691 (N_23691,N_17370,N_16922);
nand U23692 (N_23692,N_15505,N_16216);
nand U23693 (N_23693,N_18797,N_13555);
or U23694 (N_23694,N_19301,N_12406);
nand U23695 (N_23695,N_12185,N_16358);
or U23696 (N_23696,N_12651,N_15236);
nand U23697 (N_23697,N_12560,N_18316);
nand U23698 (N_23698,N_13539,N_11182);
nand U23699 (N_23699,N_12850,N_19154);
nor U23700 (N_23700,N_15812,N_16403);
or U23701 (N_23701,N_10043,N_12027);
nand U23702 (N_23702,N_14444,N_15081);
and U23703 (N_23703,N_10558,N_12855);
nor U23704 (N_23704,N_17224,N_19491);
and U23705 (N_23705,N_17819,N_15763);
nor U23706 (N_23706,N_15633,N_10371);
and U23707 (N_23707,N_11607,N_19233);
or U23708 (N_23708,N_15554,N_16820);
nor U23709 (N_23709,N_19146,N_17045);
or U23710 (N_23710,N_10952,N_15645);
xor U23711 (N_23711,N_12864,N_18262);
nand U23712 (N_23712,N_19264,N_13911);
and U23713 (N_23713,N_14777,N_19632);
and U23714 (N_23714,N_14284,N_18533);
nand U23715 (N_23715,N_14612,N_11741);
nand U23716 (N_23716,N_18360,N_19210);
nor U23717 (N_23717,N_13267,N_13294);
nor U23718 (N_23718,N_12976,N_11159);
and U23719 (N_23719,N_11692,N_19875);
or U23720 (N_23720,N_11549,N_10588);
and U23721 (N_23721,N_15215,N_11131);
and U23722 (N_23722,N_16109,N_17826);
and U23723 (N_23723,N_15572,N_14367);
nor U23724 (N_23724,N_18763,N_16710);
and U23725 (N_23725,N_18118,N_17574);
nand U23726 (N_23726,N_16565,N_12606);
nor U23727 (N_23727,N_19136,N_11900);
nor U23728 (N_23728,N_12928,N_18612);
and U23729 (N_23729,N_14391,N_14385);
nand U23730 (N_23730,N_13614,N_17044);
nor U23731 (N_23731,N_10250,N_10521);
nand U23732 (N_23732,N_11874,N_10789);
or U23733 (N_23733,N_10337,N_12700);
nor U23734 (N_23734,N_15191,N_19394);
nand U23735 (N_23735,N_16189,N_19095);
and U23736 (N_23736,N_17383,N_16137);
xnor U23737 (N_23737,N_16753,N_14903);
or U23738 (N_23738,N_17563,N_11116);
nor U23739 (N_23739,N_18746,N_17564);
nand U23740 (N_23740,N_18534,N_12847);
nor U23741 (N_23741,N_12679,N_12332);
nor U23742 (N_23742,N_14716,N_13024);
nand U23743 (N_23743,N_18438,N_12728);
or U23744 (N_23744,N_14401,N_13649);
or U23745 (N_23745,N_14732,N_17873);
and U23746 (N_23746,N_17313,N_12999);
nor U23747 (N_23747,N_18089,N_10160);
nand U23748 (N_23748,N_19451,N_18047);
and U23749 (N_23749,N_13962,N_10398);
and U23750 (N_23750,N_16479,N_12568);
nand U23751 (N_23751,N_17880,N_13852);
nor U23752 (N_23752,N_18389,N_14988);
nor U23753 (N_23753,N_13762,N_18665);
nor U23754 (N_23754,N_19313,N_19861);
and U23755 (N_23755,N_18641,N_10606);
nand U23756 (N_23756,N_11412,N_11961);
xor U23757 (N_23757,N_11301,N_12007);
nand U23758 (N_23758,N_15273,N_15546);
or U23759 (N_23759,N_14565,N_19228);
nor U23760 (N_23760,N_11674,N_16439);
and U23761 (N_23761,N_13908,N_18159);
nor U23762 (N_23762,N_18337,N_14384);
and U23763 (N_23763,N_17664,N_17251);
or U23764 (N_23764,N_10718,N_16014);
or U23765 (N_23765,N_12815,N_18273);
nand U23766 (N_23766,N_18971,N_12978);
xnor U23767 (N_23767,N_11118,N_16603);
nor U23768 (N_23768,N_15990,N_16401);
xnor U23769 (N_23769,N_14322,N_14557);
nor U23770 (N_23770,N_10240,N_13652);
and U23771 (N_23771,N_17849,N_16284);
and U23772 (N_23772,N_10985,N_19053);
nor U23773 (N_23773,N_10660,N_14813);
nor U23774 (N_23774,N_19410,N_15902);
xnor U23775 (N_23775,N_17695,N_19339);
xnor U23776 (N_23776,N_17300,N_12330);
and U23777 (N_23777,N_11463,N_10032);
xor U23778 (N_23778,N_19083,N_15416);
nand U23779 (N_23779,N_18040,N_18428);
and U23780 (N_23780,N_15875,N_15106);
or U23781 (N_23781,N_16852,N_10110);
and U23782 (N_23782,N_17816,N_16217);
or U23783 (N_23783,N_19523,N_14148);
nand U23784 (N_23784,N_17455,N_13372);
and U23785 (N_23785,N_17290,N_16963);
nor U23786 (N_23786,N_16498,N_16930);
nand U23787 (N_23787,N_17867,N_15308);
and U23788 (N_23788,N_13512,N_14436);
or U23789 (N_23789,N_10530,N_16845);
or U23790 (N_23790,N_16018,N_13687);
nor U23791 (N_23791,N_16703,N_11066);
and U23792 (N_23792,N_18610,N_10889);
nor U23793 (N_23793,N_15863,N_17742);
nand U23794 (N_23794,N_10392,N_13954);
nor U23795 (N_23795,N_10645,N_15499);
and U23796 (N_23796,N_11717,N_14899);
nor U23797 (N_23797,N_18694,N_13946);
or U23798 (N_23798,N_15014,N_11270);
or U23799 (N_23799,N_18161,N_12659);
nor U23800 (N_23800,N_19445,N_14955);
nand U23801 (N_23801,N_10759,N_12014);
nor U23802 (N_23802,N_11616,N_14179);
and U23803 (N_23803,N_11987,N_17120);
and U23804 (N_23804,N_12113,N_15053);
and U23805 (N_23805,N_13191,N_19848);
or U23806 (N_23806,N_18653,N_13509);
nor U23807 (N_23807,N_11093,N_13187);
nand U23808 (N_23808,N_18559,N_11982);
and U23809 (N_23809,N_18267,N_15233);
nor U23810 (N_23810,N_12302,N_16891);
and U23811 (N_23811,N_11991,N_16699);
and U23812 (N_23812,N_17838,N_13358);
nand U23813 (N_23813,N_11714,N_12580);
nor U23814 (N_23814,N_17554,N_16575);
or U23815 (N_23815,N_14037,N_16925);
or U23816 (N_23816,N_17749,N_12313);
nor U23817 (N_23817,N_16800,N_17725);
nand U23818 (N_23818,N_10294,N_10776);
or U23819 (N_23819,N_18979,N_19056);
nand U23820 (N_23820,N_14902,N_18512);
nand U23821 (N_23821,N_13503,N_13020);
and U23822 (N_23822,N_15512,N_18599);
and U23823 (N_23823,N_11248,N_19530);
or U23824 (N_23824,N_12414,N_19138);
or U23825 (N_23825,N_13208,N_16909);
or U23826 (N_23826,N_14965,N_19541);
xnor U23827 (N_23827,N_12004,N_11865);
or U23828 (N_23828,N_13890,N_12680);
and U23829 (N_23829,N_12303,N_10654);
xor U23830 (N_23830,N_18765,N_14233);
nor U23831 (N_23831,N_13031,N_14667);
and U23832 (N_23832,N_18498,N_13782);
xor U23833 (N_23833,N_16115,N_12834);
xor U23834 (N_23834,N_13443,N_10477);
nor U23835 (N_23835,N_15598,N_15182);
or U23836 (N_23836,N_19921,N_10790);
nor U23837 (N_23837,N_10877,N_18868);
nor U23838 (N_23838,N_12258,N_14411);
xor U23839 (N_23839,N_11597,N_10140);
or U23840 (N_23840,N_14390,N_11761);
nand U23841 (N_23841,N_12572,N_17876);
nor U23842 (N_23842,N_14682,N_19110);
nor U23843 (N_23843,N_17931,N_19337);
nor U23844 (N_23844,N_17651,N_15950);
and U23845 (N_23845,N_10113,N_11196);
nor U23846 (N_23846,N_16068,N_17474);
or U23847 (N_23847,N_19978,N_17278);
and U23848 (N_23848,N_10750,N_18698);
nor U23849 (N_23849,N_17102,N_12314);
or U23850 (N_23850,N_18695,N_11645);
nand U23851 (N_23851,N_17285,N_11896);
nand U23852 (N_23852,N_10279,N_17436);
and U23853 (N_23853,N_19202,N_17536);
nand U23854 (N_23854,N_18663,N_15327);
nor U23855 (N_23855,N_14009,N_13058);
or U23856 (N_23856,N_12464,N_12207);
and U23857 (N_23857,N_19630,N_12097);
nand U23858 (N_23858,N_16652,N_14773);
or U23859 (N_23859,N_14982,N_19222);
nor U23860 (N_23860,N_16011,N_17779);
xor U23861 (N_23861,N_11452,N_10141);
or U23862 (N_23862,N_11424,N_19789);
xor U23863 (N_23863,N_19970,N_19013);
and U23864 (N_23864,N_10189,N_16626);
or U23865 (N_23865,N_14410,N_16410);
or U23866 (N_23866,N_19962,N_16767);
or U23867 (N_23867,N_13017,N_18524);
or U23868 (N_23868,N_14653,N_15351);
nor U23869 (N_23869,N_17239,N_17164);
and U23870 (N_23870,N_18464,N_11811);
nand U23871 (N_23871,N_15377,N_16340);
and U23872 (N_23872,N_15238,N_17175);
nand U23873 (N_23873,N_14658,N_18640);
and U23874 (N_23874,N_15994,N_13141);
and U23875 (N_23875,N_12317,N_16008);
nand U23876 (N_23876,N_15700,N_18565);
nand U23877 (N_23877,N_12426,N_15056);
or U23878 (N_23878,N_10680,N_19040);
or U23879 (N_23879,N_14690,N_17671);
nor U23880 (N_23880,N_15481,N_18899);
or U23881 (N_23881,N_15853,N_11869);
and U23882 (N_23882,N_13621,N_15112);
nor U23883 (N_23883,N_12682,N_10072);
and U23884 (N_23884,N_17863,N_13754);
xor U23885 (N_23885,N_16325,N_17201);
nor U23886 (N_23886,N_15242,N_15737);
nor U23887 (N_23887,N_17542,N_16315);
nor U23888 (N_23888,N_16138,N_13000);
or U23889 (N_23889,N_16263,N_12903);
xnor U23890 (N_23890,N_16105,N_17988);
and U23891 (N_23891,N_12846,N_19681);
or U23892 (N_23892,N_14507,N_18811);
nor U23893 (N_23893,N_11032,N_18541);
or U23894 (N_23894,N_15794,N_10352);
nor U23895 (N_23895,N_18849,N_14151);
or U23896 (N_23896,N_19185,N_17145);
nand U23897 (N_23897,N_17498,N_19813);
or U23898 (N_23898,N_11345,N_18238);
and U23899 (N_23899,N_17789,N_18998);
nor U23900 (N_23900,N_11577,N_10758);
and U23901 (N_23901,N_16561,N_19184);
xor U23902 (N_23902,N_17841,N_16464);
or U23903 (N_23903,N_13709,N_14211);
nor U23904 (N_23904,N_18920,N_12768);
or U23905 (N_23905,N_17320,N_12698);
and U23906 (N_23906,N_15509,N_14237);
and U23907 (N_23907,N_18033,N_14409);
nor U23908 (N_23908,N_19644,N_12672);
nand U23909 (N_23909,N_10557,N_14735);
and U23910 (N_23910,N_18515,N_11856);
nand U23911 (N_23911,N_15962,N_19597);
or U23912 (N_23912,N_15750,N_17009);
nand U23913 (N_23913,N_13198,N_17803);
and U23914 (N_23914,N_15177,N_15040);
or U23915 (N_23915,N_12806,N_13638);
nand U23916 (N_23916,N_14033,N_18676);
nand U23917 (N_23917,N_14694,N_15969);
or U23918 (N_23918,N_14873,N_19985);
nor U23919 (N_23919,N_18119,N_10209);
and U23920 (N_23920,N_12103,N_17415);
nand U23921 (N_23921,N_17805,N_19669);
xnor U23922 (N_23922,N_15500,N_16363);
or U23923 (N_23923,N_16501,N_11243);
nand U23924 (N_23924,N_10330,N_15030);
nand U23925 (N_23925,N_18507,N_12814);
or U23926 (N_23926,N_13580,N_15251);
or U23927 (N_23927,N_14142,N_15576);
or U23928 (N_23928,N_16030,N_12199);
or U23929 (N_23929,N_15436,N_18329);
xnor U23930 (N_23930,N_17974,N_13265);
and U23931 (N_23931,N_15256,N_19769);
or U23932 (N_23932,N_12488,N_10525);
nand U23933 (N_23933,N_18454,N_10953);
or U23934 (N_23934,N_18191,N_18562);
or U23935 (N_23935,N_11534,N_10909);
nor U23936 (N_23936,N_11332,N_11767);
or U23937 (N_23937,N_14057,N_11758);
or U23938 (N_23938,N_11395,N_16448);
nor U23939 (N_23939,N_16649,N_10681);
and U23940 (N_23940,N_11897,N_16380);
xor U23941 (N_23941,N_17502,N_13420);
nand U23942 (N_23942,N_10002,N_17255);
nand U23943 (N_23943,N_10913,N_10272);
nand U23944 (N_23944,N_15791,N_12446);
nor U23945 (N_23945,N_15098,N_17254);
xor U23946 (N_23946,N_15747,N_13665);
nor U23947 (N_23947,N_15579,N_14276);
nor U23948 (N_23948,N_14166,N_13203);
or U23949 (N_23949,N_11672,N_11652);
or U23950 (N_23950,N_16765,N_14348);
and U23951 (N_23951,N_18243,N_10921);
and U23952 (N_23952,N_16136,N_13323);
nand U23953 (N_23953,N_15852,N_13530);
nand U23954 (N_23954,N_18381,N_10653);
nand U23955 (N_23955,N_17850,N_13466);
and U23956 (N_23956,N_14780,N_13291);
nand U23957 (N_23957,N_19805,N_16776);
nand U23958 (N_23958,N_15095,N_17168);
nor U23959 (N_23959,N_18568,N_12043);
nand U23960 (N_23960,N_10834,N_10801);
and U23961 (N_23961,N_14217,N_14470);
and U23962 (N_23962,N_10312,N_16434);
nor U23963 (N_23963,N_18783,N_12392);
nor U23964 (N_23964,N_15828,N_16038);
xor U23965 (N_23965,N_16060,N_12160);
nor U23966 (N_23966,N_15263,N_19251);
and U23967 (N_23967,N_10934,N_16783);
and U23968 (N_23968,N_11598,N_11772);
xor U23969 (N_23969,N_11678,N_12056);
or U23970 (N_23970,N_13971,N_15007);
xnor U23971 (N_23971,N_18476,N_13975);
or U23972 (N_23972,N_12988,N_12696);
xnor U23973 (N_23973,N_16598,N_11018);
nand U23974 (N_23974,N_12241,N_14292);
or U23975 (N_23975,N_10246,N_15504);
or U23976 (N_23976,N_10422,N_14980);
nand U23977 (N_23977,N_12275,N_11994);
or U23978 (N_23978,N_10373,N_18622);
or U23979 (N_23979,N_12208,N_15136);
or U23980 (N_23980,N_12023,N_13301);
nor U23981 (N_23981,N_19960,N_13106);
xnor U23982 (N_23982,N_19670,N_16051);
or U23983 (N_23983,N_19536,N_16148);
nor U23984 (N_23984,N_18579,N_18442);
nand U23985 (N_23985,N_10408,N_16777);
xnor U23986 (N_23986,N_18346,N_11962);
and U23987 (N_23987,N_18671,N_11906);
and U23988 (N_23988,N_14673,N_15032);
xnor U23989 (N_23989,N_12945,N_11907);
or U23990 (N_23990,N_19866,N_13507);
and U23991 (N_23991,N_10764,N_17714);
nor U23992 (N_23992,N_11596,N_15814);
or U23993 (N_23993,N_14733,N_18738);
nor U23994 (N_23994,N_11913,N_12754);
and U23995 (N_23995,N_16343,N_11935);
nor U23996 (N_23996,N_19462,N_12838);
nor U23997 (N_23997,N_14536,N_14743);
nand U23998 (N_23998,N_12237,N_10365);
or U23999 (N_23999,N_14706,N_16111);
and U24000 (N_24000,N_18880,N_15840);
nand U24001 (N_24001,N_13359,N_14267);
nor U24002 (N_24002,N_16932,N_13365);
nand U24003 (N_24003,N_13579,N_12324);
and U24004 (N_24004,N_19847,N_12297);
and U24005 (N_24005,N_13473,N_16311);
or U24006 (N_24006,N_15008,N_15076);
nor U24007 (N_24007,N_19460,N_17655);
or U24008 (N_24008,N_18319,N_16823);
xnor U24009 (N_24009,N_18053,N_19079);
xnor U24010 (N_24010,N_16317,N_16211);
nand U24011 (N_24011,N_10010,N_13505);
and U24012 (N_24012,N_19463,N_15489);
nand U24013 (N_24013,N_16888,N_11988);
or U24014 (N_24014,N_15357,N_14684);
nor U24015 (N_24015,N_15922,N_10652);
and U24016 (N_24016,N_11739,N_17915);
nand U24017 (N_24017,N_16237,N_10664);
nand U24018 (N_24018,N_11202,N_11489);
nand U24019 (N_24019,N_17682,N_13799);
nor U24020 (N_24020,N_14745,N_18291);
xnor U24021 (N_24021,N_14490,N_10014);
and U24022 (N_24022,N_11020,N_18063);
nand U24023 (N_24023,N_17694,N_16086);
nor U24024 (N_24024,N_18627,N_17334);
xor U24025 (N_24025,N_14234,N_17133);
and U24026 (N_24026,N_14458,N_11398);
or U24027 (N_24027,N_19111,N_19790);
xor U24028 (N_24028,N_17421,N_12156);
or U24029 (N_24029,N_14352,N_14228);
nand U24030 (N_24030,N_19002,N_13093);
or U24031 (N_24031,N_19975,N_13379);
nand U24032 (N_24032,N_17753,N_17139);
or U24033 (N_24033,N_12233,N_13764);
or U24034 (N_24034,N_11948,N_10937);
or U24035 (N_24035,N_10989,N_18419);
or U24036 (N_24036,N_11951,N_18093);
and U24037 (N_24037,N_10470,N_16293);
nor U24038 (N_24038,N_19459,N_18909);
or U24039 (N_24039,N_10730,N_18493);
nor U24040 (N_24040,N_15244,N_16471);
or U24041 (N_24041,N_19287,N_13482);
xnor U24042 (N_24042,N_17108,N_10701);
and U24043 (N_24043,N_17689,N_10566);
xnor U24044 (N_24044,N_18091,N_19354);
nor U24045 (N_24045,N_16409,N_13475);
nor U24046 (N_24046,N_15883,N_19834);
nor U24047 (N_24047,N_14692,N_16657);
nor U24048 (N_24048,N_12189,N_15164);
and U24049 (N_24049,N_13224,N_12791);
and U24050 (N_24050,N_12080,N_11504);
nand U24051 (N_24051,N_19130,N_18446);
and U24052 (N_24052,N_14513,N_11983);
and U24053 (N_24053,N_15761,N_18731);
and U24054 (N_24054,N_11428,N_10034);
nand U24055 (N_24055,N_15893,N_19772);
and U24056 (N_24056,N_10693,N_17930);
or U24057 (N_24057,N_13993,N_12001);
and U24058 (N_24058,N_14306,N_10683);
xor U24059 (N_24059,N_16301,N_14330);
and U24060 (N_24060,N_10484,N_12186);
or U24061 (N_24061,N_13056,N_18919);
nand U24062 (N_24062,N_17685,N_18850);
or U24063 (N_24063,N_10532,N_12254);
nand U24064 (N_24064,N_16463,N_11516);
nand U24065 (N_24065,N_12581,N_13790);
xnor U24066 (N_24066,N_14746,N_12504);
or U24067 (N_24067,N_14523,N_12776);
xor U24068 (N_24068,N_10846,N_13945);
nand U24069 (N_24069,N_14457,N_15089);
or U24070 (N_24070,N_19505,N_15102);
nand U24071 (N_24071,N_18962,N_14719);
nor U24072 (N_24072,N_14749,N_11614);
or U24073 (N_24073,N_13796,N_17158);
and U24074 (N_24074,N_19689,N_18841);
nor U24075 (N_24075,N_14279,N_15471);
nand U24076 (N_24076,N_10598,N_17090);
nand U24077 (N_24077,N_15311,N_14312);
or U24078 (N_24078,N_19223,N_18214);
nor U24079 (N_24079,N_14473,N_11792);
xor U24080 (N_24080,N_17613,N_10630);
xor U24081 (N_24081,N_17552,N_15343);
nor U24082 (N_24082,N_10019,N_10647);
nor U24083 (N_24083,N_16186,N_10344);
and U24084 (N_24084,N_10197,N_13245);
or U24085 (N_24085,N_12872,N_18965);
nor U24086 (N_24086,N_17754,N_10443);
and U24087 (N_24087,N_17081,N_14505);
nand U24088 (N_24088,N_13234,N_15528);
or U24089 (N_24089,N_17492,N_10845);
nand U24090 (N_24090,N_17967,N_12841);
nand U24091 (N_24091,N_10056,N_17970);
nand U24092 (N_24092,N_15022,N_16628);
or U24093 (N_24093,N_15735,N_16660);
xnor U24094 (N_24094,N_10173,N_14584);
or U24095 (N_24095,N_18132,N_19907);
nor U24096 (N_24096,N_19171,N_10232);
nor U24097 (N_24097,N_19428,N_10381);
nor U24098 (N_24098,N_14303,N_16304);
or U24099 (N_24099,N_19595,N_11755);
nor U24100 (N_24100,N_15861,N_17883);
xnor U24101 (N_24101,N_19873,N_19155);
nand U24102 (N_24102,N_18733,N_19306);
or U24103 (N_24103,N_16261,N_16252);
nor U24104 (N_24104,N_15132,N_16064);
nand U24105 (N_24105,N_17173,N_15954);
or U24106 (N_24106,N_15774,N_10698);
or U24107 (N_24107,N_10329,N_12034);
and U24108 (N_24108,N_15931,N_19607);
nor U24109 (N_24109,N_15302,N_16144);
or U24110 (N_24110,N_13550,N_11373);
nand U24111 (N_24111,N_17690,N_15026);
nand U24112 (N_24112,N_14427,N_15047);
nor U24113 (N_24113,N_19329,N_10319);
or U24114 (N_24114,N_11177,N_18589);
nand U24115 (N_24115,N_12353,N_14518);
xor U24116 (N_24116,N_17665,N_12362);
nor U24117 (N_24117,N_15935,N_14847);
and U24118 (N_24118,N_16398,N_12796);
nor U24119 (N_24119,N_15675,N_18215);
nand U24120 (N_24120,N_19403,N_19302);
nand U24121 (N_24121,N_15767,N_19435);
nor U24122 (N_24122,N_10608,N_19317);
and U24123 (N_24123,N_10748,N_17330);
nand U24124 (N_24124,N_16171,N_12991);
and U24125 (N_24125,N_14215,N_10621);
xnor U24126 (N_24126,N_10390,N_16720);
xnor U24127 (N_24127,N_18176,N_10073);
or U24128 (N_24128,N_18365,N_19298);
nand U24129 (N_24129,N_13213,N_12279);
or U24130 (N_24130,N_13659,N_10715);
and U24131 (N_24131,N_13699,N_14855);
or U24132 (N_24132,N_16073,N_12183);
and U24133 (N_24133,N_12621,N_12805);
and U24134 (N_24134,N_11122,N_19800);
nor U24135 (N_24135,N_18418,N_14347);
nor U24136 (N_24136,N_19716,N_16787);
or U24137 (N_24137,N_14981,N_17615);
xor U24138 (N_24138,N_14632,N_12878);
or U24139 (N_24139,N_13362,N_17756);
nor U24140 (N_24140,N_11659,N_17443);
xnor U24141 (N_24141,N_12729,N_13366);
or U24142 (N_24142,N_18547,N_17933);
or U24143 (N_24143,N_14867,N_12900);
nor U24144 (N_24144,N_14341,N_15088);
nor U24145 (N_24145,N_13584,N_16833);
nor U24146 (N_24146,N_12249,N_10370);
nand U24147 (N_24147,N_19592,N_18745);
and U24148 (N_24148,N_11140,N_11141);
xor U24149 (N_24149,N_17042,N_17852);
nor U24150 (N_24150,N_18748,N_16576);
nor U24151 (N_24151,N_19280,N_17656);
xor U24152 (N_24152,N_19984,N_14023);
xnor U24153 (N_24153,N_15440,N_16462);
or U24154 (N_24154,N_14688,N_13811);
nand U24155 (N_24155,N_16927,N_11751);
nand U24156 (N_24156,N_15771,N_19307);
and U24157 (N_24157,N_10024,N_19250);
and U24158 (N_24158,N_17331,N_12675);
or U24159 (N_24159,N_16335,N_15844);
nor U24160 (N_24160,N_11089,N_14621);
nor U24161 (N_24161,N_14960,N_14291);
or U24162 (N_24162,N_13677,N_19107);
and U24163 (N_24163,N_19131,N_10568);
or U24164 (N_24164,N_16781,N_18525);
nor U24165 (N_24165,N_15051,N_14967);
nor U24166 (N_24166,N_15166,N_19259);
nand U24167 (N_24167,N_19874,N_17071);
and U24168 (N_24168,N_11925,N_18149);
xnor U24169 (N_24169,N_16546,N_17881);
nand U24170 (N_24170,N_16549,N_15720);
nor U24171 (N_24171,N_15239,N_11738);
nand U24172 (N_24172,N_16866,N_16010);
nor U24173 (N_24173,N_18182,N_10826);
nand U24174 (N_24174,N_19236,N_13829);
or U24175 (N_24175,N_10045,N_19159);
nand U24176 (N_24176,N_15664,N_12370);
nand U24177 (N_24177,N_18485,N_15188);
xor U24178 (N_24178,N_13178,N_18487);
xor U24179 (N_24179,N_18799,N_10227);
and U24180 (N_24180,N_18270,N_19631);
nand U24181 (N_24181,N_16749,N_17728);
and U24182 (N_24182,N_17333,N_19373);
xor U24183 (N_24183,N_13625,N_14883);
nor U24184 (N_24184,N_19336,N_14019);
and U24185 (N_24185,N_16572,N_18724);
nand U24186 (N_24186,N_15667,N_19008);
nor U24187 (N_24187,N_12907,N_13392);
and U24188 (N_24188,N_15611,N_14918);
and U24189 (N_24189,N_17730,N_17571);
or U24190 (N_24190,N_10746,N_11156);
nand U24191 (N_24191,N_18287,N_13104);
xnor U24192 (N_24192,N_19781,N_10105);
and U24193 (N_24193,N_15928,N_16611);
or U24194 (N_24194,N_14461,N_13413);
and U24195 (N_24195,N_17587,N_10168);
or U24196 (N_24196,N_13220,N_15640);
or U24197 (N_24197,N_19284,N_11418);
nand U24198 (N_24198,N_12877,N_16312);
nand U24199 (N_24199,N_14856,N_17503);
and U24200 (N_24200,N_12704,N_18503);
nand U24201 (N_24201,N_17900,N_10977);
and U24202 (N_24202,N_16714,N_13128);
and U24203 (N_24203,N_10427,N_19820);
and U24204 (N_24204,N_12919,N_14386);
nor U24205 (N_24205,N_14149,N_11603);
nor U24206 (N_24206,N_11019,N_19761);
nand U24207 (N_24207,N_12149,N_18662);
nor U24208 (N_24208,N_14664,N_13715);
and U24209 (N_24209,N_13251,N_12840);
nor U24210 (N_24210,N_16732,N_13894);
nor U24211 (N_24211,N_13189,N_13999);
xnor U24212 (N_24212,N_15320,N_16133);
nor U24213 (N_24213,N_16047,N_15213);
nor U24214 (N_24214,N_14839,N_18742);
nor U24215 (N_24215,N_14810,N_18304);
nand U24216 (N_24216,N_14161,N_14644);
and U24217 (N_24217,N_17323,N_11033);
nor U24218 (N_24218,N_14787,N_17788);
or U24219 (N_24219,N_19464,N_13576);
xor U24220 (N_24220,N_19519,N_17306);
and U24221 (N_24221,N_13646,N_12495);
nor U24222 (N_24222,N_16686,N_16898);
nor U24223 (N_24223,N_14484,N_19206);
nor U24224 (N_24224,N_12486,N_15626);
nor U24225 (N_24225,N_15627,N_18906);
and U24226 (N_24226,N_19715,N_11804);
and U24227 (N_24227,N_17921,N_17898);
and U24228 (N_24228,N_14723,N_11021);
and U24229 (N_24229,N_17335,N_12705);
nor U24230 (N_24230,N_15891,N_16960);
nor U24231 (N_24231,N_18794,N_15961);
nor U24232 (N_24232,N_19578,N_16806);
xor U24233 (N_24233,N_17198,N_15398);
xor U24234 (N_24234,N_19237,N_14316);
xor U24235 (N_24235,N_15469,N_12268);
or U24236 (N_24236,N_14208,N_15202);
or U24237 (N_24237,N_16742,N_19458);
nor U24238 (N_24238,N_17361,N_18583);
nand U24239 (N_24239,N_12684,N_12960);
and U24240 (N_24240,N_15467,N_16222);
nor U24241 (N_24241,N_11923,N_11150);
nand U24242 (N_24242,N_10376,N_18741);
nand U24243 (N_24243,N_10975,N_12614);
nor U24244 (N_24244,N_14095,N_11268);
nor U24245 (N_24245,N_12812,N_17971);
nand U24246 (N_24246,N_19520,N_12664);
and U24247 (N_24247,N_12721,N_14025);
nand U24248 (N_24248,N_12974,N_15618);
nand U24249 (N_24249,N_16907,N_18017);
and U24250 (N_24250,N_10798,N_10915);
nand U24251 (N_24251,N_18198,N_13450);
and U24252 (N_24252,N_11919,N_11589);
and U24253 (N_24253,N_17594,N_17879);
or U24254 (N_24254,N_13279,N_12602);
or U24255 (N_24255,N_10192,N_10548);
or U24256 (N_24256,N_19663,N_15748);
nand U24257 (N_24257,N_11478,N_16052);
nor U24258 (N_24258,N_12517,N_13977);
nand U24259 (N_24259,N_15490,N_11870);
and U24260 (N_24260,N_16517,N_11917);
and U24261 (N_24261,N_16107,N_10054);
or U24262 (N_24262,N_16147,N_18566);
or U24263 (N_24263,N_10535,N_11147);
nor U24264 (N_24264,N_18608,N_12981);
or U24265 (N_24265,N_19643,N_14131);
nor U24266 (N_24266,N_15680,N_12073);
and U24267 (N_24267,N_14028,N_14887);
or U24268 (N_24268,N_14588,N_11108);
or U24269 (N_24269,N_15133,N_19137);
or U24270 (N_24270,N_12825,N_18758);
xor U24271 (N_24271,N_12371,N_13130);
nor U24272 (N_24272,N_14957,N_12746);
xnor U24273 (N_24273,N_10792,N_11768);
or U24274 (N_24274,N_12646,N_18115);
and U24275 (N_24275,N_13685,N_12407);
nor U24276 (N_24276,N_15326,N_12202);
or U24277 (N_24277,N_13560,N_15004);
nand U24278 (N_24278,N_11877,N_11163);
nand U24279 (N_24279,N_11501,N_17083);
nand U24280 (N_24280,N_16490,N_10773);
nor U24281 (N_24281,N_18253,N_14093);
nor U24282 (N_24282,N_19614,N_11304);
and U24283 (N_24283,N_15268,N_11253);
nor U24284 (N_24284,N_17572,N_15452);
and U24285 (N_24285,N_19531,N_14816);
nand U24286 (N_24286,N_12188,N_11742);
xor U24287 (N_24287,N_18659,N_13139);
and U24288 (N_24288,N_13151,N_19709);
and U24289 (N_24289,N_13632,N_18422);
nor U24290 (N_24290,N_11943,N_11171);
and U24291 (N_24291,N_19129,N_12076);
xnor U24292 (N_24292,N_11111,N_17296);
nand U24293 (N_24293,N_17180,N_10969);
nand U24294 (N_24294,N_16509,N_17628);
and U24295 (N_24295,N_10270,N_13819);
nor U24296 (N_24296,N_18817,N_14577);
nor U24297 (N_24297,N_18689,N_17675);
nor U24298 (N_24298,N_14254,N_15159);
nand U24299 (N_24299,N_13370,N_18955);
or U24300 (N_24300,N_10254,N_10943);
and U24301 (N_24301,N_14956,N_15220);
or U24302 (N_24302,N_16188,N_12190);
and U24303 (N_24303,N_12124,N_14771);
and U24304 (N_24304,N_11201,N_13660);
xnor U24305 (N_24305,N_10676,N_10216);
or U24306 (N_24306,N_12338,N_15121);
and U24307 (N_24307,N_12888,N_17428);
nand U24308 (N_24308,N_13070,N_15148);
nor U24309 (N_24309,N_13304,N_19819);
and U24310 (N_24310,N_16004,N_16342);
nor U24311 (N_24311,N_19659,N_16477);
nand U24312 (N_24312,N_11646,N_16764);
nand U24313 (N_24313,N_10212,N_10784);
nand U24314 (N_24314,N_17899,N_10180);
or U24315 (N_24315,N_10885,N_10225);
and U24316 (N_24316,N_16850,N_10970);
nor U24317 (N_24317,N_19453,N_10458);
nand U24318 (N_24318,N_14597,N_13478);
or U24319 (N_24319,N_15364,N_11213);
nor U24320 (N_24320,N_12813,N_12337);
nand U24321 (N_24321,N_15375,N_14851);
nand U24322 (N_24322,N_14286,N_15704);
nor U24323 (N_24323,N_13133,N_12016);
and U24324 (N_24324,N_10454,N_18674);
nor U24325 (N_24325,N_10738,N_16262);
and U24326 (N_24326,N_11132,N_17143);
nand U24327 (N_24327,N_15031,N_15069);
nand U24328 (N_24328,N_13477,N_15531);
and U24329 (N_24329,N_19885,N_16229);
nor U24330 (N_24330,N_17592,N_15530);
or U24331 (N_24331,N_12072,N_16466);
nand U24332 (N_24332,N_16619,N_17928);
or U24333 (N_24333,N_14044,N_12449);
or U24334 (N_24334,N_13750,N_15317);
and U24335 (N_24335,N_13904,N_17459);
nand U24336 (N_24336,N_18489,N_11365);
xnor U24337 (N_24337,N_10023,N_11986);
nand U24338 (N_24338,N_11353,N_12843);
and U24339 (N_24339,N_11773,N_19005);
nand U24340 (N_24340,N_19734,N_12152);
or U24341 (N_24341,N_15082,N_15850);
nor U24342 (N_24342,N_18791,N_10974);
nand U24343 (N_24343,N_10884,N_13544);
and U24344 (N_24344,N_13575,N_10848);
nor U24345 (N_24345,N_13546,N_15218);
and U24346 (N_24346,N_13412,N_15956);
nand U24347 (N_24347,N_18459,N_19799);
or U24348 (N_24348,N_16110,N_13524);
nor U24349 (N_24349,N_19966,N_19628);
nor U24350 (N_24350,N_10891,N_18585);
nand U24351 (N_24351,N_14091,N_19418);
nor U24352 (N_24352,N_15406,N_19270);
nand U24353 (N_24353,N_10793,N_18840);
and U24354 (N_24354,N_14535,N_11803);
nor U24355 (N_24355,N_17726,N_15105);
xnor U24356 (N_24356,N_14974,N_16142);
and U24357 (N_24357,N_18341,N_16690);
and U24358 (N_24358,N_16455,N_19028);
or U24359 (N_24359,N_14074,N_19795);
xnor U24360 (N_24360,N_19114,N_18661);
nand U24361 (N_24361,N_15358,N_15281);
and U24362 (N_24362,N_18960,N_10770);
or U24363 (N_24363,N_16215,N_16134);
or U24364 (N_24364,N_15212,N_10960);
or U24365 (N_24365,N_11362,N_17947);
or U24366 (N_24366,N_18305,N_17824);
or U24367 (N_24367,N_14152,N_13931);
nor U24368 (N_24368,N_14556,N_15257);
nor U24369 (N_24369,N_12683,N_13048);
nor U24370 (N_24370,N_11694,N_13205);
nand U24371 (N_24371,N_15287,N_14181);
nand U24372 (N_24372,N_12350,N_11206);
xor U24373 (N_24373,N_10519,N_10251);
nor U24374 (N_24374,N_17223,N_10309);
nand U24375 (N_24375,N_12240,N_11437);
or U24376 (N_24376,N_16928,N_17586);
nor U24377 (N_24377,N_12959,N_14503);
nand U24378 (N_24378,N_14601,N_19679);
xnor U24379 (N_24379,N_16504,N_13800);
nand U24380 (N_24380,N_15753,N_13411);
nor U24381 (N_24381,N_11461,N_14985);
or U24382 (N_24382,N_11221,N_10005);
and U24383 (N_24383,N_17199,N_12955);
nor U24384 (N_24384,N_17494,N_13289);
and U24385 (N_24385,N_12530,N_15142);
xnor U24386 (N_24386,N_12678,N_15101);
and U24387 (N_24387,N_19120,N_17463);
nor U24388 (N_24388,N_10167,N_14948);
nand U24389 (N_24389,N_16825,N_14574);
nand U24390 (N_24390,N_11239,N_16512);
nand U24391 (N_24391,N_12875,N_18771);
and U24392 (N_24392,N_15086,N_14042);
and U24393 (N_24393,N_10475,N_17096);
nor U24394 (N_24394,N_17067,N_13892);
and U24395 (N_24395,N_18012,N_16258);
or U24396 (N_24396,N_18677,N_12526);
or U24397 (N_24397,N_12743,N_17046);
or U24398 (N_24398,N_11191,N_10305);
nand U24399 (N_24399,N_18231,N_17661);
nor U24400 (N_24400,N_10230,N_15958);
or U24401 (N_24401,N_16279,N_11469);
xnor U24402 (N_24402,N_19534,N_13722);
or U24403 (N_24403,N_13463,N_14040);
nor U24404 (N_24404,N_11993,N_17232);
and U24405 (N_24405,N_19640,N_19717);
xnor U24406 (N_24406,N_14337,N_14189);
nand U24407 (N_24407,N_13656,N_11143);
nand U24408 (N_24408,N_14251,N_19586);
or U24409 (N_24409,N_19521,N_15099);
or U24410 (N_24410,N_10048,N_18087);
nor U24411 (N_24411,N_12912,N_16733);
and U24412 (N_24412,N_19826,N_17261);
or U24413 (N_24413,N_17960,N_19058);
or U24414 (N_24414,N_19257,N_18225);
and U24415 (N_24415,N_10726,N_17877);
and U24416 (N_24416,N_13955,N_17166);
and U24417 (N_24417,N_11707,N_13173);
nor U24418 (N_24418,N_19499,N_14870);
nor U24419 (N_24419,N_16525,N_18113);
nand U24420 (N_24420,N_13394,N_16306);
or U24421 (N_24421,N_19321,N_11249);
nand U24422 (N_24422,N_11381,N_14178);
or U24423 (N_24423,N_11012,N_18279);
nand U24424 (N_24424,N_12709,N_15558);
or U24425 (N_24425,N_13426,N_16088);
and U24426 (N_24426,N_11505,N_14261);
and U24427 (N_24427,N_12799,N_19039);
nand U24428 (N_24428,N_19727,N_13517);
and U24429 (N_24429,N_12286,N_17007);
or U24430 (N_24430,N_18085,N_13285);
or U24431 (N_24431,N_18189,N_19070);
and U24432 (N_24432,N_18691,N_13942);
or U24433 (N_24433,N_15324,N_13185);
or U24434 (N_24434,N_19407,N_12543);
xor U24435 (N_24435,N_13177,N_12573);
nor U24436 (N_24436,N_15480,N_16563);
nor U24437 (N_24437,N_18939,N_13960);
nand U24438 (N_24438,N_14476,N_11178);
nand U24439 (N_24439,N_17358,N_18021);
or U24440 (N_24440,N_16489,N_18405);
nor U24441 (N_24441,N_12828,N_19894);
and U24442 (N_24442,N_15487,N_12598);
or U24443 (N_24443,N_16604,N_19822);
or U24444 (N_24444,N_18448,N_16415);
nand U24445 (N_24445,N_17576,N_17833);
nand U24446 (N_24446,N_19591,N_18453);
and U24447 (N_24447,N_18011,N_11225);
xor U24448 (N_24448,N_13985,N_18996);
and U24449 (N_24449,N_14300,N_19074);
or U24450 (N_24450,N_14862,N_15178);
or U24451 (N_24451,N_18856,N_17389);
nor U24452 (N_24452,N_12382,N_12536);
nor U24453 (N_24453,N_18924,N_14314);
nand U24454 (N_24454,N_18041,N_14081);
and U24455 (N_24455,N_17195,N_11639);
and U24456 (N_24456,N_10936,N_17256);
and U24457 (N_24457,N_16728,N_17832);
or U24458 (N_24458,N_16194,N_12061);
nor U24459 (N_24459,N_18766,N_12356);
nor U24460 (N_24460,N_17072,N_12177);
nor U24461 (N_24461,N_16668,N_15652);
and U24462 (N_24462,N_12033,N_17662);
or U24463 (N_24463,N_17939,N_13849);
nand U24464 (N_24464,N_10739,N_16968);
and U24465 (N_24465,N_17487,N_15016);
or U24466 (N_24466,N_17987,N_10050);
nand U24467 (N_24467,N_14615,N_13741);
and U24468 (N_24468,N_13838,N_12765);
and U24469 (N_24469,N_16726,N_11183);
and U24470 (N_24470,N_19547,N_17328);
nand U24471 (N_24471,N_18614,N_19622);
nand U24472 (N_24472,N_12451,N_10911);
nor U24473 (N_24473,N_19621,N_18092);
or U24474 (N_24474,N_11322,N_18218);
nand U24475 (N_24475,N_15208,N_10112);
nand U24476 (N_24476,N_19493,N_17851);
and U24477 (N_24477,N_16318,N_19945);
or U24478 (N_24478,N_17039,N_17758);
xnor U24479 (N_24479,N_12163,N_10926);
nand U24480 (N_24480,N_17793,N_10544);
nand U24481 (N_24481,N_16179,N_16527);
or U24482 (N_24482,N_12442,N_15110);
nand U24483 (N_24483,N_10573,N_15983);
nand U24484 (N_24484,N_16971,N_11277);
nor U24485 (N_24485,N_13107,N_10213);
nor U24486 (N_24486,N_10781,N_18642);
nand U24487 (N_24487,N_13809,N_11618);
nand U24488 (N_24488,N_18537,N_18258);
and U24489 (N_24489,N_19594,N_14996);
nand U24490 (N_24490,N_14620,N_13557);
nor U24491 (N_24491,N_10612,N_12616);
nor U24492 (N_24492,N_14073,N_19692);
nand U24493 (N_24493,N_15334,N_15291);
nand U24494 (N_24494,N_19814,N_14475);
xnor U24495 (N_24495,N_13523,N_12336);
nor U24496 (N_24496,N_11736,N_16535);
nor U24497 (N_24497,N_14336,N_10383);
and U24498 (N_24498,N_14371,N_11954);
nor U24499 (N_24499,N_17676,N_13661);
and U24500 (N_24500,N_10284,N_18470);
nand U24501 (N_24501,N_13175,N_11931);
or U24502 (N_24502,N_14659,N_15915);
nor U24503 (N_24503,N_14175,N_13326);
and U24504 (N_24504,N_15474,N_12833);
or U24505 (N_24505,N_10405,N_18260);
nand U24506 (N_24506,N_19396,N_10961);
nor U24507 (N_24507,N_15429,N_18075);
nand U24508 (N_24508,N_12906,N_12234);
or U24509 (N_24509,N_13639,N_11370);
nand U24510 (N_24510,N_16805,N_19239);
xnor U24511 (N_24511,N_18452,N_18511);
xnor U24512 (N_24512,N_11999,N_13915);
nand U24513 (N_24513,N_12948,N_17170);
nor U24514 (N_24514,N_15232,N_12376);
nor U24515 (N_24515,N_18598,N_10620);
xnor U24516 (N_24516,N_12585,N_18883);
or U24517 (N_24517,N_16596,N_13016);
or U24518 (N_24518,N_17269,N_18236);
nand U24519 (N_24519,N_19700,N_14853);
nor U24520 (N_24520,N_16680,N_12760);
nand U24521 (N_24521,N_10563,N_15325);
and U24522 (N_24522,N_10107,N_19606);
or U24523 (N_24523,N_13884,N_13791);
nand U24524 (N_24524,N_16769,N_13195);
nand U24525 (N_24525,N_13036,N_15292);
nor U24526 (N_24526,N_14417,N_19167);
or U24527 (N_24527,N_11550,N_13439);
nor U24528 (N_24528,N_12269,N_18067);
nor U24529 (N_24529,N_10207,N_13415);
and U24530 (N_24530,N_16944,N_17134);
or U24531 (N_24531,N_17627,N_14453);
and U24532 (N_24532,N_13393,N_10963);
nand U24533 (N_24533,N_14992,N_15322);
and U24534 (N_24534,N_19612,N_13110);
or U24535 (N_24535,N_13793,N_13298);
or U24536 (N_24536,N_13541,N_18721);
and U24537 (N_24537,N_15692,N_16658);
or U24538 (N_24538,N_18197,N_18383);
or U24539 (N_24539,N_18154,N_11554);
nand U24540 (N_24540,N_19779,N_13281);
and U24541 (N_24541,N_10130,N_13776);
nand U24542 (N_24542,N_13170,N_19686);
or U24543 (N_24543,N_11256,N_13142);
nor U24544 (N_24544,N_17777,N_13204);
xor U24545 (N_24545,N_10839,N_12115);
nand U24546 (N_24546,N_18864,N_18266);
nand U24547 (N_24547,N_13719,N_16685);
nand U24548 (N_24548,N_15247,N_16814);
and U24549 (N_24549,N_19347,N_11864);
and U24550 (N_24550,N_19049,N_19956);
nand U24551 (N_24551,N_15849,N_11126);
nand U24552 (N_24552,N_13258,N_17030);
nand U24553 (N_24553,N_19935,N_17598);
nand U24554 (N_24554,N_18413,N_10651);
nand U24555 (N_24555,N_14359,N_18156);
or U24556 (N_24556,N_12715,N_15890);
nor U24557 (N_24557,N_13072,N_14413);
nand U24558 (N_24558,N_17752,N_13136);
nor U24559 (N_24559,N_16559,N_16694);
nand U24560 (N_24560,N_18248,N_19581);
nor U24561 (N_24561,N_19381,N_17314);
and U24562 (N_24562,N_12782,N_13077);
and U24563 (N_24563,N_18940,N_15153);
nand U24564 (N_24564,N_11460,N_16857);
or U24565 (N_24565,N_13256,N_13785);
nand U24566 (N_24566,N_10870,N_12990);
or U24567 (N_24567,N_19217,N_11700);
nand U24568 (N_24568,N_12060,N_12091);
and U24569 (N_24569,N_10281,N_18988);
nand U24570 (N_24570,N_18631,N_12851);
and U24571 (N_24571,N_11933,N_11593);
and U24572 (N_24572,N_16063,N_19054);
nand U24573 (N_24573,N_10833,N_18580);
xnor U24574 (N_24574,N_19997,N_13430);
xor U24575 (N_24575,N_12934,N_14983);
xnor U24576 (N_24576,N_18153,N_15592);
nand U24577 (N_24577,N_10768,N_19637);
nor U24578 (N_24578,N_10439,N_10347);
and U24579 (N_24579,N_19412,N_12473);
nand U24580 (N_24580,N_13693,N_16632);
and U24581 (N_24581,N_11307,N_14714);
or U24582 (N_24582,N_17156,N_18692);
nor U24583 (N_24583,N_19032,N_18157);
xnor U24584 (N_24584,N_14766,N_10321);
or U24585 (N_24585,N_13214,N_10829);
nor U24586 (N_24586,N_13949,N_16428);
or U24587 (N_24587,N_10070,N_14545);
and U24588 (N_24588,N_17231,N_16751);
xnor U24589 (N_24589,N_19751,N_12242);
nand U24590 (N_24590,N_12887,N_11495);
or U24591 (N_24591,N_12509,N_11476);
or U24592 (N_24592,N_19261,N_10327);
nor U24593 (N_24593,N_14196,N_17732);
nor U24594 (N_24594,N_15486,N_11732);
nand U24595 (N_24595,N_12592,N_17352);
and U24596 (N_24596,N_17736,N_12859);
and U24597 (N_24597,N_18408,N_13492);
or U24598 (N_24598,N_16986,N_18717);
and U24599 (N_24599,N_14202,N_13526);
and U24600 (N_24600,N_10333,N_19156);
and U24601 (N_24601,N_10326,N_15561);
nand U24602 (N_24602,N_18148,N_16493);
nand U24603 (N_24603,N_16629,N_15745);
nor U24604 (N_24604,N_15981,N_17092);
nor U24605 (N_24605,N_19165,N_18501);
nand U24606 (N_24606,N_16384,N_13098);
nand U24607 (N_24607,N_15373,N_16775);
nand U24608 (N_24608,N_18623,N_16892);
nand U24609 (N_24609,N_11571,N_18049);
or U24610 (N_24610,N_15204,N_14937);
nor U24611 (N_24611,N_18352,N_11892);
nor U24612 (N_24612,N_16123,N_18617);
or U24613 (N_24613,N_13221,N_15856);
nand U24614 (N_24614,N_19234,N_16081);
nor U24615 (N_24615,N_13690,N_16438);
nor U24616 (N_24616,N_14666,N_18326);
or U24617 (N_24617,N_14943,N_18761);
nor U24618 (N_24618,N_19408,N_18073);
nor U24619 (N_24619,N_11518,N_13087);
and U24620 (N_24620,N_10163,N_13921);
xor U24621 (N_24621,N_16388,N_10345);
or U24622 (N_24622,N_10832,N_16873);
and U24623 (N_24623,N_15971,N_19949);
or U24624 (N_24624,N_10059,N_18361);
xor U24625 (N_24625,N_12865,N_12962);
or U24626 (N_24626,N_17674,N_10508);
and U24627 (N_24627,N_17406,N_15458);
nand U24628 (N_24628,N_18045,N_12824);
nor U24629 (N_24629,N_10164,N_11459);
nor U24630 (N_24630,N_13019,N_13027);
nand U24631 (N_24631,N_15261,N_17400);
or U24632 (N_24632,N_11841,N_19263);
and U24633 (N_24633,N_17267,N_17638);
and U24634 (N_24634,N_18462,N_11152);
nor U24635 (N_24635,N_10488,N_17637);
and U24636 (N_24636,N_11663,N_19798);
nor U24637 (N_24637,N_12943,N_16447);
nand U24638 (N_24638,N_13035,N_12644);
nand U24639 (N_24639,N_15285,N_18995);
and U24640 (N_24640,N_13075,N_10627);
nor U24641 (N_24641,N_15061,N_10393);
xor U24642 (N_24642,N_11034,N_11292);
or U24643 (N_24643,N_16416,N_14599);
nor U24644 (N_24644,N_19046,N_11076);
nor U24645 (N_24645,N_10629,N_13732);
xnor U24646 (N_24646,N_12062,N_18046);
nand U24647 (N_24647,N_12953,N_16738);
and U24648 (N_24648,N_16482,N_19629);
nand U24649 (N_24649,N_17289,N_16739);
nand U24650 (N_24650,N_10102,N_12375);
nand U24651 (N_24651,N_15344,N_10579);
nand U24652 (N_24652,N_18016,N_12499);
nand U24653 (N_24653,N_18824,N_18963);
and U24654 (N_24654,N_15356,N_11575);
or U24655 (N_24655,N_12924,N_13143);
nor U24656 (N_24656,N_12294,N_10901);
nor U24657 (N_24657,N_10355,N_13698);
nor U24658 (N_24658,N_19667,N_12725);
xor U24659 (N_24659,N_12538,N_13119);
and U24660 (N_24660,N_11421,N_19052);
nor U24661 (N_24661,N_16772,N_14321);
nor U24662 (N_24662,N_12151,N_11950);
and U24663 (N_24663,N_17663,N_10590);
nand U24664 (N_24664,N_14986,N_12193);
nand U24665 (N_24665,N_14707,N_10063);
nor U24666 (N_24666,N_14720,N_15859);
nor U24667 (N_24667,N_14067,N_12808);
nor U24668 (N_24668,N_18700,N_17080);
and U24669 (N_24669,N_15676,N_13479);
nand U24670 (N_24670,N_13836,N_16305);
and U24671 (N_24671,N_11187,N_12172);
and U24672 (N_24672,N_14995,N_11535);
nand U24673 (N_24673,N_18964,N_13380);
nand U24674 (N_24674,N_18942,N_10788);
nor U24675 (N_24675,N_15724,N_13655);
nor U24676 (N_24676,N_11279,N_16066);
nor U24677 (N_24677,N_10656,N_12947);
or U24678 (N_24678,N_17213,N_11007);
nand U24679 (N_24679,N_11809,N_14046);
nor U24680 (N_24680,N_15387,N_15258);
and U24681 (N_24681,N_18888,N_16417);
or U24682 (N_24682,N_18293,N_16003);
nor U24683 (N_24683,N_19140,N_13761);
or U24684 (N_24684,N_10941,N_16672);
or U24685 (N_24685,N_17569,N_14324);
nor U24686 (N_24686,N_11184,N_15271);
nor U24687 (N_24687,N_18603,N_16637);
and U24688 (N_24688,N_10994,N_12645);
nor U24689 (N_24689,N_13984,N_17162);
nand U24690 (N_24690,N_17980,N_16282);
and U24691 (N_24691,N_12346,N_11867);
or U24692 (N_24692,N_15578,N_16451);
nand U24693 (N_24693,N_13748,N_11560);
nor U24694 (N_24694,N_15673,N_17483);
nand U24695 (N_24695,N_18984,N_18380);
and U24696 (N_24696,N_15732,N_16104);
or U24697 (N_24697,N_14987,N_19356);
xnor U24698 (N_24698,N_19276,N_13848);
nor U24699 (N_24699,N_10461,N_17621);
or U24700 (N_24700,N_11022,N_17616);
nor U24701 (N_24701,N_12939,N_19572);
nor U24702 (N_24702,N_11315,N_12966);
nand U24703 (N_24703,N_16581,N_14089);
nand U24704 (N_24704,N_12653,N_14657);
and U24705 (N_24705,N_10346,N_13795);
xor U24706 (N_24706,N_16789,N_18518);
nor U24707 (N_24707,N_16090,N_14509);
or U24708 (N_24708,N_19047,N_11806);
nor U24709 (N_24709,N_14232,N_12600);
or U24710 (N_24710,N_10316,N_18288);
or U24711 (N_24711,N_11989,N_18836);
nand U24712 (N_24712,N_16993,N_12260);
and U24713 (N_24713,N_10863,N_13895);
or U24714 (N_24714,N_12022,N_16496);
and U24715 (N_24715,N_18299,N_14931);
and U24716 (N_24716,N_11937,N_11375);
nand U24717 (N_24717,N_13902,N_15400);
or U24718 (N_24718,N_17624,N_15921);
xnor U24719 (N_24719,N_17262,N_10696);
xor U24720 (N_24720,N_17197,N_18759);
nand U24721 (N_24721,N_18921,N_15574);
or U24722 (N_24722,N_18278,N_19334);
or U24723 (N_24723,N_13585,N_17294);
or U24724 (N_24724,N_15706,N_17864);
or U24725 (N_24725,N_18229,N_19362);
and U24726 (N_24726,N_10946,N_14668);
or U24727 (N_24727,N_15255,N_19844);
or U24728 (N_24728,N_15341,N_11648);
and U24729 (N_24729,N_11195,N_14872);
nor U24730 (N_24730,N_12886,N_14868);
nor U24731 (N_24731,N_16173,N_14225);
nand U24732 (N_24732,N_10123,N_15321);
nor U24733 (N_24733,N_10763,N_19180);
and U24734 (N_24734,N_18318,N_13417);
nor U24735 (N_24735,N_18373,N_19712);
nand U24736 (N_24736,N_12369,N_13184);
nand U24737 (N_24737,N_19756,N_11343);
nand U24738 (N_24738,N_18374,N_10377);
xor U24739 (N_24739,N_12827,N_14404);
nor U24740 (N_24740,N_13193,N_11323);
and U24741 (N_24741,N_12218,N_13972);
and U24742 (N_24742,N_15623,N_19296);
nand U24743 (N_24743,N_11197,N_14686);
nor U24744 (N_24744,N_19089,N_10285);
or U24745 (N_24745,N_12093,N_16533);
nand U24746 (N_24746,N_15044,N_12694);
nand U24747 (N_24747,N_18300,N_17354);
nor U24748 (N_24748,N_11660,N_10607);
or U24749 (N_24749,N_15011,N_11726);
or U24750 (N_24750,N_16206,N_18992);
nor U24751 (N_24751,N_17523,N_19319);
nor U24752 (N_24752,N_14651,N_15862);
xnor U24753 (N_24753,N_15039,N_15708);
or U24754 (N_24754,N_16161,N_12610);
nor U24755 (N_24755,N_19188,N_14681);
nand U24756 (N_24756,N_12863,N_11247);
xor U24757 (N_24757,N_16404,N_13820);
xnor U24758 (N_24758,N_12583,N_11794);
and U24759 (N_24759,N_19024,N_16566);
nor U24760 (N_24760,N_17128,N_15927);
or U24761 (N_24761,N_12378,N_12687);
nor U24762 (N_24762,N_11211,N_17835);
and U24763 (N_24763,N_17235,N_10628);
nand U24764 (N_24764,N_17302,N_16324);
and U24765 (N_24765,N_19341,N_17461);
or U24766 (N_24766,N_18976,N_17340);
nor U24767 (N_24767,N_16153,N_17399);
or U24768 (N_24768,N_11318,N_12835);
nor U24769 (N_24769,N_13160,N_18643);
nor U24770 (N_24770,N_19563,N_16458);
nor U24771 (N_24771,N_16949,N_15613);
nand U24772 (N_24772,N_19923,N_10669);
or U24773 (N_24773,N_16877,N_10966);
or U24774 (N_24774,N_17153,N_12121);
nor U24775 (N_24775,N_16089,N_15975);
nor U24776 (N_24776,N_17171,N_14752);
nor U24777 (N_24777,N_11807,N_16675);
xnor U24778 (N_24778,N_12247,N_17104);
or U24779 (N_24779,N_14483,N_17008);
nor U24780 (N_24780,N_11293,N_11073);
nor U24781 (N_24781,N_18821,N_19768);
nand U24782 (N_24782,N_16524,N_17964);
xnor U24783 (N_24783,N_13780,N_17891);
and U24784 (N_24784,N_12624,N_13033);
or U24785 (N_24785,N_12987,N_13122);
nor U24786 (N_24786,N_14665,N_12724);
or U24787 (N_24787,N_12596,N_12628);
xnor U24788 (N_24788,N_12194,N_11778);
xor U24789 (N_24789,N_18669,N_14433);
nand U24790 (N_24790,N_10584,N_17519);
xor U24791 (N_24791,N_10907,N_16245);
and U24792 (N_24792,N_11967,N_11081);
and U24793 (N_24793,N_18862,N_19043);
nor U24794 (N_24794,N_18578,N_13556);
or U24795 (N_24795,N_15083,N_16114);
and U24796 (N_24796,N_15374,N_19106);
and U24797 (N_24797,N_19105,N_17446);
and U24798 (N_24798,N_14350,N_17750);
and U24799 (N_24799,N_15551,N_19627);
or U24800 (N_24800,N_17028,N_15536);
nand U24801 (N_24801,N_14061,N_18835);
and U24802 (N_24802,N_15946,N_17786);
nor U24803 (N_24803,N_11175,N_13723);
nor U24804 (N_24804,N_14354,N_12292);
or U24805 (N_24805,N_16092,N_12977);
or U24806 (N_24806,N_19439,N_12941);
and U24807 (N_24807,N_16972,N_11826);
nand U24808 (N_24808,N_16630,N_18540);
nor U24809 (N_24809,N_15241,N_16113);
nand U24810 (N_24810,N_16040,N_11231);
nor U24811 (N_24811,N_15707,N_19195);
nand U24812 (N_24812,N_17403,N_17450);
nor U24813 (N_24813,N_16087,N_18615);
nor U24814 (N_24814,N_15027,N_13700);
nor U24815 (N_24815,N_13044,N_12755);
nand U24816 (N_24816,N_11795,N_16106);
nand U24817 (N_24817,N_14298,N_17068);
xnor U24818 (N_24818,N_13135,N_12416);
or U24819 (N_24819,N_19787,N_10084);
and U24820 (N_24820,N_13531,N_18134);
or U24821 (N_24821,N_10997,N_18886);
and U24822 (N_24822,N_10586,N_17022);
and U24823 (N_24823,N_10085,N_13287);
and U24824 (N_24824,N_13869,N_17003);
nor U24825 (N_24825,N_18628,N_17013);
nor U24826 (N_24826,N_15235,N_13226);
or U24827 (N_24827,N_18581,N_13470);
and U24828 (N_24828,N_13026,N_15137);
or U24829 (N_24829,N_13465,N_16221);
or U24830 (N_24830,N_17263,N_13609);
nand U24831 (N_24831,N_15270,N_14297);
nand U24832 (N_24832,N_12701,N_11808);
or U24833 (N_24833,N_14656,N_16069);
or U24834 (N_24834,N_16100,N_12821);
and U24835 (N_24835,N_15246,N_12420);
nor U24836 (N_24836,N_17433,N_16392);
nand U24837 (N_24837,N_11918,N_14052);
and U24838 (N_24838,N_17218,N_10021);
xor U24839 (N_24839,N_11760,N_11438);
xor U24840 (N_24840,N_19674,N_11681);
or U24841 (N_24841,N_12220,N_15294);
nand U24842 (N_24842,N_14277,N_10528);
nand U24843 (N_24843,N_10416,N_11675);
nor U24844 (N_24844,N_10505,N_19759);
nand U24845 (N_24845,N_15869,N_14124);
and U24846 (N_24846,N_14863,N_14258);
xor U24847 (N_24847,N_17174,N_18710);
xor U24848 (N_24848,N_19037,N_18934);
xor U24849 (N_24849,N_12891,N_13242);
xnor U24850 (N_24850,N_13604,N_14949);
and U24851 (N_24851,N_12950,N_15207);
xnor U24852 (N_24852,N_18798,N_11016);
or U24853 (N_24853,N_10090,N_12410);
and U24854 (N_24854,N_10639,N_15900);
and U24855 (N_24855,N_16042,N_17772);
and U24856 (N_24856,N_18037,N_10184);
or U24857 (N_24857,N_15437,N_14479);
nor U24858 (N_24858,N_15339,N_13336);
nor U24859 (N_24859,N_16551,N_19685);
nor U24860 (N_24860,N_10323,N_10391);
or U24861 (N_24861,N_12326,N_11789);
and U24862 (N_24862,N_15020,N_12508);
nor U24863 (N_24863,N_18991,N_14897);
nand U24864 (N_24864,N_17543,N_19292);
and U24865 (N_24865,N_10871,N_12355);
nor U24866 (N_24866,N_16542,N_14220);
nor U24867 (N_24867,N_18716,N_13368);
nand U24868 (N_24868,N_12603,N_13354);
nand U24869 (N_24869,N_14434,N_17766);
xor U24870 (N_24870,N_12874,N_15615);
nand U24871 (N_24871,N_13270,N_12599);
nand U24872 (N_24872,N_18348,N_10879);
nand U24873 (N_24873,N_13297,N_16034);
nor U24874 (N_24874,N_19647,N_10271);
nor U24875 (N_24875,N_15851,N_14637);
and U24876 (N_24876,N_10816,N_14517);
nor U24877 (N_24877,N_15307,N_12307);
and U24878 (N_24878,N_10887,N_17309);
or U24879 (N_24879,N_17625,N_13040);
nor U24880 (N_24880,N_11224,N_12915);
and U24881 (N_24881,N_16362,N_17561);
xor U24882 (N_24882,N_15685,N_17562);
or U24883 (N_24883,N_19948,N_13459);
or U24884 (N_24884,N_12857,N_15661);
nor U24885 (N_24885,N_16239,N_16826);
or U24886 (N_24886,N_14158,N_12597);
nor U24887 (N_24887,N_17064,N_16297);
or U24888 (N_24888,N_17652,N_16896);
or U24889 (N_24889,N_18556,N_10506);
or U24890 (N_24890,N_15817,N_17858);
or U24891 (N_24891,N_11427,N_15628);
nor U24892 (N_24892,N_14190,N_13461);
nand U24893 (N_24893,N_15447,N_12735);
and U24894 (N_24894,N_14721,N_10406);
and U24895 (N_24895,N_11036,N_11862);
nor U24896 (N_24896,N_14940,N_19297);
xor U24897 (N_24897,N_17024,N_19952);
nand U24898 (N_24898,N_15280,N_18752);
nand U24899 (N_24899,N_11901,N_18486);
xor U24900 (N_24900,N_13515,N_12299);
and U24901 (N_24901,N_12327,N_12065);
nand U24902 (N_24902,N_14406,N_16249);
xor U24903 (N_24903,N_15873,N_10219);
or U24904 (N_24904,N_16938,N_11321);
and U24905 (N_24905,N_19552,N_10367);
nor U24906 (N_24906,N_10166,N_15562);
nor U24907 (N_24907,N_12266,N_15690);
nand U24908 (N_24908,N_10865,N_14197);
xnor U24909 (N_24909,N_15049,N_15433);
and U24910 (N_24910,N_19735,N_16334);
xnor U24911 (N_24911,N_14480,N_18095);
or U24912 (N_24912,N_14854,N_17747);
or U24913 (N_24913,N_15985,N_19570);
nand U24914 (N_24914,N_10908,N_15210);
nor U24915 (N_24915,N_14106,N_17882);
nor U24916 (N_24916,N_10489,N_17106);
nand U24917 (N_24917,N_15963,N_10842);
nor U24918 (N_24918,N_16407,N_18228);
or U24919 (N_24919,N_15847,N_16676);
or U24920 (N_24920,N_18102,N_15550);
and U24921 (N_24921,N_14730,N_13876);
nand U24922 (N_24922,N_19849,N_19020);
nand U24923 (N_24923,N_13233,N_14423);
nand U24924 (N_24924,N_19542,N_15448);
and U24925 (N_24925,N_12558,N_11264);
xor U24926 (N_24926,N_10196,N_15478);
and U24927 (N_24927,N_10714,N_17012);
and U24928 (N_24928,N_11003,N_15943);
or U24929 (N_24929,N_19963,N_15209);
nor U24930 (N_24930,N_19786,N_10444);
nor U24931 (N_24931,N_15511,N_12095);
nor U24932 (N_24932,N_18223,N_17465);
or U24933 (N_24933,N_18529,N_14301);
or U24934 (N_24934,N_11940,N_14147);
or U24935 (N_24935,N_13925,N_19774);
and U24936 (N_24936,N_15666,N_13572);
or U24937 (N_24937,N_19363,N_13922);
nor U24938 (N_24938,N_17057,N_10289);
nor U24939 (N_24939,N_12112,N_15046);
xnor U24940 (N_24940,N_15620,N_15390);
or U24941 (N_24941,N_15459,N_18735);
xnor U24942 (N_24942,N_18194,N_18274);
nand U24943 (N_24943,N_17681,N_12534);
and U24944 (N_24944,N_11477,N_16000);
or U24945 (N_24945,N_17761,N_15653);
nor U24946 (N_24946,N_19219,N_14070);
or U24947 (N_24947,N_17393,N_17666);
and U24948 (N_24948,N_11400,N_16713);
nand U24949 (N_24949,N_15996,N_13244);
or U24950 (N_24950,N_10754,N_11099);
nand U24951 (N_24951,N_10958,N_10469);
nor U24952 (N_24952,N_15593,N_13282);
or U24953 (N_24953,N_13355,N_10545);
nor U24954 (N_24954,N_14709,N_16840);
nand U24955 (N_24955,N_13484,N_12380);
xnor U24956 (N_24956,N_14946,N_12130);
and U24957 (N_24957,N_15514,N_11621);
nor U24958 (N_24958,N_17167,N_18550);
xor U24959 (N_24959,N_13218,N_17113);
and U24960 (N_24960,N_13123,N_17342);
nand U24961 (N_24961,N_11626,N_14323);
nand U24962 (N_24962,N_16602,N_14154);
nor U24963 (N_24963,N_10662,N_14405);
nor U24964 (N_24964,N_17154,N_17927);
nand U24965 (N_24965,N_18339,N_11952);
or U24966 (N_24966,N_19352,N_12774);
or U24967 (N_24967,N_11849,N_12155);
and U24968 (N_24968,N_19971,N_16475);
and U24969 (N_24969,N_15276,N_12810);
or U24970 (N_24970,N_17332,N_11712);
or U24971 (N_24971,N_19245,N_11561);
and U24972 (N_24972,N_13936,N_15171);
xnor U24973 (N_24973,N_18972,N_17696);
or U24974 (N_24974,N_16143,N_16094);
or U24975 (N_24975,N_12816,N_19535);
nand U24976 (N_24976,N_15160,N_15738);
or U24977 (N_24977,N_12298,N_14699);
and U24978 (N_24978,N_17095,N_15066);
nand U24979 (N_24979,N_10065,N_10791);
nand U24980 (N_24980,N_16578,N_17026);
or U24981 (N_24981,N_10678,N_17639);
xnor U24982 (N_24982,N_12349,N_14858);
nand U24983 (N_24983,N_14755,N_19057);
xnor U24984 (N_24984,N_16121,N_10649);
nand U24985 (N_24985,N_14834,N_14935);
and U24986 (N_24986,N_19496,N_18259);
nor U24987 (N_24987,N_13194,N_18521);
nor U24988 (N_24988,N_11244,N_13823);
nor U24989 (N_24989,N_13644,N_12431);
nor U24990 (N_24990,N_12116,N_17999);
nand U24991 (N_24991,N_14819,N_11599);
nand U24992 (N_24992,N_18330,N_19434);
and U24993 (N_24993,N_16746,N_11889);
nor U24994 (N_24994,N_19776,N_19852);
nand U24995 (N_24995,N_11280,N_15911);
or U24996 (N_24996,N_19198,N_19447);
nand U24997 (N_24997,N_14163,N_10830);
nand U24998 (N_24998,N_15009,N_13944);
nor U24999 (N_24999,N_15694,N_10673);
and U25000 (N_25000,N_14064,N_12003);
and U25001 (N_25001,N_13545,N_11436);
nand U25002 (N_25002,N_17896,N_14040);
nand U25003 (N_25003,N_14699,N_19256);
nor U25004 (N_25004,N_14740,N_15510);
nor U25005 (N_25005,N_18621,N_11910);
nand U25006 (N_25006,N_17436,N_11333);
nor U25007 (N_25007,N_14673,N_12008);
xnor U25008 (N_25008,N_17924,N_14507);
nor U25009 (N_25009,N_18794,N_11742);
nor U25010 (N_25010,N_10052,N_19427);
and U25011 (N_25011,N_19076,N_18742);
nor U25012 (N_25012,N_17625,N_12097);
nand U25013 (N_25013,N_18223,N_19837);
or U25014 (N_25014,N_14071,N_13451);
or U25015 (N_25015,N_17670,N_13185);
and U25016 (N_25016,N_16915,N_17631);
nand U25017 (N_25017,N_18036,N_12664);
nand U25018 (N_25018,N_18461,N_13179);
or U25019 (N_25019,N_14645,N_16086);
nor U25020 (N_25020,N_15545,N_10889);
nand U25021 (N_25021,N_18587,N_15106);
or U25022 (N_25022,N_16880,N_10049);
nor U25023 (N_25023,N_17407,N_16268);
and U25024 (N_25024,N_13966,N_12816);
nand U25025 (N_25025,N_12576,N_14677);
or U25026 (N_25026,N_19338,N_18971);
nor U25027 (N_25027,N_11736,N_16917);
and U25028 (N_25028,N_19753,N_14318);
nand U25029 (N_25029,N_12658,N_19769);
nor U25030 (N_25030,N_15899,N_11412);
nand U25031 (N_25031,N_12511,N_15027);
nor U25032 (N_25032,N_11808,N_14014);
or U25033 (N_25033,N_17465,N_17495);
or U25034 (N_25034,N_14416,N_13639);
nand U25035 (N_25035,N_17345,N_17374);
and U25036 (N_25036,N_16293,N_17208);
nand U25037 (N_25037,N_10307,N_15397);
nor U25038 (N_25038,N_16320,N_15066);
nand U25039 (N_25039,N_16120,N_19006);
or U25040 (N_25040,N_15790,N_11802);
nand U25041 (N_25041,N_10628,N_10249);
or U25042 (N_25042,N_14683,N_17711);
nand U25043 (N_25043,N_17543,N_16029);
or U25044 (N_25044,N_15247,N_14705);
nand U25045 (N_25045,N_12731,N_14034);
nand U25046 (N_25046,N_12915,N_17668);
or U25047 (N_25047,N_18528,N_12752);
or U25048 (N_25048,N_15914,N_18770);
nor U25049 (N_25049,N_16369,N_19137);
nand U25050 (N_25050,N_13283,N_12931);
and U25051 (N_25051,N_16543,N_16036);
nor U25052 (N_25052,N_10281,N_13001);
xor U25053 (N_25053,N_13311,N_15215);
nor U25054 (N_25054,N_16472,N_13363);
nor U25055 (N_25055,N_14684,N_14815);
and U25056 (N_25056,N_19122,N_10905);
nor U25057 (N_25057,N_16337,N_19241);
nand U25058 (N_25058,N_10816,N_11002);
xnor U25059 (N_25059,N_16517,N_15043);
nor U25060 (N_25060,N_13619,N_16908);
and U25061 (N_25061,N_13363,N_13261);
and U25062 (N_25062,N_14912,N_15987);
and U25063 (N_25063,N_13786,N_11097);
nand U25064 (N_25064,N_13769,N_12795);
nor U25065 (N_25065,N_11554,N_18737);
xor U25066 (N_25066,N_13336,N_12473);
nand U25067 (N_25067,N_14887,N_15840);
nand U25068 (N_25068,N_17531,N_18129);
and U25069 (N_25069,N_16310,N_14452);
nand U25070 (N_25070,N_10201,N_14428);
or U25071 (N_25071,N_15601,N_11917);
xor U25072 (N_25072,N_18888,N_18720);
nand U25073 (N_25073,N_10569,N_14253);
nand U25074 (N_25074,N_19266,N_16405);
nor U25075 (N_25075,N_12964,N_12935);
nor U25076 (N_25076,N_15927,N_11640);
xor U25077 (N_25077,N_15692,N_12103);
nand U25078 (N_25078,N_11190,N_13907);
nor U25079 (N_25079,N_19271,N_13209);
nor U25080 (N_25080,N_13096,N_15268);
nor U25081 (N_25081,N_10063,N_18391);
or U25082 (N_25082,N_19037,N_12328);
nor U25083 (N_25083,N_19795,N_18984);
nor U25084 (N_25084,N_19223,N_16169);
nand U25085 (N_25085,N_13041,N_16342);
and U25086 (N_25086,N_13854,N_16110);
nand U25087 (N_25087,N_17185,N_18762);
or U25088 (N_25088,N_13960,N_12491);
or U25089 (N_25089,N_13192,N_18309);
or U25090 (N_25090,N_16106,N_17658);
and U25091 (N_25091,N_13337,N_13220);
nand U25092 (N_25092,N_17276,N_11482);
nor U25093 (N_25093,N_13061,N_11424);
nor U25094 (N_25094,N_10205,N_19318);
nand U25095 (N_25095,N_10856,N_19807);
or U25096 (N_25096,N_13750,N_14898);
and U25097 (N_25097,N_15509,N_17601);
or U25098 (N_25098,N_15826,N_17847);
nand U25099 (N_25099,N_15980,N_10500);
xnor U25100 (N_25100,N_15382,N_19888);
nor U25101 (N_25101,N_11828,N_11025);
xor U25102 (N_25102,N_13545,N_12492);
and U25103 (N_25103,N_17280,N_19278);
xnor U25104 (N_25104,N_14576,N_14290);
nor U25105 (N_25105,N_14237,N_15638);
and U25106 (N_25106,N_16645,N_10009);
or U25107 (N_25107,N_18771,N_18974);
and U25108 (N_25108,N_10426,N_13562);
nand U25109 (N_25109,N_13315,N_13057);
nor U25110 (N_25110,N_13376,N_10831);
nor U25111 (N_25111,N_12307,N_11462);
nand U25112 (N_25112,N_16702,N_14352);
nor U25113 (N_25113,N_17832,N_10351);
nor U25114 (N_25114,N_14850,N_16106);
nor U25115 (N_25115,N_15158,N_10347);
nand U25116 (N_25116,N_12979,N_17023);
nor U25117 (N_25117,N_18126,N_11497);
xor U25118 (N_25118,N_19521,N_11927);
nor U25119 (N_25119,N_12169,N_18083);
or U25120 (N_25120,N_12826,N_19732);
or U25121 (N_25121,N_19360,N_18100);
and U25122 (N_25122,N_19484,N_19450);
or U25123 (N_25123,N_13040,N_14474);
or U25124 (N_25124,N_16493,N_15132);
or U25125 (N_25125,N_14173,N_14008);
nor U25126 (N_25126,N_19183,N_12874);
nor U25127 (N_25127,N_10790,N_12865);
and U25128 (N_25128,N_19260,N_19389);
nand U25129 (N_25129,N_14742,N_16911);
and U25130 (N_25130,N_16129,N_12296);
nand U25131 (N_25131,N_11995,N_19584);
nand U25132 (N_25132,N_18431,N_19726);
nor U25133 (N_25133,N_18552,N_10315);
nand U25134 (N_25134,N_12041,N_19901);
or U25135 (N_25135,N_14686,N_10265);
or U25136 (N_25136,N_13479,N_14107);
nand U25137 (N_25137,N_11994,N_15519);
or U25138 (N_25138,N_17133,N_17763);
and U25139 (N_25139,N_12484,N_15750);
and U25140 (N_25140,N_12184,N_10541);
nand U25141 (N_25141,N_17646,N_15178);
and U25142 (N_25142,N_12170,N_14643);
and U25143 (N_25143,N_12529,N_10741);
nor U25144 (N_25144,N_11754,N_16874);
nor U25145 (N_25145,N_19538,N_16174);
nor U25146 (N_25146,N_10117,N_18375);
nor U25147 (N_25147,N_10875,N_14101);
nor U25148 (N_25148,N_12747,N_19497);
and U25149 (N_25149,N_10482,N_17064);
or U25150 (N_25150,N_11689,N_19974);
or U25151 (N_25151,N_10656,N_17866);
and U25152 (N_25152,N_10652,N_11140);
and U25153 (N_25153,N_13114,N_10951);
or U25154 (N_25154,N_11749,N_15471);
xor U25155 (N_25155,N_17871,N_15471);
nor U25156 (N_25156,N_13072,N_19260);
nand U25157 (N_25157,N_18275,N_19520);
nor U25158 (N_25158,N_10206,N_10864);
or U25159 (N_25159,N_12178,N_10289);
nand U25160 (N_25160,N_11917,N_18802);
xor U25161 (N_25161,N_14374,N_17985);
and U25162 (N_25162,N_18298,N_18316);
nor U25163 (N_25163,N_19172,N_16096);
nor U25164 (N_25164,N_17683,N_17254);
nand U25165 (N_25165,N_16684,N_11647);
nand U25166 (N_25166,N_16101,N_18848);
and U25167 (N_25167,N_16828,N_12777);
nor U25168 (N_25168,N_19396,N_16238);
nand U25169 (N_25169,N_18379,N_18497);
or U25170 (N_25170,N_12794,N_16780);
nor U25171 (N_25171,N_11378,N_14978);
nor U25172 (N_25172,N_11200,N_16880);
nor U25173 (N_25173,N_13558,N_10385);
nand U25174 (N_25174,N_11239,N_16526);
nor U25175 (N_25175,N_18923,N_10351);
nor U25176 (N_25176,N_17604,N_17172);
and U25177 (N_25177,N_10943,N_19109);
and U25178 (N_25178,N_17373,N_19395);
and U25179 (N_25179,N_16262,N_11235);
or U25180 (N_25180,N_16291,N_16689);
xnor U25181 (N_25181,N_16165,N_10922);
or U25182 (N_25182,N_13943,N_19883);
and U25183 (N_25183,N_19213,N_14683);
nand U25184 (N_25184,N_19764,N_14611);
and U25185 (N_25185,N_17922,N_12912);
xor U25186 (N_25186,N_14449,N_12601);
nor U25187 (N_25187,N_14203,N_15257);
nor U25188 (N_25188,N_10680,N_11278);
or U25189 (N_25189,N_19072,N_13513);
nor U25190 (N_25190,N_16150,N_18990);
nand U25191 (N_25191,N_13247,N_14226);
nand U25192 (N_25192,N_19340,N_13424);
and U25193 (N_25193,N_14499,N_12680);
nor U25194 (N_25194,N_16347,N_15013);
or U25195 (N_25195,N_12039,N_10720);
or U25196 (N_25196,N_19786,N_15486);
or U25197 (N_25197,N_15176,N_13519);
nand U25198 (N_25198,N_12002,N_16234);
or U25199 (N_25199,N_12311,N_11013);
xor U25200 (N_25200,N_19141,N_19121);
nor U25201 (N_25201,N_15372,N_18095);
or U25202 (N_25202,N_18258,N_11412);
nor U25203 (N_25203,N_17287,N_15920);
or U25204 (N_25204,N_19894,N_10987);
nor U25205 (N_25205,N_19989,N_17784);
nand U25206 (N_25206,N_15158,N_11366);
or U25207 (N_25207,N_13857,N_12223);
nand U25208 (N_25208,N_16496,N_12727);
nand U25209 (N_25209,N_14016,N_13542);
nand U25210 (N_25210,N_14163,N_19526);
and U25211 (N_25211,N_13516,N_10242);
nor U25212 (N_25212,N_13959,N_19016);
xnor U25213 (N_25213,N_16402,N_15925);
and U25214 (N_25214,N_13789,N_11343);
nand U25215 (N_25215,N_12602,N_19699);
xnor U25216 (N_25216,N_18128,N_13225);
or U25217 (N_25217,N_15183,N_18521);
or U25218 (N_25218,N_19937,N_16409);
and U25219 (N_25219,N_17941,N_13721);
or U25220 (N_25220,N_11742,N_13974);
or U25221 (N_25221,N_12084,N_13003);
nand U25222 (N_25222,N_18065,N_11754);
and U25223 (N_25223,N_12279,N_13570);
nand U25224 (N_25224,N_14925,N_17546);
xor U25225 (N_25225,N_10331,N_12090);
or U25226 (N_25226,N_17731,N_10893);
nor U25227 (N_25227,N_18061,N_12456);
and U25228 (N_25228,N_15257,N_12907);
nor U25229 (N_25229,N_14743,N_13097);
nor U25230 (N_25230,N_11309,N_12080);
or U25231 (N_25231,N_15147,N_15792);
and U25232 (N_25232,N_12912,N_16553);
xnor U25233 (N_25233,N_11266,N_15695);
and U25234 (N_25234,N_14459,N_18109);
or U25235 (N_25235,N_11456,N_11024);
and U25236 (N_25236,N_11047,N_10090);
nor U25237 (N_25237,N_15652,N_10662);
nor U25238 (N_25238,N_17229,N_11394);
nand U25239 (N_25239,N_12758,N_13223);
nor U25240 (N_25240,N_16957,N_19526);
nor U25241 (N_25241,N_10343,N_15908);
or U25242 (N_25242,N_11862,N_19363);
nand U25243 (N_25243,N_19725,N_19388);
xor U25244 (N_25244,N_18346,N_16435);
nand U25245 (N_25245,N_15039,N_19289);
and U25246 (N_25246,N_10063,N_14643);
or U25247 (N_25247,N_15260,N_16001);
nand U25248 (N_25248,N_19039,N_19318);
and U25249 (N_25249,N_16834,N_16358);
and U25250 (N_25250,N_19976,N_19503);
or U25251 (N_25251,N_19533,N_17492);
xor U25252 (N_25252,N_18955,N_13170);
and U25253 (N_25253,N_15838,N_19458);
and U25254 (N_25254,N_12722,N_19312);
nor U25255 (N_25255,N_18838,N_16961);
and U25256 (N_25256,N_17113,N_19757);
nand U25257 (N_25257,N_19726,N_12829);
nor U25258 (N_25258,N_10463,N_14587);
and U25259 (N_25259,N_17259,N_17103);
nand U25260 (N_25260,N_13834,N_14644);
nand U25261 (N_25261,N_17422,N_16613);
nor U25262 (N_25262,N_12332,N_10494);
nor U25263 (N_25263,N_13505,N_10940);
nor U25264 (N_25264,N_18233,N_16706);
nand U25265 (N_25265,N_14989,N_18706);
nand U25266 (N_25266,N_14119,N_12840);
and U25267 (N_25267,N_14366,N_13107);
xor U25268 (N_25268,N_13235,N_12339);
xor U25269 (N_25269,N_12082,N_13424);
or U25270 (N_25270,N_18989,N_13991);
nand U25271 (N_25271,N_19551,N_18953);
nand U25272 (N_25272,N_19270,N_16479);
nor U25273 (N_25273,N_14613,N_17848);
and U25274 (N_25274,N_15744,N_18689);
nand U25275 (N_25275,N_15928,N_17331);
and U25276 (N_25276,N_18541,N_18992);
nor U25277 (N_25277,N_15352,N_19614);
or U25278 (N_25278,N_15523,N_10072);
xor U25279 (N_25279,N_16175,N_18877);
nand U25280 (N_25280,N_13539,N_19126);
nand U25281 (N_25281,N_11281,N_11627);
nor U25282 (N_25282,N_11436,N_16548);
nor U25283 (N_25283,N_14232,N_15100);
and U25284 (N_25284,N_17621,N_19009);
nor U25285 (N_25285,N_13344,N_17667);
nand U25286 (N_25286,N_10179,N_18060);
nor U25287 (N_25287,N_14745,N_18814);
nand U25288 (N_25288,N_16006,N_12194);
xor U25289 (N_25289,N_16956,N_10050);
nor U25290 (N_25290,N_14930,N_16498);
xor U25291 (N_25291,N_18323,N_17951);
nor U25292 (N_25292,N_19363,N_11064);
nor U25293 (N_25293,N_18513,N_10436);
nor U25294 (N_25294,N_10389,N_11298);
or U25295 (N_25295,N_16111,N_11371);
and U25296 (N_25296,N_10283,N_17787);
nor U25297 (N_25297,N_17126,N_13149);
or U25298 (N_25298,N_17373,N_15679);
nor U25299 (N_25299,N_15383,N_10842);
or U25300 (N_25300,N_11905,N_10738);
xor U25301 (N_25301,N_18789,N_10940);
nand U25302 (N_25302,N_16790,N_17130);
nor U25303 (N_25303,N_14278,N_18021);
and U25304 (N_25304,N_16645,N_17399);
nor U25305 (N_25305,N_15715,N_10003);
nand U25306 (N_25306,N_10536,N_12641);
or U25307 (N_25307,N_12269,N_17109);
and U25308 (N_25308,N_18006,N_18045);
or U25309 (N_25309,N_12387,N_11679);
or U25310 (N_25310,N_14964,N_15677);
nor U25311 (N_25311,N_13025,N_15116);
xnor U25312 (N_25312,N_11321,N_13541);
nand U25313 (N_25313,N_11060,N_17118);
nor U25314 (N_25314,N_16987,N_11899);
nand U25315 (N_25315,N_19455,N_18024);
nor U25316 (N_25316,N_14139,N_17370);
nand U25317 (N_25317,N_13404,N_11591);
nor U25318 (N_25318,N_16180,N_19040);
nor U25319 (N_25319,N_14869,N_16654);
nor U25320 (N_25320,N_11008,N_15475);
and U25321 (N_25321,N_11565,N_13511);
and U25322 (N_25322,N_13220,N_15349);
nand U25323 (N_25323,N_14437,N_19673);
nor U25324 (N_25324,N_10486,N_19360);
and U25325 (N_25325,N_19610,N_18376);
xor U25326 (N_25326,N_17289,N_15258);
and U25327 (N_25327,N_16666,N_19486);
nor U25328 (N_25328,N_17274,N_10441);
xnor U25329 (N_25329,N_14189,N_17828);
or U25330 (N_25330,N_15444,N_14314);
nand U25331 (N_25331,N_15957,N_18426);
or U25332 (N_25332,N_16574,N_12763);
or U25333 (N_25333,N_17911,N_16152);
xor U25334 (N_25334,N_12852,N_10166);
and U25335 (N_25335,N_17138,N_10386);
nand U25336 (N_25336,N_12113,N_10389);
xnor U25337 (N_25337,N_17085,N_14282);
nand U25338 (N_25338,N_14908,N_16227);
and U25339 (N_25339,N_10607,N_19697);
or U25340 (N_25340,N_14700,N_15743);
nand U25341 (N_25341,N_19162,N_19185);
and U25342 (N_25342,N_18229,N_11960);
nor U25343 (N_25343,N_14686,N_17136);
nand U25344 (N_25344,N_14987,N_13442);
or U25345 (N_25345,N_11472,N_15078);
and U25346 (N_25346,N_17976,N_16852);
or U25347 (N_25347,N_10307,N_12920);
xnor U25348 (N_25348,N_12611,N_16015);
and U25349 (N_25349,N_14715,N_11871);
nand U25350 (N_25350,N_16976,N_19553);
and U25351 (N_25351,N_11510,N_15256);
and U25352 (N_25352,N_12071,N_12097);
nor U25353 (N_25353,N_12269,N_14043);
nand U25354 (N_25354,N_12867,N_19372);
nand U25355 (N_25355,N_11539,N_19013);
and U25356 (N_25356,N_17014,N_14587);
nand U25357 (N_25357,N_18312,N_19615);
nand U25358 (N_25358,N_15465,N_12765);
nor U25359 (N_25359,N_17662,N_13073);
nor U25360 (N_25360,N_17245,N_19509);
and U25361 (N_25361,N_11644,N_16965);
or U25362 (N_25362,N_10629,N_11627);
and U25363 (N_25363,N_18616,N_11439);
nand U25364 (N_25364,N_18705,N_13617);
xor U25365 (N_25365,N_13943,N_11290);
or U25366 (N_25366,N_19399,N_15444);
nor U25367 (N_25367,N_18813,N_11722);
and U25368 (N_25368,N_14898,N_11492);
or U25369 (N_25369,N_12681,N_10668);
or U25370 (N_25370,N_11153,N_13773);
nand U25371 (N_25371,N_18682,N_14238);
nand U25372 (N_25372,N_14543,N_12846);
and U25373 (N_25373,N_12271,N_19550);
nor U25374 (N_25374,N_19985,N_11166);
nand U25375 (N_25375,N_14741,N_16715);
nor U25376 (N_25376,N_16607,N_12143);
nor U25377 (N_25377,N_14822,N_16873);
and U25378 (N_25378,N_18201,N_14165);
nand U25379 (N_25379,N_15311,N_15191);
nand U25380 (N_25380,N_16490,N_18195);
nor U25381 (N_25381,N_12391,N_12461);
nand U25382 (N_25382,N_10127,N_12023);
nor U25383 (N_25383,N_17728,N_13802);
or U25384 (N_25384,N_13498,N_14586);
and U25385 (N_25385,N_16386,N_19598);
nor U25386 (N_25386,N_10585,N_12199);
or U25387 (N_25387,N_16037,N_10417);
nor U25388 (N_25388,N_18585,N_17604);
or U25389 (N_25389,N_19147,N_13193);
or U25390 (N_25390,N_14311,N_17859);
or U25391 (N_25391,N_13714,N_12503);
or U25392 (N_25392,N_17188,N_13796);
xnor U25393 (N_25393,N_14405,N_15168);
nor U25394 (N_25394,N_19289,N_14342);
or U25395 (N_25395,N_17321,N_13260);
nand U25396 (N_25396,N_11566,N_19075);
nand U25397 (N_25397,N_17050,N_18961);
and U25398 (N_25398,N_11530,N_15895);
nor U25399 (N_25399,N_18066,N_15026);
and U25400 (N_25400,N_13211,N_16052);
nor U25401 (N_25401,N_17085,N_17291);
nand U25402 (N_25402,N_19219,N_13788);
nor U25403 (N_25403,N_15340,N_10119);
nand U25404 (N_25404,N_10832,N_19249);
nor U25405 (N_25405,N_13790,N_11595);
and U25406 (N_25406,N_14862,N_10550);
nand U25407 (N_25407,N_19809,N_13008);
nand U25408 (N_25408,N_19416,N_16239);
or U25409 (N_25409,N_12739,N_11939);
xnor U25410 (N_25410,N_19869,N_11725);
nor U25411 (N_25411,N_19934,N_12690);
or U25412 (N_25412,N_15607,N_14041);
nand U25413 (N_25413,N_19811,N_18114);
or U25414 (N_25414,N_18453,N_17203);
nand U25415 (N_25415,N_11985,N_19145);
xnor U25416 (N_25416,N_10633,N_16275);
or U25417 (N_25417,N_10433,N_17041);
nand U25418 (N_25418,N_17640,N_16448);
nor U25419 (N_25419,N_14734,N_19188);
nand U25420 (N_25420,N_10116,N_16984);
nor U25421 (N_25421,N_12568,N_13854);
nor U25422 (N_25422,N_15670,N_18412);
nor U25423 (N_25423,N_14239,N_17983);
nor U25424 (N_25424,N_13694,N_12744);
nand U25425 (N_25425,N_13909,N_16019);
nand U25426 (N_25426,N_18068,N_17496);
nand U25427 (N_25427,N_15107,N_19817);
nand U25428 (N_25428,N_13473,N_16527);
nor U25429 (N_25429,N_16950,N_13721);
nor U25430 (N_25430,N_12016,N_16449);
nand U25431 (N_25431,N_18562,N_10289);
nand U25432 (N_25432,N_18617,N_16368);
or U25433 (N_25433,N_13375,N_12980);
or U25434 (N_25434,N_10424,N_15166);
nor U25435 (N_25435,N_17377,N_12029);
nor U25436 (N_25436,N_13742,N_13675);
and U25437 (N_25437,N_13783,N_10033);
and U25438 (N_25438,N_11821,N_18518);
or U25439 (N_25439,N_16630,N_16503);
nor U25440 (N_25440,N_16521,N_18751);
or U25441 (N_25441,N_13001,N_14759);
nor U25442 (N_25442,N_12574,N_14536);
nand U25443 (N_25443,N_14562,N_19961);
xor U25444 (N_25444,N_16990,N_18334);
xnor U25445 (N_25445,N_19041,N_15442);
and U25446 (N_25446,N_10452,N_13346);
nand U25447 (N_25447,N_16806,N_16769);
and U25448 (N_25448,N_17978,N_15597);
nand U25449 (N_25449,N_14589,N_10239);
nor U25450 (N_25450,N_16266,N_14681);
and U25451 (N_25451,N_15348,N_16411);
nand U25452 (N_25452,N_17935,N_10931);
nor U25453 (N_25453,N_18701,N_10153);
or U25454 (N_25454,N_12316,N_11135);
nand U25455 (N_25455,N_13269,N_12871);
and U25456 (N_25456,N_11869,N_12924);
nor U25457 (N_25457,N_12228,N_18259);
nand U25458 (N_25458,N_14958,N_19902);
nor U25459 (N_25459,N_18056,N_17478);
xor U25460 (N_25460,N_13471,N_13753);
nand U25461 (N_25461,N_13868,N_10870);
nor U25462 (N_25462,N_11572,N_16029);
or U25463 (N_25463,N_13058,N_17358);
xor U25464 (N_25464,N_16430,N_13955);
or U25465 (N_25465,N_19955,N_19756);
nor U25466 (N_25466,N_12228,N_14833);
nand U25467 (N_25467,N_19267,N_18566);
and U25468 (N_25468,N_19813,N_11726);
or U25469 (N_25469,N_10995,N_16574);
nand U25470 (N_25470,N_13733,N_19912);
or U25471 (N_25471,N_18971,N_18956);
and U25472 (N_25472,N_13168,N_19122);
nor U25473 (N_25473,N_15168,N_17754);
and U25474 (N_25474,N_11396,N_15805);
or U25475 (N_25475,N_19115,N_15292);
or U25476 (N_25476,N_14639,N_10376);
and U25477 (N_25477,N_17672,N_15535);
nand U25478 (N_25478,N_11225,N_12385);
nand U25479 (N_25479,N_12357,N_18162);
nor U25480 (N_25480,N_14945,N_19733);
nand U25481 (N_25481,N_18838,N_11744);
or U25482 (N_25482,N_11003,N_13009);
nand U25483 (N_25483,N_19734,N_11139);
xnor U25484 (N_25484,N_13755,N_14225);
and U25485 (N_25485,N_15800,N_16970);
nor U25486 (N_25486,N_18556,N_13346);
nand U25487 (N_25487,N_14583,N_14604);
or U25488 (N_25488,N_16371,N_17532);
xor U25489 (N_25489,N_18301,N_11281);
nand U25490 (N_25490,N_14494,N_13447);
nor U25491 (N_25491,N_19992,N_14624);
or U25492 (N_25492,N_16426,N_13183);
nor U25493 (N_25493,N_13499,N_14647);
nor U25494 (N_25494,N_10628,N_12079);
nor U25495 (N_25495,N_12996,N_14152);
or U25496 (N_25496,N_15276,N_17443);
or U25497 (N_25497,N_10571,N_11298);
xnor U25498 (N_25498,N_18335,N_10397);
nand U25499 (N_25499,N_14928,N_15826);
and U25500 (N_25500,N_14758,N_16984);
and U25501 (N_25501,N_17850,N_17343);
nand U25502 (N_25502,N_13067,N_15023);
nand U25503 (N_25503,N_14095,N_16486);
xor U25504 (N_25504,N_19434,N_10920);
and U25505 (N_25505,N_15872,N_12096);
and U25506 (N_25506,N_16194,N_14336);
and U25507 (N_25507,N_16650,N_19162);
and U25508 (N_25508,N_16042,N_13140);
and U25509 (N_25509,N_17758,N_19854);
or U25510 (N_25510,N_17885,N_13668);
nor U25511 (N_25511,N_18728,N_16167);
nor U25512 (N_25512,N_19533,N_12180);
nor U25513 (N_25513,N_19487,N_11328);
and U25514 (N_25514,N_11788,N_15312);
nand U25515 (N_25515,N_16079,N_14265);
and U25516 (N_25516,N_11401,N_13367);
and U25517 (N_25517,N_11064,N_13694);
and U25518 (N_25518,N_13055,N_10571);
nand U25519 (N_25519,N_10936,N_15489);
nand U25520 (N_25520,N_18917,N_16793);
nor U25521 (N_25521,N_16197,N_12945);
nand U25522 (N_25522,N_16715,N_19026);
nor U25523 (N_25523,N_13775,N_16281);
nor U25524 (N_25524,N_17899,N_15567);
nand U25525 (N_25525,N_17853,N_11412);
nor U25526 (N_25526,N_15428,N_18735);
or U25527 (N_25527,N_19687,N_19752);
nand U25528 (N_25528,N_11109,N_17398);
nor U25529 (N_25529,N_18447,N_11886);
or U25530 (N_25530,N_17817,N_13979);
or U25531 (N_25531,N_11924,N_13346);
and U25532 (N_25532,N_10399,N_17060);
and U25533 (N_25533,N_17395,N_16601);
nand U25534 (N_25534,N_17738,N_11473);
or U25535 (N_25535,N_11791,N_17010);
and U25536 (N_25536,N_11940,N_14662);
nor U25537 (N_25537,N_10141,N_10870);
nor U25538 (N_25538,N_17401,N_19609);
and U25539 (N_25539,N_15415,N_13663);
nand U25540 (N_25540,N_19393,N_10010);
nor U25541 (N_25541,N_10520,N_17622);
or U25542 (N_25542,N_18520,N_12192);
nor U25543 (N_25543,N_13328,N_16476);
nand U25544 (N_25544,N_12075,N_16159);
nor U25545 (N_25545,N_15812,N_15062);
nand U25546 (N_25546,N_15123,N_16242);
xnor U25547 (N_25547,N_10277,N_10006);
nor U25548 (N_25548,N_14537,N_18024);
nor U25549 (N_25549,N_15087,N_10814);
and U25550 (N_25550,N_14962,N_11385);
and U25551 (N_25551,N_19761,N_15798);
and U25552 (N_25552,N_18058,N_16934);
and U25553 (N_25553,N_17878,N_10113);
or U25554 (N_25554,N_13811,N_12398);
and U25555 (N_25555,N_10677,N_16250);
or U25556 (N_25556,N_16828,N_16406);
nor U25557 (N_25557,N_13125,N_16758);
nor U25558 (N_25558,N_11609,N_17660);
or U25559 (N_25559,N_15986,N_17916);
nand U25560 (N_25560,N_11733,N_16249);
or U25561 (N_25561,N_15595,N_10417);
nor U25562 (N_25562,N_11934,N_14571);
nand U25563 (N_25563,N_14432,N_14928);
nor U25564 (N_25564,N_17203,N_14545);
nand U25565 (N_25565,N_17063,N_17039);
xor U25566 (N_25566,N_16427,N_16882);
nor U25567 (N_25567,N_18765,N_10249);
or U25568 (N_25568,N_13746,N_16811);
xor U25569 (N_25569,N_16326,N_14580);
and U25570 (N_25570,N_17412,N_19919);
nand U25571 (N_25571,N_11170,N_13424);
nor U25572 (N_25572,N_16330,N_17274);
xnor U25573 (N_25573,N_14506,N_15281);
nor U25574 (N_25574,N_10396,N_15195);
nand U25575 (N_25575,N_10664,N_13585);
or U25576 (N_25576,N_11415,N_18779);
xor U25577 (N_25577,N_11992,N_16874);
nor U25578 (N_25578,N_15021,N_14607);
or U25579 (N_25579,N_10323,N_11206);
and U25580 (N_25580,N_16606,N_11119);
and U25581 (N_25581,N_15175,N_15042);
xor U25582 (N_25582,N_19609,N_19352);
nand U25583 (N_25583,N_11224,N_10009);
xnor U25584 (N_25584,N_17992,N_18649);
nor U25585 (N_25585,N_13612,N_10978);
xor U25586 (N_25586,N_13698,N_12380);
nor U25587 (N_25587,N_18405,N_14937);
nor U25588 (N_25588,N_12826,N_18123);
xor U25589 (N_25589,N_13508,N_14334);
nand U25590 (N_25590,N_17537,N_13099);
nand U25591 (N_25591,N_18295,N_19708);
nor U25592 (N_25592,N_11385,N_15952);
nor U25593 (N_25593,N_15772,N_12625);
and U25594 (N_25594,N_11664,N_15067);
or U25595 (N_25595,N_16802,N_12789);
xnor U25596 (N_25596,N_15549,N_18356);
and U25597 (N_25597,N_17993,N_12774);
and U25598 (N_25598,N_15189,N_13196);
nor U25599 (N_25599,N_14117,N_15998);
or U25600 (N_25600,N_12811,N_16486);
nand U25601 (N_25601,N_17544,N_13849);
nor U25602 (N_25602,N_19730,N_10341);
xnor U25603 (N_25603,N_13302,N_15043);
or U25604 (N_25604,N_19253,N_14399);
or U25605 (N_25605,N_10288,N_16944);
nor U25606 (N_25606,N_17968,N_15226);
nand U25607 (N_25607,N_15631,N_16862);
or U25608 (N_25608,N_13008,N_18023);
xor U25609 (N_25609,N_12040,N_18810);
xor U25610 (N_25610,N_17707,N_17109);
nor U25611 (N_25611,N_14558,N_12109);
and U25612 (N_25612,N_18713,N_10763);
nand U25613 (N_25613,N_14650,N_17055);
and U25614 (N_25614,N_19150,N_12837);
nor U25615 (N_25615,N_19913,N_11171);
and U25616 (N_25616,N_19730,N_16924);
or U25617 (N_25617,N_18406,N_10045);
nand U25618 (N_25618,N_10357,N_13577);
or U25619 (N_25619,N_14638,N_15350);
xnor U25620 (N_25620,N_17862,N_17230);
xnor U25621 (N_25621,N_17265,N_17105);
and U25622 (N_25622,N_14048,N_13808);
or U25623 (N_25623,N_12188,N_11991);
nand U25624 (N_25624,N_18994,N_12215);
or U25625 (N_25625,N_12129,N_19125);
or U25626 (N_25626,N_11500,N_12965);
and U25627 (N_25627,N_18816,N_11378);
nor U25628 (N_25628,N_17130,N_12945);
nand U25629 (N_25629,N_17387,N_11857);
or U25630 (N_25630,N_18869,N_11377);
nor U25631 (N_25631,N_17915,N_19059);
nor U25632 (N_25632,N_11011,N_14760);
xnor U25633 (N_25633,N_13106,N_13292);
nor U25634 (N_25634,N_15169,N_17179);
nor U25635 (N_25635,N_17201,N_16232);
nor U25636 (N_25636,N_15934,N_17292);
or U25637 (N_25637,N_10259,N_19263);
and U25638 (N_25638,N_12861,N_12431);
or U25639 (N_25639,N_19360,N_17935);
nor U25640 (N_25640,N_19870,N_12260);
and U25641 (N_25641,N_13319,N_13415);
nor U25642 (N_25642,N_10424,N_12461);
xor U25643 (N_25643,N_15806,N_16131);
or U25644 (N_25644,N_14489,N_12798);
xnor U25645 (N_25645,N_18346,N_19241);
nor U25646 (N_25646,N_10017,N_17412);
xnor U25647 (N_25647,N_15931,N_12090);
xor U25648 (N_25648,N_15814,N_12218);
xnor U25649 (N_25649,N_11208,N_13586);
nand U25650 (N_25650,N_13088,N_18484);
nor U25651 (N_25651,N_15750,N_19042);
nand U25652 (N_25652,N_17487,N_15094);
nor U25653 (N_25653,N_17983,N_13758);
nand U25654 (N_25654,N_12629,N_18448);
xnor U25655 (N_25655,N_11719,N_13256);
nand U25656 (N_25656,N_12444,N_15351);
nor U25657 (N_25657,N_12932,N_14674);
nor U25658 (N_25658,N_19987,N_16063);
and U25659 (N_25659,N_14840,N_15359);
and U25660 (N_25660,N_19879,N_19522);
xnor U25661 (N_25661,N_15154,N_12335);
nor U25662 (N_25662,N_13166,N_13621);
or U25663 (N_25663,N_10576,N_16220);
nor U25664 (N_25664,N_11156,N_17341);
xor U25665 (N_25665,N_15893,N_15852);
or U25666 (N_25666,N_14433,N_18159);
nor U25667 (N_25667,N_12640,N_11480);
nand U25668 (N_25668,N_10304,N_18841);
nor U25669 (N_25669,N_16031,N_18924);
and U25670 (N_25670,N_15817,N_17977);
or U25671 (N_25671,N_13973,N_10863);
or U25672 (N_25672,N_19765,N_17743);
nand U25673 (N_25673,N_17990,N_19122);
nor U25674 (N_25674,N_11932,N_12822);
xnor U25675 (N_25675,N_14061,N_12724);
nor U25676 (N_25676,N_14901,N_10221);
and U25677 (N_25677,N_17573,N_13232);
nor U25678 (N_25678,N_15066,N_16654);
nor U25679 (N_25679,N_12304,N_13817);
nor U25680 (N_25680,N_18139,N_16141);
and U25681 (N_25681,N_12377,N_14451);
and U25682 (N_25682,N_19156,N_10262);
nor U25683 (N_25683,N_18388,N_10293);
nand U25684 (N_25684,N_17794,N_16787);
nand U25685 (N_25685,N_12389,N_16923);
nor U25686 (N_25686,N_15806,N_11432);
and U25687 (N_25687,N_13602,N_19159);
xnor U25688 (N_25688,N_11457,N_17954);
or U25689 (N_25689,N_18922,N_16178);
nand U25690 (N_25690,N_19941,N_11541);
or U25691 (N_25691,N_12977,N_15759);
or U25692 (N_25692,N_17457,N_11229);
or U25693 (N_25693,N_10763,N_14947);
or U25694 (N_25694,N_10614,N_11626);
xor U25695 (N_25695,N_10496,N_12616);
and U25696 (N_25696,N_19614,N_14722);
nor U25697 (N_25697,N_14684,N_16436);
nor U25698 (N_25698,N_18494,N_11886);
nand U25699 (N_25699,N_16798,N_15199);
and U25700 (N_25700,N_16725,N_18606);
or U25701 (N_25701,N_16679,N_11767);
and U25702 (N_25702,N_11190,N_11890);
or U25703 (N_25703,N_10486,N_10708);
nand U25704 (N_25704,N_17104,N_10285);
nand U25705 (N_25705,N_11923,N_11140);
nor U25706 (N_25706,N_13465,N_17801);
xnor U25707 (N_25707,N_12203,N_13161);
nor U25708 (N_25708,N_10815,N_18459);
nand U25709 (N_25709,N_15209,N_17103);
and U25710 (N_25710,N_14798,N_11642);
nand U25711 (N_25711,N_18002,N_10727);
nand U25712 (N_25712,N_12335,N_17420);
nor U25713 (N_25713,N_10970,N_18340);
and U25714 (N_25714,N_19461,N_15579);
nand U25715 (N_25715,N_12593,N_18879);
nand U25716 (N_25716,N_19007,N_18492);
nor U25717 (N_25717,N_16874,N_18095);
or U25718 (N_25718,N_13325,N_18875);
xnor U25719 (N_25719,N_18729,N_18865);
nand U25720 (N_25720,N_18952,N_16261);
or U25721 (N_25721,N_14247,N_17479);
or U25722 (N_25722,N_10619,N_14639);
or U25723 (N_25723,N_11713,N_17509);
or U25724 (N_25724,N_16983,N_14955);
nand U25725 (N_25725,N_14204,N_16699);
nor U25726 (N_25726,N_11763,N_14042);
nand U25727 (N_25727,N_17259,N_10430);
or U25728 (N_25728,N_17981,N_10209);
and U25729 (N_25729,N_11084,N_18174);
and U25730 (N_25730,N_18808,N_19281);
or U25731 (N_25731,N_16336,N_16183);
xnor U25732 (N_25732,N_13063,N_12644);
nand U25733 (N_25733,N_13857,N_10508);
and U25734 (N_25734,N_18931,N_19322);
or U25735 (N_25735,N_12885,N_16401);
nor U25736 (N_25736,N_18556,N_18276);
nor U25737 (N_25737,N_14632,N_12724);
nor U25738 (N_25738,N_14614,N_14871);
and U25739 (N_25739,N_13624,N_12293);
or U25740 (N_25740,N_18505,N_11245);
nand U25741 (N_25741,N_10612,N_16336);
nand U25742 (N_25742,N_14926,N_18778);
and U25743 (N_25743,N_11788,N_16271);
or U25744 (N_25744,N_16002,N_17956);
or U25745 (N_25745,N_17140,N_10522);
nand U25746 (N_25746,N_15685,N_12224);
xnor U25747 (N_25747,N_11409,N_12010);
nor U25748 (N_25748,N_17395,N_16419);
and U25749 (N_25749,N_19046,N_17771);
xor U25750 (N_25750,N_12597,N_17538);
nor U25751 (N_25751,N_13671,N_12363);
or U25752 (N_25752,N_17568,N_10858);
or U25753 (N_25753,N_16160,N_14057);
xnor U25754 (N_25754,N_12746,N_15015);
nor U25755 (N_25755,N_14857,N_14819);
nand U25756 (N_25756,N_16016,N_10310);
or U25757 (N_25757,N_19605,N_11310);
xnor U25758 (N_25758,N_13135,N_15024);
or U25759 (N_25759,N_13201,N_10189);
nand U25760 (N_25760,N_16236,N_13415);
or U25761 (N_25761,N_12914,N_11137);
nor U25762 (N_25762,N_10645,N_12769);
nor U25763 (N_25763,N_15459,N_13472);
nand U25764 (N_25764,N_19183,N_14407);
or U25765 (N_25765,N_14592,N_10192);
and U25766 (N_25766,N_11151,N_12329);
and U25767 (N_25767,N_18778,N_18810);
or U25768 (N_25768,N_15129,N_18000);
and U25769 (N_25769,N_18549,N_12094);
or U25770 (N_25770,N_15343,N_11170);
nor U25771 (N_25771,N_17911,N_10346);
nor U25772 (N_25772,N_18768,N_12588);
nor U25773 (N_25773,N_17439,N_11476);
nor U25774 (N_25774,N_12675,N_13624);
or U25775 (N_25775,N_19241,N_16800);
nand U25776 (N_25776,N_12237,N_14831);
and U25777 (N_25777,N_12965,N_17043);
nor U25778 (N_25778,N_14785,N_12008);
nor U25779 (N_25779,N_15837,N_18596);
and U25780 (N_25780,N_19859,N_13698);
nand U25781 (N_25781,N_14650,N_13446);
nor U25782 (N_25782,N_11989,N_19325);
and U25783 (N_25783,N_17512,N_11313);
and U25784 (N_25784,N_14072,N_18314);
and U25785 (N_25785,N_16996,N_16283);
xnor U25786 (N_25786,N_13885,N_18483);
or U25787 (N_25787,N_11745,N_17641);
and U25788 (N_25788,N_15316,N_16856);
and U25789 (N_25789,N_14034,N_12174);
and U25790 (N_25790,N_11641,N_15416);
nor U25791 (N_25791,N_10550,N_12924);
nor U25792 (N_25792,N_19568,N_19200);
nor U25793 (N_25793,N_15771,N_19948);
xnor U25794 (N_25794,N_16731,N_16213);
and U25795 (N_25795,N_13899,N_13388);
nor U25796 (N_25796,N_15211,N_10407);
or U25797 (N_25797,N_12257,N_12248);
nand U25798 (N_25798,N_17409,N_10826);
or U25799 (N_25799,N_14164,N_11813);
nand U25800 (N_25800,N_11087,N_11330);
nand U25801 (N_25801,N_18028,N_15535);
or U25802 (N_25802,N_12241,N_16473);
or U25803 (N_25803,N_18524,N_16362);
nor U25804 (N_25804,N_18183,N_18676);
or U25805 (N_25805,N_14310,N_11606);
xor U25806 (N_25806,N_18851,N_11284);
and U25807 (N_25807,N_19600,N_13054);
nor U25808 (N_25808,N_11432,N_15488);
and U25809 (N_25809,N_18931,N_17929);
or U25810 (N_25810,N_14648,N_16850);
xnor U25811 (N_25811,N_16073,N_12973);
nand U25812 (N_25812,N_14575,N_11926);
or U25813 (N_25813,N_12144,N_18102);
nand U25814 (N_25814,N_16504,N_13794);
and U25815 (N_25815,N_12131,N_18034);
or U25816 (N_25816,N_16679,N_18518);
or U25817 (N_25817,N_13513,N_11846);
and U25818 (N_25818,N_10267,N_10447);
and U25819 (N_25819,N_16932,N_15055);
and U25820 (N_25820,N_12305,N_19707);
xnor U25821 (N_25821,N_16674,N_13765);
or U25822 (N_25822,N_14207,N_18463);
or U25823 (N_25823,N_15301,N_19427);
or U25824 (N_25824,N_17450,N_18225);
or U25825 (N_25825,N_15787,N_15029);
nor U25826 (N_25826,N_15888,N_10300);
and U25827 (N_25827,N_15003,N_14823);
nand U25828 (N_25828,N_12860,N_14221);
nor U25829 (N_25829,N_16091,N_17538);
xor U25830 (N_25830,N_11104,N_11171);
nor U25831 (N_25831,N_12458,N_15475);
nand U25832 (N_25832,N_10900,N_18065);
and U25833 (N_25833,N_13121,N_13865);
or U25834 (N_25834,N_13222,N_14137);
xor U25835 (N_25835,N_13492,N_18887);
nand U25836 (N_25836,N_13884,N_15754);
nand U25837 (N_25837,N_15393,N_17759);
or U25838 (N_25838,N_11141,N_15585);
and U25839 (N_25839,N_16209,N_13393);
xor U25840 (N_25840,N_12205,N_16121);
and U25841 (N_25841,N_17080,N_10956);
and U25842 (N_25842,N_11600,N_14212);
nand U25843 (N_25843,N_19924,N_10755);
xor U25844 (N_25844,N_11125,N_19793);
xor U25845 (N_25845,N_19754,N_19951);
nand U25846 (N_25846,N_15783,N_12540);
and U25847 (N_25847,N_14611,N_13692);
nand U25848 (N_25848,N_16210,N_13820);
nor U25849 (N_25849,N_16235,N_19353);
or U25850 (N_25850,N_13797,N_12689);
or U25851 (N_25851,N_18333,N_18676);
and U25852 (N_25852,N_10069,N_15184);
and U25853 (N_25853,N_14616,N_13725);
or U25854 (N_25854,N_19047,N_16513);
nor U25855 (N_25855,N_11679,N_16188);
nand U25856 (N_25856,N_15677,N_12902);
nor U25857 (N_25857,N_18991,N_13342);
or U25858 (N_25858,N_11177,N_15835);
xor U25859 (N_25859,N_16084,N_15973);
nor U25860 (N_25860,N_14669,N_15286);
and U25861 (N_25861,N_19855,N_11720);
nor U25862 (N_25862,N_19040,N_17972);
and U25863 (N_25863,N_18691,N_10692);
and U25864 (N_25864,N_16677,N_14758);
xnor U25865 (N_25865,N_13781,N_14338);
or U25866 (N_25866,N_13495,N_13021);
or U25867 (N_25867,N_14100,N_10925);
nor U25868 (N_25868,N_17020,N_19033);
and U25869 (N_25869,N_18055,N_14256);
nand U25870 (N_25870,N_16154,N_19749);
xor U25871 (N_25871,N_18612,N_11851);
xor U25872 (N_25872,N_18438,N_14117);
or U25873 (N_25873,N_13442,N_12597);
or U25874 (N_25874,N_19806,N_19141);
or U25875 (N_25875,N_14303,N_17737);
and U25876 (N_25876,N_10700,N_17057);
nand U25877 (N_25877,N_12124,N_19436);
nand U25878 (N_25878,N_10413,N_18044);
and U25879 (N_25879,N_18022,N_16270);
nor U25880 (N_25880,N_17773,N_17327);
nor U25881 (N_25881,N_18741,N_11437);
and U25882 (N_25882,N_10561,N_13860);
xnor U25883 (N_25883,N_13521,N_12458);
and U25884 (N_25884,N_15110,N_17676);
nand U25885 (N_25885,N_18709,N_10009);
nor U25886 (N_25886,N_12778,N_17085);
nor U25887 (N_25887,N_19059,N_16347);
and U25888 (N_25888,N_16034,N_14112);
xnor U25889 (N_25889,N_12723,N_13200);
nand U25890 (N_25890,N_15415,N_19899);
nand U25891 (N_25891,N_19289,N_11068);
or U25892 (N_25892,N_12662,N_15537);
and U25893 (N_25893,N_15589,N_14528);
nor U25894 (N_25894,N_19634,N_17128);
or U25895 (N_25895,N_15869,N_19992);
or U25896 (N_25896,N_14000,N_16688);
nand U25897 (N_25897,N_19454,N_14407);
xor U25898 (N_25898,N_12564,N_10092);
nand U25899 (N_25899,N_16848,N_18992);
or U25900 (N_25900,N_13797,N_12842);
or U25901 (N_25901,N_18112,N_12110);
nor U25902 (N_25902,N_14850,N_18161);
or U25903 (N_25903,N_11960,N_14502);
and U25904 (N_25904,N_18842,N_12430);
and U25905 (N_25905,N_11363,N_19247);
nand U25906 (N_25906,N_12895,N_19204);
xor U25907 (N_25907,N_14613,N_19788);
nor U25908 (N_25908,N_16850,N_12882);
or U25909 (N_25909,N_14891,N_15437);
and U25910 (N_25910,N_17214,N_14291);
or U25911 (N_25911,N_17018,N_19438);
nor U25912 (N_25912,N_11951,N_15349);
or U25913 (N_25913,N_15758,N_12577);
or U25914 (N_25914,N_16877,N_19617);
nor U25915 (N_25915,N_10075,N_15671);
nor U25916 (N_25916,N_11295,N_12197);
and U25917 (N_25917,N_13284,N_16381);
nor U25918 (N_25918,N_17498,N_18539);
nand U25919 (N_25919,N_17179,N_11318);
or U25920 (N_25920,N_14389,N_14854);
nor U25921 (N_25921,N_16907,N_16939);
or U25922 (N_25922,N_19976,N_19238);
or U25923 (N_25923,N_14622,N_13623);
xnor U25924 (N_25924,N_18832,N_11424);
nand U25925 (N_25925,N_13518,N_18917);
and U25926 (N_25926,N_18004,N_19544);
or U25927 (N_25927,N_14245,N_16201);
or U25928 (N_25928,N_16130,N_12224);
or U25929 (N_25929,N_17858,N_12332);
or U25930 (N_25930,N_15147,N_18046);
nand U25931 (N_25931,N_12438,N_18288);
nand U25932 (N_25932,N_17906,N_17961);
xor U25933 (N_25933,N_11148,N_17957);
and U25934 (N_25934,N_17007,N_15163);
nand U25935 (N_25935,N_15819,N_18352);
or U25936 (N_25936,N_19783,N_11740);
nand U25937 (N_25937,N_19566,N_14923);
and U25938 (N_25938,N_16405,N_10258);
nand U25939 (N_25939,N_18628,N_18762);
nor U25940 (N_25940,N_16835,N_10908);
or U25941 (N_25941,N_19002,N_16492);
and U25942 (N_25942,N_19865,N_18649);
or U25943 (N_25943,N_18770,N_13467);
or U25944 (N_25944,N_11006,N_19819);
and U25945 (N_25945,N_15268,N_12387);
xor U25946 (N_25946,N_14170,N_18844);
and U25947 (N_25947,N_10465,N_19495);
nor U25948 (N_25948,N_13440,N_11419);
or U25949 (N_25949,N_18565,N_17493);
xnor U25950 (N_25950,N_14038,N_14824);
or U25951 (N_25951,N_13896,N_13334);
nand U25952 (N_25952,N_14491,N_10074);
nand U25953 (N_25953,N_19899,N_19104);
nor U25954 (N_25954,N_19676,N_10453);
and U25955 (N_25955,N_12052,N_19558);
and U25956 (N_25956,N_15349,N_18765);
xnor U25957 (N_25957,N_10354,N_18820);
nand U25958 (N_25958,N_18348,N_17133);
nand U25959 (N_25959,N_19179,N_17917);
or U25960 (N_25960,N_11095,N_16219);
or U25961 (N_25961,N_12136,N_19399);
or U25962 (N_25962,N_17133,N_14183);
or U25963 (N_25963,N_12223,N_14536);
nand U25964 (N_25964,N_13275,N_15337);
xnor U25965 (N_25965,N_17117,N_15034);
and U25966 (N_25966,N_11454,N_15440);
or U25967 (N_25967,N_12430,N_19144);
or U25968 (N_25968,N_16885,N_12506);
xor U25969 (N_25969,N_12584,N_17784);
and U25970 (N_25970,N_15500,N_17732);
or U25971 (N_25971,N_14457,N_12003);
and U25972 (N_25972,N_17727,N_18303);
nor U25973 (N_25973,N_17948,N_19005);
xnor U25974 (N_25974,N_18599,N_13847);
nand U25975 (N_25975,N_10454,N_10941);
and U25976 (N_25976,N_19752,N_11492);
or U25977 (N_25977,N_14830,N_16148);
and U25978 (N_25978,N_14989,N_14655);
nor U25979 (N_25979,N_19042,N_15439);
nand U25980 (N_25980,N_13033,N_16721);
and U25981 (N_25981,N_12994,N_10456);
or U25982 (N_25982,N_11053,N_11778);
xor U25983 (N_25983,N_17459,N_18007);
nor U25984 (N_25984,N_19463,N_10486);
or U25985 (N_25985,N_10625,N_15908);
nor U25986 (N_25986,N_13698,N_17183);
and U25987 (N_25987,N_13321,N_19701);
or U25988 (N_25988,N_18029,N_11503);
nand U25989 (N_25989,N_18129,N_19308);
and U25990 (N_25990,N_16506,N_12925);
and U25991 (N_25991,N_10748,N_18384);
nand U25992 (N_25992,N_11939,N_18008);
nor U25993 (N_25993,N_17432,N_11833);
nand U25994 (N_25994,N_16023,N_18933);
nor U25995 (N_25995,N_12764,N_17518);
or U25996 (N_25996,N_11678,N_10044);
or U25997 (N_25997,N_13891,N_14501);
or U25998 (N_25998,N_11070,N_18488);
nor U25999 (N_25999,N_12928,N_13603);
or U26000 (N_26000,N_13674,N_10362);
nand U26001 (N_26001,N_17863,N_15198);
or U26002 (N_26002,N_13733,N_18426);
nand U26003 (N_26003,N_14214,N_15404);
and U26004 (N_26004,N_12427,N_15751);
and U26005 (N_26005,N_10029,N_18136);
nand U26006 (N_26006,N_19492,N_15438);
nand U26007 (N_26007,N_15866,N_12606);
nor U26008 (N_26008,N_18808,N_19229);
nor U26009 (N_26009,N_17931,N_14236);
and U26010 (N_26010,N_11723,N_16550);
or U26011 (N_26011,N_15053,N_19462);
and U26012 (N_26012,N_13983,N_11483);
and U26013 (N_26013,N_11029,N_12689);
and U26014 (N_26014,N_15284,N_13585);
and U26015 (N_26015,N_12609,N_15016);
nor U26016 (N_26016,N_15598,N_18617);
or U26017 (N_26017,N_11427,N_18443);
nor U26018 (N_26018,N_16829,N_14597);
and U26019 (N_26019,N_13558,N_13212);
nor U26020 (N_26020,N_19836,N_19298);
nand U26021 (N_26021,N_16960,N_15414);
xnor U26022 (N_26022,N_17220,N_17677);
nor U26023 (N_26023,N_15011,N_17803);
nor U26024 (N_26024,N_15377,N_12484);
or U26025 (N_26025,N_16462,N_17419);
and U26026 (N_26026,N_11935,N_16250);
or U26027 (N_26027,N_15118,N_17543);
xor U26028 (N_26028,N_19074,N_10937);
or U26029 (N_26029,N_11244,N_13464);
nor U26030 (N_26030,N_14083,N_17458);
nor U26031 (N_26031,N_18098,N_17788);
nand U26032 (N_26032,N_15591,N_11080);
or U26033 (N_26033,N_18820,N_17391);
nand U26034 (N_26034,N_18606,N_14944);
nand U26035 (N_26035,N_18361,N_11958);
xnor U26036 (N_26036,N_11092,N_13486);
and U26037 (N_26037,N_10560,N_14553);
nor U26038 (N_26038,N_19610,N_18973);
nor U26039 (N_26039,N_13901,N_15547);
or U26040 (N_26040,N_12528,N_17127);
or U26041 (N_26041,N_18871,N_14197);
nor U26042 (N_26042,N_16084,N_17298);
and U26043 (N_26043,N_12225,N_10239);
nand U26044 (N_26044,N_14330,N_15239);
or U26045 (N_26045,N_13163,N_17824);
nor U26046 (N_26046,N_16572,N_11573);
or U26047 (N_26047,N_18624,N_11987);
xor U26048 (N_26048,N_12668,N_17839);
xnor U26049 (N_26049,N_16040,N_14248);
or U26050 (N_26050,N_18178,N_18365);
xor U26051 (N_26051,N_19508,N_10003);
nand U26052 (N_26052,N_13163,N_10149);
nand U26053 (N_26053,N_17027,N_16690);
xnor U26054 (N_26054,N_16439,N_14478);
nor U26055 (N_26055,N_16964,N_10136);
or U26056 (N_26056,N_16175,N_17285);
xor U26057 (N_26057,N_11167,N_13398);
nand U26058 (N_26058,N_16347,N_14508);
nand U26059 (N_26059,N_16164,N_18602);
or U26060 (N_26060,N_17147,N_11882);
and U26061 (N_26061,N_14760,N_10762);
or U26062 (N_26062,N_19689,N_13391);
nor U26063 (N_26063,N_13803,N_19032);
or U26064 (N_26064,N_10273,N_12179);
xor U26065 (N_26065,N_10600,N_11051);
xor U26066 (N_26066,N_19978,N_12826);
nor U26067 (N_26067,N_16932,N_12040);
or U26068 (N_26068,N_18144,N_10857);
xor U26069 (N_26069,N_17497,N_11373);
and U26070 (N_26070,N_14344,N_12200);
nand U26071 (N_26071,N_17837,N_17664);
nor U26072 (N_26072,N_10015,N_11294);
or U26073 (N_26073,N_18433,N_15135);
nor U26074 (N_26074,N_10325,N_11530);
and U26075 (N_26075,N_13655,N_16395);
nand U26076 (N_26076,N_17895,N_17888);
nand U26077 (N_26077,N_15024,N_18711);
and U26078 (N_26078,N_14886,N_11571);
and U26079 (N_26079,N_10387,N_10877);
and U26080 (N_26080,N_14083,N_16160);
or U26081 (N_26081,N_15617,N_12018);
nand U26082 (N_26082,N_13254,N_12609);
or U26083 (N_26083,N_19992,N_11620);
xnor U26084 (N_26084,N_19535,N_18469);
xor U26085 (N_26085,N_17877,N_12732);
nor U26086 (N_26086,N_14379,N_12524);
or U26087 (N_26087,N_10421,N_11992);
and U26088 (N_26088,N_12515,N_15008);
and U26089 (N_26089,N_18255,N_12715);
xor U26090 (N_26090,N_18471,N_18875);
and U26091 (N_26091,N_18422,N_16696);
and U26092 (N_26092,N_15448,N_11108);
nand U26093 (N_26093,N_11339,N_13760);
and U26094 (N_26094,N_15378,N_17543);
or U26095 (N_26095,N_14178,N_10460);
nand U26096 (N_26096,N_19908,N_14938);
nand U26097 (N_26097,N_15257,N_19264);
and U26098 (N_26098,N_13598,N_11345);
or U26099 (N_26099,N_18650,N_19278);
or U26100 (N_26100,N_11012,N_14761);
nand U26101 (N_26101,N_19027,N_11324);
or U26102 (N_26102,N_11135,N_11782);
or U26103 (N_26103,N_13571,N_18558);
nor U26104 (N_26104,N_15229,N_16441);
nand U26105 (N_26105,N_11681,N_10286);
nand U26106 (N_26106,N_15124,N_11431);
or U26107 (N_26107,N_11274,N_16815);
nor U26108 (N_26108,N_12557,N_17162);
or U26109 (N_26109,N_18920,N_13992);
nor U26110 (N_26110,N_14343,N_15791);
or U26111 (N_26111,N_16838,N_16986);
or U26112 (N_26112,N_16332,N_14440);
or U26113 (N_26113,N_15711,N_11279);
xnor U26114 (N_26114,N_13355,N_18527);
nand U26115 (N_26115,N_15517,N_13981);
xnor U26116 (N_26116,N_16592,N_14237);
nand U26117 (N_26117,N_18014,N_11300);
or U26118 (N_26118,N_13495,N_18675);
and U26119 (N_26119,N_16219,N_14839);
nand U26120 (N_26120,N_11309,N_15642);
or U26121 (N_26121,N_11192,N_15986);
nor U26122 (N_26122,N_14070,N_10125);
nor U26123 (N_26123,N_16716,N_14416);
nor U26124 (N_26124,N_13248,N_17268);
and U26125 (N_26125,N_10091,N_11896);
nor U26126 (N_26126,N_18234,N_10485);
nand U26127 (N_26127,N_18421,N_13222);
nor U26128 (N_26128,N_11719,N_15432);
nand U26129 (N_26129,N_13929,N_17579);
nor U26130 (N_26130,N_11082,N_17727);
nor U26131 (N_26131,N_19874,N_12132);
and U26132 (N_26132,N_18321,N_18157);
xnor U26133 (N_26133,N_19755,N_11703);
and U26134 (N_26134,N_19553,N_14084);
or U26135 (N_26135,N_10678,N_14604);
xor U26136 (N_26136,N_13901,N_10350);
or U26137 (N_26137,N_12200,N_11021);
nand U26138 (N_26138,N_17253,N_16322);
xnor U26139 (N_26139,N_13437,N_19285);
nand U26140 (N_26140,N_14853,N_16910);
nor U26141 (N_26141,N_16555,N_17242);
nor U26142 (N_26142,N_16213,N_13222);
nand U26143 (N_26143,N_18893,N_14698);
nor U26144 (N_26144,N_18817,N_14194);
nor U26145 (N_26145,N_15515,N_15004);
nand U26146 (N_26146,N_17584,N_14812);
and U26147 (N_26147,N_14972,N_11488);
or U26148 (N_26148,N_18413,N_16111);
nor U26149 (N_26149,N_19354,N_19734);
nor U26150 (N_26150,N_11586,N_13064);
xor U26151 (N_26151,N_14104,N_14637);
xnor U26152 (N_26152,N_15943,N_12010);
nor U26153 (N_26153,N_17911,N_15708);
nor U26154 (N_26154,N_19483,N_17017);
and U26155 (N_26155,N_15708,N_18092);
nor U26156 (N_26156,N_18319,N_19312);
nand U26157 (N_26157,N_19947,N_10466);
nor U26158 (N_26158,N_12515,N_18380);
nor U26159 (N_26159,N_14547,N_11113);
xnor U26160 (N_26160,N_11058,N_18128);
xor U26161 (N_26161,N_12334,N_18321);
nand U26162 (N_26162,N_12933,N_16090);
and U26163 (N_26163,N_12456,N_14702);
nand U26164 (N_26164,N_11069,N_15275);
nor U26165 (N_26165,N_14598,N_18218);
and U26166 (N_26166,N_13109,N_13166);
xor U26167 (N_26167,N_16631,N_13077);
nor U26168 (N_26168,N_15216,N_13934);
or U26169 (N_26169,N_13438,N_16280);
and U26170 (N_26170,N_15434,N_17654);
xor U26171 (N_26171,N_10053,N_18941);
nor U26172 (N_26172,N_12410,N_12667);
and U26173 (N_26173,N_17203,N_17258);
nor U26174 (N_26174,N_18671,N_11551);
nor U26175 (N_26175,N_10326,N_16795);
or U26176 (N_26176,N_12682,N_12854);
or U26177 (N_26177,N_19435,N_16222);
nand U26178 (N_26178,N_10050,N_16264);
or U26179 (N_26179,N_18885,N_17910);
nor U26180 (N_26180,N_14608,N_18609);
and U26181 (N_26181,N_12924,N_19280);
and U26182 (N_26182,N_19183,N_13075);
nor U26183 (N_26183,N_17448,N_14749);
nand U26184 (N_26184,N_14268,N_19781);
and U26185 (N_26185,N_14613,N_14593);
and U26186 (N_26186,N_16526,N_15818);
and U26187 (N_26187,N_13672,N_11949);
or U26188 (N_26188,N_13258,N_10576);
or U26189 (N_26189,N_15748,N_13022);
or U26190 (N_26190,N_16348,N_10988);
or U26191 (N_26191,N_13749,N_13897);
and U26192 (N_26192,N_11303,N_13181);
nand U26193 (N_26193,N_14670,N_16164);
nor U26194 (N_26194,N_15173,N_16813);
nor U26195 (N_26195,N_17217,N_15950);
nor U26196 (N_26196,N_19895,N_12426);
and U26197 (N_26197,N_18223,N_12970);
and U26198 (N_26198,N_10291,N_15630);
nand U26199 (N_26199,N_11465,N_16608);
or U26200 (N_26200,N_16401,N_17262);
and U26201 (N_26201,N_14508,N_17183);
and U26202 (N_26202,N_11219,N_10614);
and U26203 (N_26203,N_16209,N_16301);
or U26204 (N_26204,N_11084,N_17218);
nor U26205 (N_26205,N_13873,N_19260);
and U26206 (N_26206,N_17970,N_14314);
nor U26207 (N_26207,N_17969,N_14848);
and U26208 (N_26208,N_11868,N_15760);
and U26209 (N_26209,N_18390,N_15711);
nand U26210 (N_26210,N_13788,N_12780);
nor U26211 (N_26211,N_19915,N_14481);
xnor U26212 (N_26212,N_18251,N_19901);
and U26213 (N_26213,N_12927,N_14315);
and U26214 (N_26214,N_16596,N_17105);
or U26215 (N_26215,N_16743,N_12589);
or U26216 (N_26216,N_15279,N_11988);
and U26217 (N_26217,N_12619,N_19203);
and U26218 (N_26218,N_14858,N_13281);
or U26219 (N_26219,N_10866,N_18661);
xor U26220 (N_26220,N_15263,N_12223);
and U26221 (N_26221,N_14926,N_15613);
nor U26222 (N_26222,N_19684,N_19379);
nand U26223 (N_26223,N_12206,N_19447);
and U26224 (N_26224,N_13770,N_14280);
or U26225 (N_26225,N_16985,N_10370);
xor U26226 (N_26226,N_16099,N_16598);
or U26227 (N_26227,N_18664,N_13042);
or U26228 (N_26228,N_16599,N_15275);
nor U26229 (N_26229,N_14863,N_10102);
nand U26230 (N_26230,N_12312,N_11755);
nand U26231 (N_26231,N_13492,N_11877);
or U26232 (N_26232,N_12320,N_17055);
xor U26233 (N_26233,N_13432,N_14466);
nand U26234 (N_26234,N_13398,N_15046);
nor U26235 (N_26235,N_16882,N_15324);
nor U26236 (N_26236,N_18519,N_14852);
xor U26237 (N_26237,N_19587,N_14852);
nor U26238 (N_26238,N_17791,N_17357);
xnor U26239 (N_26239,N_15744,N_18509);
nor U26240 (N_26240,N_10210,N_12389);
nor U26241 (N_26241,N_13474,N_17626);
and U26242 (N_26242,N_14115,N_17868);
or U26243 (N_26243,N_12588,N_17351);
and U26244 (N_26244,N_11907,N_12044);
nor U26245 (N_26245,N_14844,N_14403);
nand U26246 (N_26246,N_13590,N_16166);
nor U26247 (N_26247,N_10423,N_12609);
nand U26248 (N_26248,N_16760,N_11299);
nor U26249 (N_26249,N_10801,N_18344);
nor U26250 (N_26250,N_11834,N_14498);
nor U26251 (N_26251,N_10279,N_16569);
xor U26252 (N_26252,N_16184,N_15854);
and U26253 (N_26253,N_15184,N_13970);
nor U26254 (N_26254,N_13879,N_11741);
nand U26255 (N_26255,N_14932,N_11957);
and U26256 (N_26256,N_14740,N_11771);
and U26257 (N_26257,N_11960,N_12356);
or U26258 (N_26258,N_19987,N_12579);
or U26259 (N_26259,N_18356,N_16786);
and U26260 (N_26260,N_11617,N_19599);
nor U26261 (N_26261,N_17099,N_18827);
nand U26262 (N_26262,N_13308,N_15219);
nand U26263 (N_26263,N_14765,N_10528);
xnor U26264 (N_26264,N_17846,N_11484);
nand U26265 (N_26265,N_12003,N_11334);
nor U26266 (N_26266,N_15362,N_12435);
and U26267 (N_26267,N_11498,N_14626);
nor U26268 (N_26268,N_12058,N_11028);
and U26269 (N_26269,N_18337,N_19771);
nand U26270 (N_26270,N_11329,N_14778);
nor U26271 (N_26271,N_15742,N_14828);
nand U26272 (N_26272,N_11142,N_19485);
xnor U26273 (N_26273,N_19005,N_18614);
nor U26274 (N_26274,N_15478,N_17784);
xnor U26275 (N_26275,N_10615,N_10302);
and U26276 (N_26276,N_15276,N_11462);
and U26277 (N_26277,N_19490,N_19297);
and U26278 (N_26278,N_12320,N_17899);
nor U26279 (N_26279,N_18925,N_11493);
and U26280 (N_26280,N_19472,N_11439);
and U26281 (N_26281,N_13964,N_19424);
or U26282 (N_26282,N_10793,N_16426);
and U26283 (N_26283,N_10317,N_11254);
or U26284 (N_26284,N_10745,N_16757);
and U26285 (N_26285,N_11488,N_18710);
nand U26286 (N_26286,N_15242,N_15401);
nor U26287 (N_26287,N_18964,N_18991);
or U26288 (N_26288,N_10875,N_12876);
and U26289 (N_26289,N_12048,N_17600);
or U26290 (N_26290,N_13614,N_12897);
nand U26291 (N_26291,N_14672,N_19620);
nor U26292 (N_26292,N_17746,N_13402);
nor U26293 (N_26293,N_15460,N_14592);
nor U26294 (N_26294,N_10659,N_17466);
and U26295 (N_26295,N_16711,N_11686);
and U26296 (N_26296,N_12376,N_14078);
xnor U26297 (N_26297,N_18926,N_17631);
and U26298 (N_26298,N_18465,N_10343);
nand U26299 (N_26299,N_18161,N_16142);
or U26300 (N_26300,N_14295,N_11405);
nand U26301 (N_26301,N_17350,N_18487);
or U26302 (N_26302,N_11686,N_14804);
nand U26303 (N_26303,N_18832,N_15543);
nor U26304 (N_26304,N_11407,N_16690);
or U26305 (N_26305,N_19480,N_10893);
or U26306 (N_26306,N_13752,N_14211);
nand U26307 (N_26307,N_14472,N_11228);
or U26308 (N_26308,N_13652,N_12938);
xnor U26309 (N_26309,N_18767,N_11190);
nand U26310 (N_26310,N_16387,N_17148);
nand U26311 (N_26311,N_10818,N_13133);
and U26312 (N_26312,N_14154,N_14183);
nand U26313 (N_26313,N_18841,N_14044);
nand U26314 (N_26314,N_19724,N_19995);
and U26315 (N_26315,N_16872,N_19875);
or U26316 (N_26316,N_10516,N_13214);
nor U26317 (N_26317,N_16431,N_15398);
and U26318 (N_26318,N_17199,N_10439);
and U26319 (N_26319,N_13596,N_12593);
nor U26320 (N_26320,N_15973,N_16268);
or U26321 (N_26321,N_13202,N_14007);
or U26322 (N_26322,N_16460,N_16196);
or U26323 (N_26323,N_19521,N_13441);
nand U26324 (N_26324,N_19820,N_17169);
nand U26325 (N_26325,N_17780,N_19130);
xnor U26326 (N_26326,N_14695,N_19053);
nand U26327 (N_26327,N_13445,N_16464);
and U26328 (N_26328,N_14803,N_12804);
or U26329 (N_26329,N_14110,N_12242);
and U26330 (N_26330,N_19220,N_11729);
nand U26331 (N_26331,N_12927,N_17254);
or U26332 (N_26332,N_16232,N_12673);
nand U26333 (N_26333,N_15956,N_11689);
nor U26334 (N_26334,N_11916,N_12274);
or U26335 (N_26335,N_17622,N_15850);
or U26336 (N_26336,N_17415,N_19883);
nor U26337 (N_26337,N_11260,N_19677);
nor U26338 (N_26338,N_18857,N_11531);
and U26339 (N_26339,N_13985,N_16161);
and U26340 (N_26340,N_12247,N_19854);
and U26341 (N_26341,N_15470,N_11563);
nand U26342 (N_26342,N_18722,N_17807);
or U26343 (N_26343,N_17353,N_17328);
nor U26344 (N_26344,N_19853,N_10207);
and U26345 (N_26345,N_18764,N_12797);
or U26346 (N_26346,N_14759,N_11249);
or U26347 (N_26347,N_18365,N_15339);
and U26348 (N_26348,N_16194,N_16163);
and U26349 (N_26349,N_13247,N_10441);
nor U26350 (N_26350,N_12098,N_11772);
or U26351 (N_26351,N_18409,N_19031);
nor U26352 (N_26352,N_11237,N_10779);
nand U26353 (N_26353,N_19112,N_11668);
or U26354 (N_26354,N_11736,N_13614);
and U26355 (N_26355,N_17961,N_13251);
xor U26356 (N_26356,N_16920,N_17287);
and U26357 (N_26357,N_16570,N_13573);
and U26358 (N_26358,N_12701,N_12118);
and U26359 (N_26359,N_14658,N_15692);
nand U26360 (N_26360,N_15860,N_14600);
or U26361 (N_26361,N_15314,N_17283);
xor U26362 (N_26362,N_16864,N_16807);
nand U26363 (N_26363,N_17467,N_15510);
nand U26364 (N_26364,N_10613,N_18102);
and U26365 (N_26365,N_13405,N_17574);
or U26366 (N_26366,N_11288,N_12799);
nor U26367 (N_26367,N_18921,N_10302);
or U26368 (N_26368,N_15455,N_18818);
or U26369 (N_26369,N_13439,N_18438);
xor U26370 (N_26370,N_17407,N_12002);
or U26371 (N_26371,N_10776,N_16436);
xor U26372 (N_26372,N_11527,N_12719);
nor U26373 (N_26373,N_16776,N_11146);
nand U26374 (N_26374,N_13948,N_15131);
nor U26375 (N_26375,N_18350,N_16247);
and U26376 (N_26376,N_18903,N_12888);
xnor U26377 (N_26377,N_10978,N_14834);
xnor U26378 (N_26378,N_16675,N_13609);
and U26379 (N_26379,N_17265,N_17911);
and U26380 (N_26380,N_16566,N_15336);
xnor U26381 (N_26381,N_18881,N_15556);
or U26382 (N_26382,N_17644,N_13761);
nor U26383 (N_26383,N_17650,N_14589);
or U26384 (N_26384,N_11884,N_18305);
nand U26385 (N_26385,N_11120,N_10608);
and U26386 (N_26386,N_10516,N_13940);
nor U26387 (N_26387,N_18989,N_11571);
nor U26388 (N_26388,N_16910,N_14775);
and U26389 (N_26389,N_13514,N_13322);
nand U26390 (N_26390,N_10622,N_17819);
and U26391 (N_26391,N_10277,N_11558);
xnor U26392 (N_26392,N_14238,N_16177);
nor U26393 (N_26393,N_15269,N_13581);
nor U26394 (N_26394,N_18201,N_12289);
nor U26395 (N_26395,N_18143,N_19106);
and U26396 (N_26396,N_17435,N_17980);
nor U26397 (N_26397,N_17443,N_10030);
nand U26398 (N_26398,N_13121,N_19062);
nand U26399 (N_26399,N_18024,N_19559);
and U26400 (N_26400,N_18117,N_11489);
nor U26401 (N_26401,N_19814,N_16291);
xor U26402 (N_26402,N_14683,N_13100);
or U26403 (N_26403,N_11762,N_10948);
and U26404 (N_26404,N_14875,N_13460);
nand U26405 (N_26405,N_14860,N_13809);
nand U26406 (N_26406,N_13416,N_16752);
nor U26407 (N_26407,N_14718,N_11578);
and U26408 (N_26408,N_16299,N_16023);
and U26409 (N_26409,N_13547,N_15680);
or U26410 (N_26410,N_18799,N_14406);
or U26411 (N_26411,N_15414,N_19867);
nor U26412 (N_26412,N_11398,N_18593);
nand U26413 (N_26413,N_17065,N_11348);
or U26414 (N_26414,N_13020,N_10783);
and U26415 (N_26415,N_18798,N_16198);
and U26416 (N_26416,N_12587,N_15404);
and U26417 (N_26417,N_12467,N_14696);
or U26418 (N_26418,N_18756,N_16427);
xnor U26419 (N_26419,N_15768,N_16915);
or U26420 (N_26420,N_17265,N_13306);
or U26421 (N_26421,N_16763,N_11186);
nand U26422 (N_26422,N_16869,N_18766);
xnor U26423 (N_26423,N_13265,N_13366);
nand U26424 (N_26424,N_10591,N_12649);
or U26425 (N_26425,N_17702,N_18675);
nand U26426 (N_26426,N_19502,N_15314);
and U26427 (N_26427,N_17626,N_12898);
nor U26428 (N_26428,N_19444,N_17380);
nor U26429 (N_26429,N_10249,N_10588);
or U26430 (N_26430,N_18804,N_11224);
nand U26431 (N_26431,N_12926,N_14305);
and U26432 (N_26432,N_19477,N_19402);
and U26433 (N_26433,N_19149,N_18243);
nor U26434 (N_26434,N_17995,N_13813);
nand U26435 (N_26435,N_13083,N_12494);
nor U26436 (N_26436,N_15087,N_11354);
nand U26437 (N_26437,N_12108,N_11957);
or U26438 (N_26438,N_13349,N_14042);
nor U26439 (N_26439,N_15194,N_16237);
nand U26440 (N_26440,N_12377,N_17467);
and U26441 (N_26441,N_13954,N_11849);
or U26442 (N_26442,N_19023,N_15657);
xor U26443 (N_26443,N_16596,N_14370);
xor U26444 (N_26444,N_19108,N_19553);
or U26445 (N_26445,N_16753,N_15693);
or U26446 (N_26446,N_18118,N_17779);
or U26447 (N_26447,N_15866,N_16605);
or U26448 (N_26448,N_10394,N_17753);
or U26449 (N_26449,N_18413,N_18913);
nor U26450 (N_26450,N_12028,N_15075);
or U26451 (N_26451,N_14203,N_15089);
or U26452 (N_26452,N_17346,N_13038);
nand U26453 (N_26453,N_14732,N_19268);
nor U26454 (N_26454,N_17528,N_11658);
xnor U26455 (N_26455,N_15054,N_13824);
or U26456 (N_26456,N_19222,N_12205);
nor U26457 (N_26457,N_18312,N_19959);
nand U26458 (N_26458,N_19069,N_12994);
and U26459 (N_26459,N_11234,N_10293);
or U26460 (N_26460,N_15495,N_15832);
nor U26461 (N_26461,N_18102,N_11608);
or U26462 (N_26462,N_10849,N_13132);
xnor U26463 (N_26463,N_14674,N_15937);
nor U26464 (N_26464,N_11424,N_13184);
and U26465 (N_26465,N_10029,N_11242);
xnor U26466 (N_26466,N_14310,N_16006);
nor U26467 (N_26467,N_19262,N_13161);
or U26468 (N_26468,N_11480,N_15346);
or U26469 (N_26469,N_14190,N_15275);
xnor U26470 (N_26470,N_15849,N_13171);
nand U26471 (N_26471,N_12585,N_11553);
nor U26472 (N_26472,N_17871,N_16787);
nor U26473 (N_26473,N_11555,N_14473);
nand U26474 (N_26474,N_11054,N_18465);
or U26475 (N_26475,N_14958,N_17884);
and U26476 (N_26476,N_10114,N_15288);
and U26477 (N_26477,N_19817,N_15888);
nand U26478 (N_26478,N_12291,N_10761);
nand U26479 (N_26479,N_17676,N_10818);
and U26480 (N_26480,N_14361,N_14582);
nand U26481 (N_26481,N_11744,N_14603);
nor U26482 (N_26482,N_18545,N_10087);
nand U26483 (N_26483,N_16684,N_19895);
and U26484 (N_26484,N_16159,N_13973);
nand U26485 (N_26485,N_14107,N_17600);
nor U26486 (N_26486,N_18432,N_19532);
or U26487 (N_26487,N_14519,N_15217);
and U26488 (N_26488,N_11360,N_12614);
xnor U26489 (N_26489,N_19698,N_10113);
or U26490 (N_26490,N_13614,N_10495);
or U26491 (N_26491,N_15121,N_17109);
nor U26492 (N_26492,N_13503,N_10805);
xnor U26493 (N_26493,N_15913,N_14418);
or U26494 (N_26494,N_14750,N_11703);
or U26495 (N_26495,N_14067,N_13118);
or U26496 (N_26496,N_16128,N_13035);
nor U26497 (N_26497,N_17868,N_18001);
nor U26498 (N_26498,N_12086,N_10230);
nand U26499 (N_26499,N_17438,N_16348);
and U26500 (N_26500,N_11049,N_13049);
and U26501 (N_26501,N_14533,N_12024);
nand U26502 (N_26502,N_13318,N_15335);
nand U26503 (N_26503,N_12247,N_12840);
nand U26504 (N_26504,N_12083,N_14076);
nand U26505 (N_26505,N_19812,N_19702);
xnor U26506 (N_26506,N_13286,N_14718);
nand U26507 (N_26507,N_11871,N_18277);
and U26508 (N_26508,N_12172,N_10712);
and U26509 (N_26509,N_15040,N_11005);
nand U26510 (N_26510,N_13677,N_11131);
or U26511 (N_26511,N_14717,N_11529);
nand U26512 (N_26512,N_13171,N_18380);
and U26513 (N_26513,N_13140,N_17685);
nand U26514 (N_26514,N_15109,N_10115);
nand U26515 (N_26515,N_11303,N_13592);
nand U26516 (N_26516,N_12221,N_12019);
or U26517 (N_26517,N_14548,N_16560);
or U26518 (N_26518,N_14476,N_13595);
or U26519 (N_26519,N_13334,N_10980);
nor U26520 (N_26520,N_13399,N_12649);
or U26521 (N_26521,N_10052,N_15119);
xor U26522 (N_26522,N_18528,N_17857);
nand U26523 (N_26523,N_15808,N_19526);
xor U26524 (N_26524,N_10322,N_16019);
or U26525 (N_26525,N_13556,N_19318);
and U26526 (N_26526,N_13781,N_11101);
nor U26527 (N_26527,N_17199,N_11377);
nor U26528 (N_26528,N_17656,N_17024);
xor U26529 (N_26529,N_13475,N_17254);
or U26530 (N_26530,N_16257,N_15654);
nand U26531 (N_26531,N_13508,N_11354);
and U26532 (N_26532,N_16375,N_19341);
and U26533 (N_26533,N_14765,N_19926);
and U26534 (N_26534,N_14961,N_12480);
or U26535 (N_26535,N_15498,N_16035);
and U26536 (N_26536,N_15431,N_12353);
nor U26537 (N_26537,N_19327,N_14161);
nor U26538 (N_26538,N_10118,N_10578);
nand U26539 (N_26539,N_11731,N_13894);
and U26540 (N_26540,N_17257,N_16121);
and U26541 (N_26541,N_17140,N_12423);
or U26542 (N_26542,N_12016,N_18567);
and U26543 (N_26543,N_12394,N_13207);
xnor U26544 (N_26544,N_14791,N_19912);
nor U26545 (N_26545,N_11744,N_10186);
and U26546 (N_26546,N_18588,N_12802);
xnor U26547 (N_26547,N_13705,N_15988);
nand U26548 (N_26548,N_16484,N_16448);
nor U26549 (N_26549,N_18806,N_15662);
nor U26550 (N_26550,N_12281,N_15745);
or U26551 (N_26551,N_16469,N_14236);
xnor U26552 (N_26552,N_19882,N_13904);
and U26553 (N_26553,N_11355,N_16530);
or U26554 (N_26554,N_16865,N_18974);
nor U26555 (N_26555,N_18332,N_15785);
nor U26556 (N_26556,N_19899,N_18120);
nand U26557 (N_26557,N_17367,N_11263);
nor U26558 (N_26558,N_17320,N_17629);
nor U26559 (N_26559,N_14410,N_13847);
nor U26560 (N_26560,N_10051,N_19262);
xnor U26561 (N_26561,N_12270,N_17202);
or U26562 (N_26562,N_11640,N_18337);
and U26563 (N_26563,N_15482,N_13094);
xnor U26564 (N_26564,N_19261,N_19430);
or U26565 (N_26565,N_14322,N_18959);
nor U26566 (N_26566,N_15423,N_16775);
nor U26567 (N_26567,N_10476,N_15517);
nand U26568 (N_26568,N_14602,N_17058);
and U26569 (N_26569,N_17026,N_11459);
nor U26570 (N_26570,N_12783,N_14595);
nand U26571 (N_26571,N_16557,N_10787);
nand U26572 (N_26572,N_18544,N_13391);
or U26573 (N_26573,N_17699,N_15025);
nand U26574 (N_26574,N_17079,N_10660);
and U26575 (N_26575,N_18983,N_16816);
and U26576 (N_26576,N_11373,N_12995);
or U26577 (N_26577,N_11411,N_15737);
nor U26578 (N_26578,N_15983,N_12362);
nor U26579 (N_26579,N_12872,N_14688);
nor U26580 (N_26580,N_19201,N_18105);
or U26581 (N_26581,N_15744,N_13235);
or U26582 (N_26582,N_15228,N_10677);
nand U26583 (N_26583,N_11661,N_15349);
or U26584 (N_26584,N_10124,N_10233);
and U26585 (N_26585,N_11386,N_10130);
nor U26586 (N_26586,N_14233,N_16157);
nand U26587 (N_26587,N_14221,N_19970);
nand U26588 (N_26588,N_12526,N_10039);
nor U26589 (N_26589,N_14073,N_17356);
and U26590 (N_26590,N_14522,N_16498);
nand U26591 (N_26591,N_13767,N_19324);
xnor U26592 (N_26592,N_13159,N_19461);
and U26593 (N_26593,N_12663,N_11893);
or U26594 (N_26594,N_19397,N_15195);
xnor U26595 (N_26595,N_18405,N_18693);
or U26596 (N_26596,N_16900,N_15741);
nand U26597 (N_26597,N_16238,N_19488);
nor U26598 (N_26598,N_14839,N_10766);
nand U26599 (N_26599,N_16600,N_11248);
xor U26600 (N_26600,N_15388,N_13026);
nor U26601 (N_26601,N_18952,N_16685);
and U26602 (N_26602,N_16557,N_19380);
and U26603 (N_26603,N_15844,N_10547);
nand U26604 (N_26604,N_15839,N_19805);
xnor U26605 (N_26605,N_12232,N_16550);
and U26606 (N_26606,N_11814,N_19986);
or U26607 (N_26607,N_19959,N_12881);
nand U26608 (N_26608,N_15962,N_14301);
or U26609 (N_26609,N_11053,N_15266);
or U26610 (N_26610,N_15093,N_19026);
or U26611 (N_26611,N_15290,N_19205);
or U26612 (N_26612,N_10828,N_15811);
nor U26613 (N_26613,N_12784,N_15533);
nand U26614 (N_26614,N_10131,N_15769);
nand U26615 (N_26615,N_19860,N_16518);
nand U26616 (N_26616,N_16985,N_18263);
and U26617 (N_26617,N_19187,N_14678);
or U26618 (N_26618,N_10277,N_14042);
or U26619 (N_26619,N_17719,N_12632);
nor U26620 (N_26620,N_15219,N_16000);
and U26621 (N_26621,N_17386,N_15565);
and U26622 (N_26622,N_13084,N_12129);
or U26623 (N_26623,N_16030,N_15570);
and U26624 (N_26624,N_18982,N_13079);
and U26625 (N_26625,N_10628,N_15053);
nor U26626 (N_26626,N_15183,N_10107);
nand U26627 (N_26627,N_17460,N_18160);
or U26628 (N_26628,N_14884,N_13109);
or U26629 (N_26629,N_10254,N_18828);
xnor U26630 (N_26630,N_16015,N_10668);
xnor U26631 (N_26631,N_14883,N_14752);
or U26632 (N_26632,N_15589,N_10312);
nand U26633 (N_26633,N_17912,N_17461);
and U26634 (N_26634,N_17969,N_15329);
nor U26635 (N_26635,N_19496,N_15620);
and U26636 (N_26636,N_16574,N_12980);
nand U26637 (N_26637,N_11247,N_14560);
nor U26638 (N_26638,N_18722,N_11962);
and U26639 (N_26639,N_14106,N_10464);
and U26640 (N_26640,N_15667,N_17365);
nand U26641 (N_26641,N_10591,N_16913);
or U26642 (N_26642,N_11131,N_15913);
or U26643 (N_26643,N_13487,N_12406);
or U26644 (N_26644,N_17082,N_18408);
or U26645 (N_26645,N_11865,N_16077);
and U26646 (N_26646,N_13675,N_10467);
nand U26647 (N_26647,N_11629,N_19449);
nor U26648 (N_26648,N_15785,N_13424);
or U26649 (N_26649,N_15346,N_18460);
or U26650 (N_26650,N_14089,N_17294);
and U26651 (N_26651,N_15199,N_11991);
and U26652 (N_26652,N_12817,N_12336);
or U26653 (N_26653,N_16799,N_10774);
nor U26654 (N_26654,N_18770,N_12058);
nor U26655 (N_26655,N_19172,N_18748);
nand U26656 (N_26656,N_16639,N_14139);
and U26657 (N_26657,N_12670,N_19895);
and U26658 (N_26658,N_19728,N_18410);
nand U26659 (N_26659,N_18902,N_14919);
and U26660 (N_26660,N_10523,N_19222);
nand U26661 (N_26661,N_13672,N_13155);
or U26662 (N_26662,N_10854,N_19800);
and U26663 (N_26663,N_19289,N_18792);
or U26664 (N_26664,N_13658,N_12608);
or U26665 (N_26665,N_16911,N_10420);
nor U26666 (N_26666,N_12508,N_15037);
nor U26667 (N_26667,N_18344,N_12633);
nand U26668 (N_26668,N_17328,N_16081);
or U26669 (N_26669,N_10070,N_16058);
nand U26670 (N_26670,N_12400,N_11186);
nand U26671 (N_26671,N_13798,N_11356);
and U26672 (N_26672,N_11325,N_15530);
or U26673 (N_26673,N_13601,N_10398);
nor U26674 (N_26674,N_11011,N_11055);
nor U26675 (N_26675,N_10222,N_11033);
and U26676 (N_26676,N_13733,N_11794);
and U26677 (N_26677,N_17410,N_14737);
nand U26678 (N_26678,N_11257,N_15015);
xnor U26679 (N_26679,N_19791,N_14877);
nand U26680 (N_26680,N_18332,N_16117);
or U26681 (N_26681,N_17893,N_16098);
and U26682 (N_26682,N_14406,N_18928);
nor U26683 (N_26683,N_14294,N_13146);
nor U26684 (N_26684,N_11340,N_10685);
nor U26685 (N_26685,N_14300,N_10300);
nor U26686 (N_26686,N_18087,N_11241);
nand U26687 (N_26687,N_15974,N_11019);
nor U26688 (N_26688,N_18529,N_15224);
and U26689 (N_26689,N_10473,N_14520);
and U26690 (N_26690,N_17001,N_13342);
nor U26691 (N_26691,N_16257,N_15185);
or U26692 (N_26692,N_12194,N_18946);
nand U26693 (N_26693,N_12739,N_12600);
nor U26694 (N_26694,N_14579,N_11241);
or U26695 (N_26695,N_17546,N_16300);
or U26696 (N_26696,N_14093,N_16371);
and U26697 (N_26697,N_15951,N_12149);
nor U26698 (N_26698,N_16072,N_12172);
and U26699 (N_26699,N_14658,N_19014);
or U26700 (N_26700,N_18991,N_18374);
or U26701 (N_26701,N_12598,N_10126);
nand U26702 (N_26702,N_19843,N_19889);
nor U26703 (N_26703,N_18701,N_18560);
nor U26704 (N_26704,N_18633,N_16840);
or U26705 (N_26705,N_19969,N_18490);
nor U26706 (N_26706,N_14119,N_17163);
or U26707 (N_26707,N_16599,N_15822);
nand U26708 (N_26708,N_13163,N_12262);
nand U26709 (N_26709,N_12786,N_19415);
and U26710 (N_26710,N_14187,N_16800);
and U26711 (N_26711,N_19568,N_17228);
nor U26712 (N_26712,N_10247,N_10041);
nor U26713 (N_26713,N_14538,N_17302);
or U26714 (N_26714,N_13694,N_18587);
or U26715 (N_26715,N_11501,N_10442);
nor U26716 (N_26716,N_15859,N_19829);
nor U26717 (N_26717,N_15985,N_13834);
and U26718 (N_26718,N_12090,N_14159);
or U26719 (N_26719,N_19314,N_16002);
nand U26720 (N_26720,N_14761,N_11997);
nand U26721 (N_26721,N_17069,N_17840);
xor U26722 (N_26722,N_13752,N_13853);
nand U26723 (N_26723,N_10956,N_18959);
or U26724 (N_26724,N_17867,N_13963);
nor U26725 (N_26725,N_19639,N_14485);
or U26726 (N_26726,N_10339,N_10410);
or U26727 (N_26727,N_11493,N_11923);
nor U26728 (N_26728,N_10484,N_13625);
or U26729 (N_26729,N_15528,N_15158);
or U26730 (N_26730,N_18717,N_14275);
nor U26731 (N_26731,N_13691,N_16718);
and U26732 (N_26732,N_15977,N_16025);
and U26733 (N_26733,N_17254,N_18771);
and U26734 (N_26734,N_10154,N_17018);
nand U26735 (N_26735,N_10090,N_12705);
nor U26736 (N_26736,N_15665,N_15585);
or U26737 (N_26737,N_13302,N_15191);
and U26738 (N_26738,N_17220,N_11498);
or U26739 (N_26739,N_11636,N_17500);
nor U26740 (N_26740,N_16786,N_14198);
or U26741 (N_26741,N_11314,N_12642);
or U26742 (N_26742,N_19654,N_13994);
nand U26743 (N_26743,N_11611,N_18001);
or U26744 (N_26744,N_11686,N_16544);
and U26745 (N_26745,N_15483,N_11982);
or U26746 (N_26746,N_18399,N_19023);
and U26747 (N_26747,N_11220,N_18777);
or U26748 (N_26748,N_18097,N_19960);
nor U26749 (N_26749,N_17415,N_12464);
and U26750 (N_26750,N_10636,N_13426);
or U26751 (N_26751,N_17414,N_19915);
nor U26752 (N_26752,N_12826,N_12766);
nor U26753 (N_26753,N_19674,N_18484);
nand U26754 (N_26754,N_15532,N_17052);
nand U26755 (N_26755,N_16618,N_18329);
nor U26756 (N_26756,N_11183,N_19984);
xnor U26757 (N_26757,N_18771,N_11463);
nor U26758 (N_26758,N_10423,N_18508);
nor U26759 (N_26759,N_15931,N_16761);
nand U26760 (N_26760,N_15734,N_11726);
or U26761 (N_26761,N_10301,N_15166);
nor U26762 (N_26762,N_17342,N_13005);
or U26763 (N_26763,N_13291,N_16649);
and U26764 (N_26764,N_13623,N_13955);
nor U26765 (N_26765,N_11500,N_11435);
or U26766 (N_26766,N_19337,N_14084);
nor U26767 (N_26767,N_11994,N_15065);
and U26768 (N_26768,N_16043,N_19030);
nand U26769 (N_26769,N_12490,N_10808);
and U26770 (N_26770,N_11819,N_12890);
nor U26771 (N_26771,N_17850,N_17994);
nand U26772 (N_26772,N_18106,N_10608);
xor U26773 (N_26773,N_12653,N_19612);
nand U26774 (N_26774,N_13253,N_16514);
and U26775 (N_26775,N_13636,N_18232);
nor U26776 (N_26776,N_15612,N_19843);
nor U26777 (N_26777,N_19756,N_13073);
or U26778 (N_26778,N_10811,N_11425);
and U26779 (N_26779,N_19312,N_15151);
xnor U26780 (N_26780,N_12393,N_11196);
and U26781 (N_26781,N_16058,N_10417);
nand U26782 (N_26782,N_12730,N_12737);
and U26783 (N_26783,N_19186,N_11251);
or U26784 (N_26784,N_10016,N_14645);
and U26785 (N_26785,N_12574,N_13685);
nor U26786 (N_26786,N_14507,N_10212);
nor U26787 (N_26787,N_12489,N_19427);
nand U26788 (N_26788,N_16773,N_14586);
xor U26789 (N_26789,N_10200,N_16700);
or U26790 (N_26790,N_17716,N_17825);
nor U26791 (N_26791,N_19909,N_12108);
nor U26792 (N_26792,N_10864,N_18371);
nand U26793 (N_26793,N_18309,N_15592);
nand U26794 (N_26794,N_17140,N_16356);
or U26795 (N_26795,N_19210,N_16436);
nand U26796 (N_26796,N_15201,N_17128);
nand U26797 (N_26797,N_12551,N_19433);
and U26798 (N_26798,N_13890,N_11247);
nor U26799 (N_26799,N_14524,N_13316);
and U26800 (N_26800,N_14263,N_10528);
or U26801 (N_26801,N_18597,N_17903);
nor U26802 (N_26802,N_15027,N_19998);
nand U26803 (N_26803,N_18581,N_18947);
xnor U26804 (N_26804,N_18801,N_19336);
or U26805 (N_26805,N_10347,N_17601);
xor U26806 (N_26806,N_12172,N_16523);
or U26807 (N_26807,N_13443,N_16303);
xnor U26808 (N_26808,N_12236,N_13084);
or U26809 (N_26809,N_18395,N_10344);
nor U26810 (N_26810,N_12723,N_10178);
nand U26811 (N_26811,N_13846,N_10515);
nor U26812 (N_26812,N_10543,N_19338);
nand U26813 (N_26813,N_18908,N_16034);
or U26814 (N_26814,N_14926,N_17592);
nor U26815 (N_26815,N_15052,N_14471);
and U26816 (N_26816,N_16988,N_11815);
nand U26817 (N_26817,N_13902,N_11424);
nand U26818 (N_26818,N_16733,N_19026);
nor U26819 (N_26819,N_14425,N_18608);
and U26820 (N_26820,N_17254,N_17765);
nand U26821 (N_26821,N_16638,N_12891);
and U26822 (N_26822,N_11577,N_19571);
nor U26823 (N_26823,N_16551,N_12130);
xnor U26824 (N_26824,N_18897,N_18081);
or U26825 (N_26825,N_13817,N_18758);
or U26826 (N_26826,N_15164,N_16786);
nand U26827 (N_26827,N_10542,N_18003);
and U26828 (N_26828,N_16153,N_12624);
nor U26829 (N_26829,N_13993,N_13003);
and U26830 (N_26830,N_19201,N_11779);
or U26831 (N_26831,N_16796,N_14547);
and U26832 (N_26832,N_11600,N_18389);
nor U26833 (N_26833,N_15939,N_10907);
and U26834 (N_26834,N_18863,N_18426);
or U26835 (N_26835,N_17892,N_13736);
nand U26836 (N_26836,N_15390,N_16020);
and U26837 (N_26837,N_12043,N_11554);
nand U26838 (N_26838,N_18608,N_19181);
nor U26839 (N_26839,N_11457,N_19182);
xnor U26840 (N_26840,N_18484,N_18679);
nand U26841 (N_26841,N_19551,N_14339);
and U26842 (N_26842,N_14668,N_11990);
or U26843 (N_26843,N_17625,N_14696);
nand U26844 (N_26844,N_19731,N_16388);
nor U26845 (N_26845,N_13832,N_10673);
nand U26846 (N_26846,N_12751,N_18037);
or U26847 (N_26847,N_16839,N_18600);
nand U26848 (N_26848,N_11716,N_17600);
nand U26849 (N_26849,N_19307,N_16330);
or U26850 (N_26850,N_19081,N_16977);
nand U26851 (N_26851,N_15194,N_19321);
and U26852 (N_26852,N_11807,N_19701);
nor U26853 (N_26853,N_12640,N_18783);
nand U26854 (N_26854,N_17072,N_14567);
nand U26855 (N_26855,N_15605,N_18658);
or U26856 (N_26856,N_15441,N_19706);
or U26857 (N_26857,N_12007,N_12650);
or U26858 (N_26858,N_10521,N_14195);
or U26859 (N_26859,N_13744,N_10963);
nand U26860 (N_26860,N_17721,N_15837);
nor U26861 (N_26861,N_15347,N_10212);
or U26862 (N_26862,N_14915,N_16802);
xnor U26863 (N_26863,N_12729,N_15563);
nand U26864 (N_26864,N_17590,N_19186);
xnor U26865 (N_26865,N_14686,N_13077);
or U26866 (N_26866,N_14154,N_19115);
and U26867 (N_26867,N_12297,N_15623);
or U26868 (N_26868,N_18419,N_17377);
xnor U26869 (N_26869,N_14188,N_14634);
or U26870 (N_26870,N_14386,N_10161);
nand U26871 (N_26871,N_10768,N_18365);
or U26872 (N_26872,N_19009,N_18099);
nand U26873 (N_26873,N_17345,N_13978);
nor U26874 (N_26874,N_19213,N_15280);
nor U26875 (N_26875,N_19630,N_13221);
nand U26876 (N_26876,N_10613,N_10066);
nor U26877 (N_26877,N_19240,N_16266);
xor U26878 (N_26878,N_16253,N_12240);
or U26879 (N_26879,N_12310,N_13715);
nor U26880 (N_26880,N_10810,N_17742);
and U26881 (N_26881,N_18776,N_10856);
nand U26882 (N_26882,N_19592,N_11039);
nand U26883 (N_26883,N_19975,N_12849);
nor U26884 (N_26884,N_13565,N_16855);
xnor U26885 (N_26885,N_13230,N_17923);
nor U26886 (N_26886,N_13131,N_14699);
nand U26887 (N_26887,N_15690,N_12895);
or U26888 (N_26888,N_14963,N_17301);
or U26889 (N_26889,N_17570,N_15430);
nand U26890 (N_26890,N_16734,N_14267);
nor U26891 (N_26891,N_12796,N_16071);
nor U26892 (N_26892,N_19983,N_14462);
and U26893 (N_26893,N_10477,N_17538);
and U26894 (N_26894,N_11121,N_15927);
nor U26895 (N_26895,N_17465,N_11716);
nand U26896 (N_26896,N_17887,N_16363);
or U26897 (N_26897,N_18897,N_18758);
nor U26898 (N_26898,N_13703,N_10401);
or U26899 (N_26899,N_10537,N_15325);
nor U26900 (N_26900,N_11070,N_11318);
or U26901 (N_26901,N_16284,N_12317);
nor U26902 (N_26902,N_13957,N_17185);
and U26903 (N_26903,N_12656,N_17468);
nor U26904 (N_26904,N_18793,N_12492);
or U26905 (N_26905,N_16844,N_12511);
nor U26906 (N_26906,N_17609,N_11852);
xor U26907 (N_26907,N_19317,N_16257);
and U26908 (N_26908,N_19902,N_10774);
or U26909 (N_26909,N_14805,N_18925);
or U26910 (N_26910,N_14618,N_11318);
and U26911 (N_26911,N_17987,N_10917);
nor U26912 (N_26912,N_15233,N_15526);
or U26913 (N_26913,N_12350,N_18271);
and U26914 (N_26914,N_15182,N_10551);
and U26915 (N_26915,N_15694,N_11884);
and U26916 (N_26916,N_17595,N_18192);
or U26917 (N_26917,N_11514,N_19169);
nand U26918 (N_26918,N_15531,N_16669);
or U26919 (N_26919,N_13589,N_12394);
or U26920 (N_26920,N_12030,N_19587);
xnor U26921 (N_26921,N_11100,N_13855);
nand U26922 (N_26922,N_18382,N_14448);
nor U26923 (N_26923,N_16857,N_12282);
nor U26924 (N_26924,N_14037,N_14001);
nand U26925 (N_26925,N_19070,N_19865);
nor U26926 (N_26926,N_14431,N_10918);
and U26927 (N_26927,N_13290,N_13830);
and U26928 (N_26928,N_19447,N_11030);
and U26929 (N_26929,N_14483,N_16873);
or U26930 (N_26930,N_11340,N_12917);
nor U26931 (N_26931,N_16674,N_11334);
nor U26932 (N_26932,N_14209,N_13294);
or U26933 (N_26933,N_13822,N_11379);
nor U26934 (N_26934,N_14647,N_10659);
nand U26935 (N_26935,N_15780,N_18039);
and U26936 (N_26936,N_12583,N_19265);
or U26937 (N_26937,N_10400,N_19561);
nor U26938 (N_26938,N_12237,N_15303);
nor U26939 (N_26939,N_17345,N_10975);
or U26940 (N_26940,N_10000,N_17629);
xor U26941 (N_26941,N_10354,N_12029);
nor U26942 (N_26942,N_13126,N_10734);
or U26943 (N_26943,N_13965,N_15304);
xor U26944 (N_26944,N_15929,N_11790);
or U26945 (N_26945,N_13303,N_16237);
nor U26946 (N_26946,N_12259,N_15393);
nor U26947 (N_26947,N_13328,N_19579);
and U26948 (N_26948,N_17911,N_17418);
nor U26949 (N_26949,N_16353,N_14994);
xor U26950 (N_26950,N_11689,N_16836);
nor U26951 (N_26951,N_19750,N_15329);
nand U26952 (N_26952,N_11014,N_18976);
nand U26953 (N_26953,N_14347,N_10491);
nand U26954 (N_26954,N_14036,N_10186);
nand U26955 (N_26955,N_16608,N_11178);
nor U26956 (N_26956,N_16104,N_18990);
or U26957 (N_26957,N_16049,N_14322);
nor U26958 (N_26958,N_18892,N_11460);
xor U26959 (N_26959,N_12832,N_13244);
and U26960 (N_26960,N_19024,N_16329);
or U26961 (N_26961,N_18337,N_17628);
nor U26962 (N_26962,N_16519,N_16828);
or U26963 (N_26963,N_14418,N_11466);
nor U26964 (N_26964,N_17820,N_15390);
xnor U26965 (N_26965,N_18906,N_11127);
nand U26966 (N_26966,N_11792,N_14478);
nand U26967 (N_26967,N_17527,N_14254);
and U26968 (N_26968,N_10700,N_19605);
xor U26969 (N_26969,N_16698,N_16339);
nand U26970 (N_26970,N_19678,N_16246);
and U26971 (N_26971,N_15881,N_19512);
or U26972 (N_26972,N_14203,N_14375);
nand U26973 (N_26973,N_12000,N_12750);
or U26974 (N_26974,N_16869,N_10112);
nor U26975 (N_26975,N_15485,N_14285);
or U26976 (N_26976,N_17770,N_18655);
and U26977 (N_26977,N_18066,N_19334);
nand U26978 (N_26978,N_19312,N_11603);
xnor U26979 (N_26979,N_17422,N_19874);
nand U26980 (N_26980,N_17908,N_14119);
nand U26981 (N_26981,N_17623,N_14884);
nand U26982 (N_26982,N_14303,N_17940);
nor U26983 (N_26983,N_18889,N_17447);
nor U26984 (N_26984,N_12955,N_11770);
nand U26985 (N_26985,N_10956,N_17927);
nand U26986 (N_26986,N_17844,N_10518);
nand U26987 (N_26987,N_16870,N_13750);
nand U26988 (N_26988,N_13878,N_19918);
or U26989 (N_26989,N_18194,N_12238);
xor U26990 (N_26990,N_12527,N_16325);
nand U26991 (N_26991,N_12787,N_15930);
or U26992 (N_26992,N_15320,N_19428);
and U26993 (N_26993,N_12607,N_13911);
nor U26994 (N_26994,N_11838,N_17231);
or U26995 (N_26995,N_16804,N_18719);
or U26996 (N_26996,N_12381,N_15708);
nor U26997 (N_26997,N_16858,N_13288);
nand U26998 (N_26998,N_12140,N_15898);
and U26999 (N_26999,N_17220,N_19956);
nor U27000 (N_27000,N_12291,N_11077);
nor U27001 (N_27001,N_15899,N_16473);
or U27002 (N_27002,N_11254,N_13025);
nand U27003 (N_27003,N_12006,N_18557);
xor U27004 (N_27004,N_14135,N_19279);
and U27005 (N_27005,N_10285,N_12108);
or U27006 (N_27006,N_19987,N_16023);
or U27007 (N_27007,N_19110,N_15075);
or U27008 (N_27008,N_12928,N_19274);
and U27009 (N_27009,N_13972,N_19219);
xnor U27010 (N_27010,N_16563,N_11497);
or U27011 (N_27011,N_15595,N_13236);
nor U27012 (N_27012,N_14008,N_16946);
or U27013 (N_27013,N_17583,N_18219);
or U27014 (N_27014,N_12037,N_19552);
or U27015 (N_27015,N_18317,N_12073);
nor U27016 (N_27016,N_17756,N_19121);
or U27017 (N_27017,N_12056,N_15598);
and U27018 (N_27018,N_12307,N_17393);
nand U27019 (N_27019,N_15665,N_18618);
nand U27020 (N_27020,N_13927,N_17767);
and U27021 (N_27021,N_15981,N_17603);
and U27022 (N_27022,N_12289,N_14183);
or U27023 (N_27023,N_10304,N_15788);
or U27024 (N_27024,N_19833,N_10563);
or U27025 (N_27025,N_11905,N_17659);
xnor U27026 (N_27026,N_13751,N_12235);
nand U27027 (N_27027,N_16141,N_10690);
or U27028 (N_27028,N_13769,N_11955);
nand U27029 (N_27029,N_14404,N_12458);
or U27030 (N_27030,N_16635,N_16335);
xnor U27031 (N_27031,N_12545,N_10677);
nand U27032 (N_27032,N_15872,N_14846);
and U27033 (N_27033,N_18649,N_15631);
nor U27034 (N_27034,N_12337,N_17064);
or U27035 (N_27035,N_19183,N_10425);
xor U27036 (N_27036,N_17868,N_19604);
or U27037 (N_27037,N_19906,N_11108);
nand U27038 (N_27038,N_13309,N_18851);
and U27039 (N_27039,N_18381,N_15567);
nand U27040 (N_27040,N_10364,N_19204);
nor U27041 (N_27041,N_11061,N_19216);
nor U27042 (N_27042,N_15287,N_14679);
nor U27043 (N_27043,N_19292,N_16076);
nand U27044 (N_27044,N_17878,N_12875);
or U27045 (N_27045,N_17388,N_15184);
xor U27046 (N_27046,N_13151,N_16961);
nand U27047 (N_27047,N_16733,N_14093);
or U27048 (N_27048,N_10622,N_12014);
nor U27049 (N_27049,N_12041,N_15922);
nor U27050 (N_27050,N_10727,N_19047);
nand U27051 (N_27051,N_11442,N_17312);
nor U27052 (N_27052,N_17970,N_13834);
nor U27053 (N_27053,N_12105,N_13373);
nand U27054 (N_27054,N_13286,N_10981);
and U27055 (N_27055,N_15469,N_11894);
nand U27056 (N_27056,N_13117,N_15239);
xnor U27057 (N_27057,N_19167,N_15975);
nor U27058 (N_27058,N_13629,N_13138);
nand U27059 (N_27059,N_18757,N_16101);
nor U27060 (N_27060,N_15159,N_16155);
nor U27061 (N_27061,N_10316,N_11937);
and U27062 (N_27062,N_17281,N_18682);
nand U27063 (N_27063,N_12959,N_12001);
xor U27064 (N_27064,N_10864,N_16897);
or U27065 (N_27065,N_17509,N_17279);
nor U27066 (N_27066,N_19653,N_12081);
nor U27067 (N_27067,N_19325,N_14791);
nor U27068 (N_27068,N_14612,N_12444);
nor U27069 (N_27069,N_13015,N_10621);
nand U27070 (N_27070,N_10331,N_14425);
nand U27071 (N_27071,N_10644,N_11358);
and U27072 (N_27072,N_11467,N_13023);
xor U27073 (N_27073,N_14252,N_16743);
nand U27074 (N_27074,N_16495,N_12437);
and U27075 (N_27075,N_18889,N_14187);
nand U27076 (N_27076,N_11470,N_17730);
nor U27077 (N_27077,N_18625,N_19106);
nor U27078 (N_27078,N_13526,N_19178);
and U27079 (N_27079,N_10802,N_18042);
and U27080 (N_27080,N_10746,N_11249);
and U27081 (N_27081,N_16153,N_10735);
and U27082 (N_27082,N_16790,N_18370);
and U27083 (N_27083,N_19208,N_16257);
nand U27084 (N_27084,N_16143,N_10422);
and U27085 (N_27085,N_13836,N_19552);
nand U27086 (N_27086,N_13644,N_19341);
or U27087 (N_27087,N_19448,N_14892);
nand U27088 (N_27088,N_11724,N_12598);
nor U27089 (N_27089,N_11377,N_10307);
and U27090 (N_27090,N_13372,N_10496);
and U27091 (N_27091,N_13705,N_15265);
and U27092 (N_27092,N_13953,N_17631);
and U27093 (N_27093,N_19184,N_17563);
nor U27094 (N_27094,N_10202,N_19560);
nor U27095 (N_27095,N_15059,N_18982);
nor U27096 (N_27096,N_14754,N_19267);
xnor U27097 (N_27097,N_11661,N_13887);
nor U27098 (N_27098,N_15625,N_12311);
or U27099 (N_27099,N_10552,N_12043);
nand U27100 (N_27100,N_12371,N_10519);
or U27101 (N_27101,N_11607,N_10669);
or U27102 (N_27102,N_14928,N_12917);
xor U27103 (N_27103,N_16876,N_17537);
and U27104 (N_27104,N_10180,N_19037);
nand U27105 (N_27105,N_14087,N_15882);
nor U27106 (N_27106,N_11819,N_15460);
nand U27107 (N_27107,N_12606,N_17488);
xor U27108 (N_27108,N_12431,N_14590);
nand U27109 (N_27109,N_18532,N_13649);
nand U27110 (N_27110,N_14228,N_15051);
or U27111 (N_27111,N_11311,N_11391);
xor U27112 (N_27112,N_11592,N_14295);
xor U27113 (N_27113,N_19592,N_15527);
nor U27114 (N_27114,N_17945,N_12140);
or U27115 (N_27115,N_12326,N_13129);
and U27116 (N_27116,N_13711,N_15881);
nand U27117 (N_27117,N_14782,N_13788);
nor U27118 (N_27118,N_12889,N_12842);
and U27119 (N_27119,N_19531,N_15239);
or U27120 (N_27120,N_11082,N_17996);
or U27121 (N_27121,N_19041,N_16559);
nand U27122 (N_27122,N_15986,N_17919);
nand U27123 (N_27123,N_10233,N_15948);
nor U27124 (N_27124,N_13089,N_17698);
nor U27125 (N_27125,N_18576,N_17755);
nor U27126 (N_27126,N_12300,N_11159);
nand U27127 (N_27127,N_19431,N_15287);
nand U27128 (N_27128,N_11907,N_13865);
nand U27129 (N_27129,N_12385,N_14707);
nor U27130 (N_27130,N_18479,N_13396);
nand U27131 (N_27131,N_11445,N_16293);
and U27132 (N_27132,N_19476,N_12463);
and U27133 (N_27133,N_11136,N_10702);
or U27134 (N_27134,N_13961,N_19116);
nand U27135 (N_27135,N_16986,N_11912);
nor U27136 (N_27136,N_15920,N_18236);
nor U27137 (N_27137,N_15093,N_11150);
nor U27138 (N_27138,N_18228,N_11314);
and U27139 (N_27139,N_19875,N_13320);
and U27140 (N_27140,N_12715,N_16187);
nor U27141 (N_27141,N_14325,N_11628);
nand U27142 (N_27142,N_12980,N_13467);
or U27143 (N_27143,N_14962,N_18904);
xor U27144 (N_27144,N_17176,N_17460);
or U27145 (N_27145,N_17537,N_12033);
xnor U27146 (N_27146,N_17101,N_10066);
nand U27147 (N_27147,N_12204,N_10860);
nor U27148 (N_27148,N_17907,N_18846);
or U27149 (N_27149,N_17012,N_15160);
nor U27150 (N_27150,N_11928,N_19795);
or U27151 (N_27151,N_14464,N_10891);
nor U27152 (N_27152,N_15622,N_12373);
nor U27153 (N_27153,N_13636,N_16056);
xor U27154 (N_27154,N_13486,N_16438);
or U27155 (N_27155,N_18814,N_13409);
or U27156 (N_27156,N_10435,N_15632);
nand U27157 (N_27157,N_11312,N_19541);
or U27158 (N_27158,N_12220,N_17991);
nand U27159 (N_27159,N_11719,N_15781);
xnor U27160 (N_27160,N_15973,N_16298);
nor U27161 (N_27161,N_18098,N_17950);
and U27162 (N_27162,N_14621,N_15141);
and U27163 (N_27163,N_11776,N_14321);
and U27164 (N_27164,N_19890,N_19960);
and U27165 (N_27165,N_18091,N_13252);
nor U27166 (N_27166,N_10798,N_12957);
or U27167 (N_27167,N_11342,N_16118);
nand U27168 (N_27168,N_16501,N_10900);
and U27169 (N_27169,N_14127,N_11254);
nand U27170 (N_27170,N_16085,N_16370);
xor U27171 (N_27171,N_10945,N_16768);
or U27172 (N_27172,N_16182,N_14402);
or U27173 (N_27173,N_18650,N_10170);
or U27174 (N_27174,N_10864,N_11460);
and U27175 (N_27175,N_12591,N_15155);
and U27176 (N_27176,N_17770,N_18330);
or U27177 (N_27177,N_11808,N_13020);
nor U27178 (N_27178,N_15045,N_14779);
nand U27179 (N_27179,N_13034,N_19091);
xor U27180 (N_27180,N_18722,N_16672);
nand U27181 (N_27181,N_10245,N_18384);
xnor U27182 (N_27182,N_18744,N_16643);
and U27183 (N_27183,N_14352,N_11879);
or U27184 (N_27184,N_16565,N_13171);
nand U27185 (N_27185,N_11186,N_10045);
nand U27186 (N_27186,N_16641,N_15111);
nor U27187 (N_27187,N_16252,N_13538);
or U27188 (N_27188,N_17876,N_16855);
nand U27189 (N_27189,N_17591,N_11486);
nand U27190 (N_27190,N_16283,N_10423);
nor U27191 (N_27191,N_11626,N_10400);
nand U27192 (N_27192,N_19057,N_18806);
and U27193 (N_27193,N_16467,N_15045);
xor U27194 (N_27194,N_18607,N_14429);
nand U27195 (N_27195,N_13522,N_14291);
and U27196 (N_27196,N_19220,N_15550);
nor U27197 (N_27197,N_18320,N_10720);
nand U27198 (N_27198,N_11003,N_15726);
or U27199 (N_27199,N_13765,N_19043);
or U27200 (N_27200,N_17190,N_18848);
nand U27201 (N_27201,N_14009,N_13342);
and U27202 (N_27202,N_11327,N_16494);
xnor U27203 (N_27203,N_12536,N_14887);
nor U27204 (N_27204,N_18753,N_17387);
and U27205 (N_27205,N_12779,N_19651);
and U27206 (N_27206,N_14948,N_12134);
or U27207 (N_27207,N_17194,N_11209);
and U27208 (N_27208,N_10955,N_17818);
or U27209 (N_27209,N_18267,N_12191);
nor U27210 (N_27210,N_16607,N_17122);
nor U27211 (N_27211,N_11181,N_19970);
nand U27212 (N_27212,N_11747,N_16251);
nor U27213 (N_27213,N_15920,N_19603);
nand U27214 (N_27214,N_18945,N_12305);
xnor U27215 (N_27215,N_17064,N_17464);
and U27216 (N_27216,N_19770,N_13260);
nor U27217 (N_27217,N_17166,N_18170);
or U27218 (N_27218,N_14449,N_12454);
nor U27219 (N_27219,N_17888,N_17301);
nand U27220 (N_27220,N_16640,N_17870);
or U27221 (N_27221,N_11262,N_10543);
and U27222 (N_27222,N_10712,N_16278);
xor U27223 (N_27223,N_14356,N_15380);
and U27224 (N_27224,N_14932,N_12943);
nor U27225 (N_27225,N_17011,N_11661);
and U27226 (N_27226,N_16930,N_14765);
and U27227 (N_27227,N_13892,N_18323);
nand U27228 (N_27228,N_19995,N_16259);
nand U27229 (N_27229,N_19702,N_12477);
nor U27230 (N_27230,N_16955,N_16465);
nand U27231 (N_27231,N_18567,N_15778);
and U27232 (N_27232,N_17348,N_12125);
and U27233 (N_27233,N_16817,N_13723);
nand U27234 (N_27234,N_10096,N_15918);
nor U27235 (N_27235,N_18073,N_15597);
nor U27236 (N_27236,N_18354,N_17018);
and U27237 (N_27237,N_17963,N_15898);
nand U27238 (N_27238,N_18919,N_13367);
nor U27239 (N_27239,N_19031,N_16107);
nor U27240 (N_27240,N_18100,N_16576);
and U27241 (N_27241,N_18558,N_19492);
or U27242 (N_27242,N_15936,N_17098);
or U27243 (N_27243,N_17421,N_13255);
or U27244 (N_27244,N_16186,N_10727);
or U27245 (N_27245,N_12410,N_10293);
and U27246 (N_27246,N_15276,N_13679);
or U27247 (N_27247,N_17713,N_10732);
nand U27248 (N_27248,N_14473,N_15469);
and U27249 (N_27249,N_13213,N_14957);
xor U27250 (N_27250,N_13320,N_13300);
nor U27251 (N_27251,N_10334,N_11575);
xor U27252 (N_27252,N_10419,N_18310);
or U27253 (N_27253,N_15996,N_18175);
nand U27254 (N_27254,N_15843,N_13444);
and U27255 (N_27255,N_15026,N_16743);
or U27256 (N_27256,N_14257,N_16022);
nand U27257 (N_27257,N_10232,N_16669);
and U27258 (N_27258,N_10340,N_18142);
nor U27259 (N_27259,N_18541,N_14654);
xnor U27260 (N_27260,N_16319,N_13452);
and U27261 (N_27261,N_12487,N_16746);
nor U27262 (N_27262,N_12135,N_16008);
nor U27263 (N_27263,N_16592,N_12823);
nand U27264 (N_27264,N_11393,N_17108);
and U27265 (N_27265,N_10588,N_13160);
nand U27266 (N_27266,N_11035,N_17109);
nor U27267 (N_27267,N_15977,N_10389);
nand U27268 (N_27268,N_16441,N_17395);
nor U27269 (N_27269,N_12878,N_11824);
xnor U27270 (N_27270,N_15742,N_15977);
or U27271 (N_27271,N_18863,N_14047);
nor U27272 (N_27272,N_11468,N_17030);
or U27273 (N_27273,N_18571,N_11682);
nor U27274 (N_27274,N_16020,N_14830);
and U27275 (N_27275,N_12106,N_16984);
nor U27276 (N_27276,N_12319,N_14250);
nand U27277 (N_27277,N_13173,N_19050);
xnor U27278 (N_27278,N_19021,N_11173);
nor U27279 (N_27279,N_11405,N_15844);
nand U27280 (N_27280,N_19766,N_16877);
and U27281 (N_27281,N_15862,N_18831);
or U27282 (N_27282,N_12574,N_19594);
and U27283 (N_27283,N_10089,N_11755);
or U27284 (N_27284,N_12110,N_11231);
or U27285 (N_27285,N_13249,N_13184);
or U27286 (N_27286,N_11546,N_14823);
nor U27287 (N_27287,N_16221,N_14870);
nor U27288 (N_27288,N_14300,N_12767);
nand U27289 (N_27289,N_15733,N_15396);
nand U27290 (N_27290,N_17699,N_13872);
or U27291 (N_27291,N_11986,N_19807);
nand U27292 (N_27292,N_15887,N_12520);
nor U27293 (N_27293,N_18694,N_12159);
xnor U27294 (N_27294,N_12919,N_14016);
xor U27295 (N_27295,N_18352,N_10773);
nand U27296 (N_27296,N_18977,N_19608);
and U27297 (N_27297,N_15178,N_13873);
and U27298 (N_27298,N_11888,N_18195);
or U27299 (N_27299,N_13706,N_17506);
nand U27300 (N_27300,N_14206,N_18924);
xor U27301 (N_27301,N_17771,N_13815);
and U27302 (N_27302,N_17641,N_18994);
or U27303 (N_27303,N_13338,N_16227);
or U27304 (N_27304,N_14713,N_12089);
nand U27305 (N_27305,N_14502,N_18855);
or U27306 (N_27306,N_16023,N_11728);
and U27307 (N_27307,N_17254,N_13467);
nor U27308 (N_27308,N_12268,N_16703);
nor U27309 (N_27309,N_19425,N_15875);
and U27310 (N_27310,N_17958,N_19417);
or U27311 (N_27311,N_13465,N_12464);
xnor U27312 (N_27312,N_17776,N_11229);
or U27313 (N_27313,N_12117,N_19913);
and U27314 (N_27314,N_17240,N_13973);
xnor U27315 (N_27315,N_13209,N_17052);
nand U27316 (N_27316,N_14022,N_12383);
nor U27317 (N_27317,N_14751,N_11723);
and U27318 (N_27318,N_16248,N_15446);
or U27319 (N_27319,N_14849,N_11763);
and U27320 (N_27320,N_15682,N_10888);
or U27321 (N_27321,N_14907,N_15907);
xnor U27322 (N_27322,N_14498,N_19338);
and U27323 (N_27323,N_15845,N_11933);
or U27324 (N_27324,N_11747,N_13515);
and U27325 (N_27325,N_15636,N_15087);
and U27326 (N_27326,N_11706,N_15627);
nor U27327 (N_27327,N_15016,N_16451);
nor U27328 (N_27328,N_13769,N_15914);
nand U27329 (N_27329,N_10461,N_12005);
or U27330 (N_27330,N_19745,N_18909);
nor U27331 (N_27331,N_10649,N_13322);
and U27332 (N_27332,N_15443,N_12060);
xnor U27333 (N_27333,N_10455,N_19582);
nor U27334 (N_27334,N_15233,N_14437);
xnor U27335 (N_27335,N_19097,N_19143);
or U27336 (N_27336,N_11196,N_16281);
and U27337 (N_27337,N_18828,N_19227);
nand U27338 (N_27338,N_16453,N_18024);
nand U27339 (N_27339,N_14347,N_17375);
and U27340 (N_27340,N_12252,N_10046);
nand U27341 (N_27341,N_11436,N_17969);
or U27342 (N_27342,N_19802,N_19946);
and U27343 (N_27343,N_19719,N_17550);
or U27344 (N_27344,N_11375,N_17932);
or U27345 (N_27345,N_13823,N_19648);
xor U27346 (N_27346,N_13133,N_15427);
nor U27347 (N_27347,N_12735,N_10464);
xnor U27348 (N_27348,N_18323,N_15598);
nor U27349 (N_27349,N_19835,N_17412);
nor U27350 (N_27350,N_11573,N_17229);
nand U27351 (N_27351,N_12983,N_14016);
nor U27352 (N_27352,N_12201,N_10552);
xor U27353 (N_27353,N_11434,N_10856);
or U27354 (N_27354,N_15621,N_18866);
xor U27355 (N_27355,N_11708,N_11138);
nor U27356 (N_27356,N_13178,N_11278);
nor U27357 (N_27357,N_17772,N_18909);
xnor U27358 (N_27358,N_11604,N_13452);
or U27359 (N_27359,N_18318,N_12112);
or U27360 (N_27360,N_19220,N_11077);
nor U27361 (N_27361,N_13853,N_18247);
nor U27362 (N_27362,N_19645,N_13707);
nor U27363 (N_27363,N_16604,N_10910);
xnor U27364 (N_27364,N_15900,N_10508);
nor U27365 (N_27365,N_19236,N_18001);
nand U27366 (N_27366,N_11469,N_13121);
and U27367 (N_27367,N_19868,N_12886);
nand U27368 (N_27368,N_14952,N_17409);
nor U27369 (N_27369,N_14194,N_12657);
nand U27370 (N_27370,N_18556,N_16707);
and U27371 (N_27371,N_19045,N_11930);
nor U27372 (N_27372,N_17078,N_19422);
nand U27373 (N_27373,N_19094,N_17485);
nor U27374 (N_27374,N_18885,N_16621);
or U27375 (N_27375,N_14907,N_17741);
nor U27376 (N_27376,N_10001,N_12358);
or U27377 (N_27377,N_13853,N_12881);
nand U27378 (N_27378,N_12449,N_17268);
nand U27379 (N_27379,N_19189,N_16505);
nand U27380 (N_27380,N_18621,N_12243);
nand U27381 (N_27381,N_11609,N_12676);
or U27382 (N_27382,N_19131,N_17471);
or U27383 (N_27383,N_11104,N_10457);
or U27384 (N_27384,N_15853,N_14887);
or U27385 (N_27385,N_11524,N_13806);
nor U27386 (N_27386,N_10723,N_11072);
nor U27387 (N_27387,N_18461,N_12704);
and U27388 (N_27388,N_15552,N_19877);
and U27389 (N_27389,N_14089,N_10079);
nor U27390 (N_27390,N_17973,N_14467);
and U27391 (N_27391,N_14441,N_18283);
nor U27392 (N_27392,N_16862,N_14201);
and U27393 (N_27393,N_13129,N_16344);
or U27394 (N_27394,N_12511,N_12760);
nand U27395 (N_27395,N_12096,N_15512);
nand U27396 (N_27396,N_15337,N_19938);
nor U27397 (N_27397,N_17871,N_11166);
xnor U27398 (N_27398,N_12131,N_16224);
nor U27399 (N_27399,N_10829,N_13771);
and U27400 (N_27400,N_16450,N_10718);
nor U27401 (N_27401,N_16056,N_15021);
and U27402 (N_27402,N_16468,N_12956);
and U27403 (N_27403,N_13299,N_16595);
nand U27404 (N_27404,N_11184,N_13630);
nand U27405 (N_27405,N_10035,N_12801);
and U27406 (N_27406,N_17646,N_11540);
nor U27407 (N_27407,N_19757,N_13424);
nor U27408 (N_27408,N_18902,N_12448);
nor U27409 (N_27409,N_14244,N_17359);
and U27410 (N_27410,N_14522,N_12198);
nor U27411 (N_27411,N_19800,N_10836);
or U27412 (N_27412,N_15950,N_15655);
nor U27413 (N_27413,N_15187,N_19845);
nor U27414 (N_27414,N_11095,N_16175);
and U27415 (N_27415,N_13808,N_15707);
and U27416 (N_27416,N_14638,N_13969);
nand U27417 (N_27417,N_14676,N_10303);
nor U27418 (N_27418,N_10553,N_15029);
and U27419 (N_27419,N_15192,N_16527);
and U27420 (N_27420,N_11690,N_18928);
nand U27421 (N_27421,N_11415,N_11144);
or U27422 (N_27422,N_16872,N_12117);
nor U27423 (N_27423,N_18111,N_14116);
or U27424 (N_27424,N_18188,N_14322);
nor U27425 (N_27425,N_16682,N_10248);
nand U27426 (N_27426,N_11434,N_14994);
and U27427 (N_27427,N_13121,N_14310);
nor U27428 (N_27428,N_19118,N_19972);
or U27429 (N_27429,N_15617,N_10110);
and U27430 (N_27430,N_17466,N_17834);
and U27431 (N_27431,N_16919,N_13326);
nor U27432 (N_27432,N_17374,N_19349);
and U27433 (N_27433,N_14609,N_14126);
or U27434 (N_27434,N_11728,N_19253);
nor U27435 (N_27435,N_10867,N_19833);
and U27436 (N_27436,N_17022,N_16396);
or U27437 (N_27437,N_12962,N_16734);
nor U27438 (N_27438,N_12570,N_15490);
or U27439 (N_27439,N_19972,N_19753);
nand U27440 (N_27440,N_14393,N_17547);
nor U27441 (N_27441,N_14456,N_14920);
xnor U27442 (N_27442,N_19910,N_15813);
nand U27443 (N_27443,N_16982,N_12331);
and U27444 (N_27444,N_16475,N_12129);
nand U27445 (N_27445,N_13527,N_19703);
nor U27446 (N_27446,N_11390,N_19507);
and U27447 (N_27447,N_19465,N_19209);
nand U27448 (N_27448,N_12771,N_11168);
xor U27449 (N_27449,N_19231,N_10391);
nor U27450 (N_27450,N_13102,N_19303);
or U27451 (N_27451,N_12804,N_11253);
nand U27452 (N_27452,N_18638,N_16383);
xnor U27453 (N_27453,N_19720,N_17490);
and U27454 (N_27454,N_10076,N_19631);
and U27455 (N_27455,N_10885,N_11793);
and U27456 (N_27456,N_16682,N_14501);
and U27457 (N_27457,N_17409,N_17460);
nand U27458 (N_27458,N_16005,N_18933);
nor U27459 (N_27459,N_16217,N_10306);
and U27460 (N_27460,N_12596,N_12915);
nand U27461 (N_27461,N_14711,N_19261);
or U27462 (N_27462,N_18367,N_15673);
and U27463 (N_27463,N_15671,N_14471);
nand U27464 (N_27464,N_18327,N_18740);
nand U27465 (N_27465,N_15760,N_10522);
nand U27466 (N_27466,N_12697,N_19153);
or U27467 (N_27467,N_11146,N_15332);
nor U27468 (N_27468,N_16898,N_10022);
nor U27469 (N_27469,N_14541,N_13050);
nor U27470 (N_27470,N_19746,N_14684);
nor U27471 (N_27471,N_18042,N_16305);
nor U27472 (N_27472,N_10772,N_12388);
or U27473 (N_27473,N_19303,N_11640);
and U27474 (N_27474,N_15624,N_14598);
nor U27475 (N_27475,N_18018,N_16818);
and U27476 (N_27476,N_10580,N_17831);
nand U27477 (N_27477,N_11822,N_17735);
nor U27478 (N_27478,N_12524,N_11892);
nor U27479 (N_27479,N_15739,N_16538);
nor U27480 (N_27480,N_11149,N_15476);
and U27481 (N_27481,N_16126,N_15793);
or U27482 (N_27482,N_12934,N_13137);
or U27483 (N_27483,N_11759,N_12132);
or U27484 (N_27484,N_14274,N_11654);
nand U27485 (N_27485,N_10985,N_16582);
xor U27486 (N_27486,N_12614,N_11152);
and U27487 (N_27487,N_13511,N_12823);
nand U27488 (N_27488,N_16031,N_11486);
nor U27489 (N_27489,N_15093,N_13456);
nand U27490 (N_27490,N_14970,N_17594);
nor U27491 (N_27491,N_13156,N_17794);
xnor U27492 (N_27492,N_12363,N_16478);
and U27493 (N_27493,N_16953,N_15349);
or U27494 (N_27494,N_10971,N_12786);
nor U27495 (N_27495,N_12127,N_13864);
nor U27496 (N_27496,N_14731,N_13663);
and U27497 (N_27497,N_12380,N_19968);
or U27498 (N_27498,N_11332,N_15711);
nand U27499 (N_27499,N_16909,N_17932);
or U27500 (N_27500,N_19748,N_14786);
xor U27501 (N_27501,N_12536,N_11334);
xor U27502 (N_27502,N_15640,N_17499);
nor U27503 (N_27503,N_16523,N_14234);
or U27504 (N_27504,N_18336,N_19931);
or U27505 (N_27505,N_14190,N_11420);
nor U27506 (N_27506,N_17962,N_16232);
and U27507 (N_27507,N_15397,N_10606);
nor U27508 (N_27508,N_14902,N_14310);
nor U27509 (N_27509,N_11290,N_16492);
nand U27510 (N_27510,N_14879,N_12051);
xnor U27511 (N_27511,N_19147,N_15217);
and U27512 (N_27512,N_17141,N_14435);
nand U27513 (N_27513,N_19526,N_12897);
nand U27514 (N_27514,N_15095,N_12227);
xor U27515 (N_27515,N_18526,N_16658);
or U27516 (N_27516,N_17186,N_12423);
or U27517 (N_27517,N_13342,N_12355);
nor U27518 (N_27518,N_19747,N_19770);
or U27519 (N_27519,N_10741,N_18934);
nor U27520 (N_27520,N_13528,N_13171);
nor U27521 (N_27521,N_16636,N_12965);
and U27522 (N_27522,N_15819,N_11917);
nor U27523 (N_27523,N_10812,N_14604);
and U27524 (N_27524,N_13946,N_15014);
nand U27525 (N_27525,N_18467,N_18672);
or U27526 (N_27526,N_15222,N_14210);
or U27527 (N_27527,N_17794,N_11122);
nor U27528 (N_27528,N_16538,N_19478);
and U27529 (N_27529,N_17219,N_17404);
nand U27530 (N_27530,N_17964,N_18492);
or U27531 (N_27531,N_17138,N_14279);
and U27532 (N_27532,N_16804,N_18948);
or U27533 (N_27533,N_14597,N_19096);
xnor U27534 (N_27534,N_17108,N_15321);
nand U27535 (N_27535,N_13762,N_15582);
nand U27536 (N_27536,N_18037,N_12788);
nor U27537 (N_27537,N_17464,N_17968);
xor U27538 (N_27538,N_15635,N_17049);
or U27539 (N_27539,N_14529,N_10231);
and U27540 (N_27540,N_16739,N_14330);
and U27541 (N_27541,N_12079,N_15754);
nand U27542 (N_27542,N_15540,N_13366);
or U27543 (N_27543,N_11680,N_15574);
and U27544 (N_27544,N_17581,N_18860);
nand U27545 (N_27545,N_19813,N_15175);
or U27546 (N_27546,N_10205,N_18040);
or U27547 (N_27547,N_18920,N_18150);
or U27548 (N_27548,N_14430,N_13376);
nand U27549 (N_27549,N_18679,N_17843);
xor U27550 (N_27550,N_12758,N_16829);
nor U27551 (N_27551,N_17164,N_10051);
nor U27552 (N_27552,N_13324,N_14486);
or U27553 (N_27553,N_13749,N_15231);
and U27554 (N_27554,N_13646,N_14479);
nand U27555 (N_27555,N_15027,N_10949);
nand U27556 (N_27556,N_14680,N_18433);
nor U27557 (N_27557,N_16305,N_11526);
or U27558 (N_27558,N_12099,N_11620);
or U27559 (N_27559,N_13189,N_12403);
xor U27560 (N_27560,N_12474,N_18212);
and U27561 (N_27561,N_11608,N_12278);
or U27562 (N_27562,N_12018,N_15917);
nor U27563 (N_27563,N_14550,N_10535);
nor U27564 (N_27564,N_17481,N_16797);
or U27565 (N_27565,N_11790,N_12449);
xnor U27566 (N_27566,N_10104,N_12924);
nand U27567 (N_27567,N_16467,N_13789);
and U27568 (N_27568,N_19517,N_11481);
nand U27569 (N_27569,N_10547,N_19627);
or U27570 (N_27570,N_12601,N_10291);
nor U27571 (N_27571,N_19453,N_16125);
or U27572 (N_27572,N_15418,N_18869);
and U27573 (N_27573,N_12571,N_11107);
and U27574 (N_27574,N_19929,N_12874);
or U27575 (N_27575,N_16774,N_12833);
and U27576 (N_27576,N_11035,N_19308);
and U27577 (N_27577,N_10064,N_13952);
and U27578 (N_27578,N_16325,N_14971);
or U27579 (N_27579,N_16818,N_10507);
nor U27580 (N_27580,N_17099,N_17193);
nor U27581 (N_27581,N_18167,N_14603);
or U27582 (N_27582,N_12427,N_11023);
and U27583 (N_27583,N_10887,N_13477);
nand U27584 (N_27584,N_18880,N_19920);
nor U27585 (N_27585,N_13725,N_17053);
or U27586 (N_27586,N_19777,N_10871);
nand U27587 (N_27587,N_15715,N_15402);
or U27588 (N_27588,N_11554,N_19142);
nor U27589 (N_27589,N_12722,N_15152);
nor U27590 (N_27590,N_14059,N_13440);
nand U27591 (N_27591,N_16978,N_10284);
xnor U27592 (N_27592,N_17906,N_15243);
nand U27593 (N_27593,N_16237,N_17196);
or U27594 (N_27594,N_16800,N_17209);
nand U27595 (N_27595,N_18187,N_11221);
nand U27596 (N_27596,N_15342,N_12775);
xor U27597 (N_27597,N_11994,N_13514);
xnor U27598 (N_27598,N_10299,N_13570);
nor U27599 (N_27599,N_18246,N_15847);
xnor U27600 (N_27600,N_14938,N_10917);
and U27601 (N_27601,N_12407,N_17228);
nand U27602 (N_27602,N_19190,N_10827);
or U27603 (N_27603,N_16184,N_16358);
nor U27604 (N_27604,N_14671,N_19402);
or U27605 (N_27605,N_13548,N_19310);
and U27606 (N_27606,N_18662,N_12000);
and U27607 (N_27607,N_12337,N_12670);
nor U27608 (N_27608,N_14196,N_15695);
and U27609 (N_27609,N_17482,N_16770);
nor U27610 (N_27610,N_10074,N_13858);
and U27611 (N_27611,N_13657,N_17100);
and U27612 (N_27612,N_19987,N_19637);
or U27613 (N_27613,N_17294,N_19715);
nor U27614 (N_27614,N_13820,N_13827);
and U27615 (N_27615,N_16130,N_17447);
and U27616 (N_27616,N_12095,N_10777);
or U27617 (N_27617,N_15115,N_15624);
or U27618 (N_27618,N_17253,N_18454);
nor U27619 (N_27619,N_11068,N_19644);
xnor U27620 (N_27620,N_12236,N_12958);
nor U27621 (N_27621,N_19535,N_13573);
xor U27622 (N_27622,N_10326,N_16760);
or U27623 (N_27623,N_13005,N_16973);
nand U27624 (N_27624,N_17416,N_14925);
or U27625 (N_27625,N_14442,N_17006);
nor U27626 (N_27626,N_18195,N_19691);
or U27627 (N_27627,N_18946,N_11654);
nand U27628 (N_27628,N_10149,N_11931);
nor U27629 (N_27629,N_16415,N_18563);
nand U27630 (N_27630,N_18195,N_15834);
nor U27631 (N_27631,N_10101,N_16407);
xor U27632 (N_27632,N_16091,N_10213);
or U27633 (N_27633,N_14699,N_17833);
and U27634 (N_27634,N_18962,N_10723);
nor U27635 (N_27635,N_11828,N_12793);
or U27636 (N_27636,N_14389,N_17813);
and U27637 (N_27637,N_17543,N_11597);
nor U27638 (N_27638,N_11329,N_11067);
or U27639 (N_27639,N_13776,N_10487);
nor U27640 (N_27640,N_14811,N_13042);
and U27641 (N_27641,N_15629,N_18618);
and U27642 (N_27642,N_15534,N_19972);
and U27643 (N_27643,N_14565,N_19918);
or U27644 (N_27644,N_12058,N_12396);
and U27645 (N_27645,N_19010,N_11566);
nor U27646 (N_27646,N_17377,N_12781);
nor U27647 (N_27647,N_11401,N_16412);
nand U27648 (N_27648,N_13242,N_16904);
nor U27649 (N_27649,N_12144,N_18476);
nor U27650 (N_27650,N_13995,N_17625);
nand U27651 (N_27651,N_17471,N_15966);
or U27652 (N_27652,N_12815,N_10511);
and U27653 (N_27653,N_10027,N_11181);
and U27654 (N_27654,N_15530,N_16842);
nand U27655 (N_27655,N_12048,N_16008);
nand U27656 (N_27656,N_12117,N_11560);
nand U27657 (N_27657,N_14809,N_10855);
or U27658 (N_27658,N_18139,N_17961);
nand U27659 (N_27659,N_17449,N_16775);
nor U27660 (N_27660,N_17030,N_17771);
and U27661 (N_27661,N_17731,N_19635);
or U27662 (N_27662,N_12405,N_19026);
and U27663 (N_27663,N_19883,N_10254);
nor U27664 (N_27664,N_16160,N_12144);
nand U27665 (N_27665,N_11638,N_19024);
and U27666 (N_27666,N_11753,N_17018);
or U27667 (N_27667,N_15087,N_18872);
or U27668 (N_27668,N_15711,N_10325);
nand U27669 (N_27669,N_11719,N_10804);
nor U27670 (N_27670,N_17029,N_12276);
or U27671 (N_27671,N_16739,N_17746);
or U27672 (N_27672,N_17081,N_12751);
nor U27673 (N_27673,N_11704,N_11773);
or U27674 (N_27674,N_12296,N_18181);
nand U27675 (N_27675,N_15326,N_16725);
nand U27676 (N_27676,N_13294,N_13340);
nor U27677 (N_27677,N_10919,N_14130);
and U27678 (N_27678,N_10302,N_11198);
or U27679 (N_27679,N_18895,N_12030);
nand U27680 (N_27680,N_12956,N_14662);
xor U27681 (N_27681,N_13182,N_13464);
nor U27682 (N_27682,N_12532,N_14900);
or U27683 (N_27683,N_12435,N_11171);
or U27684 (N_27684,N_12444,N_19956);
nor U27685 (N_27685,N_14289,N_13447);
nand U27686 (N_27686,N_10275,N_14540);
nand U27687 (N_27687,N_18037,N_15901);
or U27688 (N_27688,N_11284,N_14104);
or U27689 (N_27689,N_17514,N_19104);
and U27690 (N_27690,N_14856,N_13095);
nand U27691 (N_27691,N_13465,N_19594);
nand U27692 (N_27692,N_13880,N_17559);
and U27693 (N_27693,N_19611,N_13611);
and U27694 (N_27694,N_15156,N_10902);
nor U27695 (N_27695,N_10913,N_16200);
nor U27696 (N_27696,N_18717,N_18411);
or U27697 (N_27697,N_15785,N_12417);
and U27698 (N_27698,N_17431,N_12022);
and U27699 (N_27699,N_11518,N_16349);
or U27700 (N_27700,N_15126,N_17288);
and U27701 (N_27701,N_17937,N_12044);
nand U27702 (N_27702,N_13647,N_15232);
nand U27703 (N_27703,N_11762,N_10588);
or U27704 (N_27704,N_14042,N_12361);
and U27705 (N_27705,N_15497,N_14902);
and U27706 (N_27706,N_10637,N_17024);
nand U27707 (N_27707,N_12723,N_11820);
and U27708 (N_27708,N_11921,N_15851);
nor U27709 (N_27709,N_11336,N_14387);
nand U27710 (N_27710,N_14147,N_12460);
and U27711 (N_27711,N_16442,N_16048);
or U27712 (N_27712,N_14961,N_13184);
xnor U27713 (N_27713,N_10153,N_11315);
xnor U27714 (N_27714,N_14978,N_14367);
nor U27715 (N_27715,N_18337,N_18220);
or U27716 (N_27716,N_10088,N_11186);
nand U27717 (N_27717,N_13531,N_12245);
nor U27718 (N_27718,N_12189,N_19031);
nor U27719 (N_27719,N_10858,N_16865);
xor U27720 (N_27720,N_12609,N_10770);
nor U27721 (N_27721,N_12435,N_17465);
nand U27722 (N_27722,N_18903,N_16826);
or U27723 (N_27723,N_13901,N_13213);
and U27724 (N_27724,N_12441,N_11352);
and U27725 (N_27725,N_12516,N_16465);
nor U27726 (N_27726,N_13077,N_10877);
nor U27727 (N_27727,N_11375,N_13949);
and U27728 (N_27728,N_14446,N_10047);
nand U27729 (N_27729,N_12262,N_13766);
nor U27730 (N_27730,N_13285,N_12322);
and U27731 (N_27731,N_19826,N_17395);
and U27732 (N_27732,N_18368,N_15071);
or U27733 (N_27733,N_16207,N_15746);
or U27734 (N_27734,N_15859,N_17306);
or U27735 (N_27735,N_12989,N_14825);
and U27736 (N_27736,N_15066,N_16152);
or U27737 (N_27737,N_13623,N_15791);
or U27738 (N_27738,N_10523,N_13714);
xor U27739 (N_27739,N_10859,N_10646);
or U27740 (N_27740,N_10613,N_18993);
xor U27741 (N_27741,N_16916,N_18518);
and U27742 (N_27742,N_10852,N_10256);
and U27743 (N_27743,N_15499,N_11207);
or U27744 (N_27744,N_19502,N_17445);
xor U27745 (N_27745,N_15922,N_10829);
nand U27746 (N_27746,N_17731,N_16415);
and U27747 (N_27747,N_14187,N_14182);
and U27748 (N_27748,N_19573,N_19399);
and U27749 (N_27749,N_19216,N_11427);
and U27750 (N_27750,N_14734,N_11141);
nor U27751 (N_27751,N_14068,N_13879);
nor U27752 (N_27752,N_10993,N_14455);
nand U27753 (N_27753,N_10083,N_14018);
nand U27754 (N_27754,N_10310,N_18674);
and U27755 (N_27755,N_10128,N_11536);
xor U27756 (N_27756,N_13873,N_14092);
nor U27757 (N_27757,N_12081,N_15224);
and U27758 (N_27758,N_18575,N_14946);
nand U27759 (N_27759,N_17370,N_15091);
and U27760 (N_27760,N_19618,N_12093);
or U27761 (N_27761,N_16463,N_10569);
nand U27762 (N_27762,N_19248,N_13676);
nand U27763 (N_27763,N_16213,N_15606);
nand U27764 (N_27764,N_12666,N_16235);
nor U27765 (N_27765,N_10233,N_19044);
nor U27766 (N_27766,N_15397,N_13708);
nor U27767 (N_27767,N_16306,N_17035);
xor U27768 (N_27768,N_17519,N_11247);
nor U27769 (N_27769,N_12024,N_14840);
xnor U27770 (N_27770,N_17668,N_12592);
nor U27771 (N_27771,N_12749,N_10841);
or U27772 (N_27772,N_15557,N_19212);
or U27773 (N_27773,N_19787,N_16187);
and U27774 (N_27774,N_14139,N_16063);
xor U27775 (N_27775,N_15703,N_12612);
or U27776 (N_27776,N_17566,N_16186);
xor U27777 (N_27777,N_15597,N_14655);
nand U27778 (N_27778,N_12803,N_17776);
nor U27779 (N_27779,N_13145,N_17569);
nand U27780 (N_27780,N_18093,N_14009);
or U27781 (N_27781,N_18806,N_14786);
nand U27782 (N_27782,N_10048,N_18706);
nor U27783 (N_27783,N_12082,N_12530);
or U27784 (N_27784,N_15759,N_16798);
nor U27785 (N_27785,N_18569,N_19305);
nor U27786 (N_27786,N_12337,N_13876);
or U27787 (N_27787,N_14738,N_12879);
xnor U27788 (N_27788,N_17418,N_12308);
or U27789 (N_27789,N_18252,N_14667);
nand U27790 (N_27790,N_12074,N_17278);
and U27791 (N_27791,N_14992,N_13110);
nor U27792 (N_27792,N_10844,N_14452);
nand U27793 (N_27793,N_15140,N_14336);
or U27794 (N_27794,N_16098,N_15589);
nor U27795 (N_27795,N_17396,N_11865);
nor U27796 (N_27796,N_16660,N_11348);
nand U27797 (N_27797,N_17739,N_19591);
or U27798 (N_27798,N_18042,N_17492);
nor U27799 (N_27799,N_16247,N_13981);
and U27800 (N_27800,N_14791,N_11039);
nand U27801 (N_27801,N_11647,N_11489);
and U27802 (N_27802,N_15515,N_18430);
nor U27803 (N_27803,N_15372,N_15706);
or U27804 (N_27804,N_15093,N_14167);
or U27805 (N_27805,N_16193,N_13370);
and U27806 (N_27806,N_17286,N_10560);
and U27807 (N_27807,N_12880,N_17215);
and U27808 (N_27808,N_11499,N_10741);
nand U27809 (N_27809,N_17560,N_19901);
nand U27810 (N_27810,N_12470,N_12982);
and U27811 (N_27811,N_12047,N_16682);
or U27812 (N_27812,N_17635,N_12344);
and U27813 (N_27813,N_17280,N_14802);
nor U27814 (N_27814,N_11961,N_19738);
and U27815 (N_27815,N_14695,N_10394);
nand U27816 (N_27816,N_18450,N_18032);
or U27817 (N_27817,N_13917,N_18547);
and U27818 (N_27818,N_16997,N_12802);
and U27819 (N_27819,N_12156,N_14876);
nor U27820 (N_27820,N_12214,N_12254);
nor U27821 (N_27821,N_19728,N_16096);
xor U27822 (N_27822,N_14743,N_12062);
nand U27823 (N_27823,N_19561,N_10137);
nor U27824 (N_27824,N_14916,N_11349);
nor U27825 (N_27825,N_13195,N_17538);
or U27826 (N_27826,N_18420,N_11344);
nor U27827 (N_27827,N_19611,N_12962);
nand U27828 (N_27828,N_13946,N_10187);
nand U27829 (N_27829,N_12662,N_17498);
and U27830 (N_27830,N_13746,N_15372);
nor U27831 (N_27831,N_17536,N_12502);
or U27832 (N_27832,N_12035,N_17819);
nand U27833 (N_27833,N_17322,N_18493);
or U27834 (N_27834,N_16659,N_19501);
nand U27835 (N_27835,N_17520,N_17343);
and U27836 (N_27836,N_11999,N_16864);
nor U27837 (N_27837,N_14112,N_11030);
nor U27838 (N_27838,N_11411,N_15184);
and U27839 (N_27839,N_10972,N_15669);
or U27840 (N_27840,N_17569,N_19831);
or U27841 (N_27841,N_13186,N_10622);
nand U27842 (N_27842,N_13213,N_12894);
nand U27843 (N_27843,N_19490,N_13596);
or U27844 (N_27844,N_13614,N_14716);
and U27845 (N_27845,N_14311,N_15515);
nor U27846 (N_27846,N_10648,N_19462);
and U27847 (N_27847,N_15936,N_16214);
and U27848 (N_27848,N_16577,N_12188);
and U27849 (N_27849,N_14245,N_16276);
nand U27850 (N_27850,N_11754,N_15412);
and U27851 (N_27851,N_15319,N_14649);
or U27852 (N_27852,N_16318,N_15948);
and U27853 (N_27853,N_15021,N_13376);
nor U27854 (N_27854,N_10549,N_17106);
and U27855 (N_27855,N_16350,N_17258);
and U27856 (N_27856,N_16886,N_18904);
or U27857 (N_27857,N_16484,N_18643);
nor U27858 (N_27858,N_13410,N_19608);
and U27859 (N_27859,N_10476,N_12182);
nor U27860 (N_27860,N_12452,N_10424);
nor U27861 (N_27861,N_14065,N_10444);
nor U27862 (N_27862,N_16826,N_19686);
nor U27863 (N_27863,N_13723,N_18345);
or U27864 (N_27864,N_18556,N_13225);
nand U27865 (N_27865,N_12857,N_19205);
and U27866 (N_27866,N_17271,N_10980);
nand U27867 (N_27867,N_18995,N_13143);
nand U27868 (N_27868,N_17784,N_15218);
and U27869 (N_27869,N_16063,N_12305);
nand U27870 (N_27870,N_11121,N_18942);
xnor U27871 (N_27871,N_16729,N_13620);
or U27872 (N_27872,N_15734,N_16108);
or U27873 (N_27873,N_19187,N_13083);
or U27874 (N_27874,N_12674,N_14552);
and U27875 (N_27875,N_17149,N_10595);
nand U27876 (N_27876,N_10209,N_13648);
nand U27877 (N_27877,N_15693,N_18389);
and U27878 (N_27878,N_11860,N_10039);
or U27879 (N_27879,N_10081,N_11270);
nand U27880 (N_27880,N_13028,N_15194);
nor U27881 (N_27881,N_10060,N_18898);
nand U27882 (N_27882,N_15077,N_17797);
or U27883 (N_27883,N_11894,N_12217);
and U27884 (N_27884,N_17239,N_15103);
or U27885 (N_27885,N_11943,N_18863);
or U27886 (N_27886,N_11624,N_19156);
and U27887 (N_27887,N_10111,N_15724);
nand U27888 (N_27888,N_10818,N_11204);
nor U27889 (N_27889,N_13314,N_16285);
and U27890 (N_27890,N_15063,N_18908);
nand U27891 (N_27891,N_12275,N_16308);
nand U27892 (N_27892,N_15743,N_12387);
or U27893 (N_27893,N_11704,N_18293);
and U27894 (N_27894,N_10536,N_18378);
nand U27895 (N_27895,N_12582,N_12744);
and U27896 (N_27896,N_15500,N_13800);
nand U27897 (N_27897,N_19103,N_18014);
or U27898 (N_27898,N_15857,N_19516);
nor U27899 (N_27899,N_14946,N_15248);
and U27900 (N_27900,N_15956,N_11341);
or U27901 (N_27901,N_10674,N_14585);
or U27902 (N_27902,N_15293,N_10324);
or U27903 (N_27903,N_16623,N_12222);
nor U27904 (N_27904,N_11934,N_11423);
nand U27905 (N_27905,N_16524,N_12200);
xor U27906 (N_27906,N_14826,N_11084);
nor U27907 (N_27907,N_19108,N_19847);
and U27908 (N_27908,N_15010,N_17748);
nand U27909 (N_27909,N_12596,N_19063);
nand U27910 (N_27910,N_16772,N_18259);
xor U27911 (N_27911,N_14518,N_18170);
nand U27912 (N_27912,N_14562,N_17286);
nor U27913 (N_27913,N_17441,N_13743);
nor U27914 (N_27914,N_14095,N_17078);
nor U27915 (N_27915,N_13525,N_13763);
nor U27916 (N_27916,N_10742,N_15571);
xnor U27917 (N_27917,N_18442,N_14591);
or U27918 (N_27918,N_14680,N_16058);
and U27919 (N_27919,N_10793,N_18390);
nor U27920 (N_27920,N_15477,N_11806);
nor U27921 (N_27921,N_18496,N_18867);
nand U27922 (N_27922,N_10183,N_15117);
and U27923 (N_27923,N_14996,N_18056);
nor U27924 (N_27924,N_15939,N_19956);
and U27925 (N_27925,N_15451,N_17086);
or U27926 (N_27926,N_17479,N_15993);
and U27927 (N_27927,N_11715,N_10259);
nor U27928 (N_27928,N_18446,N_13007);
xnor U27929 (N_27929,N_15636,N_17582);
nor U27930 (N_27930,N_11187,N_17982);
nor U27931 (N_27931,N_14359,N_18468);
nor U27932 (N_27932,N_15071,N_16741);
nor U27933 (N_27933,N_17657,N_18074);
nand U27934 (N_27934,N_18745,N_18507);
and U27935 (N_27935,N_13304,N_11424);
nand U27936 (N_27936,N_18196,N_15469);
nor U27937 (N_27937,N_16066,N_14464);
and U27938 (N_27938,N_12231,N_13277);
nor U27939 (N_27939,N_19759,N_12180);
nand U27940 (N_27940,N_16536,N_13693);
nand U27941 (N_27941,N_13552,N_14609);
nor U27942 (N_27942,N_14187,N_10211);
nor U27943 (N_27943,N_12122,N_16675);
xnor U27944 (N_27944,N_19494,N_16526);
or U27945 (N_27945,N_15477,N_19575);
and U27946 (N_27946,N_15916,N_17011);
nor U27947 (N_27947,N_13232,N_11681);
and U27948 (N_27948,N_18731,N_18789);
and U27949 (N_27949,N_15959,N_13232);
and U27950 (N_27950,N_13103,N_10671);
nand U27951 (N_27951,N_14441,N_13347);
and U27952 (N_27952,N_16607,N_18623);
or U27953 (N_27953,N_11053,N_19348);
and U27954 (N_27954,N_14551,N_19054);
nand U27955 (N_27955,N_16312,N_11172);
and U27956 (N_27956,N_17122,N_14645);
nor U27957 (N_27957,N_18797,N_12450);
nor U27958 (N_27958,N_19561,N_13280);
nand U27959 (N_27959,N_12728,N_14785);
xnor U27960 (N_27960,N_19057,N_11265);
and U27961 (N_27961,N_11804,N_11501);
and U27962 (N_27962,N_17900,N_13599);
or U27963 (N_27963,N_16982,N_18003);
nand U27964 (N_27964,N_14691,N_18697);
nor U27965 (N_27965,N_16018,N_10590);
or U27966 (N_27966,N_17254,N_10741);
nand U27967 (N_27967,N_16877,N_19354);
or U27968 (N_27968,N_10586,N_14267);
or U27969 (N_27969,N_11081,N_10512);
xor U27970 (N_27970,N_15512,N_19425);
or U27971 (N_27971,N_11422,N_10736);
or U27972 (N_27972,N_16259,N_12671);
or U27973 (N_27973,N_15289,N_19749);
or U27974 (N_27974,N_18062,N_12944);
nand U27975 (N_27975,N_19130,N_15288);
or U27976 (N_27976,N_14944,N_18823);
and U27977 (N_27977,N_19514,N_19188);
or U27978 (N_27978,N_17962,N_11119);
nand U27979 (N_27979,N_16484,N_18431);
or U27980 (N_27980,N_10068,N_16744);
nor U27981 (N_27981,N_19733,N_12350);
xor U27982 (N_27982,N_16047,N_12963);
nor U27983 (N_27983,N_15377,N_19746);
xnor U27984 (N_27984,N_10021,N_18577);
nor U27985 (N_27985,N_16395,N_16846);
nor U27986 (N_27986,N_12814,N_12521);
or U27987 (N_27987,N_11679,N_15155);
nor U27988 (N_27988,N_10094,N_12666);
or U27989 (N_27989,N_16535,N_11808);
and U27990 (N_27990,N_15842,N_10102);
nand U27991 (N_27991,N_14582,N_14967);
nor U27992 (N_27992,N_16395,N_18154);
nor U27993 (N_27993,N_11121,N_19467);
nor U27994 (N_27994,N_17229,N_15377);
nor U27995 (N_27995,N_13518,N_15595);
nor U27996 (N_27996,N_13536,N_19872);
nand U27997 (N_27997,N_17655,N_15984);
and U27998 (N_27998,N_14073,N_10364);
or U27999 (N_27999,N_13869,N_18884);
or U28000 (N_28000,N_14369,N_13659);
and U28001 (N_28001,N_10867,N_11034);
nand U28002 (N_28002,N_13882,N_12055);
nand U28003 (N_28003,N_12189,N_19061);
or U28004 (N_28004,N_13755,N_18713);
nor U28005 (N_28005,N_18726,N_13320);
nor U28006 (N_28006,N_10404,N_13245);
or U28007 (N_28007,N_18701,N_16894);
and U28008 (N_28008,N_18532,N_11061);
and U28009 (N_28009,N_18836,N_16050);
nor U28010 (N_28010,N_16962,N_13428);
and U28011 (N_28011,N_12822,N_18236);
nand U28012 (N_28012,N_19411,N_16682);
nor U28013 (N_28013,N_13032,N_18156);
nor U28014 (N_28014,N_18779,N_16719);
nor U28015 (N_28015,N_16299,N_18318);
xor U28016 (N_28016,N_16693,N_18615);
nor U28017 (N_28017,N_12760,N_11244);
and U28018 (N_28018,N_17946,N_11931);
nor U28019 (N_28019,N_17442,N_17851);
nand U28020 (N_28020,N_17384,N_19960);
and U28021 (N_28021,N_10947,N_14205);
xor U28022 (N_28022,N_18123,N_15693);
or U28023 (N_28023,N_15629,N_12922);
nand U28024 (N_28024,N_15229,N_19385);
or U28025 (N_28025,N_18183,N_14075);
or U28026 (N_28026,N_11687,N_14840);
xor U28027 (N_28027,N_14548,N_18603);
nand U28028 (N_28028,N_13377,N_10396);
or U28029 (N_28029,N_11514,N_13478);
or U28030 (N_28030,N_19557,N_15437);
and U28031 (N_28031,N_11552,N_16370);
nand U28032 (N_28032,N_10771,N_10954);
xor U28033 (N_28033,N_16879,N_19302);
nor U28034 (N_28034,N_11081,N_11432);
and U28035 (N_28035,N_16239,N_10592);
nor U28036 (N_28036,N_12807,N_18886);
nor U28037 (N_28037,N_10222,N_18949);
xnor U28038 (N_28038,N_13197,N_11915);
and U28039 (N_28039,N_12413,N_18673);
nand U28040 (N_28040,N_17006,N_11461);
nand U28041 (N_28041,N_19717,N_13539);
nor U28042 (N_28042,N_15522,N_18143);
or U28043 (N_28043,N_18839,N_16695);
nand U28044 (N_28044,N_15732,N_13820);
and U28045 (N_28045,N_12848,N_10528);
and U28046 (N_28046,N_13905,N_18808);
or U28047 (N_28047,N_17814,N_13635);
nand U28048 (N_28048,N_10075,N_15769);
or U28049 (N_28049,N_15495,N_15262);
nor U28050 (N_28050,N_14554,N_15644);
nor U28051 (N_28051,N_18330,N_10007);
and U28052 (N_28052,N_14501,N_16724);
or U28053 (N_28053,N_10140,N_15593);
and U28054 (N_28054,N_14471,N_12840);
or U28055 (N_28055,N_13311,N_17103);
xnor U28056 (N_28056,N_11996,N_16307);
nor U28057 (N_28057,N_11986,N_13672);
or U28058 (N_28058,N_16742,N_14263);
nand U28059 (N_28059,N_13206,N_19533);
nor U28060 (N_28060,N_12017,N_13944);
or U28061 (N_28061,N_17270,N_10024);
nand U28062 (N_28062,N_14354,N_15172);
and U28063 (N_28063,N_13763,N_17352);
nor U28064 (N_28064,N_19351,N_16076);
or U28065 (N_28065,N_10001,N_11541);
nand U28066 (N_28066,N_15601,N_19077);
nand U28067 (N_28067,N_15268,N_11546);
xnor U28068 (N_28068,N_19013,N_18390);
nand U28069 (N_28069,N_11217,N_10455);
nand U28070 (N_28070,N_19302,N_14719);
nand U28071 (N_28071,N_10073,N_10706);
and U28072 (N_28072,N_15881,N_18360);
or U28073 (N_28073,N_16365,N_16105);
nand U28074 (N_28074,N_11466,N_10869);
xnor U28075 (N_28075,N_18169,N_13363);
xor U28076 (N_28076,N_19962,N_19173);
and U28077 (N_28077,N_19770,N_14600);
and U28078 (N_28078,N_13870,N_14865);
xor U28079 (N_28079,N_16583,N_19242);
nor U28080 (N_28080,N_11360,N_15019);
nor U28081 (N_28081,N_16652,N_19560);
nor U28082 (N_28082,N_11082,N_14596);
and U28083 (N_28083,N_18883,N_10705);
nand U28084 (N_28084,N_15800,N_16157);
nor U28085 (N_28085,N_19476,N_15600);
nor U28086 (N_28086,N_10108,N_10039);
or U28087 (N_28087,N_19309,N_18782);
and U28088 (N_28088,N_14918,N_11947);
or U28089 (N_28089,N_17548,N_15457);
xor U28090 (N_28090,N_16015,N_16521);
nand U28091 (N_28091,N_16703,N_14182);
and U28092 (N_28092,N_16239,N_19455);
nand U28093 (N_28093,N_18244,N_17910);
nor U28094 (N_28094,N_16883,N_17624);
nand U28095 (N_28095,N_18618,N_11285);
or U28096 (N_28096,N_10220,N_10808);
and U28097 (N_28097,N_12158,N_12896);
or U28098 (N_28098,N_17015,N_19705);
xnor U28099 (N_28099,N_16709,N_10560);
nand U28100 (N_28100,N_14550,N_16168);
and U28101 (N_28101,N_13676,N_15009);
nor U28102 (N_28102,N_17857,N_19701);
nand U28103 (N_28103,N_17742,N_16414);
nand U28104 (N_28104,N_10934,N_17562);
xor U28105 (N_28105,N_19183,N_17203);
or U28106 (N_28106,N_15120,N_18339);
or U28107 (N_28107,N_14614,N_12659);
xnor U28108 (N_28108,N_14373,N_11496);
nand U28109 (N_28109,N_16230,N_11636);
or U28110 (N_28110,N_18797,N_12575);
and U28111 (N_28111,N_11513,N_19090);
or U28112 (N_28112,N_16446,N_15023);
xnor U28113 (N_28113,N_15583,N_13878);
nor U28114 (N_28114,N_12004,N_12659);
or U28115 (N_28115,N_11209,N_18045);
nand U28116 (N_28116,N_15732,N_19427);
nand U28117 (N_28117,N_17073,N_11637);
nand U28118 (N_28118,N_15208,N_15237);
and U28119 (N_28119,N_18318,N_16352);
nand U28120 (N_28120,N_16561,N_12097);
or U28121 (N_28121,N_14909,N_16388);
xnor U28122 (N_28122,N_14042,N_17065);
or U28123 (N_28123,N_13099,N_16394);
nand U28124 (N_28124,N_14756,N_13900);
and U28125 (N_28125,N_14650,N_12507);
and U28126 (N_28126,N_17877,N_11827);
or U28127 (N_28127,N_14639,N_12946);
nor U28128 (N_28128,N_10362,N_15440);
nor U28129 (N_28129,N_17000,N_12433);
nand U28130 (N_28130,N_14088,N_12275);
or U28131 (N_28131,N_17080,N_19373);
and U28132 (N_28132,N_18774,N_11674);
xnor U28133 (N_28133,N_17561,N_16213);
nand U28134 (N_28134,N_10158,N_10409);
nand U28135 (N_28135,N_10556,N_10549);
and U28136 (N_28136,N_10366,N_17305);
nor U28137 (N_28137,N_10463,N_11949);
and U28138 (N_28138,N_15552,N_15468);
nand U28139 (N_28139,N_15955,N_16970);
nand U28140 (N_28140,N_11409,N_17956);
or U28141 (N_28141,N_13554,N_11866);
or U28142 (N_28142,N_19289,N_10273);
xor U28143 (N_28143,N_16153,N_12709);
xnor U28144 (N_28144,N_12826,N_11683);
or U28145 (N_28145,N_12951,N_10760);
and U28146 (N_28146,N_16694,N_15081);
nand U28147 (N_28147,N_19143,N_12103);
and U28148 (N_28148,N_14229,N_18551);
nor U28149 (N_28149,N_17360,N_16789);
nor U28150 (N_28150,N_11532,N_14030);
or U28151 (N_28151,N_19643,N_11375);
nor U28152 (N_28152,N_18741,N_16706);
nand U28153 (N_28153,N_11281,N_15547);
nor U28154 (N_28154,N_16511,N_13112);
xor U28155 (N_28155,N_13471,N_12009);
or U28156 (N_28156,N_16137,N_10677);
nor U28157 (N_28157,N_15897,N_19019);
xor U28158 (N_28158,N_12805,N_19689);
and U28159 (N_28159,N_18531,N_12210);
nand U28160 (N_28160,N_10499,N_11276);
or U28161 (N_28161,N_15432,N_10136);
and U28162 (N_28162,N_15867,N_19465);
nand U28163 (N_28163,N_16795,N_17717);
nor U28164 (N_28164,N_16551,N_17362);
or U28165 (N_28165,N_12791,N_18969);
nor U28166 (N_28166,N_13879,N_15270);
nand U28167 (N_28167,N_15065,N_11106);
nor U28168 (N_28168,N_19577,N_19666);
nand U28169 (N_28169,N_18860,N_10454);
or U28170 (N_28170,N_16219,N_14204);
and U28171 (N_28171,N_19876,N_12748);
nor U28172 (N_28172,N_17577,N_16955);
nor U28173 (N_28173,N_18046,N_17305);
nand U28174 (N_28174,N_16228,N_12991);
or U28175 (N_28175,N_16914,N_16548);
nand U28176 (N_28176,N_15626,N_13090);
xor U28177 (N_28177,N_10764,N_16436);
nand U28178 (N_28178,N_17610,N_10592);
nor U28179 (N_28179,N_14042,N_17296);
and U28180 (N_28180,N_14710,N_19584);
and U28181 (N_28181,N_13007,N_18241);
or U28182 (N_28182,N_19258,N_17788);
and U28183 (N_28183,N_11325,N_12995);
and U28184 (N_28184,N_16059,N_17810);
nand U28185 (N_28185,N_16323,N_19354);
and U28186 (N_28186,N_18014,N_15251);
xnor U28187 (N_28187,N_15214,N_16489);
and U28188 (N_28188,N_18141,N_17798);
and U28189 (N_28189,N_11923,N_17756);
or U28190 (N_28190,N_19086,N_17750);
nand U28191 (N_28191,N_16322,N_18310);
and U28192 (N_28192,N_12232,N_10283);
or U28193 (N_28193,N_14995,N_11817);
nor U28194 (N_28194,N_19929,N_16451);
nand U28195 (N_28195,N_16869,N_16133);
nand U28196 (N_28196,N_12298,N_13019);
nor U28197 (N_28197,N_13902,N_17714);
nor U28198 (N_28198,N_18940,N_10702);
nand U28199 (N_28199,N_13485,N_11553);
nand U28200 (N_28200,N_12195,N_15840);
and U28201 (N_28201,N_15290,N_11951);
or U28202 (N_28202,N_14528,N_11904);
or U28203 (N_28203,N_15539,N_14128);
nor U28204 (N_28204,N_19445,N_16506);
or U28205 (N_28205,N_14368,N_19980);
xnor U28206 (N_28206,N_13546,N_18971);
nand U28207 (N_28207,N_17150,N_17403);
and U28208 (N_28208,N_18491,N_19794);
and U28209 (N_28209,N_17510,N_11186);
nor U28210 (N_28210,N_11223,N_11735);
and U28211 (N_28211,N_15184,N_10702);
xnor U28212 (N_28212,N_17810,N_17533);
and U28213 (N_28213,N_18492,N_16323);
nor U28214 (N_28214,N_13372,N_17694);
or U28215 (N_28215,N_12128,N_14320);
nand U28216 (N_28216,N_13609,N_11924);
and U28217 (N_28217,N_12336,N_11928);
or U28218 (N_28218,N_17398,N_19451);
xnor U28219 (N_28219,N_12056,N_12689);
nand U28220 (N_28220,N_15489,N_14355);
nand U28221 (N_28221,N_10893,N_14623);
nand U28222 (N_28222,N_13479,N_11156);
or U28223 (N_28223,N_12011,N_13601);
xnor U28224 (N_28224,N_18224,N_18578);
nor U28225 (N_28225,N_14872,N_11812);
nor U28226 (N_28226,N_17346,N_18180);
and U28227 (N_28227,N_13359,N_11474);
and U28228 (N_28228,N_16293,N_16184);
nand U28229 (N_28229,N_13487,N_17108);
nor U28230 (N_28230,N_11171,N_15310);
nand U28231 (N_28231,N_14423,N_13889);
or U28232 (N_28232,N_15919,N_13187);
nor U28233 (N_28233,N_19494,N_19643);
and U28234 (N_28234,N_17136,N_13301);
nand U28235 (N_28235,N_11451,N_15071);
nand U28236 (N_28236,N_19908,N_10473);
and U28237 (N_28237,N_11535,N_14900);
or U28238 (N_28238,N_11246,N_16744);
and U28239 (N_28239,N_17984,N_19657);
nand U28240 (N_28240,N_14341,N_13597);
and U28241 (N_28241,N_11006,N_19780);
nor U28242 (N_28242,N_16588,N_14247);
nand U28243 (N_28243,N_18825,N_10921);
and U28244 (N_28244,N_13637,N_16183);
nor U28245 (N_28245,N_11669,N_10076);
xnor U28246 (N_28246,N_17953,N_14958);
and U28247 (N_28247,N_18284,N_15587);
nand U28248 (N_28248,N_10275,N_16425);
nand U28249 (N_28249,N_12710,N_18542);
or U28250 (N_28250,N_18342,N_13578);
nor U28251 (N_28251,N_17335,N_18399);
xor U28252 (N_28252,N_16635,N_13650);
nand U28253 (N_28253,N_10427,N_10728);
nand U28254 (N_28254,N_14105,N_15816);
or U28255 (N_28255,N_18356,N_16333);
nand U28256 (N_28256,N_11331,N_14186);
or U28257 (N_28257,N_13632,N_17957);
and U28258 (N_28258,N_19063,N_15736);
nand U28259 (N_28259,N_18926,N_18704);
or U28260 (N_28260,N_11215,N_10855);
nor U28261 (N_28261,N_15305,N_14685);
and U28262 (N_28262,N_14451,N_19158);
nor U28263 (N_28263,N_16078,N_13941);
or U28264 (N_28264,N_17587,N_10135);
nor U28265 (N_28265,N_13184,N_10668);
and U28266 (N_28266,N_16230,N_14030);
and U28267 (N_28267,N_13401,N_14708);
nand U28268 (N_28268,N_11611,N_19917);
nand U28269 (N_28269,N_18578,N_12610);
nor U28270 (N_28270,N_13279,N_12738);
nor U28271 (N_28271,N_14986,N_17463);
xor U28272 (N_28272,N_18059,N_18292);
and U28273 (N_28273,N_19657,N_18959);
xnor U28274 (N_28274,N_18165,N_15529);
nand U28275 (N_28275,N_19954,N_13229);
xor U28276 (N_28276,N_14283,N_11905);
or U28277 (N_28277,N_18520,N_16013);
nand U28278 (N_28278,N_10059,N_18708);
or U28279 (N_28279,N_15181,N_15793);
nor U28280 (N_28280,N_19441,N_17599);
and U28281 (N_28281,N_14955,N_10405);
and U28282 (N_28282,N_19704,N_11009);
and U28283 (N_28283,N_16936,N_11967);
nand U28284 (N_28284,N_19584,N_19710);
nor U28285 (N_28285,N_16111,N_13008);
nor U28286 (N_28286,N_11904,N_10587);
nor U28287 (N_28287,N_13569,N_10439);
nand U28288 (N_28288,N_17679,N_14431);
xor U28289 (N_28289,N_14603,N_18136);
or U28290 (N_28290,N_18357,N_16304);
and U28291 (N_28291,N_12544,N_18767);
xor U28292 (N_28292,N_11377,N_19993);
nor U28293 (N_28293,N_17411,N_13825);
or U28294 (N_28294,N_10356,N_10559);
or U28295 (N_28295,N_17529,N_17876);
or U28296 (N_28296,N_12234,N_17963);
nand U28297 (N_28297,N_12948,N_10098);
and U28298 (N_28298,N_13303,N_11240);
xnor U28299 (N_28299,N_10540,N_19646);
and U28300 (N_28300,N_19939,N_17682);
nand U28301 (N_28301,N_17193,N_13252);
nor U28302 (N_28302,N_13276,N_11858);
and U28303 (N_28303,N_10968,N_18492);
nand U28304 (N_28304,N_16220,N_12862);
or U28305 (N_28305,N_11353,N_14567);
xor U28306 (N_28306,N_10312,N_13895);
or U28307 (N_28307,N_14751,N_18272);
xnor U28308 (N_28308,N_13511,N_15812);
nand U28309 (N_28309,N_15135,N_11560);
xnor U28310 (N_28310,N_11168,N_13787);
nor U28311 (N_28311,N_11507,N_18005);
nor U28312 (N_28312,N_11592,N_12656);
nor U28313 (N_28313,N_10246,N_16818);
and U28314 (N_28314,N_14078,N_18943);
and U28315 (N_28315,N_17274,N_16095);
xor U28316 (N_28316,N_11005,N_18736);
or U28317 (N_28317,N_17256,N_14109);
or U28318 (N_28318,N_13933,N_18228);
nor U28319 (N_28319,N_10907,N_14642);
or U28320 (N_28320,N_14100,N_10740);
or U28321 (N_28321,N_18092,N_10269);
and U28322 (N_28322,N_11649,N_18493);
nor U28323 (N_28323,N_19827,N_10446);
or U28324 (N_28324,N_15486,N_10581);
or U28325 (N_28325,N_10697,N_13907);
nand U28326 (N_28326,N_19610,N_14304);
xnor U28327 (N_28327,N_18934,N_12889);
and U28328 (N_28328,N_16099,N_16039);
nand U28329 (N_28329,N_18272,N_16123);
or U28330 (N_28330,N_16070,N_11356);
or U28331 (N_28331,N_14229,N_15439);
and U28332 (N_28332,N_19145,N_17794);
xor U28333 (N_28333,N_18219,N_13310);
and U28334 (N_28334,N_13842,N_17632);
and U28335 (N_28335,N_10737,N_19386);
or U28336 (N_28336,N_14791,N_10296);
and U28337 (N_28337,N_17447,N_18013);
and U28338 (N_28338,N_10008,N_19068);
nand U28339 (N_28339,N_17227,N_18429);
and U28340 (N_28340,N_11068,N_12958);
or U28341 (N_28341,N_19441,N_12898);
nand U28342 (N_28342,N_17473,N_10695);
and U28343 (N_28343,N_10806,N_15726);
and U28344 (N_28344,N_11563,N_18336);
nand U28345 (N_28345,N_14250,N_13371);
nor U28346 (N_28346,N_11460,N_11179);
and U28347 (N_28347,N_11787,N_18430);
and U28348 (N_28348,N_16302,N_16891);
or U28349 (N_28349,N_15549,N_13944);
nand U28350 (N_28350,N_19574,N_18254);
nor U28351 (N_28351,N_14605,N_12400);
or U28352 (N_28352,N_12430,N_10674);
nand U28353 (N_28353,N_18201,N_17452);
nand U28354 (N_28354,N_18976,N_17706);
nand U28355 (N_28355,N_18193,N_11802);
nand U28356 (N_28356,N_16680,N_13172);
and U28357 (N_28357,N_17797,N_13768);
nor U28358 (N_28358,N_15669,N_18184);
nor U28359 (N_28359,N_14357,N_15817);
nor U28360 (N_28360,N_17011,N_13633);
nor U28361 (N_28361,N_18447,N_13948);
and U28362 (N_28362,N_12231,N_12419);
nand U28363 (N_28363,N_14994,N_17302);
nor U28364 (N_28364,N_10105,N_18604);
nand U28365 (N_28365,N_10147,N_15524);
and U28366 (N_28366,N_12145,N_17560);
or U28367 (N_28367,N_18991,N_18038);
and U28368 (N_28368,N_17926,N_17330);
xnor U28369 (N_28369,N_11733,N_11260);
nor U28370 (N_28370,N_11604,N_15365);
and U28371 (N_28371,N_12842,N_17895);
nand U28372 (N_28372,N_13301,N_17763);
nand U28373 (N_28373,N_15458,N_16269);
and U28374 (N_28374,N_17997,N_19076);
and U28375 (N_28375,N_14034,N_12488);
or U28376 (N_28376,N_17109,N_16624);
nand U28377 (N_28377,N_15620,N_19176);
or U28378 (N_28378,N_13739,N_15885);
nor U28379 (N_28379,N_13600,N_16787);
nand U28380 (N_28380,N_13340,N_12059);
nand U28381 (N_28381,N_12388,N_17539);
or U28382 (N_28382,N_19508,N_10429);
xnor U28383 (N_28383,N_18362,N_13111);
or U28384 (N_28384,N_17321,N_19988);
and U28385 (N_28385,N_18748,N_18763);
nor U28386 (N_28386,N_15752,N_13605);
nor U28387 (N_28387,N_12212,N_15426);
xor U28388 (N_28388,N_10473,N_12802);
or U28389 (N_28389,N_15779,N_14793);
and U28390 (N_28390,N_11710,N_11602);
nor U28391 (N_28391,N_14416,N_11410);
nor U28392 (N_28392,N_16810,N_15866);
nand U28393 (N_28393,N_15282,N_15848);
or U28394 (N_28394,N_15944,N_18439);
nor U28395 (N_28395,N_15611,N_11829);
xnor U28396 (N_28396,N_11248,N_12934);
or U28397 (N_28397,N_17597,N_10489);
nand U28398 (N_28398,N_19089,N_18940);
or U28399 (N_28399,N_16224,N_14544);
and U28400 (N_28400,N_19101,N_13352);
and U28401 (N_28401,N_18763,N_17822);
or U28402 (N_28402,N_15763,N_16776);
and U28403 (N_28403,N_18387,N_16831);
and U28404 (N_28404,N_10803,N_12278);
and U28405 (N_28405,N_13697,N_19215);
or U28406 (N_28406,N_11639,N_15321);
and U28407 (N_28407,N_18298,N_11496);
nand U28408 (N_28408,N_18744,N_16211);
and U28409 (N_28409,N_11094,N_15647);
or U28410 (N_28410,N_17503,N_16552);
and U28411 (N_28411,N_15109,N_17468);
and U28412 (N_28412,N_19334,N_17231);
nor U28413 (N_28413,N_16966,N_15207);
nor U28414 (N_28414,N_13217,N_11113);
nand U28415 (N_28415,N_16330,N_15915);
or U28416 (N_28416,N_18888,N_16698);
nand U28417 (N_28417,N_17375,N_12253);
nand U28418 (N_28418,N_16288,N_18982);
and U28419 (N_28419,N_18883,N_17126);
or U28420 (N_28420,N_11800,N_16836);
or U28421 (N_28421,N_19869,N_19721);
or U28422 (N_28422,N_12347,N_17943);
and U28423 (N_28423,N_10166,N_14034);
xor U28424 (N_28424,N_14637,N_10353);
nor U28425 (N_28425,N_14793,N_11819);
and U28426 (N_28426,N_14228,N_11469);
nor U28427 (N_28427,N_17651,N_12852);
xor U28428 (N_28428,N_11223,N_10417);
or U28429 (N_28429,N_10374,N_12038);
xnor U28430 (N_28430,N_17020,N_14894);
or U28431 (N_28431,N_17644,N_19779);
nor U28432 (N_28432,N_11773,N_16756);
nand U28433 (N_28433,N_18704,N_19628);
nor U28434 (N_28434,N_19551,N_12719);
nand U28435 (N_28435,N_15971,N_12146);
or U28436 (N_28436,N_10078,N_15292);
and U28437 (N_28437,N_11158,N_13124);
nand U28438 (N_28438,N_12808,N_18902);
nand U28439 (N_28439,N_16721,N_10055);
nand U28440 (N_28440,N_10346,N_15265);
nor U28441 (N_28441,N_18387,N_10971);
nand U28442 (N_28442,N_17131,N_10629);
nand U28443 (N_28443,N_16054,N_17509);
nand U28444 (N_28444,N_12889,N_10291);
and U28445 (N_28445,N_15010,N_13884);
nor U28446 (N_28446,N_12191,N_13070);
and U28447 (N_28447,N_13633,N_18442);
xor U28448 (N_28448,N_12602,N_19781);
nand U28449 (N_28449,N_11074,N_19860);
xor U28450 (N_28450,N_17451,N_13949);
and U28451 (N_28451,N_10671,N_18524);
nand U28452 (N_28452,N_17014,N_10310);
and U28453 (N_28453,N_18085,N_12480);
or U28454 (N_28454,N_12075,N_18580);
nand U28455 (N_28455,N_11615,N_13686);
or U28456 (N_28456,N_12336,N_11553);
nor U28457 (N_28457,N_14190,N_11638);
nor U28458 (N_28458,N_16223,N_16889);
or U28459 (N_28459,N_11493,N_14766);
nand U28460 (N_28460,N_17077,N_12460);
and U28461 (N_28461,N_16058,N_14226);
nand U28462 (N_28462,N_10853,N_16478);
and U28463 (N_28463,N_15564,N_19089);
or U28464 (N_28464,N_12260,N_11555);
or U28465 (N_28465,N_12770,N_10136);
nand U28466 (N_28466,N_12443,N_12461);
nand U28467 (N_28467,N_16160,N_19668);
and U28468 (N_28468,N_11509,N_19560);
xor U28469 (N_28469,N_15744,N_19971);
and U28470 (N_28470,N_14498,N_13057);
or U28471 (N_28471,N_13440,N_16964);
or U28472 (N_28472,N_18343,N_11322);
xnor U28473 (N_28473,N_12618,N_14156);
nand U28474 (N_28474,N_11047,N_11491);
xor U28475 (N_28475,N_19265,N_16735);
nor U28476 (N_28476,N_12448,N_12558);
or U28477 (N_28477,N_13406,N_13815);
or U28478 (N_28478,N_19264,N_10074);
nor U28479 (N_28479,N_15473,N_15406);
or U28480 (N_28480,N_11389,N_16935);
nand U28481 (N_28481,N_11002,N_12668);
nand U28482 (N_28482,N_11391,N_18987);
or U28483 (N_28483,N_10231,N_10206);
or U28484 (N_28484,N_10936,N_12935);
or U28485 (N_28485,N_17040,N_12061);
or U28486 (N_28486,N_13530,N_13822);
nor U28487 (N_28487,N_18699,N_17130);
and U28488 (N_28488,N_12169,N_19541);
or U28489 (N_28489,N_18121,N_14936);
nor U28490 (N_28490,N_19285,N_14992);
nand U28491 (N_28491,N_18849,N_15323);
nand U28492 (N_28492,N_19555,N_18220);
and U28493 (N_28493,N_18909,N_19243);
nor U28494 (N_28494,N_15978,N_15588);
and U28495 (N_28495,N_19695,N_16863);
xor U28496 (N_28496,N_17377,N_19915);
and U28497 (N_28497,N_14499,N_16738);
nand U28498 (N_28498,N_14309,N_10216);
nor U28499 (N_28499,N_10714,N_19946);
or U28500 (N_28500,N_19672,N_19285);
and U28501 (N_28501,N_16341,N_12655);
nand U28502 (N_28502,N_17685,N_14665);
and U28503 (N_28503,N_16520,N_14465);
or U28504 (N_28504,N_13178,N_17087);
and U28505 (N_28505,N_10511,N_17585);
or U28506 (N_28506,N_12091,N_17130);
xnor U28507 (N_28507,N_12670,N_17820);
or U28508 (N_28508,N_11594,N_13195);
or U28509 (N_28509,N_11452,N_13105);
nand U28510 (N_28510,N_11200,N_10592);
and U28511 (N_28511,N_17521,N_10387);
or U28512 (N_28512,N_15184,N_14330);
nand U28513 (N_28513,N_11905,N_16556);
nor U28514 (N_28514,N_17405,N_11552);
xnor U28515 (N_28515,N_10536,N_15959);
and U28516 (N_28516,N_17010,N_18829);
or U28517 (N_28517,N_10467,N_12771);
or U28518 (N_28518,N_10239,N_15995);
or U28519 (N_28519,N_13288,N_19673);
nand U28520 (N_28520,N_18919,N_10576);
nand U28521 (N_28521,N_10397,N_10040);
and U28522 (N_28522,N_12293,N_18019);
and U28523 (N_28523,N_16679,N_14191);
or U28524 (N_28524,N_10692,N_14528);
or U28525 (N_28525,N_18997,N_18884);
or U28526 (N_28526,N_16786,N_19109);
nor U28527 (N_28527,N_11081,N_10607);
nor U28528 (N_28528,N_18986,N_14163);
nor U28529 (N_28529,N_14201,N_14642);
nor U28530 (N_28530,N_19313,N_10519);
nor U28531 (N_28531,N_12628,N_11123);
and U28532 (N_28532,N_19804,N_10727);
and U28533 (N_28533,N_17152,N_13848);
xnor U28534 (N_28534,N_18779,N_12097);
and U28535 (N_28535,N_19852,N_15020);
and U28536 (N_28536,N_17967,N_12198);
xnor U28537 (N_28537,N_17147,N_18940);
nand U28538 (N_28538,N_12733,N_17008);
or U28539 (N_28539,N_19196,N_10726);
nand U28540 (N_28540,N_17195,N_10368);
nor U28541 (N_28541,N_15644,N_13843);
xnor U28542 (N_28542,N_16085,N_10562);
nor U28543 (N_28543,N_16350,N_12453);
and U28544 (N_28544,N_17083,N_15796);
and U28545 (N_28545,N_15119,N_18655);
and U28546 (N_28546,N_19011,N_16236);
and U28547 (N_28547,N_19239,N_18122);
nor U28548 (N_28548,N_10581,N_17879);
and U28549 (N_28549,N_13227,N_18061);
nor U28550 (N_28550,N_19439,N_18633);
and U28551 (N_28551,N_16183,N_13087);
xnor U28552 (N_28552,N_16382,N_11919);
nand U28553 (N_28553,N_17034,N_16984);
xnor U28554 (N_28554,N_11758,N_19350);
and U28555 (N_28555,N_12489,N_15858);
or U28556 (N_28556,N_16345,N_11936);
nand U28557 (N_28557,N_16398,N_11689);
nand U28558 (N_28558,N_15024,N_14355);
or U28559 (N_28559,N_14231,N_16495);
nor U28560 (N_28560,N_16646,N_15585);
or U28561 (N_28561,N_16707,N_19133);
nand U28562 (N_28562,N_12824,N_15298);
nor U28563 (N_28563,N_14031,N_19720);
nand U28564 (N_28564,N_16621,N_12594);
nand U28565 (N_28565,N_19808,N_11490);
and U28566 (N_28566,N_14156,N_12950);
nor U28567 (N_28567,N_17240,N_11071);
nor U28568 (N_28568,N_14876,N_12406);
and U28569 (N_28569,N_15772,N_15058);
nor U28570 (N_28570,N_16175,N_14605);
nor U28571 (N_28571,N_17890,N_12834);
nor U28572 (N_28572,N_12020,N_12263);
or U28573 (N_28573,N_19010,N_10868);
nand U28574 (N_28574,N_10310,N_10674);
or U28575 (N_28575,N_15145,N_14357);
xor U28576 (N_28576,N_15407,N_12144);
or U28577 (N_28577,N_10721,N_15345);
nand U28578 (N_28578,N_19648,N_11506);
and U28579 (N_28579,N_17075,N_12786);
or U28580 (N_28580,N_17798,N_10239);
nand U28581 (N_28581,N_14065,N_18995);
and U28582 (N_28582,N_11964,N_19209);
and U28583 (N_28583,N_18775,N_10298);
nor U28584 (N_28584,N_18569,N_13923);
xor U28585 (N_28585,N_15867,N_14147);
and U28586 (N_28586,N_17910,N_11665);
or U28587 (N_28587,N_17581,N_14888);
nand U28588 (N_28588,N_16508,N_17699);
or U28589 (N_28589,N_13424,N_15028);
and U28590 (N_28590,N_10782,N_10237);
nand U28591 (N_28591,N_18126,N_19965);
nand U28592 (N_28592,N_13602,N_12013);
nor U28593 (N_28593,N_14288,N_13617);
and U28594 (N_28594,N_13000,N_13257);
nand U28595 (N_28595,N_13524,N_12309);
and U28596 (N_28596,N_19213,N_12618);
nor U28597 (N_28597,N_12154,N_10748);
nand U28598 (N_28598,N_11433,N_15013);
nand U28599 (N_28599,N_10655,N_10474);
xnor U28600 (N_28600,N_19935,N_12724);
and U28601 (N_28601,N_15458,N_14650);
and U28602 (N_28602,N_11226,N_19775);
or U28603 (N_28603,N_13378,N_18367);
nor U28604 (N_28604,N_13436,N_19995);
or U28605 (N_28605,N_13495,N_19294);
or U28606 (N_28606,N_14573,N_18038);
nand U28607 (N_28607,N_14599,N_14979);
or U28608 (N_28608,N_13785,N_16799);
and U28609 (N_28609,N_18325,N_11614);
and U28610 (N_28610,N_12420,N_18446);
nand U28611 (N_28611,N_14812,N_13172);
or U28612 (N_28612,N_15763,N_19147);
nor U28613 (N_28613,N_18775,N_18852);
xnor U28614 (N_28614,N_17960,N_11467);
nor U28615 (N_28615,N_16861,N_10592);
nand U28616 (N_28616,N_19960,N_12640);
nand U28617 (N_28617,N_18284,N_11607);
nand U28618 (N_28618,N_13721,N_11124);
and U28619 (N_28619,N_19564,N_10354);
or U28620 (N_28620,N_10585,N_17108);
nor U28621 (N_28621,N_19096,N_13652);
or U28622 (N_28622,N_19337,N_13421);
nor U28623 (N_28623,N_15247,N_16531);
nor U28624 (N_28624,N_14555,N_11604);
and U28625 (N_28625,N_13583,N_11806);
and U28626 (N_28626,N_12885,N_16376);
nand U28627 (N_28627,N_14288,N_18859);
nor U28628 (N_28628,N_10455,N_13232);
and U28629 (N_28629,N_16008,N_19989);
nor U28630 (N_28630,N_12435,N_13766);
or U28631 (N_28631,N_16486,N_19817);
nand U28632 (N_28632,N_14979,N_17991);
nand U28633 (N_28633,N_19946,N_13926);
and U28634 (N_28634,N_15588,N_19706);
nor U28635 (N_28635,N_15427,N_10684);
xor U28636 (N_28636,N_19413,N_16569);
nand U28637 (N_28637,N_15964,N_11185);
nand U28638 (N_28638,N_10415,N_17348);
and U28639 (N_28639,N_19004,N_10443);
nor U28640 (N_28640,N_16698,N_16710);
or U28641 (N_28641,N_15653,N_18248);
or U28642 (N_28642,N_11573,N_11476);
and U28643 (N_28643,N_16606,N_16115);
or U28644 (N_28644,N_18599,N_18494);
nand U28645 (N_28645,N_12653,N_18978);
nor U28646 (N_28646,N_11625,N_17758);
nand U28647 (N_28647,N_17104,N_14344);
nor U28648 (N_28648,N_17928,N_18559);
xnor U28649 (N_28649,N_15615,N_14045);
and U28650 (N_28650,N_13104,N_13652);
and U28651 (N_28651,N_17953,N_12974);
nand U28652 (N_28652,N_14808,N_11249);
or U28653 (N_28653,N_10780,N_17321);
or U28654 (N_28654,N_15145,N_14611);
or U28655 (N_28655,N_16214,N_15899);
nor U28656 (N_28656,N_11286,N_13016);
xnor U28657 (N_28657,N_17582,N_16718);
or U28658 (N_28658,N_15680,N_14192);
and U28659 (N_28659,N_15065,N_18864);
and U28660 (N_28660,N_12342,N_16099);
and U28661 (N_28661,N_12220,N_12888);
nor U28662 (N_28662,N_15408,N_13400);
nand U28663 (N_28663,N_11775,N_18696);
nor U28664 (N_28664,N_16149,N_19136);
or U28665 (N_28665,N_15345,N_16438);
nor U28666 (N_28666,N_11819,N_12413);
and U28667 (N_28667,N_18193,N_15427);
nor U28668 (N_28668,N_16920,N_15016);
nor U28669 (N_28669,N_11078,N_14427);
nand U28670 (N_28670,N_14996,N_15224);
or U28671 (N_28671,N_11073,N_11866);
nor U28672 (N_28672,N_13852,N_15443);
and U28673 (N_28673,N_18323,N_14376);
and U28674 (N_28674,N_17474,N_16489);
or U28675 (N_28675,N_10546,N_19558);
nand U28676 (N_28676,N_16092,N_16665);
nand U28677 (N_28677,N_14892,N_11495);
and U28678 (N_28678,N_15182,N_19681);
nand U28679 (N_28679,N_19242,N_17055);
or U28680 (N_28680,N_14567,N_10488);
nand U28681 (N_28681,N_16461,N_12257);
nor U28682 (N_28682,N_17071,N_18456);
nor U28683 (N_28683,N_12730,N_12312);
or U28684 (N_28684,N_19478,N_18022);
or U28685 (N_28685,N_13191,N_12014);
nand U28686 (N_28686,N_15099,N_12331);
or U28687 (N_28687,N_10039,N_11286);
and U28688 (N_28688,N_16221,N_17683);
nor U28689 (N_28689,N_14729,N_10676);
or U28690 (N_28690,N_10476,N_16433);
nor U28691 (N_28691,N_15338,N_12511);
nor U28692 (N_28692,N_16311,N_10306);
nand U28693 (N_28693,N_16395,N_16152);
xnor U28694 (N_28694,N_18887,N_10724);
or U28695 (N_28695,N_19189,N_18683);
nand U28696 (N_28696,N_15708,N_12051);
nand U28697 (N_28697,N_15611,N_17108);
nor U28698 (N_28698,N_16278,N_15229);
nand U28699 (N_28699,N_19482,N_15847);
or U28700 (N_28700,N_12187,N_11287);
nand U28701 (N_28701,N_18223,N_15220);
or U28702 (N_28702,N_13012,N_11326);
nand U28703 (N_28703,N_15816,N_12989);
xor U28704 (N_28704,N_14883,N_16500);
nand U28705 (N_28705,N_14600,N_13828);
or U28706 (N_28706,N_18720,N_17112);
nand U28707 (N_28707,N_14676,N_18234);
and U28708 (N_28708,N_19473,N_11447);
nand U28709 (N_28709,N_18478,N_13081);
nand U28710 (N_28710,N_11882,N_12317);
and U28711 (N_28711,N_13000,N_13743);
xor U28712 (N_28712,N_12757,N_10897);
xor U28713 (N_28713,N_13250,N_18926);
nor U28714 (N_28714,N_11756,N_18936);
nand U28715 (N_28715,N_15849,N_16302);
nor U28716 (N_28716,N_11344,N_17529);
and U28717 (N_28717,N_11800,N_16834);
nand U28718 (N_28718,N_17468,N_13917);
nand U28719 (N_28719,N_11401,N_17418);
and U28720 (N_28720,N_14835,N_18929);
nand U28721 (N_28721,N_16708,N_18848);
or U28722 (N_28722,N_13148,N_12768);
or U28723 (N_28723,N_15567,N_17747);
nand U28724 (N_28724,N_16942,N_17917);
nor U28725 (N_28725,N_17867,N_12884);
nor U28726 (N_28726,N_12456,N_17832);
or U28727 (N_28727,N_12959,N_13597);
nand U28728 (N_28728,N_19299,N_18080);
nor U28729 (N_28729,N_11465,N_19341);
nor U28730 (N_28730,N_10754,N_18789);
xnor U28731 (N_28731,N_12574,N_18789);
or U28732 (N_28732,N_19360,N_14226);
nand U28733 (N_28733,N_12127,N_19718);
and U28734 (N_28734,N_13945,N_17886);
nor U28735 (N_28735,N_10260,N_11122);
nor U28736 (N_28736,N_16268,N_12420);
nor U28737 (N_28737,N_12808,N_11997);
xor U28738 (N_28738,N_16428,N_12656);
and U28739 (N_28739,N_15000,N_17128);
and U28740 (N_28740,N_16061,N_10692);
nor U28741 (N_28741,N_10878,N_19489);
and U28742 (N_28742,N_19140,N_18810);
nor U28743 (N_28743,N_19948,N_13008);
xnor U28744 (N_28744,N_12491,N_13967);
nand U28745 (N_28745,N_19975,N_18503);
xor U28746 (N_28746,N_17395,N_17479);
nor U28747 (N_28747,N_15426,N_17253);
or U28748 (N_28748,N_16032,N_11441);
nor U28749 (N_28749,N_13327,N_18458);
nor U28750 (N_28750,N_17593,N_18367);
or U28751 (N_28751,N_18868,N_15563);
nor U28752 (N_28752,N_11964,N_12474);
and U28753 (N_28753,N_15468,N_10003);
nand U28754 (N_28754,N_17570,N_15922);
or U28755 (N_28755,N_15104,N_17045);
and U28756 (N_28756,N_11150,N_18566);
nor U28757 (N_28757,N_14594,N_15955);
and U28758 (N_28758,N_15960,N_19622);
or U28759 (N_28759,N_14408,N_15123);
or U28760 (N_28760,N_17680,N_19006);
nor U28761 (N_28761,N_15387,N_10110);
nor U28762 (N_28762,N_13927,N_17880);
nor U28763 (N_28763,N_10294,N_14398);
or U28764 (N_28764,N_12836,N_13218);
nor U28765 (N_28765,N_11396,N_15004);
nor U28766 (N_28766,N_16873,N_16343);
or U28767 (N_28767,N_15475,N_18194);
or U28768 (N_28768,N_18417,N_14103);
or U28769 (N_28769,N_15110,N_19426);
and U28770 (N_28770,N_19097,N_11088);
and U28771 (N_28771,N_19771,N_14455);
nor U28772 (N_28772,N_11862,N_11518);
nand U28773 (N_28773,N_16033,N_16669);
and U28774 (N_28774,N_14034,N_18351);
nand U28775 (N_28775,N_12776,N_16108);
or U28776 (N_28776,N_18291,N_16906);
and U28777 (N_28777,N_11498,N_16906);
and U28778 (N_28778,N_19039,N_14513);
nand U28779 (N_28779,N_12022,N_12673);
nor U28780 (N_28780,N_17072,N_14454);
and U28781 (N_28781,N_15140,N_15070);
or U28782 (N_28782,N_18552,N_19561);
nand U28783 (N_28783,N_12347,N_11787);
or U28784 (N_28784,N_17988,N_12702);
xor U28785 (N_28785,N_10778,N_10729);
nand U28786 (N_28786,N_12188,N_12220);
or U28787 (N_28787,N_14908,N_19061);
and U28788 (N_28788,N_10204,N_13433);
nor U28789 (N_28789,N_15566,N_19167);
nor U28790 (N_28790,N_17901,N_18423);
or U28791 (N_28791,N_13720,N_13377);
nor U28792 (N_28792,N_11398,N_12914);
nor U28793 (N_28793,N_12491,N_11753);
and U28794 (N_28794,N_17219,N_18470);
and U28795 (N_28795,N_11754,N_13176);
nand U28796 (N_28796,N_12149,N_12387);
nand U28797 (N_28797,N_14987,N_11432);
nor U28798 (N_28798,N_12462,N_15794);
xor U28799 (N_28799,N_11520,N_11100);
nor U28800 (N_28800,N_17027,N_11098);
nand U28801 (N_28801,N_11516,N_10717);
nor U28802 (N_28802,N_19659,N_18254);
and U28803 (N_28803,N_18387,N_12678);
nor U28804 (N_28804,N_11479,N_12687);
nand U28805 (N_28805,N_15882,N_15731);
xor U28806 (N_28806,N_14025,N_17672);
nor U28807 (N_28807,N_12779,N_16001);
and U28808 (N_28808,N_17170,N_10514);
nand U28809 (N_28809,N_13030,N_10179);
nor U28810 (N_28810,N_15364,N_13003);
or U28811 (N_28811,N_15244,N_13620);
and U28812 (N_28812,N_12709,N_13475);
nand U28813 (N_28813,N_15288,N_16882);
and U28814 (N_28814,N_15239,N_10653);
nor U28815 (N_28815,N_13586,N_14401);
or U28816 (N_28816,N_13785,N_13456);
nor U28817 (N_28817,N_19403,N_12923);
and U28818 (N_28818,N_19476,N_17304);
nor U28819 (N_28819,N_12494,N_11877);
and U28820 (N_28820,N_15337,N_15644);
nand U28821 (N_28821,N_18509,N_10550);
and U28822 (N_28822,N_10274,N_14756);
nor U28823 (N_28823,N_14681,N_19379);
or U28824 (N_28824,N_10896,N_16571);
nor U28825 (N_28825,N_19263,N_12855);
or U28826 (N_28826,N_18544,N_16676);
or U28827 (N_28827,N_16867,N_11561);
xnor U28828 (N_28828,N_11743,N_14692);
nor U28829 (N_28829,N_18133,N_11692);
nor U28830 (N_28830,N_15982,N_11266);
or U28831 (N_28831,N_17198,N_16795);
nand U28832 (N_28832,N_16135,N_13297);
nor U28833 (N_28833,N_14289,N_19605);
and U28834 (N_28834,N_19190,N_11080);
nand U28835 (N_28835,N_17019,N_17103);
or U28836 (N_28836,N_12083,N_18178);
nand U28837 (N_28837,N_15660,N_10394);
nand U28838 (N_28838,N_16843,N_15076);
and U28839 (N_28839,N_19842,N_12697);
or U28840 (N_28840,N_17435,N_15191);
nand U28841 (N_28841,N_13870,N_12009);
nor U28842 (N_28842,N_14523,N_18942);
or U28843 (N_28843,N_15873,N_15129);
or U28844 (N_28844,N_13469,N_10769);
nor U28845 (N_28845,N_15498,N_18462);
and U28846 (N_28846,N_15764,N_13627);
or U28847 (N_28847,N_13605,N_15925);
nand U28848 (N_28848,N_11915,N_19437);
xor U28849 (N_28849,N_13173,N_18625);
and U28850 (N_28850,N_10353,N_11612);
or U28851 (N_28851,N_14861,N_12033);
or U28852 (N_28852,N_16771,N_17498);
or U28853 (N_28853,N_14043,N_10417);
or U28854 (N_28854,N_19036,N_14162);
nor U28855 (N_28855,N_10323,N_18645);
and U28856 (N_28856,N_10128,N_16254);
nor U28857 (N_28857,N_11182,N_19794);
nor U28858 (N_28858,N_16311,N_12734);
nand U28859 (N_28859,N_12481,N_12372);
nand U28860 (N_28860,N_11432,N_11497);
nor U28861 (N_28861,N_16434,N_18639);
or U28862 (N_28862,N_19419,N_19217);
and U28863 (N_28863,N_18827,N_12427);
or U28864 (N_28864,N_15669,N_16384);
or U28865 (N_28865,N_16726,N_13783);
and U28866 (N_28866,N_12102,N_17281);
nand U28867 (N_28867,N_13664,N_11826);
and U28868 (N_28868,N_17845,N_16212);
nand U28869 (N_28869,N_17215,N_10206);
nor U28870 (N_28870,N_15275,N_10757);
nand U28871 (N_28871,N_13948,N_11221);
or U28872 (N_28872,N_19106,N_11500);
nor U28873 (N_28873,N_18406,N_15039);
nor U28874 (N_28874,N_13782,N_16271);
nand U28875 (N_28875,N_14465,N_16670);
nor U28876 (N_28876,N_19164,N_13077);
nor U28877 (N_28877,N_11485,N_17732);
or U28878 (N_28878,N_14833,N_12000);
or U28879 (N_28879,N_16744,N_14631);
and U28880 (N_28880,N_12669,N_16390);
nor U28881 (N_28881,N_17317,N_10392);
or U28882 (N_28882,N_19167,N_12471);
nand U28883 (N_28883,N_14961,N_18868);
nand U28884 (N_28884,N_16627,N_16924);
or U28885 (N_28885,N_17108,N_14947);
nand U28886 (N_28886,N_16648,N_11379);
or U28887 (N_28887,N_11237,N_16166);
nor U28888 (N_28888,N_17104,N_10902);
and U28889 (N_28889,N_13841,N_11753);
or U28890 (N_28890,N_19937,N_14406);
and U28891 (N_28891,N_13423,N_13254);
or U28892 (N_28892,N_16499,N_12668);
and U28893 (N_28893,N_16565,N_13788);
nand U28894 (N_28894,N_12771,N_18098);
nand U28895 (N_28895,N_17979,N_14464);
nor U28896 (N_28896,N_15687,N_18017);
nor U28897 (N_28897,N_16347,N_13867);
nor U28898 (N_28898,N_16424,N_10161);
nand U28899 (N_28899,N_15347,N_12303);
or U28900 (N_28900,N_10477,N_17248);
and U28901 (N_28901,N_15750,N_16060);
nor U28902 (N_28902,N_10636,N_10561);
nor U28903 (N_28903,N_19679,N_16042);
and U28904 (N_28904,N_12640,N_19637);
nor U28905 (N_28905,N_15173,N_12662);
and U28906 (N_28906,N_15134,N_11879);
nand U28907 (N_28907,N_15487,N_12355);
and U28908 (N_28908,N_10649,N_18170);
nor U28909 (N_28909,N_16344,N_10982);
nand U28910 (N_28910,N_11390,N_10695);
nor U28911 (N_28911,N_18559,N_17919);
and U28912 (N_28912,N_19509,N_13748);
or U28913 (N_28913,N_16576,N_18056);
or U28914 (N_28914,N_11109,N_16718);
and U28915 (N_28915,N_12328,N_17236);
or U28916 (N_28916,N_16228,N_14829);
and U28917 (N_28917,N_14572,N_17773);
or U28918 (N_28918,N_18670,N_14546);
and U28919 (N_28919,N_11740,N_15836);
or U28920 (N_28920,N_18753,N_16776);
and U28921 (N_28921,N_17323,N_18544);
nand U28922 (N_28922,N_17551,N_11253);
nor U28923 (N_28923,N_13464,N_15458);
or U28924 (N_28924,N_10050,N_10882);
nand U28925 (N_28925,N_15291,N_13925);
or U28926 (N_28926,N_16695,N_16664);
and U28927 (N_28927,N_11318,N_19702);
nand U28928 (N_28928,N_10426,N_16808);
nor U28929 (N_28929,N_11753,N_16474);
or U28930 (N_28930,N_14826,N_16924);
xnor U28931 (N_28931,N_11896,N_10871);
and U28932 (N_28932,N_12872,N_10446);
nand U28933 (N_28933,N_19112,N_19503);
or U28934 (N_28934,N_16620,N_11043);
nor U28935 (N_28935,N_10600,N_19787);
nand U28936 (N_28936,N_18114,N_16316);
nor U28937 (N_28937,N_13897,N_18521);
nor U28938 (N_28938,N_18727,N_15364);
nand U28939 (N_28939,N_10986,N_13868);
nand U28940 (N_28940,N_10693,N_10742);
and U28941 (N_28941,N_18109,N_10541);
nand U28942 (N_28942,N_18391,N_16736);
nand U28943 (N_28943,N_19195,N_14377);
nand U28944 (N_28944,N_10971,N_12677);
nor U28945 (N_28945,N_16192,N_10792);
or U28946 (N_28946,N_18159,N_14332);
and U28947 (N_28947,N_10841,N_13317);
xnor U28948 (N_28948,N_15211,N_15683);
nor U28949 (N_28949,N_11745,N_14844);
and U28950 (N_28950,N_13778,N_17763);
xor U28951 (N_28951,N_19267,N_18630);
nor U28952 (N_28952,N_14099,N_10895);
nand U28953 (N_28953,N_15269,N_18182);
or U28954 (N_28954,N_10935,N_10698);
nand U28955 (N_28955,N_16878,N_10704);
or U28956 (N_28956,N_10186,N_12767);
nor U28957 (N_28957,N_18074,N_10916);
nand U28958 (N_28958,N_12518,N_19674);
and U28959 (N_28959,N_17196,N_19824);
nor U28960 (N_28960,N_12410,N_18396);
or U28961 (N_28961,N_19645,N_19420);
nand U28962 (N_28962,N_10527,N_12197);
nand U28963 (N_28963,N_12876,N_19831);
nand U28964 (N_28964,N_16675,N_13571);
or U28965 (N_28965,N_14820,N_14881);
or U28966 (N_28966,N_17161,N_17788);
or U28967 (N_28967,N_15610,N_15364);
or U28968 (N_28968,N_14304,N_16138);
nand U28969 (N_28969,N_11770,N_12783);
nand U28970 (N_28970,N_14105,N_19830);
nor U28971 (N_28971,N_14244,N_15446);
and U28972 (N_28972,N_13166,N_11019);
nand U28973 (N_28973,N_14325,N_15625);
nand U28974 (N_28974,N_14499,N_13755);
nand U28975 (N_28975,N_19689,N_17032);
or U28976 (N_28976,N_17291,N_19312);
xnor U28977 (N_28977,N_15400,N_10022);
and U28978 (N_28978,N_18214,N_15914);
and U28979 (N_28979,N_15962,N_10574);
or U28980 (N_28980,N_10332,N_15877);
xor U28981 (N_28981,N_15246,N_16498);
or U28982 (N_28982,N_18943,N_19577);
nor U28983 (N_28983,N_19077,N_18163);
or U28984 (N_28984,N_19373,N_13967);
xor U28985 (N_28985,N_12745,N_13296);
nor U28986 (N_28986,N_14801,N_17504);
or U28987 (N_28987,N_13043,N_10363);
xnor U28988 (N_28988,N_12321,N_16118);
nor U28989 (N_28989,N_11558,N_14545);
or U28990 (N_28990,N_10330,N_11898);
or U28991 (N_28991,N_13161,N_12133);
nand U28992 (N_28992,N_15485,N_10956);
and U28993 (N_28993,N_10776,N_10462);
or U28994 (N_28994,N_16418,N_12697);
and U28995 (N_28995,N_16785,N_17393);
nand U28996 (N_28996,N_14230,N_11274);
nor U28997 (N_28997,N_17074,N_18426);
nand U28998 (N_28998,N_12742,N_12350);
and U28999 (N_28999,N_11859,N_14754);
or U29000 (N_29000,N_15969,N_18164);
nor U29001 (N_29001,N_17100,N_18913);
nand U29002 (N_29002,N_17860,N_14956);
nand U29003 (N_29003,N_10741,N_15908);
nor U29004 (N_29004,N_12966,N_10696);
nand U29005 (N_29005,N_16894,N_12175);
or U29006 (N_29006,N_10988,N_11332);
nand U29007 (N_29007,N_11705,N_12775);
and U29008 (N_29008,N_13061,N_13703);
xor U29009 (N_29009,N_13202,N_13001);
nand U29010 (N_29010,N_11200,N_18678);
and U29011 (N_29011,N_19025,N_10098);
or U29012 (N_29012,N_15937,N_14107);
or U29013 (N_29013,N_15254,N_13596);
nand U29014 (N_29014,N_18266,N_17180);
nand U29015 (N_29015,N_18154,N_12655);
or U29016 (N_29016,N_12823,N_10756);
or U29017 (N_29017,N_17809,N_17393);
xor U29018 (N_29018,N_11620,N_13025);
and U29019 (N_29019,N_17972,N_15987);
and U29020 (N_29020,N_11280,N_14735);
or U29021 (N_29021,N_17113,N_17801);
and U29022 (N_29022,N_19323,N_15792);
or U29023 (N_29023,N_18569,N_14961);
nor U29024 (N_29024,N_13556,N_14429);
nand U29025 (N_29025,N_14021,N_13873);
nand U29026 (N_29026,N_13481,N_15986);
nand U29027 (N_29027,N_12767,N_17579);
nor U29028 (N_29028,N_13439,N_12344);
nand U29029 (N_29029,N_18226,N_18618);
or U29030 (N_29030,N_19212,N_12050);
xnor U29031 (N_29031,N_13333,N_10681);
nor U29032 (N_29032,N_10295,N_11681);
xor U29033 (N_29033,N_16951,N_18134);
and U29034 (N_29034,N_18608,N_19275);
or U29035 (N_29035,N_12426,N_19978);
and U29036 (N_29036,N_12578,N_13274);
and U29037 (N_29037,N_17066,N_13401);
nand U29038 (N_29038,N_15087,N_15190);
nor U29039 (N_29039,N_11851,N_15058);
nand U29040 (N_29040,N_14376,N_18878);
nand U29041 (N_29041,N_16179,N_13885);
nor U29042 (N_29042,N_12404,N_11711);
or U29043 (N_29043,N_11277,N_18692);
nand U29044 (N_29044,N_15126,N_16507);
and U29045 (N_29045,N_15025,N_10889);
nor U29046 (N_29046,N_19836,N_17271);
nand U29047 (N_29047,N_16884,N_12753);
nor U29048 (N_29048,N_11040,N_16356);
nor U29049 (N_29049,N_14309,N_19234);
xnor U29050 (N_29050,N_17547,N_10456);
nand U29051 (N_29051,N_16935,N_12217);
nor U29052 (N_29052,N_14290,N_10611);
or U29053 (N_29053,N_14068,N_13999);
and U29054 (N_29054,N_11459,N_11597);
nor U29055 (N_29055,N_17982,N_15291);
and U29056 (N_29056,N_15312,N_17245);
nor U29057 (N_29057,N_13739,N_10410);
xnor U29058 (N_29058,N_11371,N_12587);
nand U29059 (N_29059,N_10893,N_14804);
nand U29060 (N_29060,N_14005,N_11456);
xor U29061 (N_29061,N_14838,N_12499);
nor U29062 (N_29062,N_16109,N_18375);
nand U29063 (N_29063,N_10567,N_18581);
nand U29064 (N_29064,N_16223,N_11604);
and U29065 (N_29065,N_17157,N_17534);
and U29066 (N_29066,N_13854,N_11566);
nand U29067 (N_29067,N_15665,N_17551);
nor U29068 (N_29068,N_12356,N_14857);
nand U29069 (N_29069,N_13109,N_15811);
or U29070 (N_29070,N_14778,N_14079);
or U29071 (N_29071,N_17595,N_18407);
or U29072 (N_29072,N_17418,N_13127);
nand U29073 (N_29073,N_13604,N_17050);
nand U29074 (N_29074,N_18013,N_12038);
or U29075 (N_29075,N_12339,N_19966);
nand U29076 (N_29076,N_17688,N_16533);
nor U29077 (N_29077,N_14993,N_10688);
or U29078 (N_29078,N_15337,N_16198);
nor U29079 (N_29079,N_13359,N_17422);
and U29080 (N_29080,N_16797,N_18097);
nor U29081 (N_29081,N_11542,N_13097);
and U29082 (N_29082,N_19257,N_10381);
nand U29083 (N_29083,N_18778,N_17502);
nor U29084 (N_29084,N_11194,N_18958);
or U29085 (N_29085,N_12957,N_11355);
and U29086 (N_29086,N_17515,N_17903);
nor U29087 (N_29087,N_10546,N_12185);
nor U29088 (N_29088,N_12040,N_15278);
xnor U29089 (N_29089,N_18672,N_19247);
xnor U29090 (N_29090,N_15495,N_14990);
nand U29091 (N_29091,N_17437,N_10838);
or U29092 (N_29092,N_16597,N_11272);
xor U29093 (N_29093,N_16136,N_16577);
and U29094 (N_29094,N_19768,N_17405);
nand U29095 (N_29095,N_16586,N_14553);
or U29096 (N_29096,N_12501,N_18836);
nor U29097 (N_29097,N_11187,N_13565);
nor U29098 (N_29098,N_16427,N_14573);
or U29099 (N_29099,N_13172,N_13092);
and U29100 (N_29100,N_13754,N_12030);
nand U29101 (N_29101,N_18100,N_13855);
nor U29102 (N_29102,N_14360,N_10355);
nor U29103 (N_29103,N_13485,N_17050);
nor U29104 (N_29104,N_15322,N_15912);
nor U29105 (N_29105,N_13729,N_16519);
or U29106 (N_29106,N_13234,N_12257);
or U29107 (N_29107,N_11042,N_16999);
nand U29108 (N_29108,N_13664,N_19687);
nand U29109 (N_29109,N_16445,N_17850);
nand U29110 (N_29110,N_13421,N_18145);
and U29111 (N_29111,N_14051,N_18170);
nand U29112 (N_29112,N_17384,N_13501);
xor U29113 (N_29113,N_15439,N_14210);
nand U29114 (N_29114,N_10679,N_14654);
and U29115 (N_29115,N_15459,N_12166);
xnor U29116 (N_29116,N_13191,N_11069);
and U29117 (N_29117,N_15683,N_10503);
nand U29118 (N_29118,N_19360,N_14330);
and U29119 (N_29119,N_10572,N_17136);
nor U29120 (N_29120,N_17336,N_17237);
and U29121 (N_29121,N_19361,N_19443);
nand U29122 (N_29122,N_10803,N_13832);
or U29123 (N_29123,N_18533,N_19363);
nand U29124 (N_29124,N_13444,N_12726);
nand U29125 (N_29125,N_18618,N_12867);
nand U29126 (N_29126,N_10470,N_12972);
or U29127 (N_29127,N_14991,N_16477);
and U29128 (N_29128,N_19549,N_18562);
nor U29129 (N_29129,N_15411,N_19434);
and U29130 (N_29130,N_10661,N_15857);
nor U29131 (N_29131,N_19106,N_11015);
and U29132 (N_29132,N_14793,N_11998);
or U29133 (N_29133,N_16096,N_15994);
nand U29134 (N_29134,N_13915,N_16064);
nor U29135 (N_29135,N_10580,N_11967);
or U29136 (N_29136,N_10662,N_17594);
and U29137 (N_29137,N_14417,N_19211);
nor U29138 (N_29138,N_15864,N_14994);
nor U29139 (N_29139,N_18939,N_16005);
and U29140 (N_29140,N_16852,N_11767);
or U29141 (N_29141,N_11458,N_15306);
or U29142 (N_29142,N_17411,N_19518);
and U29143 (N_29143,N_10141,N_17656);
and U29144 (N_29144,N_11744,N_11141);
nor U29145 (N_29145,N_13499,N_16566);
xnor U29146 (N_29146,N_13633,N_12745);
and U29147 (N_29147,N_17302,N_13435);
or U29148 (N_29148,N_19423,N_13078);
or U29149 (N_29149,N_13365,N_19271);
and U29150 (N_29150,N_18299,N_14121);
and U29151 (N_29151,N_17690,N_18709);
and U29152 (N_29152,N_15547,N_11674);
nand U29153 (N_29153,N_15597,N_13283);
or U29154 (N_29154,N_14718,N_12730);
nand U29155 (N_29155,N_19859,N_11959);
or U29156 (N_29156,N_11798,N_17786);
and U29157 (N_29157,N_12217,N_15383);
nor U29158 (N_29158,N_13787,N_10527);
xor U29159 (N_29159,N_15049,N_14586);
and U29160 (N_29160,N_13666,N_19552);
nand U29161 (N_29161,N_13430,N_16956);
and U29162 (N_29162,N_10379,N_17922);
and U29163 (N_29163,N_18828,N_19096);
or U29164 (N_29164,N_12316,N_15332);
and U29165 (N_29165,N_18254,N_19446);
nand U29166 (N_29166,N_15709,N_16226);
nand U29167 (N_29167,N_10994,N_15629);
nand U29168 (N_29168,N_13705,N_17085);
and U29169 (N_29169,N_16928,N_15960);
and U29170 (N_29170,N_13568,N_19422);
nor U29171 (N_29171,N_16697,N_16954);
and U29172 (N_29172,N_14948,N_13999);
nand U29173 (N_29173,N_11502,N_17345);
and U29174 (N_29174,N_15465,N_18382);
or U29175 (N_29175,N_18120,N_16371);
or U29176 (N_29176,N_14698,N_11140);
nor U29177 (N_29177,N_14345,N_12354);
or U29178 (N_29178,N_18716,N_15302);
or U29179 (N_29179,N_15804,N_13056);
and U29180 (N_29180,N_16747,N_16356);
and U29181 (N_29181,N_14289,N_17190);
nor U29182 (N_29182,N_19174,N_15367);
nor U29183 (N_29183,N_19522,N_12568);
and U29184 (N_29184,N_13922,N_16264);
nand U29185 (N_29185,N_19366,N_19430);
nor U29186 (N_29186,N_13915,N_19939);
nand U29187 (N_29187,N_16924,N_18942);
nand U29188 (N_29188,N_11605,N_16624);
nand U29189 (N_29189,N_13116,N_19168);
nor U29190 (N_29190,N_11665,N_11406);
nand U29191 (N_29191,N_11573,N_18988);
and U29192 (N_29192,N_17183,N_12131);
or U29193 (N_29193,N_12756,N_17789);
nand U29194 (N_29194,N_12633,N_17367);
and U29195 (N_29195,N_16364,N_12149);
or U29196 (N_29196,N_13485,N_12100);
or U29197 (N_29197,N_15870,N_12291);
xnor U29198 (N_29198,N_14246,N_12225);
and U29199 (N_29199,N_12172,N_19829);
nor U29200 (N_29200,N_13829,N_15253);
nand U29201 (N_29201,N_12725,N_13552);
nand U29202 (N_29202,N_15238,N_17319);
nor U29203 (N_29203,N_10970,N_18840);
nor U29204 (N_29204,N_12960,N_19754);
nor U29205 (N_29205,N_17347,N_16927);
nor U29206 (N_29206,N_18342,N_14319);
xnor U29207 (N_29207,N_18874,N_10781);
nand U29208 (N_29208,N_14469,N_19839);
nor U29209 (N_29209,N_11873,N_11268);
or U29210 (N_29210,N_12404,N_13870);
nand U29211 (N_29211,N_11810,N_12385);
and U29212 (N_29212,N_12585,N_18727);
or U29213 (N_29213,N_19486,N_13236);
nor U29214 (N_29214,N_17277,N_19441);
xor U29215 (N_29215,N_19224,N_16763);
and U29216 (N_29216,N_18910,N_18637);
or U29217 (N_29217,N_19137,N_11652);
nor U29218 (N_29218,N_10264,N_16736);
and U29219 (N_29219,N_18953,N_13620);
nor U29220 (N_29220,N_16297,N_18464);
and U29221 (N_29221,N_14705,N_10822);
and U29222 (N_29222,N_17683,N_17215);
nor U29223 (N_29223,N_14710,N_17199);
or U29224 (N_29224,N_13756,N_13972);
and U29225 (N_29225,N_14483,N_17403);
or U29226 (N_29226,N_12070,N_12817);
nor U29227 (N_29227,N_16677,N_11213);
nand U29228 (N_29228,N_12389,N_12179);
nor U29229 (N_29229,N_10657,N_10237);
nand U29230 (N_29230,N_16122,N_13463);
nand U29231 (N_29231,N_13279,N_16643);
and U29232 (N_29232,N_19687,N_17397);
and U29233 (N_29233,N_15811,N_18043);
xor U29234 (N_29234,N_14724,N_16635);
or U29235 (N_29235,N_11042,N_18681);
xnor U29236 (N_29236,N_11922,N_19899);
and U29237 (N_29237,N_10573,N_17361);
nor U29238 (N_29238,N_14712,N_19799);
nor U29239 (N_29239,N_15290,N_19016);
nand U29240 (N_29240,N_17424,N_12759);
xnor U29241 (N_29241,N_13277,N_18296);
nor U29242 (N_29242,N_17340,N_12416);
or U29243 (N_29243,N_19605,N_16752);
nand U29244 (N_29244,N_15110,N_19702);
nand U29245 (N_29245,N_10799,N_17562);
or U29246 (N_29246,N_15934,N_13826);
nand U29247 (N_29247,N_14140,N_17723);
nand U29248 (N_29248,N_18741,N_17576);
or U29249 (N_29249,N_19293,N_18260);
or U29250 (N_29250,N_13408,N_18697);
nor U29251 (N_29251,N_10966,N_18940);
or U29252 (N_29252,N_18389,N_10343);
or U29253 (N_29253,N_10373,N_18664);
xnor U29254 (N_29254,N_11732,N_10259);
or U29255 (N_29255,N_14208,N_16403);
nor U29256 (N_29256,N_10305,N_15457);
and U29257 (N_29257,N_17947,N_12252);
xor U29258 (N_29258,N_12738,N_11876);
or U29259 (N_29259,N_10984,N_14633);
nor U29260 (N_29260,N_16953,N_14030);
nor U29261 (N_29261,N_19704,N_16026);
nand U29262 (N_29262,N_10899,N_19806);
nor U29263 (N_29263,N_10909,N_12643);
or U29264 (N_29264,N_11364,N_19997);
nor U29265 (N_29265,N_13001,N_16888);
and U29266 (N_29266,N_11940,N_16083);
and U29267 (N_29267,N_11603,N_17577);
xnor U29268 (N_29268,N_19415,N_16725);
xor U29269 (N_29269,N_17042,N_11877);
nand U29270 (N_29270,N_17235,N_10064);
nor U29271 (N_29271,N_15559,N_18882);
nor U29272 (N_29272,N_13810,N_12929);
nand U29273 (N_29273,N_18082,N_13370);
nor U29274 (N_29274,N_17649,N_10042);
xor U29275 (N_29275,N_12395,N_10607);
nor U29276 (N_29276,N_18244,N_12030);
nor U29277 (N_29277,N_13938,N_10619);
and U29278 (N_29278,N_14037,N_15115);
nor U29279 (N_29279,N_12171,N_17104);
or U29280 (N_29280,N_15634,N_12088);
and U29281 (N_29281,N_15318,N_18669);
or U29282 (N_29282,N_18255,N_14382);
nor U29283 (N_29283,N_18126,N_14376);
nand U29284 (N_29284,N_16545,N_12897);
or U29285 (N_29285,N_18149,N_12132);
and U29286 (N_29286,N_12403,N_19872);
or U29287 (N_29287,N_11969,N_10355);
or U29288 (N_29288,N_17749,N_15974);
nor U29289 (N_29289,N_10562,N_13107);
and U29290 (N_29290,N_18733,N_10662);
and U29291 (N_29291,N_18865,N_17581);
xor U29292 (N_29292,N_17753,N_12926);
or U29293 (N_29293,N_14302,N_18320);
xor U29294 (N_29294,N_18641,N_14734);
and U29295 (N_29295,N_14560,N_19535);
or U29296 (N_29296,N_19858,N_13896);
or U29297 (N_29297,N_18598,N_18047);
nand U29298 (N_29298,N_16827,N_14238);
nor U29299 (N_29299,N_11924,N_18689);
or U29300 (N_29300,N_10221,N_14036);
or U29301 (N_29301,N_17984,N_12821);
nand U29302 (N_29302,N_18979,N_16075);
and U29303 (N_29303,N_14366,N_12296);
or U29304 (N_29304,N_19313,N_13841);
or U29305 (N_29305,N_16729,N_15236);
nor U29306 (N_29306,N_17251,N_16873);
and U29307 (N_29307,N_16513,N_12791);
and U29308 (N_29308,N_12029,N_15673);
nand U29309 (N_29309,N_13155,N_17158);
nand U29310 (N_29310,N_15932,N_10488);
nor U29311 (N_29311,N_10506,N_12996);
and U29312 (N_29312,N_16140,N_15994);
nand U29313 (N_29313,N_11845,N_18380);
nor U29314 (N_29314,N_15128,N_16451);
nand U29315 (N_29315,N_15757,N_19883);
nand U29316 (N_29316,N_18831,N_12011);
or U29317 (N_29317,N_13178,N_15949);
or U29318 (N_29318,N_16168,N_17719);
nand U29319 (N_29319,N_11833,N_16167);
nand U29320 (N_29320,N_12303,N_12729);
nand U29321 (N_29321,N_10866,N_11916);
xor U29322 (N_29322,N_11191,N_12404);
and U29323 (N_29323,N_10731,N_13836);
nor U29324 (N_29324,N_12480,N_11844);
or U29325 (N_29325,N_10320,N_13238);
nor U29326 (N_29326,N_15379,N_18880);
nor U29327 (N_29327,N_10887,N_11651);
and U29328 (N_29328,N_14713,N_19728);
nor U29329 (N_29329,N_19236,N_14187);
nand U29330 (N_29330,N_12135,N_15358);
xnor U29331 (N_29331,N_12147,N_15306);
or U29332 (N_29332,N_19047,N_16733);
or U29333 (N_29333,N_10385,N_12139);
or U29334 (N_29334,N_19431,N_12066);
nand U29335 (N_29335,N_13698,N_13067);
or U29336 (N_29336,N_13792,N_10993);
nor U29337 (N_29337,N_14289,N_11567);
nand U29338 (N_29338,N_14832,N_18185);
or U29339 (N_29339,N_13899,N_15279);
nor U29340 (N_29340,N_17943,N_15098);
nand U29341 (N_29341,N_14808,N_17313);
xor U29342 (N_29342,N_13633,N_11134);
nor U29343 (N_29343,N_18014,N_15665);
nor U29344 (N_29344,N_12446,N_14798);
nand U29345 (N_29345,N_16693,N_19922);
xor U29346 (N_29346,N_11705,N_16627);
nand U29347 (N_29347,N_13015,N_13800);
nand U29348 (N_29348,N_19500,N_12623);
nand U29349 (N_29349,N_16671,N_16769);
or U29350 (N_29350,N_12706,N_19833);
and U29351 (N_29351,N_14421,N_13356);
and U29352 (N_29352,N_11975,N_11445);
nor U29353 (N_29353,N_14804,N_13026);
or U29354 (N_29354,N_17665,N_19378);
or U29355 (N_29355,N_13218,N_12092);
or U29356 (N_29356,N_18092,N_14425);
and U29357 (N_29357,N_15351,N_16461);
nor U29358 (N_29358,N_17986,N_13293);
or U29359 (N_29359,N_19450,N_10520);
or U29360 (N_29360,N_13409,N_11712);
nor U29361 (N_29361,N_17721,N_10086);
nor U29362 (N_29362,N_15606,N_13922);
and U29363 (N_29363,N_14793,N_15091);
and U29364 (N_29364,N_18167,N_12670);
or U29365 (N_29365,N_13273,N_15818);
and U29366 (N_29366,N_12629,N_11949);
xor U29367 (N_29367,N_16144,N_15216);
or U29368 (N_29368,N_11313,N_16295);
nand U29369 (N_29369,N_18302,N_14509);
xnor U29370 (N_29370,N_14385,N_12529);
xor U29371 (N_29371,N_15255,N_14468);
xor U29372 (N_29372,N_15334,N_10353);
nand U29373 (N_29373,N_15884,N_12535);
and U29374 (N_29374,N_18245,N_16093);
nor U29375 (N_29375,N_13659,N_12701);
nand U29376 (N_29376,N_17007,N_18894);
or U29377 (N_29377,N_16766,N_14376);
or U29378 (N_29378,N_13995,N_16039);
nand U29379 (N_29379,N_17935,N_15606);
nor U29380 (N_29380,N_19531,N_14771);
and U29381 (N_29381,N_17901,N_12528);
and U29382 (N_29382,N_15404,N_14851);
nand U29383 (N_29383,N_16665,N_18962);
or U29384 (N_29384,N_18113,N_15555);
or U29385 (N_29385,N_16246,N_16679);
nand U29386 (N_29386,N_14149,N_18804);
nand U29387 (N_29387,N_14648,N_10930);
nand U29388 (N_29388,N_11310,N_15548);
and U29389 (N_29389,N_12306,N_15765);
or U29390 (N_29390,N_15921,N_17655);
nor U29391 (N_29391,N_13762,N_18689);
nor U29392 (N_29392,N_15847,N_16445);
nand U29393 (N_29393,N_16420,N_11062);
or U29394 (N_29394,N_10243,N_15269);
nand U29395 (N_29395,N_18237,N_14136);
and U29396 (N_29396,N_18715,N_19009);
nand U29397 (N_29397,N_16813,N_13142);
nor U29398 (N_29398,N_11537,N_18345);
nand U29399 (N_29399,N_16373,N_10865);
or U29400 (N_29400,N_12032,N_12051);
nor U29401 (N_29401,N_19199,N_18757);
or U29402 (N_29402,N_17489,N_19149);
nor U29403 (N_29403,N_16513,N_14352);
and U29404 (N_29404,N_14649,N_13527);
or U29405 (N_29405,N_11496,N_14043);
and U29406 (N_29406,N_10501,N_10625);
and U29407 (N_29407,N_10315,N_18139);
nand U29408 (N_29408,N_16584,N_12671);
or U29409 (N_29409,N_10324,N_10653);
xor U29410 (N_29410,N_17743,N_18503);
and U29411 (N_29411,N_11608,N_10763);
nand U29412 (N_29412,N_16486,N_13166);
or U29413 (N_29413,N_11503,N_17243);
xor U29414 (N_29414,N_13478,N_18782);
or U29415 (N_29415,N_16222,N_10217);
nor U29416 (N_29416,N_17423,N_14303);
or U29417 (N_29417,N_17860,N_12819);
or U29418 (N_29418,N_15574,N_14032);
or U29419 (N_29419,N_18994,N_14127);
or U29420 (N_29420,N_10479,N_16751);
nand U29421 (N_29421,N_19594,N_12688);
xor U29422 (N_29422,N_14421,N_11408);
or U29423 (N_29423,N_18649,N_10274);
nor U29424 (N_29424,N_16627,N_14237);
or U29425 (N_29425,N_10125,N_10195);
or U29426 (N_29426,N_11887,N_19867);
or U29427 (N_29427,N_17132,N_17021);
or U29428 (N_29428,N_12028,N_19650);
and U29429 (N_29429,N_14501,N_18631);
or U29430 (N_29430,N_18931,N_17535);
nor U29431 (N_29431,N_16000,N_19605);
nand U29432 (N_29432,N_17662,N_12909);
nand U29433 (N_29433,N_18542,N_10595);
or U29434 (N_29434,N_14351,N_18490);
nor U29435 (N_29435,N_12901,N_14622);
nor U29436 (N_29436,N_12024,N_11124);
nand U29437 (N_29437,N_14122,N_19133);
and U29438 (N_29438,N_12356,N_15022);
and U29439 (N_29439,N_16861,N_15087);
nand U29440 (N_29440,N_11739,N_17655);
or U29441 (N_29441,N_17550,N_16882);
nand U29442 (N_29442,N_13693,N_11350);
and U29443 (N_29443,N_13621,N_17790);
or U29444 (N_29444,N_12225,N_11936);
xor U29445 (N_29445,N_15628,N_16315);
and U29446 (N_29446,N_17130,N_19059);
or U29447 (N_29447,N_15319,N_15568);
and U29448 (N_29448,N_17720,N_18893);
nand U29449 (N_29449,N_13809,N_16409);
and U29450 (N_29450,N_12168,N_18310);
and U29451 (N_29451,N_15739,N_15643);
nand U29452 (N_29452,N_12314,N_18026);
nand U29453 (N_29453,N_14677,N_19892);
nor U29454 (N_29454,N_14975,N_10344);
or U29455 (N_29455,N_11362,N_16548);
nor U29456 (N_29456,N_18614,N_14806);
and U29457 (N_29457,N_15785,N_18054);
nand U29458 (N_29458,N_15797,N_13574);
nor U29459 (N_29459,N_10971,N_15026);
xnor U29460 (N_29460,N_11317,N_11250);
nor U29461 (N_29461,N_19913,N_16129);
nand U29462 (N_29462,N_14688,N_10859);
or U29463 (N_29463,N_13959,N_19043);
nand U29464 (N_29464,N_15964,N_13288);
xnor U29465 (N_29465,N_10206,N_17794);
nor U29466 (N_29466,N_10825,N_17935);
or U29467 (N_29467,N_16483,N_10152);
xor U29468 (N_29468,N_15911,N_10508);
or U29469 (N_29469,N_14026,N_19364);
xnor U29470 (N_29470,N_12191,N_14014);
and U29471 (N_29471,N_10397,N_19251);
nor U29472 (N_29472,N_16469,N_12039);
xnor U29473 (N_29473,N_12226,N_12174);
nand U29474 (N_29474,N_10679,N_16574);
nand U29475 (N_29475,N_17337,N_10689);
and U29476 (N_29476,N_13103,N_10890);
nor U29477 (N_29477,N_15870,N_16429);
and U29478 (N_29478,N_14321,N_12473);
and U29479 (N_29479,N_14199,N_12705);
nor U29480 (N_29480,N_17792,N_12917);
nor U29481 (N_29481,N_19945,N_17517);
nor U29482 (N_29482,N_16452,N_10647);
or U29483 (N_29483,N_11102,N_12285);
nand U29484 (N_29484,N_16685,N_10170);
nand U29485 (N_29485,N_19519,N_13875);
nand U29486 (N_29486,N_11927,N_12410);
and U29487 (N_29487,N_10653,N_10777);
or U29488 (N_29488,N_12436,N_10660);
nand U29489 (N_29489,N_19899,N_16058);
nor U29490 (N_29490,N_10150,N_12424);
nor U29491 (N_29491,N_17928,N_19210);
nor U29492 (N_29492,N_16129,N_17309);
and U29493 (N_29493,N_16904,N_18771);
and U29494 (N_29494,N_10048,N_19980);
xor U29495 (N_29495,N_12965,N_10401);
xor U29496 (N_29496,N_11793,N_16431);
or U29497 (N_29497,N_15220,N_17133);
nor U29498 (N_29498,N_13628,N_11590);
and U29499 (N_29499,N_19560,N_15778);
and U29500 (N_29500,N_13698,N_17767);
xnor U29501 (N_29501,N_12569,N_11166);
xnor U29502 (N_29502,N_15651,N_14120);
nor U29503 (N_29503,N_11378,N_17448);
and U29504 (N_29504,N_11910,N_13453);
and U29505 (N_29505,N_13970,N_10459);
nor U29506 (N_29506,N_12331,N_12715);
nor U29507 (N_29507,N_19171,N_17198);
xor U29508 (N_29508,N_18202,N_11332);
or U29509 (N_29509,N_14237,N_10102);
and U29510 (N_29510,N_12625,N_15777);
xnor U29511 (N_29511,N_10589,N_10162);
or U29512 (N_29512,N_18917,N_18813);
nand U29513 (N_29513,N_11717,N_12145);
nand U29514 (N_29514,N_15248,N_11287);
nor U29515 (N_29515,N_10780,N_16745);
or U29516 (N_29516,N_14389,N_19174);
nor U29517 (N_29517,N_17809,N_12100);
or U29518 (N_29518,N_18040,N_18933);
nor U29519 (N_29519,N_15964,N_15129);
xor U29520 (N_29520,N_19288,N_17141);
and U29521 (N_29521,N_11258,N_15608);
and U29522 (N_29522,N_14722,N_18150);
and U29523 (N_29523,N_13234,N_12388);
and U29524 (N_29524,N_18358,N_16604);
xnor U29525 (N_29525,N_17331,N_17271);
or U29526 (N_29526,N_18996,N_12516);
nand U29527 (N_29527,N_13156,N_17971);
nor U29528 (N_29528,N_12167,N_12681);
or U29529 (N_29529,N_13579,N_13773);
and U29530 (N_29530,N_19182,N_17393);
nor U29531 (N_29531,N_14087,N_14313);
and U29532 (N_29532,N_17208,N_15842);
or U29533 (N_29533,N_15489,N_14311);
or U29534 (N_29534,N_18436,N_15933);
and U29535 (N_29535,N_18709,N_13500);
or U29536 (N_29536,N_18872,N_14072);
nor U29537 (N_29537,N_10913,N_13061);
or U29538 (N_29538,N_15442,N_12560);
xnor U29539 (N_29539,N_15239,N_11899);
and U29540 (N_29540,N_17757,N_13221);
nor U29541 (N_29541,N_12769,N_10950);
or U29542 (N_29542,N_13552,N_17097);
xnor U29543 (N_29543,N_11162,N_14131);
nor U29544 (N_29544,N_12316,N_15221);
nand U29545 (N_29545,N_11208,N_15963);
nand U29546 (N_29546,N_16380,N_10956);
and U29547 (N_29547,N_19414,N_19968);
nor U29548 (N_29548,N_19312,N_16906);
or U29549 (N_29549,N_12642,N_14148);
and U29550 (N_29550,N_18450,N_14107);
and U29551 (N_29551,N_18594,N_16064);
or U29552 (N_29552,N_19918,N_13933);
nor U29553 (N_29553,N_15925,N_12327);
or U29554 (N_29554,N_15807,N_15843);
xor U29555 (N_29555,N_15143,N_14495);
xnor U29556 (N_29556,N_18070,N_17445);
xor U29557 (N_29557,N_14806,N_12235);
nand U29558 (N_29558,N_11233,N_10660);
or U29559 (N_29559,N_11771,N_16677);
and U29560 (N_29560,N_10321,N_15940);
and U29561 (N_29561,N_16027,N_11692);
and U29562 (N_29562,N_19802,N_12421);
nor U29563 (N_29563,N_19770,N_11882);
xnor U29564 (N_29564,N_16997,N_11147);
nand U29565 (N_29565,N_16680,N_11261);
nand U29566 (N_29566,N_15196,N_17533);
or U29567 (N_29567,N_12721,N_12368);
or U29568 (N_29568,N_19256,N_17346);
nor U29569 (N_29569,N_14579,N_12275);
or U29570 (N_29570,N_17052,N_10721);
and U29571 (N_29571,N_18836,N_10678);
nand U29572 (N_29572,N_15235,N_16248);
and U29573 (N_29573,N_18686,N_19367);
xnor U29574 (N_29574,N_18722,N_11801);
nand U29575 (N_29575,N_19692,N_18820);
and U29576 (N_29576,N_11379,N_10567);
and U29577 (N_29577,N_10155,N_12464);
or U29578 (N_29578,N_13765,N_18782);
xnor U29579 (N_29579,N_18868,N_17856);
and U29580 (N_29580,N_18384,N_13310);
nand U29581 (N_29581,N_15194,N_11381);
nor U29582 (N_29582,N_17258,N_19627);
and U29583 (N_29583,N_10833,N_15892);
nor U29584 (N_29584,N_14803,N_14782);
and U29585 (N_29585,N_19104,N_17000);
and U29586 (N_29586,N_16632,N_13956);
nor U29587 (N_29587,N_18729,N_17061);
nor U29588 (N_29588,N_18728,N_10327);
nor U29589 (N_29589,N_14084,N_14942);
and U29590 (N_29590,N_18188,N_10488);
nand U29591 (N_29591,N_14049,N_13639);
and U29592 (N_29592,N_14613,N_17311);
nand U29593 (N_29593,N_15114,N_10337);
or U29594 (N_29594,N_12921,N_15674);
nor U29595 (N_29595,N_12509,N_19111);
or U29596 (N_29596,N_11379,N_14015);
nor U29597 (N_29597,N_11868,N_14817);
or U29598 (N_29598,N_16034,N_14802);
and U29599 (N_29599,N_17189,N_13368);
and U29600 (N_29600,N_10487,N_10991);
nor U29601 (N_29601,N_19319,N_12017);
nand U29602 (N_29602,N_11518,N_13118);
or U29603 (N_29603,N_16363,N_18403);
nor U29604 (N_29604,N_12041,N_15130);
xor U29605 (N_29605,N_10295,N_10141);
nand U29606 (N_29606,N_16803,N_16792);
nor U29607 (N_29607,N_17181,N_11713);
and U29608 (N_29608,N_18580,N_17246);
and U29609 (N_29609,N_16278,N_10934);
or U29610 (N_29610,N_16045,N_13625);
nor U29611 (N_29611,N_15750,N_14248);
xnor U29612 (N_29612,N_14889,N_11173);
nand U29613 (N_29613,N_12404,N_19057);
nor U29614 (N_29614,N_17432,N_14055);
nand U29615 (N_29615,N_12484,N_12094);
and U29616 (N_29616,N_10795,N_11916);
and U29617 (N_29617,N_18863,N_19535);
and U29618 (N_29618,N_10001,N_17162);
nor U29619 (N_29619,N_18295,N_15540);
and U29620 (N_29620,N_16083,N_15109);
nor U29621 (N_29621,N_13428,N_12412);
nor U29622 (N_29622,N_10130,N_18393);
and U29623 (N_29623,N_16564,N_11091);
or U29624 (N_29624,N_18070,N_19633);
nand U29625 (N_29625,N_12342,N_12259);
and U29626 (N_29626,N_10009,N_12613);
xnor U29627 (N_29627,N_17112,N_13291);
and U29628 (N_29628,N_16353,N_17409);
and U29629 (N_29629,N_11815,N_12127);
and U29630 (N_29630,N_14289,N_16719);
xnor U29631 (N_29631,N_16432,N_19772);
and U29632 (N_29632,N_14990,N_10424);
nor U29633 (N_29633,N_19375,N_14858);
nand U29634 (N_29634,N_19385,N_10436);
nand U29635 (N_29635,N_10547,N_17183);
nand U29636 (N_29636,N_18497,N_12436);
nor U29637 (N_29637,N_17112,N_12213);
xnor U29638 (N_29638,N_15500,N_16750);
and U29639 (N_29639,N_11513,N_11750);
and U29640 (N_29640,N_10542,N_18349);
nor U29641 (N_29641,N_15495,N_11881);
nor U29642 (N_29642,N_15922,N_17897);
nand U29643 (N_29643,N_13722,N_13309);
xnor U29644 (N_29644,N_15989,N_17819);
xor U29645 (N_29645,N_14015,N_18500);
xor U29646 (N_29646,N_16359,N_14815);
xnor U29647 (N_29647,N_18134,N_13011);
nand U29648 (N_29648,N_19836,N_12487);
nand U29649 (N_29649,N_11738,N_11516);
nor U29650 (N_29650,N_15616,N_19910);
or U29651 (N_29651,N_12963,N_12820);
and U29652 (N_29652,N_18770,N_19480);
or U29653 (N_29653,N_15804,N_17844);
xnor U29654 (N_29654,N_12980,N_19029);
nor U29655 (N_29655,N_18896,N_18972);
nand U29656 (N_29656,N_17070,N_15840);
nor U29657 (N_29657,N_10748,N_13418);
nand U29658 (N_29658,N_19068,N_14750);
nand U29659 (N_29659,N_18562,N_13036);
nand U29660 (N_29660,N_10173,N_14771);
xnor U29661 (N_29661,N_17064,N_15263);
xor U29662 (N_29662,N_18917,N_18181);
and U29663 (N_29663,N_18706,N_14680);
nand U29664 (N_29664,N_14355,N_11044);
nor U29665 (N_29665,N_16981,N_12896);
or U29666 (N_29666,N_16620,N_17699);
or U29667 (N_29667,N_14564,N_19250);
nor U29668 (N_29668,N_14231,N_15988);
nand U29669 (N_29669,N_16141,N_11373);
nand U29670 (N_29670,N_13054,N_16044);
nand U29671 (N_29671,N_16711,N_12864);
nand U29672 (N_29672,N_17941,N_10816);
and U29673 (N_29673,N_16683,N_14706);
nand U29674 (N_29674,N_11992,N_13099);
xor U29675 (N_29675,N_15448,N_19325);
or U29676 (N_29676,N_17919,N_13518);
xnor U29677 (N_29677,N_14635,N_14596);
nand U29678 (N_29678,N_15754,N_12752);
and U29679 (N_29679,N_16910,N_17934);
nor U29680 (N_29680,N_19639,N_16121);
or U29681 (N_29681,N_12715,N_12538);
xnor U29682 (N_29682,N_12805,N_18436);
nor U29683 (N_29683,N_10580,N_12909);
nor U29684 (N_29684,N_14036,N_14407);
and U29685 (N_29685,N_15119,N_19774);
nand U29686 (N_29686,N_12880,N_16479);
or U29687 (N_29687,N_17015,N_15919);
or U29688 (N_29688,N_16304,N_10709);
nor U29689 (N_29689,N_11676,N_15730);
nor U29690 (N_29690,N_15563,N_16302);
xnor U29691 (N_29691,N_14902,N_15052);
or U29692 (N_29692,N_12094,N_16494);
xor U29693 (N_29693,N_13649,N_12913);
and U29694 (N_29694,N_15037,N_19376);
or U29695 (N_29695,N_11006,N_14966);
and U29696 (N_29696,N_14175,N_10658);
xnor U29697 (N_29697,N_10321,N_18034);
or U29698 (N_29698,N_10541,N_11139);
xnor U29699 (N_29699,N_15490,N_14615);
nor U29700 (N_29700,N_17909,N_16153);
nor U29701 (N_29701,N_17479,N_15210);
or U29702 (N_29702,N_19985,N_13963);
and U29703 (N_29703,N_17512,N_10855);
nand U29704 (N_29704,N_19965,N_12673);
xor U29705 (N_29705,N_15042,N_19002);
nand U29706 (N_29706,N_17911,N_10316);
or U29707 (N_29707,N_19734,N_18827);
and U29708 (N_29708,N_10727,N_10814);
nand U29709 (N_29709,N_12498,N_13403);
and U29710 (N_29710,N_10900,N_18210);
or U29711 (N_29711,N_19415,N_19692);
and U29712 (N_29712,N_10537,N_15554);
xor U29713 (N_29713,N_11407,N_13855);
or U29714 (N_29714,N_19330,N_16493);
nor U29715 (N_29715,N_17203,N_13697);
or U29716 (N_29716,N_17489,N_18206);
xnor U29717 (N_29717,N_15776,N_16398);
and U29718 (N_29718,N_10527,N_12175);
nand U29719 (N_29719,N_17758,N_14227);
or U29720 (N_29720,N_13014,N_16749);
and U29721 (N_29721,N_11591,N_13493);
nand U29722 (N_29722,N_16191,N_12018);
or U29723 (N_29723,N_11239,N_12634);
nand U29724 (N_29724,N_17508,N_13849);
nor U29725 (N_29725,N_13655,N_13358);
and U29726 (N_29726,N_10457,N_16967);
and U29727 (N_29727,N_10060,N_17859);
nor U29728 (N_29728,N_16427,N_15294);
nand U29729 (N_29729,N_18914,N_18783);
and U29730 (N_29730,N_10137,N_11527);
xor U29731 (N_29731,N_11225,N_16255);
and U29732 (N_29732,N_11824,N_15303);
and U29733 (N_29733,N_13733,N_15932);
or U29734 (N_29734,N_12695,N_11943);
xor U29735 (N_29735,N_11617,N_15070);
or U29736 (N_29736,N_11501,N_19160);
and U29737 (N_29737,N_19127,N_15973);
or U29738 (N_29738,N_19353,N_14520);
and U29739 (N_29739,N_10009,N_12599);
and U29740 (N_29740,N_10833,N_12206);
nand U29741 (N_29741,N_18169,N_18736);
and U29742 (N_29742,N_12833,N_10427);
xor U29743 (N_29743,N_11533,N_14765);
or U29744 (N_29744,N_16293,N_19808);
and U29745 (N_29745,N_19408,N_12785);
nand U29746 (N_29746,N_14827,N_19994);
nor U29747 (N_29747,N_16000,N_19292);
and U29748 (N_29748,N_18212,N_18734);
nor U29749 (N_29749,N_16074,N_12351);
nor U29750 (N_29750,N_15433,N_13371);
nor U29751 (N_29751,N_17747,N_19038);
nor U29752 (N_29752,N_16431,N_14567);
and U29753 (N_29753,N_15563,N_11655);
or U29754 (N_29754,N_12845,N_17995);
nor U29755 (N_29755,N_10569,N_10548);
and U29756 (N_29756,N_16702,N_19693);
nor U29757 (N_29757,N_16645,N_16002);
or U29758 (N_29758,N_18626,N_13364);
or U29759 (N_29759,N_18010,N_18059);
or U29760 (N_29760,N_15259,N_14885);
xor U29761 (N_29761,N_18095,N_18471);
or U29762 (N_29762,N_16288,N_16672);
or U29763 (N_29763,N_10183,N_15915);
nor U29764 (N_29764,N_18666,N_13605);
and U29765 (N_29765,N_18171,N_18964);
or U29766 (N_29766,N_19384,N_16723);
nor U29767 (N_29767,N_10210,N_19062);
or U29768 (N_29768,N_12330,N_11524);
or U29769 (N_29769,N_10485,N_18652);
nand U29770 (N_29770,N_13321,N_15001);
nor U29771 (N_29771,N_11023,N_10114);
or U29772 (N_29772,N_17862,N_10053);
or U29773 (N_29773,N_16604,N_15286);
and U29774 (N_29774,N_15514,N_18203);
or U29775 (N_29775,N_18098,N_10758);
and U29776 (N_29776,N_10750,N_19930);
or U29777 (N_29777,N_11793,N_13429);
and U29778 (N_29778,N_19926,N_10103);
nor U29779 (N_29779,N_15357,N_13577);
or U29780 (N_29780,N_16806,N_17238);
xor U29781 (N_29781,N_16689,N_13211);
nand U29782 (N_29782,N_18388,N_12682);
and U29783 (N_29783,N_17600,N_15214);
and U29784 (N_29784,N_15493,N_10766);
and U29785 (N_29785,N_13318,N_15197);
or U29786 (N_29786,N_15948,N_15629);
nor U29787 (N_29787,N_14847,N_11767);
nor U29788 (N_29788,N_16518,N_10329);
nor U29789 (N_29789,N_13447,N_10287);
and U29790 (N_29790,N_14578,N_12059);
xnor U29791 (N_29791,N_17569,N_10051);
and U29792 (N_29792,N_12344,N_19712);
and U29793 (N_29793,N_17531,N_14937);
and U29794 (N_29794,N_11073,N_14114);
and U29795 (N_29795,N_13131,N_13613);
nor U29796 (N_29796,N_19307,N_12295);
or U29797 (N_29797,N_10028,N_15289);
xor U29798 (N_29798,N_11905,N_14510);
xor U29799 (N_29799,N_17914,N_13773);
and U29800 (N_29800,N_19940,N_18071);
or U29801 (N_29801,N_19590,N_10172);
or U29802 (N_29802,N_17538,N_18420);
or U29803 (N_29803,N_16901,N_13087);
and U29804 (N_29804,N_13714,N_12035);
xnor U29805 (N_29805,N_10613,N_19858);
or U29806 (N_29806,N_15077,N_12355);
or U29807 (N_29807,N_14989,N_12341);
nand U29808 (N_29808,N_14894,N_13347);
nor U29809 (N_29809,N_15930,N_16710);
nor U29810 (N_29810,N_19033,N_14569);
and U29811 (N_29811,N_13682,N_19679);
xnor U29812 (N_29812,N_18703,N_11428);
nand U29813 (N_29813,N_15889,N_12839);
xnor U29814 (N_29814,N_15781,N_17847);
nand U29815 (N_29815,N_17756,N_14430);
nor U29816 (N_29816,N_12092,N_18272);
and U29817 (N_29817,N_12439,N_14583);
nor U29818 (N_29818,N_11518,N_14300);
nand U29819 (N_29819,N_17697,N_12369);
nand U29820 (N_29820,N_14161,N_15121);
and U29821 (N_29821,N_10872,N_14201);
nor U29822 (N_29822,N_10175,N_16869);
and U29823 (N_29823,N_10604,N_18111);
nor U29824 (N_29824,N_19768,N_18022);
xnor U29825 (N_29825,N_13679,N_11351);
nand U29826 (N_29826,N_18377,N_10599);
nor U29827 (N_29827,N_16368,N_18358);
nand U29828 (N_29828,N_12469,N_13745);
or U29829 (N_29829,N_16261,N_14226);
or U29830 (N_29830,N_12793,N_14344);
and U29831 (N_29831,N_13926,N_19664);
nor U29832 (N_29832,N_14512,N_10961);
or U29833 (N_29833,N_10753,N_18005);
and U29834 (N_29834,N_19036,N_11378);
xnor U29835 (N_29835,N_14968,N_16807);
and U29836 (N_29836,N_18226,N_16782);
nand U29837 (N_29837,N_19623,N_11150);
nand U29838 (N_29838,N_13809,N_18559);
nand U29839 (N_29839,N_16655,N_17631);
nor U29840 (N_29840,N_15178,N_15650);
xor U29841 (N_29841,N_17877,N_10720);
or U29842 (N_29842,N_16061,N_12338);
nor U29843 (N_29843,N_14285,N_19771);
nor U29844 (N_29844,N_11788,N_16329);
and U29845 (N_29845,N_17344,N_19614);
nor U29846 (N_29846,N_12250,N_11304);
nand U29847 (N_29847,N_16468,N_12182);
and U29848 (N_29848,N_10572,N_15543);
and U29849 (N_29849,N_11195,N_14268);
and U29850 (N_29850,N_19826,N_17796);
nor U29851 (N_29851,N_19445,N_14557);
xnor U29852 (N_29852,N_10663,N_15611);
nand U29853 (N_29853,N_13136,N_14676);
nor U29854 (N_29854,N_10227,N_19920);
nand U29855 (N_29855,N_13291,N_18450);
and U29856 (N_29856,N_16973,N_19570);
nand U29857 (N_29857,N_14765,N_14925);
nor U29858 (N_29858,N_13433,N_13642);
nand U29859 (N_29859,N_19568,N_19412);
and U29860 (N_29860,N_15785,N_16137);
or U29861 (N_29861,N_15379,N_18501);
or U29862 (N_29862,N_16493,N_13091);
or U29863 (N_29863,N_12498,N_11872);
nor U29864 (N_29864,N_17418,N_10620);
nor U29865 (N_29865,N_12847,N_13428);
nor U29866 (N_29866,N_19089,N_14001);
nor U29867 (N_29867,N_19174,N_10719);
or U29868 (N_29868,N_17702,N_16995);
nor U29869 (N_29869,N_18818,N_13054);
or U29870 (N_29870,N_17207,N_18303);
nor U29871 (N_29871,N_19819,N_19522);
or U29872 (N_29872,N_12190,N_14478);
xor U29873 (N_29873,N_14966,N_18924);
xnor U29874 (N_29874,N_10882,N_15580);
nand U29875 (N_29875,N_19866,N_18065);
and U29876 (N_29876,N_12001,N_10522);
or U29877 (N_29877,N_17189,N_18815);
or U29878 (N_29878,N_12127,N_12832);
and U29879 (N_29879,N_17353,N_18965);
or U29880 (N_29880,N_16546,N_19475);
or U29881 (N_29881,N_17988,N_11151);
and U29882 (N_29882,N_14730,N_16305);
nand U29883 (N_29883,N_17348,N_12849);
nand U29884 (N_29884,N_13684,N_14542);
and U29885 (N_29885,N_14855,N_11192);
nor U29886 (N_29886,N_10050,N_13176);
nor U29887 (N_29887,N_13606,N_11430);
or U29888 (N_29888,N_17033,N_17337);
nor U29889 (N_29889,N_17432,N_17245);
nor U29890 (N_29890,N_12611,N_11194);
nand U29891 (N_29891,N_11194,N_14295);
nor U29892 (N_29892,N_12539,N_19967);
or U29893 (N_29893,N_16637,N_10050);
and U29894 (N_29894,N_19219,N_18285);
nand U29895 (N_29895,N_13473,N_16894);
nor U29896 (N_29896,N_12232,N_11117);
or U29897 (N_29897,N_13336,N_19072);
nor U29898 (N_29898,N_16770,N_16352);
nand U29899 (N_29899,N_15244,N_16114);
nor U29900 (N_29900,N_15402,N_10322);
or U29901 (N_29901,N_18080,N_18833);
nand U29902 (N_29902,N_11024,N_18025);
nor U29903 (N_29903,N_13062,N_11998);
nor U29904 (N_29904,N_14091,N_14035);
nand U29905 (N_29905,N_14727,N_14704);
or U29906 (N_29906,N_10766,N_10189);
nand U29907 (N_29907,N_12666,N_18925);
or U29908 (N_29908,N_17512,N_18717);
nor U29909 (N_29909,N_16255,N_18052);
nand U29910 (N_29910,N_18843,N_13350);
nand U29911 (N_29911,N_18597,N_12196);
or U29912 (N_29912,N_18688,N_14255);
nor U29913 (N_29913,N_12158,N_11734);
nand U29914 (N_29914,N_19390,N_16675);
and U29915 (N_29915,N_14856,N_10142);
or U29916 (N_29916,N_15392,N_11566);
nor U29917 (N_29917,N_17931,N_15722);
xor U29918 (N_29918,N_18409,N_13270);
nand U29919 (N_29919,N_15727,N_16748);
xnor U29920 (N_29920,N_16250,N_17252);
nor U29921 (N_29921,N_11112,N_16798);
and U29922 (N_29922,N_13639,N_18404);
xor U29923 (N_29923,N_19680,N_13010);
xnor U29924 (N_29924,N_11425,N_10827);
or U29925 (N_29925,N_19332,N_18780);
xor U29926 (N_29926,N_11285,N_11561);
and U29927 (N_29927,N_10543,N_12715);
or U29928 (N_29928,N_11780,N_14310);
or U29929 (N_29929,N_17877,N_12935);
and U29930 (N_29930,N_18280,N_16073);
xnor U29931 (N_29931,N_14879,N_16597);
or U29932 (N_29932,N_15743,N_17455);
and U29933 (N_29933,N_18864,N_14371);
or U29934 (N_29934,N_18808,N_10123);
and U29935 (N_29935,N_19636,N_10568);
nand U29936 (N_29936,N_18532,N_18891);
nand U29937 (N_29937,N_19188,N_16600);
or U29938 (N_29938,N_17591,N_16188);
xnor U29939 (N_29939,N_13497,N_17435);
nor U29940 (N_29940,N_11017,N_10833);
and U29941 (N_29941,N_19387,N_19294);
or U29942 (N_29942,N_15005,N_11153);
xor U29943 (N_29943,N_11079,N_12650);
nor U29944 (N_29944,N_18465,N_17142);
xnor U29945 (N_29945,N_14713,N_10159);
nor U29946 (N_29946,N_18088,N_10762);
xnor U29947 (N_29947,N_14297,N_16351);
nor U29948 (N_29948,N_17378,N_15189);
xnor U29949 (N_29949,N_13049,N_15883);
or U29950 (N_29950,N_11510,N_19020);
and U29951 (N_29951,N_12472,N_16042);
and U29952 (N_29952,N_10595,N_18280);
nor U29953 (N_29953,N_10831,N_16916);
or U29954 (N_29954,N_18036,N_14347);
and U29955 (N_29955,N_18338,N_11326);
nand U29956 (N_29956,N_10698,N_13377);
or U29957 (N_29957,N_18857,N_17579);
or U29958 (N_29958,N_13551,N_13746);
and U29959 (N_29959,N_12599,N_15198);
nor U29960 (N_29960,N_17635,N_16285);
nand U29961 (N_29961,N_15951,N_11090);
or U29962 (N_29962,N_19286,N_16299);
xnor U29963 (N_29963,N_17620,N_13007);
nand U29964 (N_29964,N_17900,N_16577);
nand U29965 (N_29965,N_14498,N_14122);
or U29966 (N_29966,N_12774,N_19697);
nand U29967 (N_29967,N_16417,N_15927);
or U29968 (N_29968,N_13214,N_17774);
nand U29969 (N_29969,N_17958,N_18157);
or U29970 (N_29970,N_15800,N_16053);
nand U29971 (N_29971,N_13719,N_16828);
and U29972 (N_29972,N_18023,N_15073);
xor U29973 (N_29973,N_17688,N_18794);
nor U29974 (N_29974,N_15642,N_11403);
nor U29975 (N_29975,N_15369,N_13031);
nor U29976 (N_29976,N_11273,N_17818);
nor U29977 (N_29977,N_16119,N_15535);
and U29978 (N_29978,N_11225,N_19049);
or U29979 (N_29979,N_12969,N_18353);
nand U29980 (N_29980,N_13842,N_18562);
and U29981 (N_29981,N_19186,N_17966);
nand U29982 (N_29982,N_13083,N_17758);
nand U29983 (N_29983,N_17159,N_12806);
or U29984 (N_29984,N_10527,N_18512);
nand U29985 (N_29985,N_19403,N_12930);
and U29986 (N_29986,N_18814,N_17199);
or U29987 (N_29987,N_19240,N_14642);
nor U29988 (N_29988,N_11093,N_14942);
xor U29989 (N_29989,N_14321,N_16540);
or U29990 (N_29990,N_15378,N_14015);
and U29991 (N_29991,N_17831,N_18055);
xnor U29992 (N_29992,N_13352,N_13693);
nor U29993 (N_29993,N_14038,N_13216);
or U29994 (N_29994,N_18517,N_12387);
and U29995 (N_29995,N_13544,N_10401);
nor U29996 (N_29996,N_19293,N_15122);
and U29997 (N_29997,N_13827,N_16318);
nand U29998 (N_29998,N_18811,N_10651);
and U29999 (N_29999,N_11904,N_19495);
nand U30000 (N_30000,N_20864,N_24143);
nor U30001 (N_30001,N_22582,N_22005);
xor U30002 (N_30002,N_26099,N_23740);
xor U30003 (N_30003,N_24031,N_29236);
nand U30004 (N_30004,N_29065,N_25213);
and U30005 (N_30005,N_21989,N_25730);
or U30006 (N_30006,N_29959,N_22464);
nand U30007 (N_30007,N_27348,N_20777);
nand U30008 (N_30008,N_24771,N_23592);
nand U30009 (N_30009,N_24321,N_24435);
and U30010 (N_30010,N_28346,N_26441);
nor U30011 (N_30011,N_25170,N_24171);
or U30012 (N_30012,N_20394,N_29406);
or U30013 (N_30013,N_22669,N_23892);
nand U30014 (N_30014,N_26855,N_26561);
nor U30015 (N_30015,N_25562,N_22156);
nor U30016 (N_30016,N_26872,N_21173);
and U30017 (N_30017,N_22419,N_23824);
nand U30018 (N_30018,N_27048,N_27550);
or U30019 (N_30019,N_28895,N_27758);
and U30020 (N_30020,N_28562,N_20423);
nor U30021 (N_30021,N_26152,N_22110);
and U30022 (N_30022,N_28422,N_26764);
xnor U30023 (N_30023,N_26058,N_26140);
or U30024 (N_30024,N_29573,N_20428);
nor U30025 (N_30025,N_22345,N_28545);
xor U30026 (N_30026,N_20845,N_25135);
or U30027 (N_30027,N_27116,N_24496);
nor U30028 (N_30028,N_21135,N_25534);
nor U30029 (N_30029,N_23861,N_22214);
and U30030 (N_30030,N_25846,N_28388);
nand U30031 (N_30031,N_25982,N_20364);
nand U30032 (N_30032,N_20384,N_25996);
or U30033 (N_30033,N_26292,N_24599);
or U30034 (N_30034,N_27586,N_21198);
or U30035 (N_30035,N_25939,N_29451);
or U30036 (N_30036,N_21064,N_29498);
and U30037 (N_30037,N_28696,N_24233);
or U30038 (N_30038,N_29361,N_23919);
nand U30039 (N_30039,N_20708,N_20935);
and U30040 (N_30040,N_24533,N_20096);
xnor U30041 (N_30041,N_26647,N_22797);
xnor U30042 (N_30042,N_29612,N_25073);
and U30043 (N_30043,N_22097,N_28808);
or U30044 (N_30044,N_21971,N_25734);
nor U30045 (N_30045,N_27402,N_28238);
xnor U30046 (N_30046,N_23601,N_23034);
or U30047 (N_30047,N_24107,N_26601);
xnor U30048 (N_30048,N_24932,N_21422);
and U30049 (N_30049,N_22776,N_25098);
or U30050 (N_30050,N_23556,N_22642);
nor U30051 (N_30051,N_26911,N_29393);
nor U30052 (N_30052,N_29534,N_26821);
nor U30053 (N_30053,N_25858,N_25684);
or U30054 (N_30054,N_25610,N_23220);
nand U30055 (N_30055,N_28482,N_23706);
or U30056 (N_30056,N_25201,N_21102);
nor U30057 (N_30057,N_25943,N_23090);
xor U30058 (N_30058,N_25778,N_20284);
or U30059 (N_30059,N_21851,N_23494);
nand U30060 (N_30060,N_24073,N_27946);
and U30061 (N_30061,N_29006,N_27942);
nor U30062 (N_30062,N_21654,N_28927);
nor U30063 (N_30063,N_23149,N_22966);
or U30064 (N_30064,N_24589,N_29033);
nor U30065 (N_30065,N_22268,N_25083);
nand U30066 (N_30066,N_22896,N_23820);
nor U30067 (N_30067,N_20083,N_27441);
nor U30068 (N_30068,N_23839,N_27042);
or U30069 (N_30069,N_26384,N_28530);
and U30070 (N_30070,N_20163,N_24736);
xor U30071 (N_30071,N_24060,N_26507);
nor U30072 (N_30072,N_27807,N_25782);
nand U30073 (N_30073,N_29081,N_26347);
nand U30074 (N_30074,N_29435,N_22031);
nor U30075 (N_30075,N_22876,N_29003);
nand U30076 (N_30076,N_26961,N_20258);
nand U30077 (N_30077,N_29744,N_24817);
and U30078 (N_30078,N_26592,N_23719);
and U30079 (N_30079,N_20850,N_29248);
or U30080 (N_30080,N_23735,N_23732);
or U30081 (N_30081,N_22518,N_28386);
nand U30082 (N_30082,N_21900,N_20216);
nor U30083 (N_30083,N_21044,N_25474);
and U30084 (N_30084,N_25513,N_21586);
and U30085 (N_30085,N_28431,N_27543);
nor U30086 (N_30086,N_24306,N_24159);
nor U30087 (N_30087,N_22880,N_21000);
or U30088 (N_30088,N_23041,N_28925);
or U30089 (N_30089,N_24330,N_22298);
nand U30090 (N_30090,N_27400,N_20797);
nor U30091 (N_30091,N_26653,N_27151);
nor U30092 (N_30092,N_27768,N_21772);
or U30093 (N_30093,N_25161,N_24219);
and U30094 (N_30094,N_25922,N_27983);
nand U30095 (N_30095,N_24680,N_26915);
nand U30096 (N_30096,N_27438,N_29778);
or U30097 (N_30097,N_28838,N_24299);
nand U30098 (N_30098,N_25061,N_22159);
xor U30099 (N_30099,N_26771,N_29490);
and U30100 (N_30100,N_29019,N_22125);
nor U30101 (N_30101,N_22674,N_26499);
and U30102 (N_30102,N_27347,N_22833);
xnor U30103 (N_30103,N_23874,N_21888);
nand U30104 (N_30104,N_27104,N_23607);
or U30105 (N_30105,N_20499,N_26382);
nand U30106 (N_30106,N_27740,N_28297);
and U30107 (N_30107,N_29521,N_27839);
nand U30108 (N_30108,N_20734,N_23176);
and U30109 (N_30109,N_20771,N_20564);
nand U30110 (N_30110,N_22272,N_29815);
or U30111 (N_30111,N_28789,N_28986);
nor U30112 (N_30112,N_20370,N_22150);
xor U30113 (N_30113,N_24075,N_25623);
or U30114 (N_30114,N_22511,N_28836);
and U30115 (N_30115,N_23665,N_20642);
and U30116 (N_30116,N_21860,N_25791);
or U30117 (N_30117,N_28210,N_22531);
and U30118 (N_30118,N_23903,N_28662);
and U30119 (N_30119,N_29888,N_28454);
or U30120 (N_30120,N_23125,N_27761);
and U30121 (N_30121,N_24058,N_24994);
nor U30122 (N_30122,N_20086,N_22057);
and U30123 (N_30123,N_24696,N_24510);
xnor U30124 (N_30124,N_22229,N_21255);
and U30125 (N_30125,N_25501,N_26097);
nand U30126 (N_30126,N_29046,N_26091);
nand U30127 (N_30127,N_22529,N_28471);
and U30128 (N_30128,N_25404,N_25181);
or U30129 (N_30129,N_27567,N_24894);
or U30130 (N_30130,N_27140,N_29314);
or U30131 (N_30131,N_24838,N_24292);
or U30132 (N_30132,N_26278,N_20616);
nor U30133 (N_30133,N_23274,N_29224);
nor U30134 (N_30134,N_26583,N_23539);
and U30135 (N_30135,N_23112,N_28244);
xor U30136 (N_30136,N_27650,N_23777);
or U30137 (N_30137,N_21861,N_23587);
xor U30138 (N_30138,N_28447,N_29858);
nor U30139 (N_30139,N_23760,N_26526);
nand U30140 (N_30140,N_23875,N_26195);
and U30141 (N_30141,N_23517,N_29769);
and U30142 (N_30142,N_24478,N_23991);
and U30143 (N_30143,N_28220,N_24447);
or U30144 (N_30144,N_27606,N_26324);
nand U30145 (N_30145,N_29589,N_23940);
nor U30146 (N_30146,N_28743,N_26669);
nand U30147 (N_30147,N_25936,N_26129);
and U30148 (N_30148,N_22019,N_23351);
nor U30149 (N_30149,N_23202,N_26286);
xor U30150 (N_30150,N_25882,N_28682);
or U30151 (N_30151,N_29975,N_21548);
nor U30152 (N_30152,N_21870,N_28164);
or U30153 (N_30153,N_26831,N_23636);
nand U30154 (N_30154,N_20154,N_22738);
nor U30155 (N_30155,N_26030,N_24236);
nor U30156 (N_30156,N_23158,N_24432);
nor U30157 (N_30157,N_24032,N_29917);
or U30158 (N_30158,N_20871,N_21645);
nand U30159 (N_30159,N_21566,N_23217);
and U30160 (N_30160,N_25875,N_22020);
or U30161 (N_30161,N_22842,N_21287);
nor U30162 (N_30162,N_23659,N_24665);
nor U30163 (N_30163,N_21349,N_25008);
or U30164 (N_30164,N_26791,N_23431);
or U30165 (N_30165,N_28401,N_26790);
nor U30166 (N_30166,N_24551,N_28765);
nand U30167 (N_30167,N_29181,N_21774);
or U30168 (N_30168,N_23726,N_27244);
nor U30169 (N_30169,N_28189,N_28661);
nor U30170 (N_30170,N_26722,N_21823);
nand U30171 (N_30171,N_26267,N_24747);
or U30172 (N_30172,N_25461,N_28591);
and U30173 (N_30173,N_21767,N_28292);
or U30174 (N_30174,N_20013,N_20067);
and U30175 (N_30175,N_26355,N_21021);
nand U30176 (N_30176,N_20140,N_27082);
nor U30177 (N_30177,N_27050,N_22258);
and U30178 (N_30178,N_29558,N_25191);
nor U30179 (N_30179,N_29556,N_28116);
xnor U30180 (N_30180,N_23397,N_25207);
nand U30181 (N_30181,N_22651,N_26554);
nor U30182 (N_30182,N_25374,N_28278);
nor U30183 (N_30183,N_20362,N_23260);
and U30184 (N_30184,N_27750,N_24459);
and U30185 (N_30185,N_24648,N_23970);
nand U30186 (N_30186,N_20298,N_25384);
xor U30187 (N_30187,N_22432,N_27692);
or U30188 (N_30188,N_28827,N_29501);
and U30189 (N_30189,N_22625,N_26459);
nand U30190 (N_30190,N_25937,N_26198);
xnor U30191 (N_30191,N_26861,N_25650);
nand U30192 (N_30192,N_24986,N_22507);
and U30193 (N_30193,N_26241,N_29675);
nor U30194 (N_30194,N_26128,N_25375);
nand U30195 (N_30195,N_26811,N_28197);
nand U30196 (N_30196,N_20452,N_28865);
nand U30197 (N_30197,N_29184,N_20409);
nand U30198 (N_30198,N_27753,N_25547);
or U30199 (N_30199,N_21483,N_23802);
nand U30200 (N_30200,N_24652,N_25362);
nor U30201 (N_30201,N_20730,N_22777);
nor U30202 (N_30202,N_22112,N_28603);
and U30203 (N_30203,N_28188,N_25783);
nand U30204 (N_30204,N_23000,N_29814);
nand U30205 (N_30205,N_22162,N_27812);
nor U30206 (N_30206,N_28525,N_24526);
nor U30207 (N_30207,N_24416,N_28203);
and U30208 (N_30208,N_24429,N_23146);
nor U30209 (N_30209,N_24616,N_21477);
or U30210 (N_30210,N_25327,N_23506);
or U30211 (N_30211,N_26598,N_21754);
nor U30212 (N_30212,N_20002,N_21098);
nor U30213 (N_30213,N_22163,N_26815);
nor U30214 (N_30214,N_26137,N_27667);
or U30215 (N_30215,N_29353,N_29131);
nor U30216 (N_30216,N_22058,N_22506);
or U30217 (N_30217,N_29791,N_29156);
or U30218 (N_30218,N_23532,N_22590);
xor U30219 (N_30219,N_21023,N_21384);
or U30220 (N_30220,N_28050,N_28908);
or U30221 (N_30221,N_29378,N_27882);
nor U30222 (N_30222,N_21040,N_29264);
or U30223 (N_30223,N_21435,N_28380);
or U30224 (N_30224,N_26644,N_21273);
nand U30225 (N_30225,N_23855,N_24572);
xor U30226 (N_30226,N_22557,N_23114);
nor U30227 (N_30227,N_21148,N_28398);
or U30228 (N_30228,N_21095,N_28163);
nand U30229 (N_30229,N_28598,N_27461);
nor U30230 (N_30230,N_24353,N_23646);
nor U30231 (N_30231,N_25838,N_29690);
nand U30232 (N_30232,N_21981,N_23213);
xnor U30233 (N_30233,N_28452,N_23942);
nor U30234 (N_30234,N_27844,N_29162);
nand U30235 (N_30235,N_20030,N_28449);
and U30236 (N_30236,N_23411,N_21522);
and U30237 (N_30237,N_24647,N_23708);
or U30238 (N_30238,N_29740,N_28034);
and U30239 (N_30239,N_26652,N_28156);
nand U30240 (N_30240,N_25226,N_27407);
xnor U30241 (N_30241,N_22332,N_29047);
and U30242 (N_30242,N_23884,N_21270);
and U30243 (N_30243,N_20749,N_29271);
and U30244 (N_30244,N_27000,N_24492);
xor U30245 (N_30245,N_23704,N_26699);
and U30246 (N_30246,N_28759,N_21138);
nand U30247 (N_30247,N_23574,N_24221);
nand U30248 (N_30248,N_25480,N_20210);
or U30249 (N_30249,N_29332,N_29043);
nand U30250 (N_30250,N_26689,N_24815);
nand U30251 (N_30251,N_23547,N_25358);
nor U30252 (N_30252,N_29736,N_27950);
and U30253 (N_30253,N_23782,N_26211);
and U30254 (N_30254,N_20443,N_24948);
xnor U30255 (N_30255,N_23712,N_21049);
nor U30256 (N_30256,N_23598,N_21608);
or U30257 (N_30257,N_21022,N_27536);
nor U30258 (N_30258,N_24776,N_25107);
nor U30259 (N_30259,N_26929,N_21394);
and U30260 (N_30260,N_20925,N_26639);
and U30261 (N_30261,N_29066,N_26970);
xnor U30262 (N_30262,N_21511,N_29565);
nand U30263 (N_30263,N_27747,N_24020);
nor U30264 (N_30264,N_25920,N_28772);
and U30265 (N_30265,N_29242,N_28778);
and U30266 (N_30266,N_25023,N_23421);
nor U30267 (N_30267,N_24093,N_25261);
nand U30268 (N_30268,N_28932,N_22362);
nand U30269 (N_30269,N_23196,N_29255);
nand U30270 (N_30270,N_27309,N_25842);
nand U30271 (N_30271,N_23182,N_25526);
nand U30272 (N_30272,N_29277,N_22976);
nand U30273 (N_30273,N_24226,N_29036);
xnor U30274 (N_30274,N_23252,N_24110);
or U30275 (N_30275,N_25238,N_22450);
nor U30276 (N_30276,N_24423,N_26479);
and U30277 (N_30277,N_23905,N_29459);
and U30278 (N_30278,N_29627,N_22364);
and U30279 (N_30279,N_24452,N_29203);
xnor U30280 (N_30280,N_25126,N_26112);
nand U30281 (N_30281,N_21735,N_22698);
or U30282 (N_30282,N_25906,N_23923);
nor U30283 (N_30283,N_23657,N_26510);
nand U30284 (N_30284,N_22011,N_29202);
or U30285 (N_30285,N_21020,N_24298);
or U30286 (N_30286,N_20208,N_21815);
and U30287 (N_30287,N_26700,N_27580);
and U30288 (N_30288,N_21336,N_25607);
nand U30289 (N_30289,N_27446,N_29848);
nor U30290 (N_30290,N_28839,N_22818);
nor U30291 (N_30291,N_26794,N_20908);
or U30292 (N_30292,N_24770,N_26356);
nor U30293 (N_30293,N_22591,N_20100);
nor U30294 (N_30294,N_29404,N_25378);
and U30295 (N_30295,N_28185,N_22356);
and U30296 (N_30296,N_21622,N_20119);
and U30297 (N_30297,N_23168,N_28068);
xnor U30298 (N_30298,N_23248,N_29391);
xor U30299 (N_30299,N_27097,N_20141);
nand U30300 (N_30300,N_20690,N_25114);
nor U30301 (N_30301,N_21380,N_28355);
nand U30302 (N_30302,N_26664,N_27191);
nor U30303 (N_30303,N_21504,N_29645);
xnor U30304 (N_30304,N_26317,N_29390);
or U30305 (N_30305,N_28924,N_25244);
and U30306 (N_30306,N_20201,N_22923);
nor U30307 (N_30307,N_29630,N_22664);
nand U30308 (N_30308,N_26345,N_23552);
nor U30309 (N_30309,N_20227,N_25401);
or U30310 (N_30310,N_20514,N_22472);
nor U30311 (N_30311,N_26687,N_28991);
nand U30312 (N_30312,N_20230,N_24205);
or U30313 (N_30313,N_23464,N_23145);
nor U30314 (N_30314,N_24843,N_27113);
nor U30315 (N_30315,N_28524,N_22448);
and U30316 (N_30316,N_22746,N_23658);
nor U30317 (N_30317,N_21263,N_27486);
nand U30318 (N_30318,N_28055,N_20464);
or U30319 (N_30319,N_21634,N_22391);
nor U30320 (N_30320,N_29567,N_25494);
or U30321 (N_30321,N_28004,N_24398);
nand U30322 (N_30322,N_25835,N_22510);
nor U30323 (N_30323,N_21330,N_22887);
or U30324 (N_30324,N_28118,N_25265);
or U30325 (N_30325,N_23586,N_21493);
and U30326 (N_30326,N_22694,N_27656);
xnor U30327 (N_30327,N_23354,N_27867);
and U30328 (N_30328,N_23046,N_20557);
or U30329 (N_30329,N_21862,N_28053);
xor U30330 (N_30330,N_24793,N_24713);
nand U30331 (N_30331,N_22139,N_29083);
nand U30332 (N_30332,N_21375,N_23073);
or U30333 (N_30333,N_20235,N_22868);
nor U30334 (N_30334,N_26176,N_27816);
xnor U30335 (N_30335,N_26302,N_26081);
nand U30336 (N_30336,N_29399,N_21628);
nor U30337 (N_30337,N_25080,N_29885);
xnor U30338 (N_30338,N_21975,N_28726);
nand U30339 (N_30339,N_23976,N_20901);
nor U30340 (N_30340,N_23364,N_20073);
nor U30341 (N_30341,N_21651,N_28635);
nor U30342 (N_30342,N_22329,N_28922);
nand U30343 (N_30343,N_22645,N_24612);
nor U30344 (N_30344,N_26725,N_29631);
xnor U30345 (N_30345,N_21010,N_21990);
and U30346 (N_30346,N_23858,N_22589);
and U30347 (N_30347,N_23885,N_21026);
or U30348 (N_30348,N_26545,N_27832);
nor U30349 (N_30349,N_29327,N_20937);
and U30350 (N_30350,N_27852,N_21415);
nand U30351 (N_30351,N_25393,N_28445);
and U30352 (N_30352,N_29087,N_21429);
or U30353 (N_30353,N_23384,N_21234);
or U30354 (N_30354,N_28243,N_24878);
xnor U30355 (N_30355,N_27004,N_28944);
and U30356 (N_30356,N_29145,N_20739);
nand U30357 (N_30357,N_29527,N_27017);
and U30358 (N_30358,N_28280,N_27282);
nor U30359 (N_30359,N_27681,N_28742);
or U30360 (N_30360,N_23171,N_24136);
nor U30361 (N_30361,N_29074,N_20881);
and U30362 (N_30362,N_27639,N_29237);
and U30363 (N_30363,N_29032,N_27566);
nand U30364 (N_30364,N_20459,N_24170);
and U30365 (N_30365,N_26000,N_27170);
nand U30366 (N_30366,N_24968,N_24576);
and U30367 (N_30367,N_21322,N_29654);
nand U30368 (N_30368,N_27871,N_23295);
nand U30369 (N_30369,N_23850,N_24714);
or U30370 (N_30370,N_25595,N_27440);
and U30371 (N_30371,N_22971,N_21379);
nor U30372 (N_30372,N_24208,N_28550);
nand U30373 (N_30373,N_28785,N_25037);
nor U30374 (N_30374,N_23424,N_29106);
xor U30375 (N_30375,N_29983,N_27019);
nand U30376 (N_30376,N_20205,N_23830);
and U30377 (N_30377,N_29564,N_23512);
nor U30378 (N_30378,N_27202,N_28056);
nor U30379 (N_30379,N_29441,N_22787);
nor U30380 (N_30380,N_25168,N_20065);
nand U30381 (N_30381,N_26440,N_20190);
and U30382 (N_30382,N_25019,N_24070);
or U30383 (N_30383,N_29135,N_29999);
and U30384 (N_30384,N_22614,N_22183);
nor U30385 (N_30385,N_21746,N_24748);
nand U30386 (N_30386,N_22990,N_25692);
and U30387 (N_30387,N_20214,N_23150);
and U30388 (N_30388,N_27063,N_24643);
nor U30389 (N_30389,N_25465,N_21866);
nor U30390 (N_30390,N_23249,N_24690);
xnor U30391 (N_30391,N_23635,N_22858);
xor U30392 (N_30392,N_27916,N_20244);
nand U30393 (N_30393,N_29951,N_25340);
nor U30394 (N_30394,N_23501,N_21366);
xnor U30395 (N_30395,N_28484,N_26006);
or U30396 (N_30396,N_26280,N_23151);
or U30397 (N_30397,N_20849,N_24787);
xnor U30398 (N_30398,N_23133,N_25252);
or U30399 (N_30399,N_20462,N_26281);
nand U30400 (N_30400,N_20390,N_20614);
or U30401 (N_30401,N_29365,N_27077);
xnor U30402 (N_30402,N_25487,N_27966);
and U30403 (N_30403,N_27061,N_24707);
nand U30404 (N_30404,N_21052,N_27940);
nand U30405 (N_30405,N_25407,N_26523);
nand U30406 (N_30406,N_28822,N_22279);
and U30407 (N_30407,N_25097,N_29863);
or U30408 (N_30408,N_22978,N_29424);
nor U30409 (N_30409,N_21442,N_28767);
nand U30410 (N_30410,N_29217,N_24051);
nand U30411 (N_30411,N_20544,N_28310);
and U30412 (N_30412,N_25026,N_26276);
nor U30413 (N_30413,N_24630,N_20355);
nor U30414 (N_30414,N_26110,N_23037);
and U30415 (N_30415,N_24792,N_27030);
and U30416 (N_30416,N_29721,N_23823);
or U30417 (N_30417,N_21820,N_23952);
nor U30418 (N_30418,N_23811,N_20639);
or U30419 (N_30419,N_20874,N_29673);
nand U30420 (N_30420,N_21489,N_24923);
or U30421 (N_30421,N_29011,N_26165);
nand U30422 (N_30422,N_25036,N_24715);
or U30423 (N_30423,N_28340,N_26336);
or U30424 (N_30424,N_24308,N_29045);
or U30425 (N_30425,N_24626,N_29127);
nand U30426 (N_30426,N_25893,N_21706);
nand U30427 (N_30427,N_28930,N_21213);
nand U30428 (N_30428,N_29345,N_24061);
and U30429 (N_30429,N_22027,N_28311);
and U30430 (N_30430,N_28366,N_28649);
and U30431 (N_30431,N_27835,N_26673);
nand U30432 (N_30432,N_29840,N_24590);
and U30433 (N_30433,N_27258,N_23045);
xnor U30434 (N_30434,N_26388,N_29280);
nand U30435 (N_30435,N_24198,N_27653);
xnor U30436 (N_30436,N_28949,N_23257);
nor U30437 (N_30437,N_24040,N_21082);
nand U30438 (N_30438,N_29770,N_29057);
nand U30439 (N_30439,N_23767,N_23882);
nand U30440 (N_30440,N_22793,N_26067);
nand U30441 (N_30441,N_28744,N_29086);
and U30442 (N_30442,N_25593,N_24834);
and U30443 (N_30443,N_28899,N_20082);
and U30444 (N_30444,N_26953,N_24274);
nor U30445 (N_30445,N_28493,N_23081);
nand U30446 (N_30446,N_23910,N_26167);
and U30447 (N_30447,N_24337,N_22455);
or U30448 (N_30448,N_26621,N_29766);
or U30449 (N_30449,N_26579,N_28901);
and U30450 (N_30450,N_24230,N_22543);
nand U30451 (N_30451,N_22046,N_26977);
and U30452 (N_30452,N_28667,N_20166);
nand U30453 (N_30453,N_27603,N_23367);
nand U30454 (N_30454,N_27222,N_23455);
or U30455 (N_30455,N_25289,N_28605);
and U30456 (N_30456,N_21530,N_28085);
or U30457 (N_30457,N_24798,N_21982);
nand U30458 (N_30458,N_29444,N_26896);
and U30459 (N_30459,N_27573,N_29750);
nor U30460 (N_30460,N_29454,N_22704);
or U30461 (N_30461,N_22227,N_29215);
nand U30462 (N_30462,N_25787,N_23068);
nand U30463 (N_30463,N_26981,N_29680);
nand U30464 (N_30464,N_25283,N_28089);
nand U30465 (N_30465,N_26581,N_22265);
and U30466 (N_30466,N_28779,N_27630);
nor U30467 (N_30467,N_23054,N_25216);
nand U30468 (N_30468,N_20556,N_27519);
nor U30469 (N_30469,N_20916,N_22906);
and U30470 (N_30470,N_22242,N_24538);
nand U30471 (N_30471,N_28896,N_28463);
nand U30472 (N_30472,N_28523,N_22071);
nor U30473 (N_30473,N_27500,N_25549);
or U30474 (N_30474,N_27276,N_26363);
and U30475 (N_30475,N_21441,N_22555);
and U30476 (N_30476,N_25856,N_27840);
nand U30477 (N_30477,N_25245,N_28968);
nand U30478 (N_30478,N_28905,N_21535);
or U30479 (N_30479,N_29640,N_22686);
nand U30480 (N_30480,N_23689,N_29330);
nand U30481 (N_30481,N_22556,N_21512);
or U30482 (N_30482,N_29165,N_26162);
nor U30483 (N_30483,N_27138,N_23938);
nand U30484 (N_30484,N_28975,N_22323);
or U30485 (N_30485,N_22598,N_20759);
or U30486 (N_30486,N_27450,N_26352);
or U30487 (N_30487,N_26224,N_24546);
or U30488 (N_30488,N_24644,N_23661);
and U30489 (N_30489,N_26287,N_21373);
or U30490 (N_30490,N_24741,N_28641);
nor U30491 (N_30491,N_25738,N_23616);
or U30492 (N_30492,N_25218,N_29284);
nand U30493 (N_30493,N_22250,N_23934);
nor U30494 (N_30494,N_28228,N_22185);
nand U30495 (N_30495,N_27147,N_25538);
xor U30496 (N_30496,N_27876,N_27128);
or U30497 (N_30497,N_29201,N_27674);
and U30498 (N_30498,N_25255,N_21955);
xor U30499 (N_30499,N_20552,N_23617);
nand U30500 (N_30500,N_20213,N_28751);
or U30501 (N_30501,N_26304,N_20961);
nand U30502 (N_30502,N_21621,N_28065);
nand U30503 (N_30503,N_25206,N_28096);
and U30504 (N_30504,N_26826,N_25975);
nand U30505 (N_30505,N_29553,N_20570);
or U30506 (N_30506,N_27306,N_20832);
nor U30507 (N_30507,N_21850,N_25724);
or U30508 (N_30508,N_23626,N_27843);
nand U30509 (N_30509,N_21035,N_26731);
and U30510 (N_30510,N_27130,N_21763);
xnor U30511 (N_30511,N_20246,N_24318);
nand U30512 (N_30512,N_25524,N_21632);
xor U30513 (N_30513,N_28417,N_29496);
nand U30514 (N_30514,N_23893,N_27891);
xor U30515 (N_30515,N_24606,N_24362);
or U30516 (N_30516,N_24117,N_23605);
xor U30517 (N_30517,N_20615,N_29533);
nand U30518 (N_30518,N_23419,N_24368);
and U30519 (N_30519,N_23828,N_22341);
nor U30520 (N_30520,N_22231,N_23630);
or U30521 (N_30521,N_23692,N_25442);
or U30522 (N_30522,N_26717,N_20300);
nand U30523 (N_30523,N_27102,N_29267);
xnor U30524 (N_30524,N_20179,N_20887);
nor U30525 (N_30525,N_26916,N_24509);
or U30526 (N_30526,N_23966,N_25125);
xnor U30527 (N_30527,N_23988,N_28009);
nand U30528 (N_30528,N_27417,N_25752);
or U30529 (N_30529,N_21297,N_26031);
nor U30530 (N_30530,N_24495,N_28464);
nor U30531 (N_30531,N_20132,N_24698);
or U30532 (N_30532,N_20497,N_20207);
or U30533 (N_30533,N_24413,N_29849);
and U30534 (N_30534,N_28387,N_26438);
nor U30535 (N_30535,N_22220,N_24939);
xor U30536 (N_30536,N_21737,N_26825);
nor U30537 (N_30537,N_29285,N_27547);
nor U30538 (N_30538,N_20037,N_24767);
nor U30539 (N_30539,N_20003,N_22226);
and U30540 (N_30540,N_27958,N_29337);
nand U30541 (N_30541,N_29315,N_20704);
nor U30542 (N_30542,N_21633,N_25837);
nand U30543 (N_30543,N_22705,N_22964);
xor U30544 (N_30544,N_25700,N_26709);
or U30545 (N_30545,N_26570,N_24681);
and U30546 (N_30546,N_26696,N_26188);
or U30547 (N_30547,N_27028,N_21251);
nor U30548 (N_30548,N_28602,N_20040);
nand U30549 (N_30549,N_22111,N_20211);
nor U30550 (N_30550,N_25355,N_27939);
nand U30551 (N_30551,N_23043,N_22509);
nor U30552 (N_30552,N_26918,N_28906);
nand U30553 (N_30553,N_25770,N_20289);
or U30554 (N_30554,N_20633,N_20480);
nor U30555 (N_30555,N_29827,N_20990);
nor U30556 (N_30556,N_24177,N_27411);
or U30557 (N_30557,N_24844,N_24842);
nor U30558 (N_30558,N_24216,N_29350);
or U30559 (N_30559,N_27722,N_26475);
and U30560 (N_30560,N_20099,N_20836);
nand U30561 (N_30561,N_27903,N_22264);
nand U30562 (N_30562,N_27524,N_28415);
or U30563 (N_30563,N_27088,N_20993);
and U30564 (N_30564,N_26425,N_28689);
and U30565 (N_30565,N_27877,N_28337);
nand U30566 (N_30566,N_29082,N_26159);
nand U30567 (N_30567,N_22766,N_22186);
and U30568 (N_30568,N_21570,N_26930);
nand U30569 (N_30569,N_23835,N_27884);
and U30570 (N_30570,N_21128,N_29466);
and U30571 (N_30571,N_25172,N_28306);
and U30572 (N_30572,N_20987,N_28222);
or U30573 (N_30573,N_28877,N_24141);
and U30574 (N_30574,N_21264,N_28900);
and U30575 (N_30575,N_28377,N_29767);
nor U30576 (N_30576,N_29913,N_28128);
nor U30577 (N_30577,N_22814,N_29832);
and U30578 (N_30578,N_21261,N_27729);
xor U30579 (N_30579,N_22918,N_23759);
nor U30580 (N_30580,N_29898,N_23999);
nand U30581 (N_30581,N_26884,N_22171);
and U30582 (N_30582,N_22679,N_29772);
or U30583 (N_30583,N_29905,N_22930);
nand U30584 (N_30584,N_22260,N_24067);
nand U30585 (N_30585,N_27013,N_26530);
and U30586 (N_30586,N_23460,N_26203);
and U30587 (N_30587,N_27106,N_25645);
and U30588 (N_30588,N_20979,N_22382);
xor U30589 (N_30589,N_20021,N_20192);
nand U30590 (N_30590,N_26420,N_29803);
and U30591 (N_30591,N_24933,N_21702);
nand U30592 (N_30592,N_24685,N_25137);
or U30593 (N_30593,N_29470,N_27196);
nand U30594 (N_30594,N_22015,N_29241);
and U30595 (N_30595,N_25344,N_26988);
or U30596 (N_30596,N_25560,N_29638);
nor U30597 (N_30597,N_24004,N_29954);
and U30598 (N_30598,N_25763,N_22866);
xor U30599 (N_30599,N_24397,N_21601);
nand U30600 (N_30600,N_28989,N_23353);
nand U30601 (N_30601,N_22563,N_25686);
or U30602 (N_30602,N_28296,N_25681);
nor U30603 (N_30603,N_24901,N_27819);
xnor U30604 (N_30604,N_29275,N_27745);
and U30605 (N_30605,N_25689,N_26898);
nand U30606 (N_30606,N_20193,N_25728);
xor U30607 (N_30607,N_26655,N_26643);
nor U30608 (N_30608,N_25493,N_21614);
nand U30609 (N_30609,N_20029,N_24824);
nor U30610 (N_30610,N_27397,N_21226);
or U30611 (N_30611,N_20125,N_29112);
and U30612 (N_30612,N_27521,N_20041);
nor U30613 (N_30613,N_27231,N_29157);
and U30614 (N_30614,N_26919,N_26150);
nand U30615 (N_30615,N_26237,N_23205);
nor U30616 (N_30616,N_23810,N_20375);
nor U30617 (N_30617,N_24440,N_28078);
nand U30618 (N_30618,N_25944,N_28308);
nor U30619 (N_30619,N_29266,N_22819);
xnor U30620 (N_30620,N_26248,N_22962);
and U30621 (N_30621,N_20657,N_28397);
or U30622 (N_30622,N_27322,N_20343);
or U30623 (N_30623,N_22379,N_21527);
nor U30624 (N_30624,N_25410,N_21507);
nand U30625 (N_30625,N_25693,N_20670);
nand U30626 (N_30626,N_29161,N_25162);
nor U30627 (N_30627,N_20280,N_23678);
nor U30628 (N_30628,N_25478,N_26402);
xor U30629 (N_30629,N_21929,N_24427);
nand U30630 (N_30630,N_23377,N_26692);
and U30631 (N_30631,N_20187,N_24252);
xnor U30632 (N_30632,N_21333,N_22259);
and U30633 (N_30633,N_29054,N_29023);
nor U30634 (N_30634,N_21948,N_24563);
nor U30635 (N_30635,N_28258,N_26103);
nor U30636 (N_30636,N_26715,N_25926);
or U30637 (N_30637,N_22985,N_20275);
or U30638 (N_30638,N_26395,N_22633);
nand U30639 (N_30639,N_28304,N_24243);
and U30640 (N_30640,N_22428,N_22079);
nand U30641 (N_30641,N_28629,N_28934);
and U30642 (N_30642,N_27240,N_28969);
nand U30643 (N_30643,N_29613,N_22177);
or U30644 (N_30644,N_26539,N_25486);
or U30645 (N_30645,N_22013,N_25637);
nor U30646 (N_30646,N_22276,N_23457);
or U30647 (N_30647,N_25923,N_20441);
nand U30648 (N_30648,N_23647,N_28695);
nand U30649 (N_30649,N_20649,N_29287);
nand U30650 (N_30650,N_23947,N_26451);
and U30651 (N_30651,N_23662,N_25514);
nor U30652 (N_30652,N_24201,N_24725);
nand U30653 (N_30653,N_20372,N_22418);
xor U30654 (N_30654,N_27087,N_26011);
nand U30655 (N_30655,N_21771,N_23591);
nor U30656 (N_30656,N_21146,N_24981);
and U30657 (N_30657,N_25809,N_23674);
and U30658 (N_30658,N_25777,N_29950);
or U30659 (N_30659,N_27168,N_22012);
nand U30660 (N_30660,N_27162,N_25707);
nor U30661 (N_30661,N_21120,N_26079);
nor U30662 (N_30662,N_20425,N_27990);
nor U30663 (N_30663,N_26903,N_26672);
and U30664 (N_30664,N_29873,N_24527);
or U30665 (N_30665,N_29194,N_21085);
or U30666 (N_30666,N_28697,N_26803);
or U30667 (N_30667,N_24248,N_25253);
nor U30668 (N_30668,N_28363,N_27645);
nor U30669 (N_30669,N_21712,N_29820);
nor U30670 (N_30670,N_23879,N_22039);
nand U30671 (N_30671,N_20102,N_25812);
nor U30672 (N_30672,N_25091,N_29336);
nor U30673 (N_30673,N_23982,N_22794);
nand U30674 (N_30674,N_22465,N_29549);
nand U30675 (N_30675,N_25330,N_27419);
nand U30676 (N_30676,N_29037,N_25232);
xor U30677 (N_30677,N_27669,N_29354);
and U30678 (N_30678,N_23599,N_23025);
xnor U30679 (N_30679,N_28917,N_29641);
or U30680 (N_30680,N_25917,N_25697);
nor U30681 (N_30681,N_20078,N_27715);
nand U30682 (N_30682,N_24483,N_24710);
nor U30683 (N_30683,N_23688,N_28980);
nor U30684 (N_30684,N_24673,N_25336);
and U30685 (N_30685,N_28950,N_27954);
or U30686 (N_30686,N_27993,N_25371);
xor U30687 (N_30687,N_27952,N_25490);
nor U30688 (N_30688,N_25750,N_26610);
and U30689 (N_30689,N_29587,N_21912);
and U30690 (N_30690,N_25470,N_24246);
and U30691 (N_30691,N_24972,N_21999);
nor U30692 (N_30692,N_28826,N_29058);
or U30693 (N_30693,N_21817,N_22042);
and U30694 (N_30694,N_27895,N_25776);
and U30695 (N_30695,N_29696,N_23160);
and U30696 (N_30696,N_20861,N_22325);
nor U30697 (N_30697,N_29782,N_21500);
nand U30698 (N_30698,N_24030,N_23483);
and U30699 (N_30699,N_29528,N_21296);
nand U30700 (N_30700,N_24348,N_20374);
and U30701 (N_30701,N_23660,N_28574);
xnor U30702 (N_30702,N_28617,N_20701);
or U30703 (N_30703,N_29828,N_29442);
and U30704 (N_30704,N_20264,N_27994);
nand U30705 (N_30705,N_28218,N_20168);
nand U30706 (N_30706,N_29799,N_24780);
xnor U30707 (N_30707,N_29576,N_23637);
and U30708 (N_30708,N_25994,N_21047);
and U30709 (N_30709,N_26034,N_21872);
or U30710 (N_30710,N_23467,N_29291);
and U30711 (N_30711,N_29618,N_29269);
and U30712 (N_30712,N_28520,N_21439);
or U30713 (N_30713,N_24354,N_21424);
and U30714 (N_30714,N_25764,N_23631);
xnor U30715 (N_30715,N_24729,N_25998);
and U30716 (N_30716,N_20854,N_23404);
xnor U30717 (N_30717,N_26379,N_27200);
and U30718 (N_30718,N_29824,N_25145);
nand U30719 (N_30719,N_27356,N_22789);
or U30720 (N_30720,N_24836,N_21560);
nand U30721 (N_30721,N_27855,N_28459);
or U30722 (N_30722,N_29326,N_26587);
xor U30723 (N_30723,N_25086,N_27626);
nand U30724 (N_30724,N_25075,N_28212);
or U30725 (N_30725,N_20888,N_23918);
nand U30726 (N_30726,N_20733,N_26119);
and U30727 (N_30727,N_27841,N_28780);
nand U30728 (N_30728,N_20506,N_20266);
or U30729 (N_30729,N_28375,N_25096);
or U30730 (N_30730,N_24135,N_21019);
or U30731 (N_30731,N_29172,N_27770);
nand U30732 (N_30732,N_28655,N_20540);
xor U30733 (N_30733,N_21642,N_29642);
nand U30734 (N_30734,N_23936,N_29439);
or U30735 (N_30735,N_25970,N_20225);
nor U30736 (N_30736,N_21863,N_27338);
nand U30737 (N_30737,N_25954,N_24323);
xnor U30738 (N_30738,N_29025,N_29520);
and U30739 (N_30739,N_23681,N_21551);
or U30740 (N_30740,N_21308,N_25397);
nor U30741 (N_30741,N_27615,N_20273);
or U30742 (N_30742,N_25815,N_27505);
nor U30743 (N_30743,N_25793,N_20754);
and U30744 (N_30744,N_28007,N_22050);
or U30745 (N_30745,N_23596,N_22409);
xnor U30746 (N_30746,N_24082,N_22728);
nand U30747 (N_30747,N_21951,N_26987);
or U30748 (N_30748,N_29836,N_23653);
or U30749 (N_30749,N_28384,N_28730);
or U30750 (N_30750,N_20000,N_29288);
nand U30751 (N_30751,N_28028,N_25182);
and U30752 (N_30752,N_22532,N_26743);
and U30753 (N_30753,N_22467,N_20800);
or U30754 (N_30754,N_22851,N_24593);
and U30755 (N_30755,N_25351,N_20151);
or U30756 (N_30756,N_24392,N_22198);
xor U30757 (N_30757,N_22319,N_26646);
xnor U30758 (N_30758,N_24909,N_20114);
nand U30759 (N_30759,N_25625,N_25376);
nand U30760 (N_30760,N_27429,N_22730);
nor U30761 (N_30761,N_27269,N_23346);
or U30762 (N_30762,N_25733,N_27410);
nor U30763 (N_30763,N_27034,N_20766);
nand U30764 (N_30764,N_21048,N_24488);
nand U30765 (N_30765,N_23259,N_27694);
nand U30766 (N_30766,N_27941,N_20722);
nor U30767 (N_30767,N_22151,N_29537);
or U30768 (N_30768,N_27250,N_29140);
and U30769 (N_30769,N_27336,N_27036);
and U30770 (N_30770,N_26677,N_23785);
nand U30771 (N_30771,N_27251,N_20194);
or U30772 (N_30772,N_23356,N_23853);
nor U30773 (N_30773,N_23258,N_23793);
or U30774 (N_30774,N_23435,N_21684);
and U30775 (N_30775,N_20809,N_22173);
or U30776 (N_30776,N_25116,N_27066);
nor U30777 (N_30777,N_24085,N_24409);
nor U30778 (N_30778,N_25576,N_29952);
and U30779 (N_30779,N_20142,N_20798);
nand U30780 (N_30780,N_27628,N_23526);
and U30781 (N_30781,N_23790,N_21711);
xnor U30782 (N_30782,N_25160,N_24706);
nand U30783 (N_30783,N_26258,N_22599);
xnor U30784 (N_30784,N_27727,N_26989);
or U30785 (N_30785,N_29029,N_21831);
and U30786 (N_30786,N_25677,N_20430);
nor U30787 (N_30787,N_21802,N_24858);
and U30788 (N_30788,N_22678,N_29469);
or U30789 (N_30789,N_21433,N_23312);
or U30790 (N_30790,N_21805,N_23901);
nand U30791 (N_30791,N_25010,N_21109);
nor U30792 (N_30792,N_22068,N_25790);
and U30793 (N_30793,N_28575,N_29480);
and U30794 (N_30794,N_21549,N_27980);
nor U30795 (N_30795,N_28832,N_28137);
nor U30796 (N_30796,N_28374,N_25239);
or U30797 (N_30797,N_22924,N_20787);
nand U30798 (N_30798,N_27921,N_21867);
nand U30799 (N_30799,N_28783,N_27266);
or U30800 (N_30800,N_21879,N_21363);
nor U30801 (N_30801,N_28555,N_25638);
and U30802 (N_30802,N_21525,N_22892);
nor U30803 (N_30803,N_25300,N_20302);
nor U30804 (N_30804,N_22179,N_20843);
or U30805 (N_30805,N_27796,N_24985);
xor U30806 (N_30806,N_27763,N_23175);
nor U30807 (N_30807,N_20404,N_21314);
and U30808 (N_30808,N_27648,N_22190);
nor U30809 (N_30809,N_28506,N_26505);
nor U30810 (N_30810,N_29821,N_28819);
nand U30811 (N_30811,N_22752,N_22817);
nor U30812 (N_30812,N_20233,N_26761);
or U30813 (N_30813,N_28115,N_28669);
nor U30814 (N_30814,N_27108,N_22921);
and U30815 (N_30815,N_25006,N_29958);
or U30816 (N_30816,N_21731,N_29777);
or U30817 (N_30817,N_24559,N_20317);
or U30818 (N_30818,N_20191,N_22998);
nor U30819 (N_30819,N_27273,N_23224);
nor U30820 (N_30820,N_25113,N_21166);
nor U30821 (N_30821,N_21042,N_20547);
nor U30822 (N_30822,N_24178,N_22367);
nand U30823 (N_30823,N_21970,N_27902);
nor U30824 (N_30824,N_24104,N_24852);
nor U30825 (N_30825,N_23102,N_29715);
nand U30826 (N_30826,N_24621,N_27766);
and U30827 (N_30827,N_23981,N_28119);
and U30828 (N_30828,N_20687,N_21638);
xnor U30829 (N_30829,N_27911,N_20933);
nor U30830 (N_30830,N_21773,N_26435);
nor U30831 (N_30831,N_23426,N_28853);
xor U30832 (N_30832,N_27593,N_20116);
and U30833 (N_30833,N_27541,N_21705);
or U30834 (N_30834,N_26623,N_21810);
and U30835 (N_30835,N_24346,N_29126);
nor U30836 (N_30836,N_26002,N_20376);
or U30837 (N_30837,N_24066,N_23335);
nor U30838 (N_30838,N_23776,N_27621);
nand U30839 (N_30839,N_26076,N_28548);
nand U30840 (N_30840,N_29166,N_25765);
xor U30841 (N_30841,N_26775,N_27607);
nor U30842 (N_30842,N_29197,N_24167);
nand U30843 (N_30843,N_23950,N_23585);
nor U30844 (N_30844,N_28320,N_22783);
nor U30845 (N_30845,N_22586,N_23563);
and U30846 (N_30846,N_24785,N_27131);
xor U30847 (N_30847,N_28170,N_20115);
and U30848 (N_30848,N_25680,N_27225);
and U30849 (N_30849,N_29735,N_21495);
or U30850 (N_30850,N_22750,N_27686);
or U30851 (N_30851,N_28921,N_28162);
and U30852 (N_30852,N_27714,N_20414);
and U30853 (N_30853,N_29415,N_22378);
xnor U30854 (N_30854,N_28776,N_29940);
nor U30855 (N_30855,N_28107,N_20989);
and U30856 (N_30856,N_24307,N_21799);
xnor U30857 (N_30857,N_23890,N_24378);
nand U30858 (N_30858,N_26560,N_28123);
and U30859 (N_30859,N_23768,N_27713);
nand U30860 (N_30860,N_22741,N_29700);
nand U30861 (N_30861,N_29195,N_24097);
and U30862 (N_30862,N_21640,N_22195);
nand U30863 (N_30863,N_22342,N_21976);
nor U30864 (N_30864,N_26925,N_28994);
nand U30865 (N_30865,N_26564,N_20220);
or U30866 (N_30866,N_24349,N_20095);
and U30867 (N_30867,N_27931,N_27447);
or U30868 (N_30868,N_28870,N_22836);
nand U30869 (N_30869,N_26456,N_24523);
and U30870 (N_30870,N_24998,N_23247);
and U30871 (N_30871,N_24041,N_22197);
xnor U30872 (N_30872,N_22519,N_28342);
nor U30873 (N_30873,N_24500,N_28941);
or U30874 (N_30874,N_20304,N_23801);
nor U30875 (N_30875,N_28233,N_21229);
nor U30876 (N_30876,N_21956,N_23652);
and U30877 (N_30877,N_26556,N_28435);
and U30878 (N_30878,N_20138,N_26712);
nand U30879 (N_30879,N_22363,N_26434);
nand U30880 (N_30880,N_21848,N_21846);
or U30881 (N_30881,N_27974,N_21252);
and U30882 (N_30882,N_28045,N_26219);
or U30883 (N_30883,N_25732,N_26542);
and U30884 (N_30884,N_29877,N_21928);
and U30885 (N_30885,N_26992,N_24261);
nand U30886 (N_30886,N_29748,N_23369);
nand U30887 (N_30887,N_27111,N_20555);
or U30888 (N_30888,N_24743,N_26502);
nor U30889 (N_30889,N_20886,N_27490);
and U30890 (N_30890,N_24585,N_27451);
nand U30891 (N_30891,N_21615,N_29002);
nor U30892 (N_30892,N_26437,N_27037);
or U30893 (N_30893,N_25186,N_28284);
nand U30894 (N_30894,N_26346,N_28597);
nor U30895 (N_30895,N_22727,N_24188);
nand U30896 (N_30896,N_24111,N_26177);
and U30897 (N_30897,N_28632,N_29341);
and U30898 (N_30898,N_25820,N_27935);
or U30899 (N_30899,N_20471,N_25949);
and U30900 (N_30900,N_20591,N_29467);
nand U30901 (N_30901,N_25429,N_25074);
nor U30902 (N_30902,N_22157,N_20767);
nand U30903 (N_30903,N_20957,N_29578);
nor U30904 (N_30904,N_21859,N_21046);
nand U30905 (N_30905,N_22486,N_26513);
and U30906 (N_30906,N_29996,N_22369);
or U30907 (N_30907,N_26770,N_29150);
nor U30908 (N_30908,N_22142,N_24668);
or U30909 (N_30909,N_23718,N_29016);
nand U30910 (N_30910,N_23549,N_24232);
nor U30911 (N_30911,N_29909,N_26191);
nand U30912 (N_30912,N_29548,N_25139);
nand U30913 (N_30913,N_20735,N_23867);
nand U30914 (N_30914,N_21393,N_24536);
and U30915 (N_30915,N_23625,N_20009);
nor U30916 (N_30916,N_26983,N_20835);
xnor U30917 (N_30917,N_25250,N_22102);
nor U30918 (N_30918,N_29125,N_21946);
nand U30919 (N_30919,N_22515,N_20674);
or U30920 (N_30920,N_23383,N_21838);
nor U30921 (N_30921,N_20450,N_27600);
nor U30922 (N_30922,N_23870,N_20180);
nand U30923 (N_30923,N_20270,N_20596);
or U30924 (N_30924,N_26186,N_24379);
nor U30925 (N_30925,N_20109,N_22885);
nor U30926 (N_30926,N_28198,N_20543);
or U30927 (N_30927,N_20248,N_29426);
nand U30928 (N_30928,N_24598,N_22388);
and U30929 (N_30929,N_21563,N_26262);
nor U30930 (N_30930,N_26029,N_29273);
nor U30931 (N_30931,N_25847,N_23497);
nor U30932 (N_30932,N_27464,N_21553);
and U30933 (N_30933,N_25556,N_27976);
xnor U30934 (N_30934,N_22132,N_21644);
or U30935 (N_30935,N_28169,N_22435);
xnor U30936 (N_30936,N_28019,N_25150);
nand U30937 (N_30937,N_20062,N_23032);
nand U30938 (N_30938,N_27209,N_22993);
or U30939 (N_30939,N_28231,N_20820);
xnor U30940 (N_30940,N_20139,N_24347);
or U30941 (N_30941,N_26407,N_29850);
xor U30942 (N_30942,N_27366,N_24667);
nor U30943 (N_30943,N_22773,N_29953);
nand U30944 (N_30944,N_21230,N_27742);
nor U30945 (N_30945,N_24520,N_23784);
and U30946 (N_30946,N_28092,N_29990);
nand U30947 (N_30947,N_27233,N_21398);
and U30948 (N_30948,N_23581,N_20562);
nand U30949 (N_30949,N_21271,N_24207);
nand U30950 (N_30950,N_28782,N_22981);
or U30951 (N_30951,N_24457,N_26680);
or U30952 (N_30952,N_22936,N_21072);
or U30953 (N_30953,N_22305,N_21700);
xnor U30954 (N_30954,N_22583,N_29729);
or U30955 (N_30955,N_26854,N_28527);
xor U30956 (N_30956,N_26424,N_23300);
nand U30957 (N_30957,N_29357,N_29098);
xor U30958 (N_30958,N_20929,N_22085);
nor U30959 (N_30959,N_24615,N_24271);
or U30960 (N_30960,N_22853,N_25176);
and U30961 (N_30961,N_27247,N_23119);
nand U30962 (N_30962,N_26907,N_28806);
or U30963 (N_30963,N_21005,N_20217);
nand U30964 (N_30964,N_20365,N_23697);
and U30965 (N_30965,N_27099,N_23529);
and U30966 (N_30966,N_25735,N_21268);
or U30967 (N_30967,N_20483,N_28769);
or U30968 (N_30968,N_20655,N_25816);
nand U30969 (N_30969,N_21891,N_22635);
xnor U30970 (N_30970,N_27144,N_22129);
xnor U30971 (N_30971,N_28577,N_29557);
and U30972 (N_30972,N_29204,N_21589);
nor U30973 (N_30973,N_23069,N_27712);
nor U30974 (N_30974,N_28326,N_20966);
or U30975 (N_30975,N_24490,N_22007);
and U30976 (N_30976,N_29523,N_25611);
or U30977 (N_30977,N_20903,N_28547);
or U30978 (N_30978,N_28571,N_24065);
nor U30979 (N_30979,N_26205,N_28026);
nor U30980 (N_30980,N_29887,N_29808);
or U30981 (N_30981,N_23214,N_23250);
and U30982 (N_30982,N_26799,N_29771);
nand U30983 (N_30983,N_20036,N_29724);
or U30984 (N_30984,N_20523,N_26886);
nor U30985 (N_30985,N_23641,N_21655);
nand U30986 (N_30986,N_22209,N_29021);
xor U30987 (N_30987,N_24660,N_28580);
xnor U30988 (N_30988,N_25169,N_24212);
and U30989 (N_30989,N_23111,N_28872);
nor U30990 (N_30990,N_22307,N_21257);
xnor U30991 (N_30991,N_26100,N_21053);
nor U30992 (N_30992,N_24876,N_25462);
nand U30993 (N_30993,N_23116,N_29116);
nor U30994 (N_30994,N_22212,N_22394);
and U30995 (N_30995,N_23430,N_28738);
and U30996 (N_30996,N_22168,N_26102);
and U30997 (N_30997,N_22606,N_25264);
nor U30998 (N_30998,N_28286,N_28929);
nor U30999 (N_30999,N_24254,N_28209);
and U31000 (N_31000,N_21931,N_26967);
and U31001 (N_31001,N_24028,N_21749);
nand U31002 (N_31002,N_27340,N_29017);
nand U31003 (N_31003,N_27969,N_28219);
and U31004 (N_31004,N_24934,N_20202);
nor U31005 (N_31005,N_22516,N_28875);
and U31006 (N_31006,N_29238,N_23019);
xnor U31007 (N_31007,N_23624,N_28746);
or U31008 (N_31008,N_21678,N_29506);
nand U31009 (N_31009,N_22512,N_25270);
and U31010 (N_31010,N_26265,N_29968);
or U31011 (N_31011,N_27563,N_24275);
nand U31012 (N_31012,N_22601,N_24052);
or U31013 (N_31013,N_24036,N_21137);
nand U31014 (N_31014,N_27083,N_26196);
nor U31015 (N_31015,N_26494,N_21501);
nand U31016 (N_31016,N_20301,N_20129);
xor U31017 (N_31017,N_29308,N_22283);
nand U31018 (N_31018,N_28013,N_27716);
nor U31019 (N_31019,N_29810,N_28749);
nor U31020 (N_31020,N_29304,N_21602);
and U31021 (N_31021,N_22397,N_28585);
and U31022 (N_31022,N_29614,N_20044);
and U31023 (N_31023,N_27800,N_24560);
nor U31024 (N_31024,N_28274,N_28359);
nor U31025 (N_31025,N_26371,N_26710);
nand U31026 (N_31026,N_25212,N_22347);
xor U31027 (N_31027,N_25360,N_20056);
nand U31028 (N_31028,N_22024,N_28918);
nor U31029 (N_31029,N_26616,N_21240);
nor U31030 (N_31030,N_24278,N_20943);
or U31031 (N_31031,N_21231,N_28294);
and U31032 (N_31032,N_29387,N_24807);
nand U31033 (N_31033,N_23894,N_25015);
or U31034 (N_31034,N_27609,N_22236);
or U31035 (N_31035,N_28223,N_23292);
and U31036 (N_31036,N_28325,N_20997);
or U31037 (N_31037,N_20597,N_26651);
and U31038 (N_31038,N_22952,N_29392);
nor U31039 (N_31039,N_28804,N_20958);
xnor U31040 (N_31040,N_21789,N_28664);
and U31041 (N_31041,N_23307,N_22023);
nor U31042 (N_31042,N_22032,N_24297);
nor U31043 (N_31043,N_27046,N_24687);
nor U31044 (N_31044,N_28288,N_28569);
nand U31045 (N_31045,N_23080,N_20826);
and U31046 (N_31046,N_25916,N_29214);
xor U31047 (N_31047,N_20382,N_21222);
or U31048 (N_31048,N_25333,N_23004);
nor U31049 (N_31049,N_28911,N_26056);
and U31050 (N_31050,N_21370,N_20685);
nand U31051 (N_31051,N_21066,N_28752);
xnor U31052 (N_31052,N_28133,N_25924);
or U31053 (N_31053,N_20121,N_26634);
nor U31054 (N_31054,N_26445,N_21423);
nor U31055 (N_31055,N_26756,N_29425);
nand U31056 (N_31056,N_21492,N_21719);
nand U31057 (N_31057,N_25656,N_21460);
nor U31058 (N_31058,N_28849,N_28111);
nor U31059 (N_31059,N_20696,N_21184);
nor U31060 (N_31060,N_28270,N_20532);
xnor U31061 (N_31061,N_28518,N_23187);
nor U31062 (N_31062,N_26969,N_22520);
and U31063 (N_31063,N_27423,N_23725);
xnor U31064 (N_31064,N_25328,N_23374);
or U31065 (N_31065,N_25452,N_23123);
nor U31066 (N_31066,N_28857,N_24674);
nor U31067 (N_31067,N_29947,N_22224);
or U31068 (N_31068,N_29376,N_26955);
and U31069 (N_31069,N_21303,N_27587);
or U31070 (N_31070,N_20148,N_28104);
nand U31071 (N_31071,N_25320,N_26917);
and U31072 (N_31072,N_26923,N_20410);
nor U31073 (N_31073,N_26013,N_23242);
xnor U31074 (N_31074,N_24731,N_29519);
or U31075 (N_31075,N_20057,N_28492);
and U31076 (N_31076,N_25124,N_28942);
and U31077 (N_31077,N_25449,N_28718);
and U31078 (N_31078,N_25604,N_25368);
nor U31079 (N_31079,N_28350,N_24417);
and U31080 (N_31080,N_29379,N_27156);
xor U31081 (N_31081,N_21041,N_23189);
nand U31082 (N_31082,N_26204,N_20624);
xor U31083 (N_31083,N_21150,N_24571);
or U31084 (N_31084,N_22103,N_23006);
or U31085 (N_31085,N_20159,N_20111);
and U31086 (N_31086,N_21626,N_28404);
and U31087 (N_31087,N_29509,N_27146);
or U31088 (N_31088,N_29966,N_24334);
nor U31089 (N_31089,N_22775,N_20593);
nor U31090 (N_31090,N_26252,N_29938);
and U31091 (N_31091,N_27139,N_27631);
and U31092 (N_31092,N_23492,N_25840);
nor U31093 (N_31093,N_20239,N_28358);
and U31094 (N_31094,N_27227,N_27142);
nor U31095 (N_31095,N_27389,N_22593);
nand U31096 (N_31096,N_22547,N_28619);
nand U31097 (N_31097,N_21177,N_21167);
or U31098 (N_31098,N_28946,N_24862);
nor U31099 (N_31099,N_20879,N_24587);
nand U31100 (N_31100,N_22886,N_21533);
or U31101 (N_31101,N_26077,N_21612);
xor U31102 (N_31102,N_26657,N_23849);
nand U31103 (N_31103,N_26492,N_25952);
nor U31104 (N_31104,N_25582,N_24945);
nand U31105 (N_31105,N_20035,N_28333);
and U31106 (N_31106,N_23925,N_20087);
nand U31107 (N_31107,N_27284,N_24101);
nor U31108 (N_31108,N_23974,N_29093);
xnor U31109 (N_31109,N_24820,N_28314);
and U31110 (N_31110,N_27062,N_20417);
nand U31111 (N_31111,N_27158,N_24826);
nor U31112 (N_31112,N_25586,N_22568);
nand U31113 (N_31113,N_22470,N_28437);
or U31114 (N_31114,N_20502,N_20952);
nor U31115 (N_31115,N_22361,N_28959);
and U31116 (N_31116,N_24173,N_25522);
and U31117 (N_31117,N_22530,N_26273);
nor U31118 (N_31118,N_27730,N_23063);
or U31119 (N_31119,N_25193,N_22812);
or U31120 (N_31120,N_23456,N_25950);
or U31121 (N_31121,N_25105,N_24019);
or U31122 (N_31122,N_28868,N_26613);
nand U31123 (N_31123,N_24463,N_29388);
nand U31124 (N_31124,N_21488,N_29676);
or U31125 (N_31125,N_27478,N_28933);
or U31126 (N_31126,N_28720,N_23104);
nor U31127 (N_31127,N_22637,N_22218);
nand U31128 (N_31128,N_22499,N_25079);
nor U31129 (N_31129,N_24304,N_24890);
or U31130 (N_31130,N_26784,N_22128);
and U31131 (N_31131,N_29321,N_20870);
or U31132 (N_31132,N_22908,N_29371);
or U31133 (N_31133,N_28882,N_20454);
xnor U31134 (N_31134,N_29707,N_20250);
and U31135 (N_31135,N_22113,N_29749);
nand U31136 (N_31136,N_27904,N_22213);
nor U31137 (N_31137,N_28867,N_26487);
and U31138 (N_31138,N_26341,N_21011);
xor U31139 (N_31139,N_27608,N_22376);
nand U31140 (N_31140,N_23067,N_20113);
and U31141 (N_31141,N_23695,N_27912);
nor U31142 (N_31142,N_23011,N_29063);
xnor U31143 (N_31143,N_24290,N_22178);
nor U31144 (N_31144,N_24946,N_28250);
or U31145 (N_31145,N_25237,N_27658);
and U31146 (N_31146,N_21649,N_23061);
or U31147 (N_31147,N_28419,N_21957);
nor U31148 (N_31148,N_29812,N_21677);
or U31149 (N_31149,N_20714,N_28426);
nand U31150 (N_31150,N_24619,N_22137);
or U31151 (N_31151,N_20736,N_26064);
nand U31152 (N_31152,N_23783,N_23929);
or U31153 (N_31153,N_26786,N_25672);
nand U31154 (N_31154,N_20059,N_22955);
or U31155 (N_31155,N_26812,N_27811);
and U31156 (N_31156,N_25627,N_26339);
or U31157 (N_31157,N_29292,N_27186);
and U31158 (N_31158,N_24568,N_22334);
xnor U31159 (N_31159,N_23634,N_25719);
nor U31160 (N_31160,N_22712,N_26574);
xnor U31161 (N_31161,N_23756,N_22251);
and U31162 (N_31162,N_27215,N_28636);
and U31163 (N_31163,N_22622,N_21580);
nor U31164 (N_31164,N_22500,N_26261);
nor U31165 (N_31165,N_26457,N_29518);
or U31166 (N_31166,N_27382,N_26490);
xnor U31167 (N_31167,N_20688,N_21277);
nand U31168 (N_31168,N_20110,N_20859);
nor U31169 (N_31169,N_26589,N_26593);
nor U31170 (N_31170,N_24839,N_25454);
and U31171 (N_31171,N_25919,N_27588);
xnor U31172 (N_31172,N_21961,N_29461);
or U31173 (N_31173,N_21937,N_20810);
nand U31174 (N_31174,N_22327,N_24900);
or U31175 (N_31175,N_23716,N_21913);
and U31176 (N_31176,N_26004,N_22638);
or U31177 (N_31177,N_20803,N_25204);
or U31178 (N_31178,N_20071,N_23135);
or U31179 (N_31179,N_27489,N_23565);
or U31180 (N_31180,N_28488,N_28051);
or U31181 (N_31181,N_27344,N_22891);
and U31182 (N_31182,N_20960,N_26693);
nand U31183 (N_31183,N_28568,N_25347);
nor U31184 (N_31184,N_24046,N_29333);
xor U31185 (N_31185,N_20445,N_26320);
nand U31186 (N_31186,N_25127,N_28316);
nor U31187 (N_31187,N_29319,N_21455);
nand U31188 (N_31188,N_29191,N_22763);
nor U31189 (N_31189,N_22043,N_29764);
and U31190 (N_31190,N_29859,N_21579);
nand U31191 (N_31191,N_22407,N_27571);
and U31192 (N_31192,N_25706,N_28237);
nand U31193 (N_31193,N_24530,N_24466);
nand U31194 (N_31194,N_29693,N_28328);
nand U31195 (N_31195,N_23309,N_20342);
or U31196 (N_31196,N_22166,N_27015);
nor U31197 (N_31197,N_27123,N_27611);
nor U31198 (N_31198,N_27885,N_29738);
xor U31199 (N_31199,N_29920,N_29219);
nand U31200 (N_31200,N_23553,N_21312);
or U31201 (N_31201,N_20938,N_20053);
and U31202 (N_31202,N_22587,N_28341);
nor U31203 (N_31203,N_26489,N_20158);
or U31204 (N_31204,N_20784,N_20097);
nand U31205 (N_31205,N_23305,N_27388);
nor U31206 (N_31206,N_26024,N_23165);
or U31207 (N_31207,N_28309,N_26935);
nor U31208 (N_31208,N_25762,N_23417);
nand U31209 (N_31209,N_20360,N_29864);
nand U31210 (N_31210,N_26134,N_25544);
or U31211 (N_31211,N_28234,N_24617);
nand U31212 (N_31212,N_27597,N_22521);
and U31213 (N_31213,N_29381,N_27485);
and U31214 (N_31214,N_24486,N_23142);
xnor U31215 (N_31215,N_20118,N_29447);
or U31216 (N_31216,N_28046,N_25198);
and U31217 (N_31217,N_21063,N_23222);
and U31218 (N_31218,N_28072,N_28313);
and U31219 (N_31219,N_27548,N_25158);
nand U31220 (N_31220,N_28940,N_23593);
or U31221 (N_31221,N_27471,N_21032);
nand U31222 (N_31222,N_25977,N_22117);
and U31223 (N_31223,N_27027,N_28161);
and U31224 (N_31224,N_21450,N_21168);
nor U31225 (N_31225,N_24833,N_26518);
and U31226 (N_31226,N_20918,N_28528);
nand U31227 (N_31227,N_22861,N_22641);
nand U31228 (N_31228,N_24937,N_23709);
nand U31229 (N_31229,N_29660,N_21598);
and U31230 (N_31230,N_25388,N_24718);
xnor U31231 (N_31231,N_21051,N_24350);
nor U31232 (N_31232,N_23555,N_22977);
and U31233 (N_31233,N_22424,N_21179);
nand U31234 (N_31234,N_29505,N_25467);
nor U31235 (N_31235,N_28596,N_27436);
nand U31236 (N_31236,N_26508,N_20906);
xor U31237 (N_31237,N_29896,N_23436);
xnor U31238 (N_31238,N_25390,N_24682);
nand U31239 (N_31239,N_27264,N_26844);
or U31240 (N_31240,N_20666,N_26802);
and U31241 (N_31241,N_23479,N_21054);
and U31242 (N_31242,N_26830,N_20519);
nor U31243 (N_31243,N_27551,N_22446);
and U31244 (N_31244,N_28589,N_27706);
or U31245 (N_31245,N_26359,N_29030);
nand U31246 (N_31246,N_24701,N_24800);
nand U31247 (N_31247,N_27951,N_26882);
nand U31248 (N_31248,N_27552,N_27422);
and U31249 (N_31249,N_21883,N_21698);
and U31250 (N_31250,N_20010,N_29347);
and U31251 (N_31251,N_29666,N_26627);
nand U31252 (N_31252,N_24158,N_27542);
and U31253 (N_31253,N_20522,N_24650);
or U31254 (N_31254,N_20602,N_21059);
nor U31255 (N_31255,N_22748,N_27691);
nand U31256 (N_31256,N_25353,N_23201);
nand U31257 (N_31257,N_20146,N_29623);
nor U31258 (N_31258,N_27502,N_28038);
and U31259 (N_31259,N_25532,N_27889);
nor U31260 (N_31260,N_29153,N_22018);
xnor U31261 (N_31261,N_26391,N_22567);
and U31262 (N_31262,N_29230,N_20383);
or U31263 (N_31263,N_25251,N_29449);
and U31264 (N_31264,N_26534,N_20005);
nor U31265 (N_31265,N_29373,N_23724);
xor U31266 (N_31266,N_29432,N_26048);
nand U31267 (N_31267,N_27875,N_26117);
nor U31268 (N_31268,N_28347,N_27594);
and U31269 (N_31269,N_23538,N_29468);
nor U31270 (N_31270,N_23183,N_22815);
and U31271 (N_31271,N_28495,N_27689);
xor U31272 (N_31272,N_21395,N_29055);
nor U31273 (N_31273,N_24906,N_22890);
and U31274 (N_31274,N_25383,N_25194);
nand U31275 (N_31275,N_22541,N_24281);
nor U31276 (N_31276,N_27731,N_24197);
or U31277 (N_31277,N_20717,N_28192);
nor U31278 (N_31278,N_28859,N_20860);
nand U31279 (N_31279,N_27604,N_22045);
xnor U31280 (N_31280,N_23638,N_27828);
and U31281 (N_31281,N_25365,N_20080);
or U31282 (N_31282,N_21097,N_25909);
and U31283 (N_31283,N_21979,N_28633);
nand U31284 (N_31284,N_20574,N_25725);
nor U31285 (N_31285,N_21934,N_26251);
or U31286 (N_31286,N_23216,N_23342);
nor U31287 (N_31287,N_22967,N_20622);
nand U31288 (N_31288,N_20131,N_24196);
nor U31289 (N_31289,N_21755,N_28160);
nand U31290 (N_31290,N_24657,N_28856);
nand U31291 (N_31291,N_26720,N_26483);
and U31292 (N_31292,N_23866,N_25363);
or U31293 (N_31293,N_20631,N_20513);
xnor U31294 (N_31294,N_22739,N_29530);
nor U31295 (N_31295,N_28674,N_22808);
nand U31296 (N_31296,N_24089,N_22869);
nor U31297 (N_31297,N_28265,N_28961);
nand U31298 (N_31298,N_20281,N_27310);
or U31299 (N_31299,N_26335,N_25418);
nand U31300 (N_31300,N_26850,N_29453);
and U31301 (N_31301,N_21083,N_25121);
or U31302 (N_31302,N_22940,N_23212);
or U31303 (N_31303,N_27554,N_29257);
or U31304 (N_31304,N_26573,N_28953);
nand U31305 (N_31305,N_23710,N_21412);
nor U31306 (N_31306,N_22313,N_25272);
xnor U31307 (N_31307,N_25709,N_23044);
nand U31308 (N_31308,N_29433,N_24420);
and U31309 (N_31309,N_22422,N_29122);
nand U31310 (N_31310,N_23164,N_22749);
xor U31311 (N_31311,N_20149,N_24134);
or U31312 (N_31312,N_21065,N_27635);
and U31313 (N_31313,N_26867,N_20387);
nand U31314 (N_31314,N_23649,N_23386);
nand U31315 (N_31315,N_27781,N_24720);
and U31316 (N_31316,N_28367,N_29992);
xor U31317 (N_31317,N_20165,N_26512);
xnor U31318 (N_31318,N_29251,N_29758);
and U31319 (N_31319,N_29911,N_23370);
nor U31320 (N_31320,N_25579,N_22901);
or U31321 (N_31321,N_26940,N_28073);
nand U31322 (N_31322,N_21381,N_21337);
or U31323 (N_31323,N_25831,N_21088);
nand U31324 (N_31324,N_24411,N_29064);
nand U31325 (N_31325,N_21290,N_29684);
and U31326 (N_31326,N_29050,N_27598);
nor U31327 (N_31327,N_22796,N_20197);
nand U31328 (N_31328,N_24582,N_26309);
or U31329 (N_31329,N_28634,N_25737);
and U31330 (N_31330,N_28125,N_23352);
nor U31331 (N_31331,N_28887,N_22548);
nand U31332 (N_31332,N_20412,N_23385);
nand U31333 (N_31333,N_20720,N_25933);
nand U31334 (N_31334,N_24125,N_25403);
nand U31335 (N_31335,N_25851,N_26496);
nand U31336 (N_31336,N_27636,N_28491);
and U31337 (N_31337,N_23355,N_25523);
and U31338 (N_31338,N_27183,N_22737);
xnor U31339 (N_31339,N_24959,N_26426);
and U31340 (N_31340,N_21588,N_20811);
nand U31341 (N_31341,N_23920,N_22115);
xnor U31342 (N_31342,N_25337,N_21671);
or U31343 (N_31343,N_23477,N_21208);
nand U31344 (N_31344,N_28958,N_23514);
nand U31345 (N_31345,N_26040,N_20752);
nor U31346 (N_31346,N_28414,N_26772);
nand U31347 (N_31347,N_21401,N_29290);
xnor U31348 (N_31348,N_20904,N_23105);
nor U31349 (N_31349,N_22210,N_28609);
or U31350 (N_31350,N_21768,N_28850);
or U31351 (N_31351,N_24294,N_25188);
or U31352 (N_31352,N_21110,N_25761);
and U31353 (N_31353,N_23434,N_23832);
and U31354 (N_31354,N_27863,N_20917);
and U31355 (N_31355,N_24328,N_23755);
and U31356 (N_31356,N_28372,N_26232);
or U31357 (N_31357,N_29619,N_25553);
nor U31358 (N_31358,N_23391,N_22974);
xor U31359 (N_31359,N_21555,N_23548);
nand U31360 (N_31360,N_27076,N_22040);
xnor U31361 (N_31361,N_27733,N_23505);
nor U31362 (N_31362,N_24424,N_26491);
nand U31363 (N_31363,N_20296,N_24365);
nand U31364 (N_31364,N_24989,N_24952);
nor U31365 (N_31365,N_27293,N_22792);
xnor U31366 (N_31366,N_27720,N_25269);
or U31367 (N_31367,N_20793,N_23279);
nor U31368 (N_31368,N_27494,N_27465);
nand U31369 (N_31369,N_20847,N_21265);
and U31370 (N_31370,N_20440,N_28473);
nor U31371 (N_31371,N_20738,N_27792);
or U31372 (N_31372,N_24819,N_27643);
nor U31373 (N_31373,N_23699,N_28938);
and U31374 (N_31374,N_24186,N_22340);
and U31375 (N_31375,N_29817,N_21186);
and U31376 (N_31376,N_20429,N_27782);
nand U31377 (N_31377,N_26374,N_23495);
nor U31378 (N_31378,N_20768,N_25497);
and U31379 (N_31379,N_27760,N_21298);
nor U31380 (N_31380,N_21962,N_27893);
xnor U31381 (N_31381,N_24237,N_26019);
and U31382 (N_31382,N_24451,N_29568);
and U31383 (N_31383,N_26168,N_22034);
and U31384 (N_31384,N_23632,N_26557);
or U31385 (N_31385,N_29245,N_26266);
xor U31386 (N_31386,N_21115,N_22907);
and U31387 (N_31387,N_22956,N_29995);
and U31388 (N_31388,N_20548,N_21721);
or U31389 (N_31389,N_20538,N_22067);
nor U31390 (N_31390,N_24762,N_21254);
or U31391 (N_31391,N_21285,N_25517);
or U31392 (N_31392,N_25059,N_29904);
nand U31393 (N_31393,N_27749,N_20638);
xor U31394 (N_31394,N_24545,N_22658);
and U31395 (N_31395,N_27672,N_25873);
and U31396 (N_31396,N_27457,N_23389);
nor U31397 (N_31397,N_22055,N_22838);
nand U31398 (N_31398,N_24074,N_27967);
or U31399 (N_31399,N_20866,N_23031);
nand U31400 (N_31400,N_24921,N_20763);
nor U31401 (N_31401,N_23804,N_23743);
nor U31402 (N_31402,N_22275,N_23595);
nand U31403 (N_31403,N_27361,N_22731);
and U31404 (N_31404,N_28037,N_21235);
nand U31405 (N_31405,N_27242,N_24874);
and U31406 (N_31406,N_25415,N_21445);
nand U31407 (N_31407,N_23128,N_23198);
or U31408 (N_31408,N_27908,N_25900);
or U31409 (N_31409,N_26136,N_23509);
and U31410 (N_31410,N_27031,N_21425);
and U31411 (N_31411,N_26952,N_28299);
and U31412 (N_31412,N_26515,N_25921);
and U31413 (N_31413,N_23545,N_28920);
or U31414 (N_31414,N_29972,N_25561);
nand U31415 (N_31415,N_20345,N_26035);
and U31416 (N_31416,N_28187,N_29307);
nor U31417 (N_31417,N_28136,N_27592);
and U31418 (N_31418,N_20672,N_28533);
nand U31419 (N_31419,N_20728,N_23939);
nand U31420 (N_31420,N_22351,N_27531);
or U31421 (N_31421,N_24489,N_28971);
or U31422 (N_31422,N_26838,N_23193);
or U31423 (N_31423,N_21723,N_28521);
nor U31424 (N_31424,N_25177,N_26401);
nor U31425 (N_31425,N_23805,N_28998);
and U31426 (N_31426,N_23998,N_21262);
nand U31427 (N_31427,N_26370,N_23267);
nor U31428 (N_31428,N_22339,N_22254);
nand U31429 (N_31429,N_22784,N_29601);
or U31430 (N_31430,N_29809,N_23733);
nand U31431 (N_31431,N_22009,N_25385);
nor U31432 (N_31432,N_25948,N_23612);
nor U31433 (N_31433,N_27110,N_26991);
or U31434 (N_31434,N_29348,N_21195);
or U31435 (N_31435,N_21743,N_23338);
nor U31436 (N_31436,N_23609,N_27562);
xnor U31437 (N_31437,N_25382,N_28624);
nor U31438 (N_31438,N_22820,N_28031);
nand U31439 (N_31439,N_22761,N_23002);
nor U31440 (N_31440,N_27117,N_29819);
nand U31441 (N_31441,N_28732,N_25243);
and U31442 (N_31442,N_29160,N_21539);
and U31443 (N_31443,N_22126,N_28207);
and U31444 (N_31444,N_24395,N_25584);
and U31445 (N_31445,N_27274,N_25356);
nor U31446 (N_31446,N_21714,N_24355);
nor U31447 (N_31447,N_21770,N_24848);
nor U31448 (N_31448,N_21617,N_29993);
xnor U31449 (N_31449,N_25807,N_27558);
or U31450 (N_31450,N_23572,N_29563);
and U31451 (N_31451,N_26599,N_20668);
nand U31452 (N_31452,N_26944,N_23629);
or U31453 (N_31453,N_23814,N_21728);
and U31454 (N_31454,N_23444,N_25242);
nand U31455 (N_31455,N_23365,N_22322);
nor U31456 (N_31456,N_21532,N_27192);
and U31457 (N_31457,N_21404,N_20498);
or U31458 (N_31458,N_23243,N_25138);
and U31459 (N_31459,N_26143,N_22080);
nor U31460 (N_31460,N_23817,N_29260);
or U31461 (N_31461,N_22717,N_25367);
nand U31462 (N_31462,N_29756,N_29511);
and U31463 (N_31463,N_28201,N_25366);
nor U31464 (N_31464,N_29965,N_20050);
nand U31465 (N_31465,N_25228,N_20331);
nand U31466 (N_31466,N_27301,N_28645);
and U31467 (N_31467,N_23569,N_23713);
nor U31468 (N_31468,N_22788,N_26600);
nand U31469 (N_31469,N_23926,N_21142);
xor U31470 (N_31470,N_24436,N_20188);
or U31471 (N_31471,N_24239,N_22596);
xor U31472 (N_31472,N_29437,N_29363);
nand U31473 (N_31473,N_20309,N_26965);
xnor U31474 (N_31474,N_23476,N_28143);
nand U31475 (N_31475,N_29853,N_25447);
nor U31476 (N_31476,N_20448,N_20265);
nor U31477 (N_31477,N_29532,N_23441);
and U31478 (N_31478,N_22437,N_25694);
nor U31479 (N_31479,N_20731,N_24327);
xnor U31480 (N_31480,N_20819,N_23745);
or U31481 (N_31481,N_23329,N_23340);
nor U31482 (N_31482,N_29577,N_28796);
nand U31483 (N_31483,N_28542,N_20449);
nor U31484 (N_31484,N_21408,N_22410);
nor U31485 (N_31485,N_20521,N_20262);
and U31486 (N_31486,N_24863,N_23272);
and U31487 (N_31487,N_29489,N_25540);
nor U31488 (N_31488,N_24795,N_24671);
and U31489 (N_31489,N_20976,N_20636);
and U31490 (N_31490,N_26230,N_21552);
nand U31491 (N_31491,N_28565,N_25653);
or U31492 (N_31492,N_27569,N_28892);
and U31493 (N_31493,N_20389,N_20589);
and U31494 (N_31494,N_20586,N_23035);
nor U31495 (N_31495,N_22207,N_29121);
nand U31496 (N_31496,N_23521,N_23840);
nand U31497 (N_31497,N_24183,N_29398);
and U31498 (N_31498,N_28902,N_28748);
nor U31499 (N_31499,N_21227,N_24279);
or U31500 (N_31500,N_23780,N_23753);
nor U31501 (N_31501,N_24001,N_22884);
or U31502 (N_31502,N_27589,N_24116);
nand U31503 (N_31503,N_23844,N_25131);
nor U31504 (N_31504,N_29765,N_23326);
or U31505 (N_31505,N_24068,N_28052);
nor U31506 (N_31506,N_25335,N_22600);
nand U31507 (N_31507,N_24345,N_22534);
or U31508 (N_31508,N_21775,N_23382);
or U31509 (N_31509,N_24960,N_26984);
or U31510 (N_31510,N_25993,N_26737);
nand U31511 (N_31511,N_23167,N_24596);
xnor U31512 (N_31512,N_28016,N_23558);
and U31513 (N_31513,N_21076,N_24263);
nor U31514 (N_31514,N_29889,N_23230);
nand U31515 (N_31515,N_29882,N_29899);
nand U31516 (N_31516,N_24565,N_25354);
nand U31517 (N_31517,N_25892,N_29278);
nor U31518 (N_31518,N_22822,N_25179);
and U31519 (N_31519,N_24542,N_22181);
or U31520 (N_31520,N_28631,N_20599);
nor U31521 (N_31521,N_24738,N_28194);
or U31522 (N_31522,N_27454,N_26087);
and U31523 (N_31523,N_22087,N_20106);
or U31524 (N_31524,N_26748,N_28734);
nor U31525 (N_31525,N_21896,N_22468);
and U31526 (N_31526,N_25884,N_21427);
nand U31527 (N_31527,N_22053,N_23429);
nand U31528 (N_31528,N_20947,N_23454);
or U31529 (N_31529,N_23608,N_29028);
nand U31530 (N_31530,N_24213,N_29048);
xor U31531 (N_31531,N_24702,N_26982);
nand U31532 (N_31532,N_20640,N_22451);
nor U31533 (N_31533,N_22569,N_27239);
and U31534 (N_31534,N_24976,N_22546);
nand U31535 (N_31535,N_26752,N_27927);
and U31536 (N_31536,N_20549,N_29686);
or U31537 (N_31537,N_20198,N_23619);
nor U31538 (N_31538,N_24997,N_23611);
nor U31539 (N_31539,N_27143,N_27596);
and U31540 (N_31540,N_23458,N_24726);
nand U31541 (N_31541,N_20105,N_28625);
or U31542 (N_31542,N_24268,N_23748);
nor U31543 (N_31543,N_24461,N_21520);
or U31544 (N_31544,N_20268,N_29948);
nor U31545 (N_31545,N_21798,N_21901);
and U31546 (N_31546,N_29091,N_20385);
nand U31547 (N_31547,N_29794,N_24677);
or U31548 (N_31548,N_29226,N_23781);
nand U31549 (N_31549,N_25753,N_26682);
and U31550 (N_31550,N_25318,N_21217);
nor U31551 (N_31551,N_22368,N_20011);
and U31552 (N_31552,N_21939,N_21174);
and U31553 (N_31553,N_25102,N_20269);
nor U31554 (N_31554,N_20535,N_29880);
and U31555 (N_31555,N_22154,N_23161);
xnor U31556 (N_31556,N_24916,N_28005);
or U31557 (N_31557,N_27530,N_28193);
and U31558 (N_31558,N_23264,N_26615);
and U31559 (N_31559,N_27058,N_21459);
and U31560 (N_31560,N_29420,N_29227);
or U31561 (N_31561,N_29395,N_23670);
and U31562 (N_31562,N_23297,N_21977);
nand U31563 (N_31563,N_28705,N_20256);
and U31564 (N_31564,N_24477,N_22474);
and U31565 (N_31565,N_26606,N_20055);
and U31566 (N_31566,N_26055,N_29507);
and U31567 (N_31567,N_21995,N_28891);
and U31568 (N_31568,N_24967,N_28546);
nand U31569 (N_31569,N_23912,N_21154);
or U31570 (N_31570,N_22810,N_29989);
or U31571 (N_31571,N_29130,N_24880);
nand U31572 (N_31572,N_25925,N_20229);
or U31573 (N_31573,N_23003,N_21171);
and U31574 (N_31574,N_24931,N_27924);
nor U31575 (N_31575,N_22093,N_22937);
nand U31576 (N_31576,N_21131,N_26660);
or U31577 (N_31577,N_28956,N_22999);
xor U31578 (N_31578,N_23403,N_25727);
nand U31579 (N_31579,N_22282,N_28190);
xor U31580 (N_31580,N_20839,N_26017);
nor U31581 (N_31581,N_21479,N_25654);
nand U31582 (N_31582,N_24487,N_27556);
nor U31583 (N_31583,N_26575,N_28964);
and U31584 (N_31584,N_25683,N_26028);
or U31585 (N_31585,N_27682,N_20122);
or U31586 (N_31586,N_26173,N_22969);
and U31587 (N_31587,N_24539,N_26810);
nor U31588 (N_31588,N_20136,N_27853);
xnor U31589 (N_31589,N_22983,N_25666);
nand U31590 (N_31590,N_25432,N_23275);
and U31591 (N_31591,N_25548,N_22270);
or U31592 (N_31592,N_22083,N_21272);
nand U31593 (N_31593,N_28879,N_26865);
nor U31594 (N_31594,N_23406,N_28700);
nor U31595 (N_31595,N_21932,N_26841);
xor U31596 (N_31596,N_23322,N_21561);
nand U31597 (N_31597,N_20437,N_24282);
xor U31598 (N_31598,N_26533,N_29967);
nand U31599 (N_31599,N_21748,N_29105);
and U31600 (N_31600,N_22735,N_20988);
and U31601 (N_31601,N_23527,N_25974);
xor U31602 (N_31602,N_23130,N_28126);
nand U31603 (N_31603,N_28990,N_29143);
nor U31604 (N_31604,N_23524,N_25369);
nor U31605 (N_31605,N_27416,N_26711);
or U31606 (N_31606,N_27482,N_25247);
nand U31607 (N_31607,N_28348,N_27703);
and U31608 (N_31608,N_29414,N_28529);
nor U31609 (N_31609,N_23597,N_26210);
nand U31610 (N_31610,N_23542,N_24467);
or U31611 (N_31611,N_20711,N_25668);
and U31612 (N_31612,N_27813,N_20941);
and U31613 (N_31613,N_28831,N_26163);
or U31614 (N_31614,N_22493,N_25020);
or U31615 (N_31615,N_24209,N_25563);
and U31616 (N_31616,N_21907,N_21606);
and U31617 (N_31617,N_25569,N_28370);
nor U31618 (N_31618,N_25427,N_28714);
nor U31619 (N_31619,N_21238,N_23941);
and U31620 (N_31620,N_23086,N_28086);
nor U31621 (N_31621,N_21360,N_28777);
or U31622 (N_31622,N_29902,N_20573);
nor U31623 (N_31623,N_20012,N_27809);
or U31624 (N_31624,N_26776,N_20812);
nand U31625 (N_31625,N_25669,N_29205);
xor U31626 (N_31626,N_27298,N_21777);
nor U31627 (N_31627,N_28254,N_24917);
nand U31628 (N_31628,N_21892,N_22243);
or U31629 (N_31629,N_26755,N_28851);
or U31630 (N_31630,N_24672,N_24172);
nand U31631 (N_31631,N_24856,N_25322);
or U31632 (N_31632,N_26200,N_28590);
or U31633 (N_31633,N_27024,N_28174);
and U31634 (N_31634,N_22863,N_21067);
or U31635 (N_31635,N_23357,N_29510);
or U31636 (N_31636,N_27345,N_25655);
or U31637 (N_31637,N_25646,N_22628);
or U31638 (N_31638,N_24575,N_23478);
xor U31639 (N_31639,N_21376,N_24180);
xor U31640 (N_31640,N_20470,N_27228);
nand U31641 (N_31641,N_25409,N_26096);
and U31642 (N_31642,N_25078,N_25024);
and U31643 (N_31643,N_25568,N_21657);
or U31644 (N_31644,N_24156,N_29703);
nor U31645 (N_31645,N_24473,N_20875);
or U31646 (N_31646,N_21409,N_21538);
nand U31647 (N_31647,N_23559,N_28247);
nor U31648 (N_31648,N_21335,N_29147);
nand U31649 (N_31649,N_23017,N_25271);
xnor U31650 (N_31650,N_25406,N_25740);
or U31651 (N_31651,N_26506,N_25444);
and U31652 (N_31652,N_20824,N_26378);
nor U31653 (N_31653,N_22116,N_23774);
nor U31654 (N_31654,N_27112,N_28845);
nor U31655 (N_31655,N_25726,N_22433);
and U31656 (N_31656,N_25863,N_23334);
nor U31657 (N_31657,N_21889,N_29070);
and U31658 (N_31658,N_20241,N_21420);
nand U31659 (N_31659,N_21744,N_24242);
nor U31660 (N_31660,N_25592,N_22082);
or U31661 (N_31661,N_28121,N_28741);
xnor U31662 (N_31662,N_25968,N_26197);
or U31663 (N_31663,N_24284,N_26625);
xor U31664 (N_31664,N_21778,N_24238);
nor U31665 (N_31665,N_26883,N_22502);
or U31666 (N_31666,N_26125,N_25278);
or U31667 (N_31667,N_26853,N_20934);
xor U31668 (N_31668,N_25133,N_21591);
nor U31669 (N_31669,N_26301,N_22321);
xnor U31670 (N_31670,N_25868,N_28253);
xnor U31671 (N_31671,N_27207,N_22762);
nand U31672 (N_31672,N_24797,N_22623);
and U31673 (N_31673,N_22004,N_27354);
or U31674 (N_31674,N_23106,N_25199);
and U31675 (N_31675,N_22665,N_27476);
nor U31676 (N_31676,N_25951,N_27283);
xor U31677 (N_31677,N_28158,N_20363);
and U31678 (N_31678,N_25321,N_29822);
and U31679 (N_31679,N_22565,N_24512);
and U31680 (N_31680,N_28502,N_20931);
or U31681 (N_31681,N_21668,N_22487);
and U31682 (N_31682,N_28539,N_24244);
xnor U31683 (N_31683,N_24144,N_22722);
xor U31684 (N_31684,N_21084,N_28428);
nor U31685 (N_31685,N_22772,N_25464);
nand U31686 (N_31686,N_24154,N_22834);
nand U31687 (N_31687,N_25789,N_25032);
nor U31688 (N_31688,N_20460,N_20495);
and U31689 (N_31689,N_29982,N_23562);
and U31690 (N_31690,N_24896,N_20539);
and U31691 (N_31691,N_24184,N_23420);
and U31692 (N_31692,N_23948,N_22091);
xnor U31693 (N_31693,N_26995,N_27767);
nand U31694 (N_31694,N_22191,N_27224);
nand U31695 (N_31695,N_23739,N_21386);
or U31696 (N_31696,N_28841,N_22400);
and U31697 (N_31697,N_28433,N_26837);
and U31698 (N_31698,N_27053,N_20652);
or U31699 (N_31699,N_26765,N_26993);
and U31700 (N_31700,N_23838,N_22375);
xor U31701 (N_31701,N_26350,N_24225);
nor U31702 (N_31702,N_20223,N_25070);
nand U31703 (N_31703,N_24750,N_29592);
or U31704 (N_31704,N_23951,N_26957);
nor U31705 (N_31705,N_23236,N_26848);
xnor U31706 (N_31706,N_27033,N_21221);
nand U31707 (N_31707,N_29719,N_21960);
or U31708 (N_31708,N_21908,N_25361);
or U31709 (N_31709,N_27396,N_29231);
xnor U31710 (N_31710,N_21482,N_25042);
or U31711 (N_31711,N_20721,N_21458);
nor U31712 (N_31712,N_25788,N_24818);
or U31713 (N_31713,N_28178,N_24534);
nor U31714 (N_31714,N_22070,N_21116);
nor U31715 (N_31715,N_21874,N_23944);
nor U31716 (N_31716,N_29486,N_20890);
xor U31717 (N_31717,N_29916,N_28438);
nor U31718 (N_31718,N_28451,N_28719);
and U31719 (N_31719,N_24521,N_25972);
and U31720 (N_31720,N_27663,N_28098);
xnor U31721 (N_31721,N_23773,N_20334);
nor U31722 (N_31722,N_25860,N_26454);
and U31723 (N_31723,N_20677,N_29908);
and U31724 (N_31724,N_22723,N_23675);
nand U31725 (N_31725,N_22634,N_23381);
xnor U31726 (N_31726,N_24431,N_26433);
or U31727 (N_31727,N_21856,N_27707);
or U31728 (N_31728,N_25210,N_20478);
and U31729 (N_31729,N_26179,N_25986);
nor U31730 (N_31730,N_27583,N_28728);
nor U31731 (N_31731,N_28349,N_26980);
xor U31732 (N_31732,N_26393,N_20117);
nor U31733 (N_31733,N_25712,N_24120);
nand U31734 (N_31734,N_26960,N_20515);
nor U31735 (N_31735,N_21690,N_20294);
nand U31736 (N_31736,N_22016,N_23962);
or U31737 (N_31737,N_20015,N_23868);
or U31738 (N_31738,N_22689,N_28248);
or U31739 (N_31739,N_24941,N_29079);
or U31740 (N_31740,N_20671,N_29482);
nor U31741 (N_31741,N_20553,N_25888);
and U31742 (N_31742,N_20520,N_20613);
nor U31743 (N_31743,N_21811,N_24930);
and U31744 (N_31744,N_21658,N_24708);
or U31745 (N_31745,N_26427,N_23091);
xnor U31746 (N_31746,N_27303,N_29562);
or U31747 (N_31747,N_29265,N_26423);
or U31748 (N_31748,N_21241,N_24468);
nand U31749 (N_31749,N_25236,N_23551);
xor U31750 (N_31750,N_23615,N_29570);
and U31751 (N_31751,N_22411,N_26661);
and U31752 (N_31752,N_25028,N_22871);
nor U31753 (N_31753,N_28184,N_28405);
and U31754 (N_31754,N_25667,N_27302);
nand U31755 (N_31755,N_26453,N_22655);
nand U31756 (N_31756,N_28319,N_25864);
and U31757 (N_31757,N_27213,N_29535);
and U31758 (N_31758,N_22244,N_29829);
or U31759 (N_31759,N_23734,N_27364);
or U31760 (N_31760,N_28458,N_29602);
and U31761 (N_31761,N_28795,N_20985);
and U31762 (N_31762,N_28120,N_21295);
nor U31763 (N_31763,N_20038,N_26151);
and U31764 (N_31764,N_22199,N_28871);
nand U31765 (N_31765,N_28093,N_23304);
and U31766 (N_31766,N_27677,N_25504);
nand U31767 (N_31767,N_21006,N_21315);
xnor U31768 (N_31768,N_28722,N_26323);
and U31769 (N_31769,N_28063,N_28660);
nor U31770 (N_31770,N_28657,N_20878);
and U31771 (N_31771,N_24845,N_28793);
or U31772 (N_31772,N_27272,N_28792);
xnor U31773 (N_31773,N_22536,N_20883);
xor U31774 (N_31774,N_25596,N_22219);
nor U31775 (N_31775,N_27549,N_20899);
nor U31776 (N_31776,N_20756,N_22706);
nand U31777 (N_31777,N_26902,N_25065);
or U31778 (N_31778,N_23983,N_26874);
or U31779 (N_31779,N_22514,N_24912);
nor U31780 (N_31780,N_26635,N_27834);
or U31781 (N_31781,N_24954,N_25600);
xor U31782 (N_31782,N_26259,N_21157);
or U31783 (N_31783,N_21447,N_24679);
nand U31784 (N_31784,N_27933,N_23568);
or U31785 (N_31785,N_22544,N_25613);
nor U31786 (N_31786,N_28217,N_26795);
nand U31787 (N_31787,N_28321,N_21201);
nand U31788 (N_31788,N_24266,N_20780);
or U31789 (N_31789,N_23655,N_25004);
and U31790 (N_31790,N_20349,N_20173);
xnor U31791 (N_31791,N_28332,N_27962);
or U31792 (N_31792,N_21785,N_29136);
nor U31793 (N_31793,N_20900,N_27057);
and U31794 (N_31794,N_28498,N_26315);
and U31795 (N_31795,N_25570,N_27936);
and U31796 (N_31796,N_24191,N_21106);
nor U31797 (N_31797,N_23977,N_23481);
and U31798 (N_31798,N_28425,N_23984);
or U31799 (N_31799,N_29937,N_28814);
nand U31800 (N_31800,N_26249,N_20042);
xnor U31801 (N_31801,N_27285,N_26104);
and U31802 (N_31802,N_29742,N_22308);
nand U31803 (N_31803,N_26832,N_28626);
and U31804 (N_31804,N_29192,N_29436);
xor U31805 (N_31805,N_27886,N_24390);
nor U31806 (N_31806,N_26571,N_26734);
and U31807 (N_31807,N_28456,N_25622);
nand U31808 (N_31808,N_21302,N_20406);
nor U31809 (N_31809,N_20411,N_20724);
nand U31810 (N_31810,N_23490,N_22030);
nor U31811 (N_31811,N_29957,N_23215);
and U31812 (N_31812,N_24309,N_22003);
and U31813 (N_31813,N_23129,N_25841);
nor U31814 (N_31814,N_25551,N_29648);
nand U31815 (N_31815,N_28361,N_24875);
nor U31816 (N_31816,N_23134,N_26290);
nand U31817 (N_31817,N_29149,N_27762);
nor U31818 (N_31818,N_20238,N_26974);
and U31819 (N_31819,N_24256,N_23177);
nand U31820 (N_31820,N_20637,N_27774);
nor U31821 (N_31821,N_24721,N_29410);
or U31822 (N_31822,N_25577,N_24453);
nor U31823 (N_31823,N_21159,N_23299);
nor U31824 (N_31824,N_25531,N_24109);
nor U31825 (N_31825,N_24071,N_22390);
xnor U31826 (N_31826,N_20867,N_26419);
or U31827 (N_31827,N_23273,N_28345);
nand U31828 (N_31828,N_27468,N_22309);
nor U31829 (N_31829,N_26044,N_29142);
nand U31830 (N_31830,N_21428,N_20872);
xor U31831 (N_31831,N_21935,N_24084);
nand U31832 (N_31832,N_25528,N_24140);
nor U31833 (N_31833,N_20335,N_25844);
nor U31834 (N_31834,N_24645,N_25602);
xor U31835 (N_31835,N_29872,N_20130);
nand U31836 (N_31836,N_29297,N_24929);
or U31837 (N_31837,N_23282,N_22676);
nand U31838 (N_31838,N_22175,N_20852);
xnor U31839 (N_31839,N_29878,N_26766);
and U31840 (N_31840,N_22314,N_23543);
nor U31841 (N_31841,N_25005,N_27532);
or U31842 (N_31842,N_29096,N_21509);
nor U31843 (N_31843,N_24375,N_21542);
nand U31844 (N_31844,N_22196,N_28910);
and U31845 (N_31845,N_24227,N_24927);
nor U31846 (N_31846,N_27008,N_27595);
or U31847 (N_31847,N_23298,N_28787);
nand U31848 (N_31848,N_23139,N_24578);
nand U31849 (N_31849,N_25315,N_24695);
nor U31850 (N_31850,N_20725,N_22296);
nor U31851 (N_31851,N_21857,N_27212);
nor U31852 (N_31852,N_29356,N_24342);
and U31853 (N_31853,N_29508,N_29939);
nand U31854 (N_31854,N_27335,N_28353);
and U31855 (N_31855,N_24000,N_25428);
nand U31856 (N_31856,N_21001,N_29148);
or U31857 (N_31857,N_25414,N_25507);
nand U31858 (N_31858,N_28010,N_20981);
nor U31859 (N_31859,N_29798,N_23442);
xor U31860 (N_31860,N_20590,N_29986);
xnor U31861 (N_31861,N_21577,N_29443);
nand U31862 (N_31862,N_28775,N_28030);
nor U31863 (N_31863,N_23915,N_25463);
and U31864 (N_31864,N_22285,N_23826);
xor U31865 (N_31865,N_22496,N_21750);
nor U31866 (N_31866,N_29581,N_24811);
and U31867 (N_31867,N_28334,N_25642);
and U31868 (N_31868,N_24166,N_27430);
nor U31869 (N_31869,N_20299,N_21550);
nand U31870 (N_31870,N_20723,N_27460);
nand U31871 (N_31871,N_26477,N_27084);
nor U31872 (N_31872,N_29789,N_23190);
nand U31873 (N_31873,N_20143,N_20024);
nor U31874 (N_31874,N_20956,N_29886);
or U31875 (N_31875,N_27380,N_25855);
and U31876 (N_31876,N_25268,N_27847);
or U31877 (N_31877,N_25736,N_29487);
xor U31878 (N_31878,N_23184,N_23255);
and U31879 (N_31879,N_29555,N_23682);
or U31880 (N_31880,N_27230,N_25609);
xnor U31881 (N_31881,N_26603,N_20776);
nor U31882 (N_31882,N_24712,N_26185);
xor U31883 (N_31883,N_23088,N_24594);
nor U31884 (N_31884,N_28421,N_24403);
xnor U31885 (N_31885,N_26400,N_20373);
nand U31886 (N_31886,N_23276,N_24755);
and U31887 (N_31887,N_29302,N_27350);
nor U31888 (N_31888,N_28561,N_20444);
nor U31889 (N_31889,N_20841,N_21416);
or U31890 (N_31890,N_29697,N_29210);
or U31891 (N_31891,N_27204,N_28966);
nand U31892 (N_31892,N_29552,N_21075);
or U31893 (N_31893,N_25057,N_25233);
nand U31894 (N_31894,N_25578,N_25310);
nor U31895 (N_31895,N_26146,N_29208);
and U31896 (N_31896,N_26787,N_21091);
xor U31897 (N_31897,N_20664,N_21382);
and U31898 (N_31898,N_29383,N_27109);
nand U31899 (N_31899,N_20204,N_23677);
or U31900 (N_31900,N_27363,N_20361);
nand U31901 (N_31901,N_27769,N_22961);
nor U31902 (N_31902,N_26736,N_23148);
nand U31903 (N_31903,N_22533,N_25589);
nor U31904 (N_31904,N_24910,N_29293);
nor U31905 (N_31905,N_24313,N_28236);
or U31906 (N_31906,N_29600,N_26263);
nand U31907 (N_31907,N_27226,N_29428);
nand U31908 (N_31908,N_20350,N_21784);
xor U31909 (N_31909,N_29094,N_27193);
nor U31910 (N_31910,N_24809,N_22306);
and U31911 (N_31911,N_21819,N_25292);
and U31912 (N_31912,N_24017,N_27771);
or U31913 (N_31913,N_24868,N_29051);
nor U31914 (N_31914,N_25590,N_27487);
nand U31915 (N_31915,N_27326,N_26214);
nand U31916 (N_31916,N_28874,N_26785);
or U31917 (N_31917,N_24240,N_26979);
and U31918 (N_31918,N_26548,N_21068);
and U31919 (N_31919,N_22550,N_25364);
or U31920 (N_31920,N_25839,N_21367);
nand U31921 (N_31921,N_25263,N_29022);
and U31922 (N_31922,N_27052,N_27047);
nor U31923 (N_31923,N_27152,N_25588);
and U31924 (N_31924,N_26654,N_21845);
or U31925 (N_31925,N_25717,N_26366);
and U31926 (N_31926,N_25767,N_23979);
and U31927 (N_31927,N_21329,N_28061);
or U31928 (N_31928,N_25400,N_24611);
or U31929 (N_31929,N_23876,N_25865);
and U31930 (N_31930,N_25225,N_21361);
nand U31931 (N_31931,N_25911,N_21094);
nor U31932 (N_31932,N_23980,N_23325);
nor U31933 (N_31933,N_20660,N_20936);
nand U31934 (N_31934,N_23141,N_24045);
and U31935 (N_31935,N_22957,N_25854);
nor U31936 (N_31936,N_25935,N_25227);
nand U31937 (N_31937,N_24505,N_26127);
nand U31938 (N_31938,N_20667,N_24970);
xor U31939 (N_31939,N_26313,N_21942);
xor U31940 (N_31940,N_28047,N_27211);
and U31941 (N_31941,N_23337,N_28960);
and U31942 (N_31942,N_20276,N_28003);
or U31943 (N_31943,N_20108,N_22235);
or U31944 (N_31944,N_21964,N_21787);
xnor U31945 (N_31945,N_20610,N_22703);
nand U31946 (N_31946,N_24730,N_22813);
nand U31947 (N_31947,N_21788,N_22421);
or U31948 (N_31948,N_27105,N_21220);
nor U31949 (N_31949,N_22771,N_24955);
and U31950 (N_31950,N_21356,N_29464);
and U31951 (N_31951,N_29616,N_24498);
xnor U31952 (N_31952,N_22301,N_20744);
or U31953 (N_31953,N_20399,N_28260);
or U31954 (N_31954,N_21827,N_23137);
xnor U31955 (N_31955,N_25466,N_27409);
nor U31956 (N_31956,N_27248,N_28675);
nand U31957 (N_31957,N_26462,N_20442);
and U31958 (N_31958,N_21536,N_20027);
and U31959 (N_31959,N_28088,N_27135);
nor U31960 (N_31960,N_25053,N_26642);
nor U31961 (N_31961,N_26342,N_28809);
xnor U31962 (N_31962,N_28173,N_26446);
nor U31963 (N_31963,N_21824,N_29495);
and U31964 (N_31964,N_23311,N_21461);
xnor U31965 (N_31965,N_29024,N_26749);
nor U31966 (N_31966,N_28854,N_24884);
or U31967 (N_31967,N_20020,N_28522);
or U31968 (N_31968,N_22438,N_25317);
xor U31969 (N_31969,N_26285,N_22075);
xor U31970 (N_31970,N_28844,N_20814);
xnor U31971 (N_31971,N_23644,N_25372);
nand U31972 (N_31972,N_25443,N_23261);
xor U31973 (N_31973,N_20932,N_29984);
xor U31974 (N_31974,N_28343,N_22164);
nand U31975 (N_31975,N_26025,N_25187);
nor U31976 (N_31976,N_29635,N_24200);
or U31977 (N_31977,N_21332,N_20028);
and U31978 (N_31978,N_23577,N_25319);
nor U31979 (N_31979,N_26892,N_22963);
and U31980 (N_31980,N_21497,N_22076);
xor U31981 (N_31981,N_25357,N_21855);
xor U31982 (N_31982,N_28365,N_26758);
nor U31983 (N_31983,N_24387,N_25947);
or U31984 (N_31984,N_26170,N_21629);
or U31985 (N_31985,N_20940,N_25825);
nor U31986 (N_31986,N_23313,N_20407);
and U31987 (N_31987,N_21294,N_27176);
or U31988 (N_31988,N_22670,N_28642);
nand U31989 (N_31989,N_29211,N_27470);
or U31990 (N_31990,N_26380,N_23089);
or U31991 (N_31991,N_21038,N_25505);
and U31992 (N_31992,N_22130,N_29062);
nor U31993 (N_31993,N_23156,N_21604);
or U31994 (N_31994,N_22488,N_20098);
and U31995 (N_31995,N_25099,N_25502);
or U31996 (N_31996,N_28000,N_26845);
nand U31997 (N_31997,N_29927,N_26577);
nand U31998 (N_31998,N_28750,N_20427);
and U31999 (N_31999,N_23651,N_21639);
xnor U32000 (N_32000,N_24121,N_25806);
and U32001 (N_32001,N_29183,N_23179);
or U32002 (N_32002,N_22571,N_21898);
or U32003 (N_32003,N_21170,N_26217);
and U32004 (N_32004,N_24825,N_21073);
or U32005 (N_32005,N_25631,N_24964);
or U32006 (N_32006,N_22059,N_23827);
and U32007 (N_32007,N_22029,N_26522);
or U32008 (N_32008,N_20134,N_22734);
nor U32009 (N_32009,N_21372,N_23930);
nand U32010 (N_32010,N_20123,N_24132);
and U32011 (N_32011,N_21307,N_23336);
and U32012 (N_32012,N_26094,N_21343);
nor U32013 (N_32013,N_28581,N_25962);
or U32014 (N_32014,N_24247,N_22124);
and U32015 (N_32015,N_27948,N_22584);
nor U32016 (N_32016,N_21792,N_22426);
and U32017 (N_32017,N_29554,N_29041);
nor U32018 (N_32018,N_21664,N_25014);
nor U32019 (N_32019,N_23897,N_27039);
nor U32020 (N_32020,N_21926,N_21015);
and U32021 (N_32021,N_23803,N_26406);
nand U32022 (N_32022,N_25288,N_20465);
nand U32023 (N_32023,N_28487,N_21403);
nor U32024 (N_32024,N_24494,N_24602);
nor U32025 (N_32025,N_22002,N_23854);
or U32026 (N_32026,N_23350,N_24535);
and U32027 (N_32027,N_27384,N_25877);
nand U32028 (N_32028,N_21776,N_25436);
or U32029 (N_32029,N_29919,N_26057);
and U32030 (N_32030,N_24335,N_29154);
nand U32031 (N_32031,N_26973,N_23448);
nand U32032 (N_32032,N_29934,N_29513);
and U32033 (N_32033,N_24662,N_29678);
nand U32034 (N_32034,N_29971,N_23407);
or U32035 (N_32035,N_23945,N_22133);
or U32036 (N_32036,N_22666,N_22643);
or U32037 (N_32037,N_28916,N_20516);
nand U32038 (N_32038,N_26464,N_21902);
nand U32039 (N_32039,N_20446,N_24861);
nor U32040 (N_32040,N_23623,N_28110);
and U32041 (N_32041,N_21465,N_21969);
and U32042 (N_32042,N_25426,N_28381);
and U32043 (N_32043,N_20542,N_29933);
or U32044 (N_32044,N_21147,N_21111);
nand U32045 (N_32045,N_29421,N_22312);
and U32046 (N_32046,N_26294,N_25546);
xnor U32047 (N_32047,N_23795,N_27172);
nor U32048 (N_32048,N_27751,N_24013);
xor U32049 (N_32049,N_26942,N_26421);
or U32050 (N_32050,N_20340,N_25756);
and U32051 (N_32051,N_24316,N_21431);
and U32052 (N_32052,N_24522,N_25009);
nor U32053 (N_32053,N_26649,N_20287);
nand U32054 (N_32054,N_23192,N_26697);
nor U32055 (N_32055,N_21089,N_25907);
nor U32056 (N_32056,N_20070,N_20882);
and U32057 (N_32057,N_24950,N_24384);
or U32058 (N_32058,N_23321,N_28099);
xnor U32059 (N_32059,N_29377,N_21008);
or U32060 (N_32060,N_27120,N_21793);
or U32061 (N_32061,N_20779,N_23359);
nand U32062 (N_32062,N_26208,N_25045);
nand U32063 (N_32063,N_23960,N_28599);
nor U32064 (N_32064,N_23294,N_21796);
nor U32065 (N_32065,N_29895,N_26240);
xor U32066 (N_32066,N_25813,N_28706);
nand U32067 (N_32067,N_23969,N_29985);
nor U32068 (N_32068,N_24663,N_22615);
or U32069 (N_32069,N_20075,N_27959);
nand U32070 (N_32070,N_22859,N_24581);
and U32071 (N_32071,N_26873,N_25630);
nor U32072 (N_32072,N_24393,N_28995);
or U32073 (N_32073,N_27122,N_25132);
nand U32074 (N_32074,N_29101,N_23650);
and U32075 (N_32075,N_22895,N_28799);
xor U32076 (N_32076,N_27791,N_25025);
or U32077 (N_32077,N_22237,N_23928);
or U32078 (N_32078,N_22216,N_25392);
and U32079 (N_32079,N_26386,N_21334);
nor U32080 (N_32080,N_27564,N_28517);
xnor U32081 (N_32081,N_24889,N_26192);
xnor U32082 (N_32082,N_28300,N_26154);
nand U32083 (N_32083,N_20377,N_23584);
or U32084 (N_32084,N_22155,N_22463);
nor U32085 (N_32085,N_27888,N_27091);
nand U32086 (N_32086,N_21448,N_23888);
nand U32087 (N_32087,N_22189,N_25267);
nor U32088 (N_32088,N_28216,N_21033);
or U32089 (N_32089,N_26733,N_21305);
nand U32090 (N_32090,N_20848,N_26084);
nand U32091 (N_32091,N_24476,N_24181);
nand U32092 (N_32092,N_28717,N_26959);
nand U32093 (N_32093,N_24369,N_23056);
nor U32094 (N_32094,N_22041,N_28516);
nand U32095 (N_32095,N_25559,N_21945);
and U32096 (N_32096,N_28124,N_20402);
nand U32097 (N_32097,N_23390,N_25163);
nand U32098 (N_32098,N_21319,N_21625);
nor U32099 (N_32099,N_22577,N_20675);
nand U32100 (N_32100,N_29340,N_22897);
nand U32101 (N_32101,N_28947,N_27075);
or U32102 (N_32102,N_27370,N_20251);
nand U32103 (N_32103,N_20426,N_27570);
nand U32104 (N_32104,N_23847,N_22457);
nand U32105 (N_32105,N_24462,N_25768);
nor U32106 (N_32106,N_29652,N_22630);
xnor U32107 (N_32107,N_25956,N_24482);
and U32108 (N_32108,N_21864,N_26007);
xnor U32109 (N_32109,N_29018,N_24969);
and U32110 (N_32110,N_23439,N_21670);
and U32111 (N_32111,N_25041,N_26008);
or U32112 (N_32112,N_22828,N_27263);
nor U32113 (N_32113,N_23157,N_25458);
or U32114 (N_32114,N_27290,N_21736);
nand U32115 (N_32115,N_25473,N_29611);
nor U32116 (N_32116,N_23973,N_23880);
nor U32117 (N_32117,N_22098,N_27435);
nand U32118 (N_32118,N_20189,N_25016);
nor U32119 (N_32119,N_20743,N_21873);
nor U32120 (N_32120,N_28468,N_23348);
or U32121 (N_32121,N_24855,N_29634);
or U32122 (N_32122,N_20971,N_29546);
or U32123 (N_32123,N_20970,N_20473);
nand U32124 (N_32124,N_29730,N_29894);
nand U32125 (N_32125,N_26666,N_28699);
nand U32126 (N_32126,N_21547,N_22287);
or U32127 (N_32127,N_23680,N_20325);
xnor U32128 (N_32128,N_25934,N_22273);
nand U32129 (N_32129,N_28873,N_29384);
nor U32130 (N_32130,N_28142,N_28803);
xnor U32131 (N_32131,N_20755,N_26641);
nand U32132 (N_32132,N_28740,N_21524);
nor U32133 (N_32133,N_29124,N_23833);
nand U32134 (N_32134,N_24699,N_20458);
nand U32135 (N_32135,N_22592,N_26922);
or U32136 (N_32136,N_20745,N_23286);
and U32137 (N_32137,N_27199,N_21984);
or U32138 (N_32138,N_23544,N_22010);
and U32139 (N_32139,N_25106,N_26349);
nor U32140 (N_32140,N_27662,N_26544);
or U32141 (N_32141,N_29316,N_23174);
nor U32142 (N_32142,N_23330,N_20224);
nor U32143 (N_32143,N_22572,N_25430);
xnor U32144 (N_32144,N_21123,N_25685);
nand U32145 (N_32145,N_20327,N_20991);
and U32146 (N_32146,N_25698,N_26729);
or U32147 (N_32147,N_29823,N_26932);
nand U32148 (N_32148,N_20778,N_29311);
nand U32149 (N_32149,N_27999,N_27737);
xor U32150 (N_32150,N_23789,N_29256);
or U32151 (N_32151,N_21436,N_23741);
nor U32152 (N_32152,N_24735,N_28368);
nor U32153 (N_32153,N_28275,N_27404);
nor U32154 (N_32154,N_20356,N_20160);
and U32155 (N_32155,N_26964,N_21444);
nor U32156 (N_32156,N_21151,N_27845);
or U32157 (N_32157,N_26488,N_28327);
xnor U32158 (N_32158,N_25254,N_29785);
and U32159 (N_32159,N_21944,N_20090);
nand U32160 (N_32160,N_28259,N_24077);
nor U32161 (N_32161,N_29132,N_24014);
or U32162 (N_32162,N_28952,N_20914);
nand U32163 (N_32163,N_24118,N_28357);
and U32164 (N_32164,N_20567,N_28936);
nor U32165 (N_32165,N_27334,N_21499);
or U32166 (N_32166,N_21663,N_22037);
and U32167 (N_32167,N_26819,N_21096);
nor U32168 (N_32168,N_23465,N_27318);
xor U32169 (N_32169,N_29339,N_22141);
nand U32170 (N_32170,N_21624,N_27136);
or U32171 (N_32171,N_26975,N_27339);
nor U32172 (N_32172,N_25424,N_25769);
or U32173 (N_32173,N_27900,N_29151);
or U32174 (N_32174,N_20393,N_20126);
nor U32175 (N_32175,N_27369,N_29090);
nand U32176 (N_32176,N_20507,N_28196);
nand U32177 (N_32177,N_29664,N_22239);
xor U32178 (N_32178,N_21992,N_28095);
and U32179 (N_32179,N_27513,N_28441);
nor U32180 (N_32180,N_21613,N_21650);
or U32181 (N_32181,N_23462,N_22588);
or U32182 (N_32182,N_28686,N_29746);
xor U32183 (N_32183,N_20678,N_26679);
nand U32184 (N_32184,N_21452,N_21753);
and U32185 (N_32185,N_29342,N_28762);
nor U32186 (N_32186,N_24259,N_20565);
and U32187 (N_32187,N_24255,N_28430);
or U32188 (N_32188,N_21397,N_26073);
or U32189 (N_32189,N_25164,N_23121);
or U32190 (N_32190,N_28909,N_20043);
nand U32191 (N_32191,N_20033,N_22261);
xnor U32192 (N_32192,N_26357,N_25912);
or U32193 (N_32193,N_24103,N_29582);
and U32194 (N_32194,N_23132,N_21172);
nor U32195 (N_32195,N_26847,N_26254);
nor U32196 (N_32196,N_23360,N_20172);
and U32197 (N_32197,N_29572,N_28883);
nor U32198 (N_32198,N_20700,N_22230);
nand U32199 (N_32199,N_27824,N_23550);
nor U32200 (N_32200,N_25710,N_28582);
and U32201 (N_32201,N_24033,N_26404);
or U32202 (N_32202,N_25983,N_28687);
nor U32203 (N_32203,N_21572,N_28586);
or U32204 (N_32204,N_27395,N_29987);
or U32205 (N_32205,N_21090,N_23909);
nor U32206 (N_32206,N_27501,N_22255);
nand U32207 (N_32207,N_20920,N_29598);
or U32208 (N_32208,N_24918,N_24711);
or U32209 (N_32209,N_22657,N_20321);
nand U32210 (N_32210,N_26503,N_28907);
nor U32211 (N_32211,N_21567,N_22204);
xnor U32212 (N_32212,N_23408,N_29928);
nand U32213 (N_32213,N_27568,N_26963);
and U32214 (N_32214,N_29646,N_22795);
nand U32215 (N_32215,N_28745,N_20488);
nand U32216 (N_32216,N_24415,N_27472);
and U32217 (N_32217,N_25178,N_23117);
nor U32218 (N_32218,N_20503,N_25103);
xor U32219 (N_32219,N_25673,N_28083);
nor U32220 (N_32220,N_27637,N_28135);
or U32221 (N_32221,N_29918,N_24879);
nand U32222 (N_32222,N_25729,N_28263);
nor U32223 (N_32223,N_25759,N_24873);
and U32224 (N_32224,N_28018,N_27638);
nand U32225 (N_32225,N_27311,N_24165);
nor U32226 (N_32226,N_25999,N_25435);
nand U32227 (N_32227,N_21725,N_20910);
nand U32228 (N_32228,N_26909,N_26016);
nor U32229 (N_32229,N_24029,N_26759);
or U32230 (N_32230,N_22120,N_22607);
and U32231 (N_32231,N_20651,N_28679);
xor U32232 (N_32232,N_26640,N_23314);
and U32233 (N_32233,N_24965,N_21250);
xor U32234 (N_32234,N_23499,N_28379);
nand U32235 (N_32235,N_23188,N_27700);
and U32236 (N_32236,N_26418,N_28043);
nor U32237 (N_32237,N_29955,N_26514);
nor U32238 (N_32238,N_22878,N_22904);
nand U32239 (N_32239,N_29963,N_22328);
and U32240 (N_32240,N_24195,N_26121);
or U32241 (N_32241,N_23968,N_22475);
and U32242 (N_32242,N_28352,N_22061);
nand U32243 (N_32243,N_28338,N_21162);
nor U32244 (N_32244,N_26298,N_24402);
xor U32245 (N_32245,N_22344,N_29906);
or U32246 (N_32246,N_24692,N_23633);
nand U32247 (N_32247,N_25678,N_24059);
nand U32248 (N_32248,N_27281,N_23618);
nand U32249 (N_32249,N_24437,N_24133);
nor U32250 (N_32250,N_22089,N_27444);
and U32251 (N_32251,N_29644,N_27654);
and U32252 (N_32252,N_26367,N_23393);
nor U32253 (N_32253,N_29429,N_29111);
and U32254 (N_32254,N_20181,N_26108);
or U32255 (N_32255,N_28858,N_29177);
xnor U32256 (N_32256,N_20245,N_24408);
and U32257 (N_32257,N_28443,N_20357);
nand U32258 (N_32258,N_27262,N_28768);
and U32259 (N_32259,N_23594,N_26943);
nor U32260 (N_32260,N_22960,N_26620);
nand U32261 (N_32261,N_20646,N_22872);
nand U32262 (N_32262,N_24822,N_21794);
and U32263 (N_32263,N_22006,N_23280);
and U32264 (N_32264,N_23564,N_29988);
or U32265 (N_32265,N_27856,N_21816);
nor U32266 (N_32266,N_20558,N_29259);
or U32267 (N_32267,N_22537,N_26582);
nor U32268 (N_32268,N_24821,N_24315);
nor U32269 (N_32269,N_21341,N_22473);
nand U32270 (N_32270,N_29220,N_29734);
or U32271 (N_32271,N_20928,N_29334);
or U32272 (N_32272,N_23296,N_27783);
xor U32273 (N_32273,N_25001,N_22028);
nand U32274 (N_32274,N_29804,N_28594);
xnor U32275 (N_32275,N_20472,N_21828);
nor U32276 (N_32276,N_20806,N_28820);
or U32277 (N_32277,N_26158,N_27849);
or U32278 (N_32278,N_20762,N_25058);
nor U32279 (N_32279,N_27810,N_25827);
and U32280 (N_32280,N_23656,N_27319);
nand U32281 (N_32281,N_21473,N_26333);
nor U32282 (N_32282,N_23209,N_25601);
and U32283 (N_32283,N_26299,N_25313);
and U32284 (N_32284,N_21244,N_28413);
nor U32285 (N_32285,N_27977,N_21133);
and U32286 (N_32286,N_28289,N_28429);
nand U32287 (N_32287,N_29034,N_26396);
xor U32288 (N_32288,N_25805,N_26881);
or U32289 (N_32289,N_24966,N_23707);
nor U32290 (N_32290,N_28039,N_27544);
nand U32291 (N_32291,N_22785,N_22316);
nand U32292 (N_32292,N_21007,N_29317);
or U32293 (N_32293,N_26461,N_29270);
and U32294 (N_32294,N_29040,N_22233);
and U32295 (N_32295,N_27934,N_21605);
nand U32296 (N_32296,N_20973,N_25445);
nor U32297 (N_32297,N_20524,N_23953);
nor U32298 (N_32298,N_20894,N_24168);
xnor U32299 (N_32299,N_26851,N_22346);
or U32300 (N_32300,N_22905,N_25165);
nor U32301 (N_32301,N_22916,N_28962);
and U32302 (N_32302,N_26053,N_28754);
or U32303 (N_32303,N_29753,N_29038);
xor U32304 (N_32304,N_27963,N_26431);
nand U32305 (N_32305,N_25459,N_29691);
nor U32306 (N_32306,N_24091,N_26074);
nor U32307 (N_32307,N_20676,N_23405);
nand U32308 (N_32308,N_21914,N_27879);
or U32309 (N_32309,N_28798,N_21808);
nand U32310 (N_32310,N_24658,N_21695);
and U32311 (N_32311,N_25852,N_27445);
nand U32312 (N_32312,N_25334,N_28442);
or U32313 (N_32313,N_28680,N_26250);
nor U32314 (N_32314,N_27150,N_24802);
and U32315 (N_32315,N_25140,N_29364);
nor U32316 (N_32316,N_21346,N_25701);
nand U32317 (N_32317,N_26086,N_23961);
and U32318 (N_32318,N_23074,N_23092);
nor U32319 (N_32319,N_25498,N_21206);
or U32320 (N_32320,N_28761,N_24122);
nand U32321 (N_32321,N_28863,N_22169);
or U32322 (N_32322,N_26003,N_26608);
nand U32323 (N_32323,N_22933,N_23504);
and U32324 (N_32324,N_28420,N_28685);
nor U32325 (N_32325,N_26334,N_21344);
or U32326 (N_32326,N_26807,N_27540);
and U32327 (N_32327,N_22469,N_27169);
or U32328 (N_32328,N_23109,N_28408);
and U32329 (N_32329,N_23186,N_26778);
or U32330 (N_32330,N_23083,N_24339);
nor U32331 (N_32331,N_20536,N_28262);
xor U32332 (N_32332,N_21897,N_22324);
and U32333 (N_32333,N_20939,N_23959);
nor U32334 (N_32334,N_23946,N_23050);
or U32335 (N_32335,N_25857,N_26392);
and U32336 (N_32336,N_27090,N_25249);
or U32337 (N_32337,N_24441,N_21688);
and U32338 (N_32338,N_21543,N_27328);
and U32339 (N_32339,N_24130,N_22482);
xor U32340 (N_32340,N_23515,N_22804);
or U32341 (N_32341,N_25499,N_25044);
nand U32342 (N_32342,N_26527,N_27089);
xnor U32343 (N_32343,N_20457,N_21715);
nor U32344 (N_32344,N_21833,N_28501);
and U32345 (N_32345,N_23914,N_24926);
or U32346 (N_32346,N_28815,N_26773);
nand U32347 (N_32347,N_20737,N_27870);
nand U32348 (N_32348,N_25324,N_28549);
and U32349 (N_32349,N_25515,N_27561);
or U32350 (N_32350,N_20781,N_25704);
nor U32351 (N_32351,N_28866,N_22824);
xor U32352 (N_32352,N_21514,N_21369);
nor U32353 (N_32353,N_23792,N_26703);
nand U32354 (N_32354,N_21941,N_27926);
and U32355 (N_32355,N_26562,N_29323);
or U32356 (N_32356,N_23557,N_21849);
and U32357 (N_32357,N_24837,N_23927);
nand U32358 (N_32358,N_26636,N_25987);
nand U32359 (N_32359,N_26497,N_29417);
nand U32360 (N_32360,N_23992,N_26602);
and U32361 (N_32361,N_21599,N_21092);
nor U32362 (N_32362,N_24508,N_27780);
nand U32363 (N_32363,N_29233,N_26051);
nand U32364 (N_32364,N_23869,N_25115);
nor U32365 (N_32365,N_25946,N_28014);
and U32366 (N_32366,N_23816,N_23908);
nand U32367 (N_32367,N_21152,N_25482);
or U32368 (N_32368,N_25295,N_25234);
nor U32369 (N_32369,N_28558,N_27492);
nand U32370 (N_32370,N_29865,N_22049);
or U32371 (N_32371,N_21786,N_25535);
nor U32372 (N_32372,N_21130,N_26705);
and U32373 (N_32373,N_29595,N_25095);
nand U32374 (N_32374,N_29499,N_22573);
nand U32375 (N_32375,N_28972,N_23284);
nor U32376 (N_32376,N_22033,N_26829);
nand U32377 (N_32377,N_27327,N_26683);
or U32378 (N_32378,N_21875,N_23694);
nor U32379 (N_32379,N_26221,N_21192);
or U32380 (N_32380,N_23461,N_25304);
nand U32381 (N_32381,N_22288,N_29005);
nand U32382 (N_32382,N_20336,N_21055);
xor U32383 (N_32383,N_29298,N_25291);
and U32384 (N_32384,N_22404,N_27986);
and U32385 (N_32385,N_22429,N_22987);
nand U32386 (N_32386,N_23859,N_20378);
nor U32387 (N_32387,N_22476,N_27484);
nor U32388 (N_32388,N_25422,N_25231);
nor U32389 (N_32389,N_21840,N_26174);
and U32390 (N_32390,N_26387,N_25985);
nor U32391 (N_32391,N_25995,N_26864);
and U32392 (N_32392,N_26843,N_24220);
nand U32393 (N_32393,N_20773,N_24869);
nand U32394 (N_32394,N_26469,N_29412);
or U32395 (N_32395,N_22140,N_24370);
xor U32396 (N_32396,N_23065,N_24189);
nand U32397 (N_32397,N_23263,N_25471);
nand U32398 (N_32398,N_27491,N_26656);
and U32399 (N_32399,N_26676,N_25468);
nor U32400 (N_32400,N_27831,N_20492);
nor U32401 (N_32401,N_20545,N_22767);
nor U32402 (N_32402,N_22677,N_26751);
or U32403 (N_32403,N_26912,N_28378);
or U32404 (N_32404,N_23843,N_27216);
or U32405 (N_32405,N_26330,N_27218);
or U32406 (N_32406,N_20107,N_22054);
or U32407 (N_32407,N_28060,N_21852);
and U32408 (N_32408,N_27620,N_25122);
and U32409 (N_32409,N_21619,N_24430);
and U32410 (N_32410,N_20079,N_27794);
and U32411 (N_32411,N_24556,N_26408);
or U32412 (N_32412,N_25745,N_22292);
xor U32413 (N_32413,N_23339,N_28573);
nor U32414 (N_32414,N_27777,N_25260);
and U32415 (N_32415,N_27913,N_26038);
and U32416 (N_32416,N_24301,N_21809);
nor U32417 (N_32417,N_22701,N_29372);
xor U32418 (N_32418,N_22721,N_27171);
and U32419 (N_32419,N_23471,N_20694);
and U32420 (N_32420,N_25721,N_21136);
or U32421 (N_32421,N_27007,N_20434);
nand U32422 (N_32422,N_28704,N_26994);
xor U32423 (N_32423,N_24624,N_21620);
nor U32424 (N_32424,N_27220,N_20255);
nand U32425 (N_32425,N_27965,N_28951);
or U32426 (N_32426,N_24742,N_26289);
and U32427 (N_32427,N_26931,N_23113);
nand U32428 (N_32428,N_21676,N_22617);
and U32429 (N_32429,N_24112,N_24895);
xnor U32430 (N_32430,N_22222,N_20805);
nor U32431 (N_32431,N_23013,N_21028);
nand U32432 (N_32432,N_27984,N_21733);
nor U32433 (N_32433,N_23131,N_28183);
nand U32434 (N_32434,N_22501,N_23836);
nand U32435 (N_32435,N_23723,N_25437);
nand U32436 (N_32436,N_26052,N_28855);
nor U32437 (N_32437,N_28225,N_21832);
nor U32438 (N_32438,N_27516,N_29722);
and U32439 (N_32439,N_29168,N_28861);
and U32440 (N_32440,N_25312,N_22280);
and U32441 (N_32441,N_24618,N_26698);
and U32442 (N_32442,N_23554,N_24517);
and U32443 (N_32443,N_29013,N_24740);
nand U32444 (N_32444,N_26763,N_29831);
nand U32445 (N_32445,N_29743,N_21443);
nand U32446 (N_32446,N_23873,N_26088);
nand U32447 (N_32447,N_24364,N_29193);
nor U32448 (N_32448,N_28612,N_29879);
nor U32449 (N_32449,N_24357,N_28608);
and U32450 (N_32450,N_22225,N_24942);
and U32451 (N_32451,N_22380,N_29583);
and U32452 (N_32452,N_26130,N_28540);
nand U32453 (N_32453,N_22480,N_26122);
xnor U32454 (N_32454,N_21757,N_27026);
nor U32455 (N_32455,N_21340,N_27121);
and U32456 (N_32456,N_26190,N_27641);
nor U32457 (N_32457,N_23468,N_25349);
xnor U32458 (N_32458,N_28457,N_22724);
nor U32459 (N_32459,N_23310,N_28914);
xnor U32460 (N_32460,N_28637,N_21652);
nand U32461 (N_32461,N_23578,N_26894);
or U32462 (N_32462,N_28199,N_22621);
xor U32463 (N_32463,N_27360,N_27148);
and U32464 (N_32464,N_24956,N_21153);
and U32465 (N_32465,N_25348,N_29620);
nor U32466 (N_32466,N_21756,N_27869);
and U32467 (N_32467,N_23487,N_29324);
or U32468 (N_32468,N_20791,N_23997);
nand U32469 (N_32469,N_28538,N_27292);
or U32470 (N_32470,N_24733,N_29942);
or U32471 (N_32471,N_27997,N_24169);
nor U32472 (N_32472,N_24341,N_28138);
or U32473 (N_32473,N_29295,N_29394);
nand U32474 (N_32474,N_28146,N_24722);
nand U32475 (N_32475,N_27851,N_29647);
nand U32476 (N_32476,N_28082,N_28036);
and U32477 (N_32477,N_22932,N_26586);
or U32478 (N_32478,N_28450,N_26895);
nand U32479 (N_32479,N_24105,N_20145);
or U32480 (N_32480,N_26788,N_21169);
nor U32481 (N_32481,N_23001,N_22386);
or U32482 (N_32482,N_29282,N_25903);
and U32483 (N_32483,N_25931,N_23453);
nand U32484 (N_32484,N_26381,N_28703);
nor U32485 (N_32485,N_20775,N_22928);
nor U32486 (N_32486,N_29610,N_25626);
nor U32487 (N_32487,N_28335,N_29915);
nor U32488 (N_32488,N_21025,N_29970);
nor U32489 (N_32489,N_22855,N_29580);
or U32490 (N_32490,N_29943,N_21662);
xnor U32491 (N_32491,N_20554,N_21966);
nor U32492 (N_32492,N_20474,N_20509);
nor U32493 (N_32493,N_28103,N_24336);
or U32494 (N_32494,N_24734,N_22299);
and U32495 (N_32495,N_23985,N_23154);
xnor U32496 (N_32496,N_25849,N_28677);
xnor U32497 (N_32497,N_22392,N_28354);
xnor U32498 (N_32498,N_22696,N_22646);
nand U32499 (N_32499,N_28663,N_26227);
nor U32500 (N_32500,N_24637,N_22182);
xor U32501 (N_32501,N_29061,N_25574);
or U32502 (N_32502,N_23507,N_28786);
nand U32503 (N_32503,N_28461,N_24139);
nor U32504 (N_32504,N_27456,N_26868);
nand U32505 (N_32505,N_26900,N_22954);
nor U32506 (N_32506,N_28181,N_29732);
nand U32507 (N_32507,N_21122,N_22656);
nor U32508 (N_32508,N_23473,N_29301);
nand U32509 (N_32509,N_21878,N_29305);
and U32510 (N_32510,N_26645,N_24374);
and U32511 (N_32511,N_25826,N_20692);
nand U32512 (N_32512,N_21139,N_29687);
nand U32513 (N_32513,N_22396,N_22188);
nor U32514 (N_32514,N_26905,N_24717);
nand U32515 (N_32515,N_23118,N_22894);
or U32516 (N_32516,N_27988,N_21697);
nand U32517 (N_32517,N_21703,N_25434);
nand U32518 (N_32518,N_24422,N_26585);
and U32519 (N_32519,N_22415,N_25652);
or U32520 (N_32520,N_22147,N_25038);
and U32521 (N_32521,N_29229,N_29175);
nand U32522 (N_32522,N_24497,N_21918);
xor U32523 (N_32523,N_28683,N_27085);
and U32524 (N_32524,N_28816,N_22943);
nor U32525 (N_32525,N_24344,N_21895);
or U32526 (N_32526,N_25420,N_28147);
nand U32527 (N_32527,N_25389,N_27493);
nand U32528 (N_32528,N_20517,N_25708);
nand U32529 (N_32529,N_26362,N_20206);
and U32530 (N_32530,N_25872,N_24925);
or U32531 (N_32531,N_22934,N_20352);
and U32532 (N_32532,N_27698,N_27838);
and U32533 (N_32533,N_27378,N_27223);
or U32534 (N_32534,N_26242,N_28755);
and U32535 (N_32535,N_25801,N_24324);
or U32536 (N_32536,N_20665,N_28472);
nand U32537 (N_32537,N_23573,N_22585);
nand U32538 (N_32538,N_20635,N_25541);
and U32539 (N_32539,N_24704,N_24439);
nor U32540 (N_32540,N_29787,N_20351);
nor U32541 (N_32541,N_28904,N_27337);
and U32542 (N_32542,N_23238,N_23231);
nand U32543 (N_32543,N_29973,N_26537);
nor U32544 (N_32544,N_24628,N_21722);
and U32545 (N_32545,N_22443,N_24474);
or U32546 (N_32546,N_28611,N_25866);
and U32547 (N_32547,N_27752,N_25557);
and U32548 (N_32548,N_26027,N_29775);
nor U32549 (N_32549,N_20533,N_29826);
xor U32550 (N_32550,N_25352,N_27837);
or U32551 (N_32551,N_27815,N_22688);
nor U32552 (N_32552,N_21963,N_26906);
and U32553 (N_32553,N_28881,N_27187);
xor U32554 (N_32554,N_20898,N_24951);
or U32555 (N_32555,N_28512,N_29462);
nor U32556 (N_32556,N_20764,N_24854);
or U32557 (N_32557,N_23379,N_21194);
nor U32558 (N_32558,N_25580,N_23432);
or U32559 (N_32559,N_28955,N_25329);
or U32560 (N_32560,N_24218,N_22245);
or U32561 (N_32561,N_27793,N_25760);
and U32562 (N_32562,N_24419,N_20157);
or U32563 (N_32563,N_25679,N_27453);
or U32564 (N_32564,N_20439,N_25412);
nand U32565 (N_32565,N_27651,N_21506);
nor U32566 (N_32566,N_21921,N_25117);
and U32567 (N_32567,N_21759,N_21418);
xor U32568 (N_32568,N_23290,N_25914);
nor U32569 (N_32569,N_20261,N_20494);
nand U32570 (N_32570,N_21301,N_28256);
nand U32571 (N_32571,N_27134,N_21256);
and U32572 (N_32572,N_24217,N_27279);
and U32573 (N_32573,N_21943,N_25585);
nor U32574 (N_32574,N_20954,N_21417);
nand U32575 (N_32575,N_26495,N_29397);
nand U32576 (N_32576,N_29430,N_29102);
or U32577 (N_32577,N_21972,N_27697);
and U32578 (N_32578,N_27671,N_29725);
and U32579 (N_32579,N_23099,N_27801);
and U32580 (N_32580,N_24768,N_21726);
or U32581 (N_32581,N_27961,N_21611);
nand U32582 (N_32582,N_25742,N_27577);
nand U32583 (N_32583,N_23059,N_24286);
nand U32584 (N_32584,N_23395,N_20702);
nor U32585 (N_32585,N_22690,N_28817);
nand U32586 (N_32586,N_26706,N_29344);
nand U32587 (N_32587,N_22310,N_20912);
and U32588 (N_32588,N_23022,N_28177);
or U32589 (N_32589,N_22427,N_28967);
nand U32590 (N_32590,N_20632,N_26724);
nand U32591 (N_32591,N_28448,N_21983);
or U32592 (N_32592,N_24775,N_27775);
or U32593 (N_32593,N_27652,N_23606);
or U32594 (N_32594,N_28271,N_27860);
nand U32595 (N_32595,N_22123,N_22284);
or U32596 (N_32596,N_24745,N_20758);
or U32597 (N_32597,N_21985,N_27257);
and U32598 (N_32598,N_28475,N_27510);
or U32599 (N_32599,N_28576,N_26394);
or U32600 (N_32600,N_29626,N_29306);
nand U32601 (N_32601,N_22203,N_24829);
and U32602 (N_32602,N_21178,N_22405);
or U32603 (N_32603,N_27232,N_23009);
nand U32604 (N_32604,N_23103,N_29503);
xor U32605 (N_32605,N_24841,N_26590);
or U32606 (N_32606,N_28285,N_29077);
nor U32607 (N_32607,N_27503,N_24772);
xor U32608 (N_32608,N_29768,N_20915);
and U32609 (N_32609,N_25635,N_24524);
nand U32610 (N_32610,N_27610,N_23614);
and U32611 (N_32611,N_29182,N_23971);
or U32612 (N_32612,N_26740,N_22221);
nand U32613 (N_32613,N_24102,N_29494);
and U32614 (N_32614,N_22849,N_26101);
nand U32615 (N_32615,N_21410,N_24666);
nor U32616 (N_32616,N_20493,N_29525);
nand U32617 (N_32617,N_25967,N_22240);
and U32618 (N_32618,N_26131,N_27020);
or U32619 (N_32619,N_21144,N_29912);
nor U32620 (N_32620,N_21269,N_22620);
nand U32621 (N_32621,N_24062,N_29042);
and U32622 (N_32622,N_21607,N_25963);
xor U32623 (N_32623,N_28211,N_23363);
nand U32624 (N_32624,N_25301,N_24008);
or U32625 (N_32625,N_29457,N_22138);
nor U32626 (N_32626,N_20243,N_24470);
and U32627 (N_32627,N_20598,N_21801);
or U32628 (N_32628,N_21466,N_20176);
nor U32629 (N_32629,N_22640,N_24025);
nand U32630 (N_32630,N_24634,N_27124);
and U32631 (N_32631,N_28913,N_20999);
and U32632 (N_32632,N_27386,N_23097);
nand U32633 (N_32633,N_28937,N_26226);
and U32634 (N_32634,N_25758,N_27316);
nor U32635 (N_32635,N_22958,N_22917);
and U32636 (N_32636,N_24241,N_21545);
nand U32637 (N_32637,N_26222,N_20453);
or U32638 (N_32638,N_25938,N_21730);
xor U32639 (N_32639,N_22081,N_22903);
nand U32640 (N_32640,N_29945,N_28017);
nand U32641 (N_32641,N_28628,N_20942);
nand U32642 (N_32642,N_23277,N_24805);
nor U32643 (N_32643,N_25309,N_27115);
nand U32644 (N_32644,N_28948,N_29636);
or U32645 (N_32645,N_22022,N_29841);
and U32646 (N_32646,N_20203,N_28587);
or U32647 (N_32647,N_28057,N_24591);
or U32648 (N_32648,N_22554,N_23221);
and U32649 (N_32649,N_29651,N_22317);
and U32650 (N_32650,N_25047,N_27979);
nor U32651 (N_32651,N_22847,N_20307);
and U32652 (N_32652,N_27412,N_21769);
xor U32653 (N_32653,N_21081,N_28644);
nand U32654 (N_32654,N_26312,N_26948);
or U32655 (N_32655,N_24049,N_24115);
nor U32656 (N_32656,N_29400,N_24160);
or U32657 (N_32657,N_22278,N_28015);
nor U32658 (N_32658,N_22096,N_22449);
and U32659 (N_32659,N_24042,N_24812);
nor U32660 (N_32660,N_22094,N_27675);
and U32661 (N_32661,N_22211,N_21260);
or U32662 (N_32662,N_26256,N_22161);
nand U32663 (N_32663,N_29445,N_20975);
xnor U32664 (N_32664,N_25281,N_28108);
nor U32665 (N_32665,N_23412,N_26746);
nand U32666 (N_32666,N_22558,N_25200);
nand U32667 (N_32667,N_26890,N_21320);
nand U32668 (N_32668,N_26607,N_22714);
nor U32669 (N_32669,N_23602,N_25647);
nor U32670 (N_32670,N_26361,N_23978);
nor U32671 (N_32671,N_21364,N_20463);
xnor U32672 (N_32672,N_25134,N_21876);
nor U32673 (N_32673,N_23737,N_24386);
nand U32674 (N_32674,N_24176,N_25146);
xnor U32675 (N_32675,N_25705,N_29632);
or U32676 (N_32676,N_24514,N_22782);
and U32677 (N_32677,N_23671,N_27432);
nor U32678 (N_32678,N_21200,N_27189);
or U32679 (N_32679,N_21910,N_26780);
or U32680 (N_32680,N_24622,N_27375);
and U32681 (N_32681,N_25747,N_24048);
or U32682 (N_32682,N_25690,N_25508);
and U32683 (N_32683,N_28279,N_22726);
and U32684 (N_32684,N_23126,N_29763);
nand U32685 (N_32685,N_27391,N_24558);
nand U32686 (N_32686,N_26365,N_25520);
and U32687 (N_32687,N_22864,N_24963);
and U32688 (N_32688,N_26114,N_27982);
nor U32689 (N_32689,N_22997,N_21672);
and U32690 (N_32690,N_29604,N_22692);
and U32691 (N_32691,N_22736,N_29944);
or U32692 (N_32692,N_29325,N_28025);
xor U32693 (N_32693,N_27998,N_27949);
and U32694 (N_32694,N_26813,N_23856);
nand U32695 (N_32695,N_27973,N_21163);
nor U32696 (N_32696,N_22335,N_28566);
or U32697 (N_32697,N_21814,N_27624);
and U32698 (N_32698,N_21180,N_25050);
xor U32699 (N_32699,N_22875,N_28444);
nor U32700 (N_32700,N_23416,N_25180);
nand U32701 (N_32701,N_25984,N_22374);
nor U32702 (N_32702,N_21402,N_24940);
and U32703 (N_32703,N_24573,N_22844);
or U32704 (N_32704,N_23392,N_28113);
and U32705 (N_32705,N_26834,N_22206);
nand U32706 (N_32706,N_20135,N_22205);
or U32707 (N_32707,N_22001,N_24506);
nor U32708 (N_32708,N_28774,N_29146);
nor U32709 (N_32709,N_20807,N_24018);
or U32710 (N_32710,N_27234,N_25440);
xor U32711 (N_32711,N_21882,N_27217);
nor U32712 (N_32712,N_25779,N_23576);
nor U32713 (N_32713,N_29907,N_24383);
and U32714 (N_32714,N_29104,N_26741);
and U32715 (N_32715,N_24153,N_27157);
nand U32716 (N_32716,N_25969,N_23345);
nand U32717 (N_32717,N_27909,N_25408);
nor U32718 (N_32718,N_22148,N_28800);
nand U32719 (N_32719,N_21554,N_29733);
and U32720 (N_32720,N_27919,N_20435);
and U32721 (N_32721,N_27991,N_29004);
nand U32722 (N_32722,N_27405,N_24688);
nor U32723 (N_32723,N_20603,N_20292);
or U32724 (N_32724,N_20772,N_26257);
nor U32725 (N_32725,N_22399,N_22065);
nand U32726 (N_32726,N_29434,N_24779);
or U32727 (N_32727,N_23621,N_21119);
and U32728 (N_32728,N_28029,N_28643);
nor U32729 (N_32729,N_22929,N_22348);
or U32730 (N_32730,N_28402,N_29313);
nor U32731 (N_32731,N_29012,N_23765);
nor U32732 (N_32732,N_22072,N_27127);
nand U32733 (N_32733,N_20277,N_23366);
and U32734 (N_32734,N_28084,N_24016);
and U32735 (N_32735,N_22699,N_21378);
nor U32736 (N_32736,N_25853,N_26481);
nor U32737 (N_32737,N_26416,N_26910);
nor U32738 (N_32738,N_29668,N_28885);
nand U32739 (N_32739,N_27365,N_21247);
and U32740 (N_32740,N_24553,N_29474);
nor U32741 (N_32741,N_28230,N_29352);
nor U32742 (N_32742,N_27670,N_24164);
nor U32743 (N_32743,N_22576,N_24974);
and U32744 (N_32744,N_24649,N_22074);
nor U32745 (N_32745,N_24789,N_25282);
or U32746 (N_32746,N_24305,N_27462);
nor U32747 (N_32747,N_23223,N_29008);
nand U32748 (N_32748,N_23446,N_26476);
nand U32749 (N_32749,N_23480,N_20368);
nor U32750 (N_32750,N_23071,N_24095);
nor U32751 (N_32751,N_28978,N_27883);
or U32752 (N_32752,N_29413,N_27785);
nor U32753 (N_32753,N_27305,N_26565);
nor U32754 (N_32754,N_21917,N_28439);
xnor U32755 (N_32755,N_29683,N_20366);
nand U32756 (N_32756,N_27374,N_22330);
or U32757 (N_32757,N_28186,N_22801);
and U32758 (N_32758,N_23589,N_26726);
nor U32759 (N_32759,N_21745,N_27312);
nand U32760 (N_32760,N_20923,N_20303);
nand U32761 (N_32761,N_22008,N_25731);
and U32762 (N_32762,N_23518,N_26228);
nand U32763 (N_32763,N_28864,N_25908);
nor U32764 (N_32764,N_21903,N_25898);
and U32765 (N_32765,N_29261,N_20419);
nand U32766 (N_32766,N_22263,N_25331);
nor U32767 (N_32767,N_21351,N_29593);
and U32768 (N_32768,N_29716,N_24603);
and U32769 (N_32769,N_22700,N_25798);
or U32770 (N_32770,N_23519,N_27092);
or U32771 (N_32771,N_26535,N_26471);
nand U32772 (N_32772,N_22355,N_26757);
nor U32773 (N_32773,N_24211,N_27504);
nand U32774 (N_32774,N_28848,N_25068);
xor U32775 (N_32775,N_24549,N_22170);
nand U32776 (N_32776,N_25670,N_27297);
xor U32777 (N_32777,N_29385,N_24377);
nor U32778 (N_32778,N_23500,N_21058);
and U32779 (N_32779,N_27894,N_20645);
nor U32780 (N_32780,N_27009,N_27425);
or U32781 (N_32781,N_28117,N_24372);
and U32782 (N_32782,N_21973,N_27616);
nor U32783 (N_32783,N_22753,N_20046);
or U32784 (N_32784,N_25817,N_28079);
nor U32785 (N_32785,N_25082,N_25277);
and U32786 (N_32786,N_21616,N_23283);
and U32787 (N_32787,N_24835,N_24961);
nand U32788 (N_32788,N_22454,N_20949);
and U32789 (N_32789,N_23475,N_29159);
or U32790 (N_32790,N_26493,N_25167);
or U32791 (N_32791,N_28407,N_23600);
or U32792 (N_32792,N_20178,N_26888);
nor U32793 (N_32793,N_26750,N_26871);
or U32794 (N_32794,N_24810,N_25960);
nand U32795 (N_32795,N_27802,N_29780);
and U32796 (N_32796,N_20604,N_24050);
nor U32797 (N_32797,N_24485,N_25566);
nor U32798 (N_32798,N_27249,N_21564);
or U32799 (N_32799,N_27119,N_25722);
nand U32800 (N_32800,N_29409,N_20568);
and U32801 (N_32801,N_20587,N_27373);
or U32802 (N_32802,N_22575,N_29139);
xor U32803 (N_32803,N_21595,N_29258);
nand U32804 (N_32804,N_21325,N_22064);
xor U32805 (N_32805,N_20438,N_22104);
xor U32806 (N_32806,N_26480,N_21686);
nor U32807 (N_32807,N_23413,N_28756);
nand U32808 (N_32808,N_29628,N_29402);
and U32809 (N_32809,N_20761,N_27975);
and U32810 (N_32810,N_25450,N_21680);
and U32811 (N_32811,N_24885,N_22408);
nand U32812 (N_32812,N_26624,N_21113);
or U32813 (N_32813,N_20072,N_24846);
nor U32814 (N_32814,N_27296,N_23094);
nor U32815 (N_32815,N_26685,N_24380);
nor U32816 (N_32816,N_27182,N_22745);
or U32817 (N_32817,N_23254,N_23060);
or U32818 (N_32818,N_29129,N_20231);
or U32819 (N_32819,N_20371,N_27463);
nand U32820 (N_32820,N_28058,N_21546);
nand U32821 (N_32821,N_24975,N_29761);
nor U32822 (N_32822,N_26036,N_22948);
nor U32823 (N_32823,N_29976,N_24401);
nand U32824 (N_32824,N_25118,N_23253);
and U32825 (N_32825,N_21557,N_28462);
and U32826 (N_32826,N_29930,N_23872);
or U32827 (N_32827,N_23690,N_23648);
or U32828 (N_32828,N_29545,N_26082);
and U32829 (N_32829,N_29662,N_25222);
and U32830 (N_32830,N_26509,N_22848);
nand U32831 (N_32831,N_24675,N_26368);
xor U32832 (N_32832,N_21284,N_24438);
or U32833 (N_32833,N_22295,N_26032);
xnor U32834 (N_32834,N_20709,N_22835);
and U32835 (N_32835,N_21679,N_20828);
and U32836 (N_32836,N_29478,N_21797);
or U32837 (N_32837,N_21916,N_29073);
and U32838 (N_32838,N_27717,N_22143);
and U32839 (N_32839,N_29946,N_28151);
nand U32840 (N_32840,N_26798,N_22200);
and U32841 (N_32841,N_29072,N_24471);
xnor U32842 (N_32842,N_22953,N_21486);
or U32843 (N_32843,N_28040,N_24790);
or U32844 (N_32844,N_21457,N_28647);
xor U32845 (N_32845,N_29110,N_29608);
or U32846 (N_32846,N_26155,N_29921);
and U32847 (N_32847,N_26968,N_24777);
or U32848 (N_32848,N_23516,N_28876);
nor U32849 (N_32849,N_23819,N_26042);
and U32850 (N_32850,N_21868,N_21405);
or U32851 (N_32851,N_24037,N_20706);
xor U32852 (N_32852,N_22716,N_20750);
or U32853 (N_32853,N_26814,N_23301);
xor U32854 (N_32854,N_20856,N_23484);
nor U32855 (N_32855,N_20403,N_25174);
nand U32856 (N_32856,N_27408,N_26858);
nand U32857 (N_32857,N_25350,N_29688);
or U32858 (N_32858,N_27414,N_27917);
or U32859 (N_32859,N_20611,N_21835);
or U32860 (N_32860,N_25743,N_25659);
nand U32861 (N_32861,N_22911,N_29599);
or U32862 (N_32862,N_20312,N_26572);
or U32863 (N_32863,N_28639,N_21707);
xor U32864 (N_32864,N_20088,N_24515);
or U32865 (N_32865,N_22768,N_20391);
or U32866 (N_32866,N_26092,N_23525);
and U32867 (N_32867,N_27915,N_25156);
or U32868 (N_32868,N_25067,N_21729);
or U32869 (N_32869,N_21219,N_25886);
or U32870 (N_32870,N_21437,N_22337);
and U32871 (N_32871,N_26293,N_23895);
nand U32872 (N_32872,N_22618,N_28712);
or U32873 (N_32873,N_24513,N_29922);
and U32874 (N_32874,N_26954,N_28889);
and U32875 (N_32875,N_23332,N_26690);
nor U32876 (N_32876,N_22343,N_21958);
nor U32877 (N_32877,N_26369,N_27945);
nor U32878 (N_32878,N_28205,N_23042);
xor U32879 (N_32879,N_22935,N_24566);
nand U32880 (N_32880,N_29119,N_21306);
or U32881 (N_32881,N_24138,N_21997);
nand U32882 (N_32882,N_25241,N_29774);
and U32883 (N_32883,N_26161,N_22441);
and U32884 (N_32884,N_21661,N_21923);
nand U32885 (N_32885,N_20489,N_22909);
nand U32886 (N_32886,N_22232,N_21641);
nand U32887 (N_32887,N_21311,N_28048);
nor U32888 (N_32888,N_26207,N_29695);
nand U32889 (N_32889,N_25932,N_25845);
or U32890 (N_32890,N_26465,N_21618);
nand U32891 (N_32891,N_21118,N_20601);
and U32892 (N_32892,N_28382,N_26153);
nor U32893 (N_32893,N_24157,N_25664);
nand U32894 (N_32894,N_23047,N_25030);
and U32895 (N_32895,N_27265,N_22732);
nor U32896 (N_32896,N_25108,N_22047);
xnor U32897 (N_32897,N_28075,N_28416);
nand U32898 (N_32898,N_27582,N_22508);
or U32899 (N_32899,N_23078,N_23218);
nor U32900 (N_32900,N_21920,N_29591);
nor U32901 (N_32901,N_24314,N_23028);
and U32902 (N_32902,N_20858,N_22513);
and U32903 (N_32903,N_28713,N_23211);
nand U32904 (N_32904,N_24258,N_28302);
and U32905 (N_32905,N_26059,N_28001);
xnor U32906 (N_32906,N_29702,N_29609);
nor U32907 (N_32907,N_27803,N_24185);
nand U32908 (N_32908,N_27321,N_21924);
and U32909 (N_32909,N_25896,N_29416);
xnor U32910 (N_32910,N_21165,N_27533);
and U32911 (N_32911,N_23610,N_20974);
or U32912 (N_32912,N_21603,N_29844);
or U32913 (N_32913,N_26525,N_27195);
xnor U32914 (N_32914,N_28673,N_26046);
or U32915 (N_32915,N_26797,N_29854);
and U32916 (N_32916,N_20323,N_20008);
or U32917 (N_32917,N_27406,N_24295);
or U32918 (N_32918,N_27095,N_26595);
nand U32919 (N_32919,N_25572,N_22350);
nand U32920 (N_32920,N_27579,N_24898);
and U32921 (N_32921,N_28241,N_24697);
nand U32922 (N_32922,N_23762,N_25997);
or U32923 (N_32923,N_29650,N_28276);
or U32924 (N_32924,N_23664,N_22353);
nand U32925 (N_32925,N_28894,N_24202);
nand U32926 (N_32926,N_26111,N_28862);
and U32927 (N_32927,N_20579,N_25394);
nand U32928 (N_32928,N_21211,N_24532);
nor U32929 (N_32929,N_26331,N_22090);
nor U32930 (N_32930,N_20686,N_25314);
or U32931 (N_32931,N_22682,N_29781);
or U32932 (N_32932,N_20047,N_29834);
nand U32933 (N_32933,N_27288,N_23076);
and U32934 (N_32934,N_27275,N_27452);
or U32935 (N_32935,N_27858,N_24935);
or U32936 (N_32936,N_25308,N_20963);
nor U32937 (N_32937,N_26739,N_22927);
and U32938 (N_32938,N_26223,N_25823);
nor U32939 (N_32939,N_25529,N_20501);
or U32940 (N_32940,N_24540,N_25345);
nand U32941 (N_32941,N_27680,N_21836);
xor U32942 (N_32942,N_25902,N_28707);
nor U32943 (N_32943,N_22552,N_29539);
nand U32944 (N_32944,N_25431,N_26377);
or U32945 (N_32945,N_21936,N_21739);
or U32946 (N_32946,N_27401,N_22267);
or U32947 (N_32947,N_23178,N_20582);
and U32948 (N_32948,N_27433,N_26704);
or U32949 (N_32949,N_24607,N_20789);
or U32950 (N_32950,N_26095,N_29825);
nand U32951 (N_32951,N_22304,N_22580);
and U32952 (N_32952,N_24012,N_25676);
and U32953 (N_32953,N_23714,N_24601);
nor U32954 (N_32954,N_29994,N_28392);
nand U32955 (N_32955,N_25142,N_28715);
nor U32956 (N_32956,N_25000,N_23566);
nor U32957 (N_32957,N_25699,N_27687);
and U32958 (N_32958,N_21383,N_26828);
and U32959 (N_32959,N_24765,N_25110);
nand U32960 (N_32960,N_27507,N_23343);
or U32961 (N_32961,N_25491,N_28627);
nand U32962 (N_32962,N_23582,N_27506);
nor U32963 (N_32963,N_26398,N_27243);
and U32964 (N_32964,N_21018,N_21114);
and U32965 (N_32965,N_21190,N_22609);
or U32966 (N_32966,N_22479,N_26123);
and U32967 (N_32967,N_20156,N_29843);
or U32968 (N_32968,N_20528,N_28993);
nand U32969 (N_32969,N_21590,N_20808);
nand U32970 (N_32970,N_29170,N_22972);
nand U32971 (N_32971,N_26668,N_29713);
or U32972 (N_32972,N_20234,N_25093);
nand U32973 (N_32973,N_24245,N_26243);
nand U32974 (N_32974,N_28648,N_28811);
nand U32975 (N_32975,N_28807,N_29718);
or U32976 (N_32976,N_22160,N_20605);
or U32977 (N_32977,N_24027,N_20969);
and U32978 (N_32978,N_29405,N_21034);
and U32979 (N_32979,N_26567,N_20968);
nor U32980 (N_32980,N_23842,N_27576);
or U32981 (N_32981,N_29891,N_22758);
nor U32982 (N_32982,N_29243,N_28842);
nand U32983 (N_32983,N_27744,N_26297);
nor U32984 (N_32984,N_20644,N_29961);
xor U32985 (N_32985,N_20431,N_25484);
nand U32986 (N_32986,N_27678,N_21300);
xor U32987 (N_32987,N_23331,N_24850);
or U32988 (N_32988,N_25629,N_21558);
and U32989 (N_32989,N_25229,N_22770);
xnor U32990 (N_32990,N_27074,N_27901);
nor U32991 (N_32991,N_29027,N_23729);
nor U32992 (N_32992,N_27014,N_25691);
nor U32993 (N_32993,N_22165,N_28336);
and U32994 (N_32994,N_22403,N_27368);
and U32995 (N_32995,N_25123,N_22528);
or U32996 (N_32996,N_22680,N_20237);
nand U32997 (N_32997,N_23396,N_28499);
or U32998 (N_32998,N_20416,N_22136);
nand U32999 (N_32999,N_25930,N_25773);
nand U33000 (N_33000,N_24766,N_28131);
and U33001 (N_33001,N_27255,N_29876);
or U33002 (N_33002,N_22595,N_26234);
xnor U33003 (N_33003,N_21087,N_24569);
or U33004 (N_33004,N_21188,N_28893);
xor U33005 (N_33005,N_21585,N_22452);
and U33006 (N_33006,N_24988,N_21764);
nor U33007 (N_33007,N_23622,N_24614);
nor U33008 (N_33008,N_22253,N_21291);
and U33009 (N_33009,N_21660,N_21795);
and U33010 (N_33010,N_20770,N_23715);
and U33011 (N_33011,N_24625,N_22086);
and U33012 (N_33012,N_28200,N_24924);
nand U33013 (N_33013,N_21537,N_27757);
and U33014 (N_33014,N_26501,N_21396);
or U33015 (N_33015,N_25453,N_27726);
nand U33016 (N_33016,N_23744,N_20169);
or U33017 (N_33017,N_27153,N_24830);
nand U33018 (N_33018,N_25663,N_20982);
or U33019 (N_33019,N_27103,N_29279);
nand U33020 (N_33020,N_27539,N_28583);
and U33021 (N_33021,N_26284,N_24128);
or U33022 (N_33022,N_22720,N_28303);
and U33023 (N_33023,N_26429,N_25643);
and U33024 (N_33024,N_23522,N_24484);
nor U33025 (N_33025,N_23818,N_24231);
nand U33026 (N_33026,N_24443,N_29099);
nand U33027 (N_33027,N_20884,N_22626);
and U33028 (N_33028,N_20257,N_22458);
or U33029 (N_33029,N_20765,N_21717);
xor U33030 (N_33030,N_29502,N_25034);
and U33031 (N_33031,N_25012,N_21101);
nor U33032 (N_33032,N_27857,N_24982);
xnor U33033 (N_33033,N_27059,N_29723);
nor U33034 (N_33034,N_20486,N_22461);
or U33035 (N_33035,N_29962,N_22026);
nand U33036 (N_33036,N_27721,N_25214);
nand U33037 (N_33037,N_20022,N_25618);
and U33038 (N_33038,N_28396,N_29343);
nand U33039 (N_33039,N_28615,N_27968);
xnor U33040 (N_33040,N_26846,N_29997);
nor U33041 (N_33041,N_29936,N_27060);
xnor U33042 (N_33042,N_28505,N_20842);
nand U33043 (N_33043,N_22416,N_28572);
nor U33044 (N_33044,N_26540,N_21359);
nand U33045 (N_33045,N_22986,N_23887);
nor U33046 (N_33046,N_29463,N_24038);
nor U33047 (N_33047,N_29685,N_20623);
or U33048 (N_33048,N_21140,N_23513);
and U33049 (N_33049,N_21494,N_24550);
and U33050 (N_33050,N_25475,N_27702);
nor U33051 (N_33051,N_25387,N_29656);
nand U33052 (N_33052,N_28897,N_22862);
nand U33053 (N_33053,N_26804,N_22938);
nor U33054 (N_33054,N_22358,N_24654);
or U33055 (N_33055,N_27280,N_22602);
or U33056 (N_33056,N_23935,N_23085);
xnor U33057 (N_33057,N_26519,N_20846);
or U33058 (N_33058,N_20314,N_28614);
nor U33059 (N_33059,N_22889,N_22522);
and U33060 (N_33060,N_24584,N_22256);
and U33061 (N_33061,N_20844,N_24057);
nand U33062 (N_33062,N_20103,N_27880);
nand U33063 (N_33063,N_22336,N_23143);
or U33064 (N_33064,N_28105,N_20170);
nor U33065 (N_33065,N_26879,N_20662);
nor U33066 (N_33066,N_28984,N_28653);
and U33067 (N_33067,N_20926,N_26716);
xnor U33068 (N_33068,N_27125,N_23409);
or U33069 (N_33069,N_22673,N_29167);
or U33070 (N_33070,N_29488,N_21696);
or U33071 (N_33071,N_27032,N_28139);
nor U33072 (N_33072,N_26166,N_25386);
xnor U33073 (N_33073,N_23400,N_27661);
or U33074 (N_33074,N_29190,N_21581);
and U33075 (N_33075,N_26020,N_27605);
and U33076 (N_33076,N_27956,N_27878);
and U33077 (N_33077,N_25192,N_27725);
or U33078 (N_33078,N_24999,N_23410);
nor U33079 (N_33079,N_28282,N_25890);
or U33080 (N_33080,N_28041,N_26708);
nor U33081 (N_33081,N_29625,N_26468);
nor U33082 (N_33082,N_26836,N_28903);
or U33083 (N_33083,N_28351,N_27943);
nor U33084 (N_33084,N_25017,N_26010);
and U33085 (N_33085,N_21310,N_28020);
nand U33086 (N_33086,N_29956,N_27848);
or U33087 (N_33087,N_24872,N_26175);
xnor U33088 (N_33088,N_20479,N_23232);
nand U33089 (N_33089,N_21125,N_25889);
or U33090 (N_33090,N_27129,N_28226);
or U33091 (N_33091,N_20621,N_23449);
and U33092 (N_33092,N_23640,N_21432);
nand U33093 (N_33093,N_20504,N_28486);
and U33094 (N_33094,N_28091,N_28563);
and U33095 (N_33095,N_27372,N_23206);
and U33096 (N_33096,N_24751,N_24609);
and U33097 (N_33097,N_24382,N_21057);
and U33098 (N_33098,N_24310,N_22549);
or U33099 (N_33099,N_27260,N_20831);
and U33100 (N_33100,N_29335,N_24816);
nand U33101 (N_33101,N_29362,N_22756);
and U33102 (N_33102,N_29978,N_27194);
nand U33103 (N_33103,N_22854,N_24655);
nand U33104 (N_33104,N_20566,N_20684);
nor U33105 (N_33105,N_28035,N_24857);
nor U33106 (N_33106,N_28784,N_24249);
xnor U33107 (N_33107,N_25195,N_29663);
nor U33108 (N_33108,N_23669,N_25634);
or U33109 (N_33109,N_26300,N_23036);
nand U33110 (N_33110,N_21877,N_22417);
and U33111 (N_33111,N_24273,N_20726);
or U33112 (N_33112,N_23954,N_27080);
and U33113 (N_33113,N_22106,N_22228);
nor U33114 (N_33114,N_28939,N_20757);
xor U33115 (N_33115,N_20405,N_22778);
and U33116 (N_33116,N_26141,N_25063);
nor U33117 (N_33117,N_26958,N_26584);
and U33118 (N_33118,N_27864,N_26060);
nor U33119 (N_33119,N_28172,N_20922);
or U33120 (N_33120,N_21925,N_25739);
xnor U33121 (N_33121,N_28213,N_25928);
or U33122 (N_33122,N_20527,N_21104);
and U33123 (N_33123,N_21471,N_27399);
xnor U33124 (N_33124,N_24592,N_22489);
nor U33125 (N_33125,N_25702,N_28277);
and U33126 (N_33126,N_25527,N_28579);
nand U33127 (N_33127,N_24320,N_20682);
and U33128 (N_33128,N_20959,N_24761);
or U33129 (N_33129,N_23451,N_25594);
and U33130 (N_33130,N_26452,N_26876);
or U33131 (N_33131,N_22192,N_27673);
nand U33132 (N_33132,N_26849,N_25373);
and U33133 (N_33133,N_25766,N_21578);
nand U33134 (N_33134,N_21938,N_24610);
and U33135 (N_33135,N_25196,N_27174);
nor U33136 (N_33136,N_20559,N_24356);
nand U33137 (N_33137,N_21259,N_29813);
or U33138 (N_33138,N_25423,N_24472);
and U33139 (N_33139,N_20546,N_25741);
or U33140 (N_33140,N_27918,N_26678);
nand U33141 (N_33141,N_22246,N_22612);
nor U33142 (N_33142,N_24943,N_21600);
or U33143 (N_33143,N_26702,N_24190);
nor U33144 (N_33144,N_27403,N_29712);
and U33145 (N_33145,N_23204,N_23172);
and U33146 (N_33146,N_20627,N_26887);
and U33147 (N_33147,N_26990,N_21880);
or U33148 (N_33148,N_21699,N_24778);
nand U33149 (N_33149,N_27989,N_29479);
or U33150 (N_33150,N_29516,N_21389);
and U33151 (N_33151,N_27602,N_21534);
nand U33152 (N_33152,N_28758,N_26869);
nand U33153 (N_33153,N_22830,N_25821);
or U33154 (N_33154,N_22774,N_24229);
nor U33155 (N_33155,N_23964,N_21803);
or U33156 (N_33156,N_29561,N_21357);
nand U33157 (N_33157,N_28339,N_29816);
nor U33158 (N_33158,N_27349,N_25049);
nor U33159 (N_33159,N_26403,N_23051);
nand U33160 (N_33160,N_27617,N_28531);
nor U33161 (N_33161,N_29407,N_24406);
nand U33162 (N_33162,N_22504,N_28044);
and U33163 (N_33163,N_25658,N_26409);
or U33164 (N_33164,N_20354,N_20541);
and U33165 (N_33165,N_24206,N_25152);
nand U33166 (N_33166,N_26817,N_26199);
nor U33167 (N_33167,N_24096,N_23937);
nand U33168 (N_33168,N_25100,N_25311);
nand U33169 (N_33169,N_22919,N_20946);
or U33170 (N_33170,N_23015,N_23493);
or U33171 (N_33171,N_21994,N_25325);
nand U33172 (N_33172,N_28690,N_27198);
nand U33173 (N_33173,N_29860,N_27907);
xor U33174 (N_33174,N_25455,N_24331);
and U33175 (N_33175,N_25339,N_21129);
nand U33176 (N_33176,N_29187,N_25874);
xnor U33177 (N_33177,N_22823,N_20967);
nand U33178 (N_33178,N_20182,N_22744);
and U33179 (N_33179,N_25413,N_23425);
xnor U33180 (N_33180,N_21783,N_23437);
and U33181 (N_33181,N_24288,N_28731);
nand U33182 (N_33182,N_21596,N_29117);
nand U33183 (N_33183,N_20855,N_26182);
or U33184 (N_33184,N_20992,N_20316);
and U33185 (N_33185,N_23533,N_25785);
nand U33186 (N_33186,N_29741,N_24763);
and U33187 (N_33187,N_24100,N_28272);
nor U33188 (N_33188,N_26744,N_27591);
xnor U33189 (N_33189,N_29225,N_24757);
nand U33190 (N_33190,N_22146,N_21665);
or U33191 (N_33191,N_23488,N_27923);
and U33192 (N_33192,N_20512,N_25550);
and U33193 (N_33193,N_26338,N_26870);
nor U33194 (N_33194,N_23107,N_26467);
nand U33195 (N_33195,N_28943,N_21475);
nor U33196 (N_33196,N_20219,N_29299);
or U33197 (N_33197,N_29446,N_23018);
and U33198 (N_33198,N_27005,N_20481);
or U33199 (N_33199,N_23746,N_28410);
or U33200 (N_33200,N_24623,N_29141);
or U33201 (N_33201,N_29477,N_29209);
or U33202 (N_33202,N_28324,N_22816);
xnor U33203 (N_33203,N_20332,N_21967);
nand U33204 (N_33204,N_28926,N_21491);
xnor U33205 (N_33205,N_23570,N_23414);
or U33206 (N_33206,N_23727,N_20729);
nor U33207 (N_33207,N_23087,N_26665);
or U33208 (N_33208,N_28503,N_22988);
nand U33209 (N_33209,N_22073,N_21718);
or U33210 (N_33210,N_21839,N_23995);
nand U33211 (N_33211,N_26187,N_22713);
or U33212 (N_33212,N_27333,N_22826);
and U33213 (N_33213,N_26071,N_28011);
nand U33214 (N_33214,N_24920,N_29088);
nand U33215 (N_33215,N_29382,N_24993);
or U33216 (N_33216,N_23772,N_27699);
and U33217 (N_33217,N_26823,N_21016);
or U33218 (N_33218,N_23140,N_28981);
or U33219 (N_33219,N_20212,N_20200);
and U33220 (N_33220,N_29133,N_25211);
xnor U33221 (N_33221,N_26065,N_25959);
or U33222 (N_33222,N_25483,N_28923);
nor U33223 (N_33223,N_29786,N_22109);
or U33224 (N_33224,N_27210,N_23055);
or U33225 (N_33225,N_27599,N_27126);
nand U33226 (N_33226,N_20572,N_24864);
nor U33227 (N_33227,N_21841,N_29757);
and U33228 (N_33228,N_29792,N_25488);
or U33229 (N_33229,N_24414,N_26316);
or U33230 (N_33230,N_26878,N_21390);
nand U33231 (N_33231,N_27206,N_23754);
and U33232 (N_33232,N_25525,N_23180);
or U33233 (N_33233,N_25303,N_27529);
or U33234 (N_33234,N_27081,N_20226);
or U33235 (N_33235,N_20500,N_23049);
xor U33236 (N_33236,N_20147,N_24583);
and U33237 (N_33237,N_25171,N_20608);
or U33238 (N_33238,N_24709,N_27133);
xnor U33239 (N_33239,N_29158,N_29851);
xnor U33240 (N_33240,N_27413,N_20526);
and U33241 (N_33241,N_26782,N_22014);
nand U33242 (N_33242,N_28957,N_29234);
xor U33243 (N_33243,N_23199,N_29755);
or U33244 (N_33244,N_23219,N_23237);
nor U33245 (N_33245,N_27644,N_22153);
nand U33246 (N_33246,N_27640,N_20137);
and U33247 (N_33247,N_25901,N_21762);
nand U33248 (N_33248,N_28364,N_27779);
nor U33249 (N_33249,N_26184,N_20680);
nand U33250 (N_33250,N_28578,N_23822);
or U33251 (N_33251,N_20039,N_29672);
xor U33252 (N_33252,N_22092,N_29869);
nor U33253 (N_33253,N_26485,N_27821);
nand U33254 (N_33254,N_28638,N_25341);
or U33255 (N_33255,N_25290,N_22603);
nor U33256 (N_33256,N_22942,N_23271);
nor U33257 (N_33257,N_26105,N_24678);
nand U33258 (N_33258,N_26442,N_28400);
nand U33259 (N_33259,N_26694,N_24562);
nor U33260 (N_33260,N_20195,N_28650);
nand U33261 (N_33261,N_20320,N_22695);
xnor U33262 (N_33262,N_28999,N_29481);
xor U33263 (N_33263,N_20802,N_20689);
and U33264 (N_33264,N_26109,N_29862);
nor U33265 (N_33265,N_20346,N_25377);
nand U33266 (N_33266,N_20877,N_29569);
nand U33267 (N_33267,N_20326,N_20081);
nor U33268 (N_33268,N_25396,N_22395);
and U33269 (N_33269,N_23528,N_29801);
xnor U33270 (N_33270,N_24605,N_21107);
and U33271 (N_33271,N_29138,N_21503);
nand U33272 (N_33272,N_29107,N_27897);
nand U33273 (N_33273,N_27528,N_23315);
or U33274 (N_33274,N_20648,N_21708);
and U33275 (N_33275,N_26563,N_24996);
or U33276 (N_33276,N_26862,N_27175);
nand U33277 (N_33277,N_29802,N_26422);
and U33278 (N_33278,N_23791,N_21202);
nand U33279 (N_33279,N_23474,N_20324);
nand U33280 (N_33280,N_20001,N_21480);
or U33281 (N_33281,N_29128,N_24400);
nand U33282 (N_33282,N_27666,N_21328);
and U33283 (N_33283,N_23144,N_21780);
or U33284 (N_33284,N_20919,N_23751);
nor U33285 (N_33285,N_20150,N_27612);
or U33286 (N_33286,N_20184,N_21216);
xor U33287 (N_33287,N_26041,N_24913);
nand U33288 (N_33288,N_24270,N_25472);
nor U33289 (N_33289,N_21571,N_24774);
and U33290 (N_33290,N_21716,N_22485);
and U33291 (N_33291,N_20896,N_26949);
nor U33292 (N_33292,N_24983,N_22193);
or U33293 (N_33293,N_27235,N_23039);
or U33294 (N_33294,N_29837,N_24794);
nand U33295 (N_33295,N_24373,N_26216);
nor U33296 (N_33296,N_27166,N_21843);
nand U33297 (N_33297,N_23987,N_29709);
nand U33298 (N_33298,N_29366,N_24579);
or U33299 (N_33299,N_25166,N_29868);
xor U33300 (N_33300,N_27331,N_21191);
and U33301 (N_33301,N_29596,N_27114);
nand U33302 (N_33302,N_29874,N_23362);
and U33303 (N_33303,N_20607,N_26466);
or U33304 (N_33304,N_21253,N_24851);
and U33305 (N_33305,N_20885,N_27267);
and U33306 (N_33306,N_23531,N_20388);
or U33307 (N_33307,N_21905,N_26473);
nor U33308 (N_33308,N_22303,N_20829);
nand U33309 (N_33309,N_23324,N_20816);
xnor U33310 (N_33310,N_21392,N_28646);
nand U33311 (N_33311,N_28544,N_20274);
or U33312 (N_33312,N_26626,N_24276);
nor U33313 (N_33313,N_25624,N_23913);
and U33314 (N_33314,N_26149,N_23124);
and U33315 (N_33315,N_27426,N_23289);
nand U33316 (N_33316,N_21682,N_22291);
nor U33317 (N_33317,N_21233,N_22725);
xnor U33318 (N_33318,N_20876,N_27657);
nand U33319 (N_33319,N_28054,N_20790);
or U33320 (N_33320,N_25802,N_25649);
nor U33321 (N_33321,N_27040,N_20796);
nand U33322 (N_33322,N_25477,N_22991);
xor U33323 (N_33323,N_27314,N_22608);
nor U33324 (N_33324,N_26591,N_28554);
or U33325 (N_33325,N_25294,N_27613);
and U33326 (N_33326,N_20077,N_28702);
or U33327 (N_33327,N_26172,N_22431);
nor U33328 (N_33328,N_28622,N_23766);
xnor U33329 (N_33329,N_22542,N_25018);
or U33330 (N_33330,N_22331,N_24786);
or U33331 (N_33331,N_21239,N_25915);
or U33332 (N_33332,N_29594,N_21321);
nor U33333 (N_33333,N_20124,N_27145);
and U33334 (N_33334,N_29522,N_26662);
xor U33335 (N_33335,N_29322,N_27718);
or U33336 (N_33336,N_26180,N_23466);
or U33337 (N_33337,N_23007,N_22989);
or U33338 (N_33338,N_29541,N_24853);
nor U33339 (N_33339,N_21299,N_22913);
xor U33340 (N_33340,N_28182,N_27992);
nor U33341 (N_33341,N_23169,N_28130);
nand U33342 (N_33342,N_26852,N_21203);
nor U33343 (N_33343,N_29847,N_22099);
nand U33344 (N_33344,N_21523,N_27866);
and U33345 (N_33345,N_24977,N_22434);
xnor U33346 (N_33346,N_28723,N_26385);
or U33347 (N_33347,N_20964,N_29458);
nor U33348 (N_33348,N_27315,N_21258);
xor U33349 (N_33349,N_25076,N_24871);
and U33350 (N_33350,N_24063,N_29657);
or U33351 (N_33351,N_29103,N_26777);
or U33352 (N_33352,N_22524,N_26399);
and U33353 (N_33353,N_20505,N_26996);
or U33354 (N_33354,N_27625,N_23643);
nand U33355 (N_33355,N_29263,N_21316);
and U33356 (N_33356,N_29491,N_26215);
or U33357 (N_33357,N_21327,N_22715);
nand U33358 (N_33358,N_20609,N_29300);
nand U33359 (N_33359,N_22377,N_20792);
nand U33360 (N_33360,N_26553,N_28021);
and U33361 (N_33361,N_27575,N_23440);
nor U33362 (N_33362,N_21468,N_24460);
nor U33363 (N_33363,N_26604,N_28710);
xnor U33364 (N_33364,N_27618,N_22176);
xnor U33365 (N_33365,N_25495,N_20023);
nand U33366 (N_33366,N_23319,N_21214);
and U33367 (N_33367,N_29543,N_25223);
xor U33368 (N_33368,N_20741,N_25980);
or U33369 (N_33369,N_24428,N_26047);
nor U33370 (N_33370,N_29080,N_27098);
or U33371 (N_33371,N_28252,N_24548);
nor U33372 (N_33372,N_29076,N_23686);
or U33373 (N_33373,N_26430,N_23808);
nand U33374 (N_33374,N_20487,N_28812);
nand U33375 (N_33375,N_21869,N_20260);
xnor U33376 (N_33376,N_21886,N_25297);
nand U33377 (N_33377,N_25485,N_28129);
nor U33378 (N_33378,N_27100,N_26169);
nor U33379 (N_33379,N_28312,N_27208);
nor U33380 (N_33380,N_20185,N_21469);
nand U33381 (N_33381,N_26632,N_21631);
xor U33382 (N_33382,N_29010,N_21352);
nand U33383 (N_33383,N_23108,N_25043);
or U33384 (N_33384,N_29779,N_25894);
and U33385 (N_33385,N_23943,N_26271);
or U33386 (N_33386,N_29174,N_20892);
xnor U33387 (N_33387,N_24865,N_23203);
nand U33388 (N_33388,N_26023,N_28847);
or U33389 (N_33389,N_25792,N_22644);
nand U33390 (N_33390,N_27690,N_22430);
nor U33391 (N_33391,N_22931,N_21822);
or U33392 (N_33392,N_26686,N_20953);
nor U33393 (N_33393,N_22158,N_22829);
nor U33394 (N_33394,N_29560,N_22398);
nand U33395 (N_33395,N_27043,N_24161);
xor U33396 (N_33396,N_27355,N_29272);
and U33397 (N_33397,N_20353,N_22000);
or U33398 (N_33398,N_27330,N_20699);
nor U33399 (N_33399,N_24749,N_20550);
xor U33400 (N_33400,N_29795,N_28485);
and U33401 (N_33401,N_28281,N_22832);
and U33402 (N_33402,N_28965,N_28996);
nor U33403 (N_33403,N_20242,N_20569);
nor U33404 (N_33404,N_20673,N_26730);
nor U33405 (N_33405,N_28149,N_23799);
xnor U33406 (N_33406,N_24641,N_26450);
or U33407 (N_33407,N_23627,N_21100);
and U33408 (N_33408,N_27574,N_20719);
and U33409 (N_33409,N_20369,N_23860);
nor U33410 (N_33410,N_28494,N_20496);
and U33411 (N_33411,N_26458,N_28513);
nand U33412 (N_33412,N_22297,N_21865);
nand U33413 (N_33413,N_23012,N_27511);
or U33414 (N_33414,N_25039,N_20747);
nor U33415 (N_33415,N_22610,N_25870);
nand U33416 (N_33416,N_20834,N_29100);
nor U33417 (N_33417,N_23561,N_28453);
nor U33418 (N_33418,N_20313,N_21031);
nand U33419 (N_33419,N_21800,N_21720);
and U33420 (N_33420,N_22021,N_25571);
nand U33421 (N_33421,N_20869,N_23917);
nand U33422 (N_33422,N_22447,N_27137);
nand U33423 (N_33423,N_28166,N_20641);
nor U33424 (N_33424,N_28616,N_22747);
and U33425 (N_33425,N_21086,N_21904);
and U33426 (N_33426,N_28390,N_29472);
nand U33427 (N_33427,N_25257,N_21281);
xnor U33428 (N_33428,N_27526,N_28446);
nand U33429 (N_33429,N_24187,N_26472);
nor U33430 (N_33430,N_28195,N_25338);
nand U33431 (N_33431,N_21519,N_21885);
and U33432 (N_33432,N_21365,N_25273);
and U33433 (N_33433,N_25771,N_23485);
or U33434 (N_33434,N_20732,N_23775);
nor U33435 (N_33435,N_29114,N_23155);
and U33436 (N_33436,N_28490,N_20085);
nand U33437 (N_33437,N_21573,N_28688);
nand U33438 (N_33438,N_25287,N_22968);
or U33439 (N_33439,N_21160,N_28087);
nand U33440 (N_33440,N_27647,N_25457);
nand U33441 (N_33441,N_23163,N_24098);
nor U33442 (N_33442,N_20291,N_20955);
xor U33443 (N_33443,N_22389,N_25621);
nor U33444 (N_33444,N_25829,N_21467);
nor U33445 (N_33445,N_23323,N_20595);
nand U33446 (N_33446,N_28802,N_23990);
and U33447 (N_33447,N_22318,N_22950);
nand U33448 (N_33448,N_28362,N_22648);
and U33449 (N_33449,N_22387,N_20016);
nor U33450 (N_33450,N_28983,N_24264);
nor U33451 (N_33451,N_24922,N_28024);
nand U33452 (N_33452,N_22912,N_28436);
and U33453 (N_33453,N_21245,N_20104);
or U33454 (N_33454,N_22856,N_22687);
nand U33455 (N_33455,N_23281,N_20339);
nand U33456 (N_33456,N_26816,N_21012);
nor U33457 (N_33457,N_27987,N_29788);
or U33458 (N_33458,N_24265,N_20895);
or U33459 (N_33459,N_26348,N_23691);
and U33460 (N_33460,N_29575,N_26809);
and U33461 (N_33461,N_24481,N_20177);
and U33462 (N_33462,N_27320,N_28394);
and U33463 (N_33463,N_22187,N_26005);
or U33464 (N_33464,N_23469,N_24897);
xnor U33465 (N_33465,N_29737,N_26713);
or U33466 (N_33466,N_27995,N_27141);
nor U33467 (N_33467,N_23347,N_21531);
nand U33468 (N_33468,N_25141,N_21947);
and U33469 (N_33469,N_29009,N_21099);
xnor U33470 (N_33470,N_26397,N_20101);
and U33471 (N_33471,N_28551,N_22523);
xnor U33472 (N_33472,N_24758,N_24543);
nor U33473 (N_33473,N_24888,N_28006);
nor U33474 (N_33474,N_23210,N_24877);
or U33475 (N_33475,N_27299,N_25545);
and U33476 (N_33476,N_21738,N_24442);
or U33477 (N_33477,N_23098,N_28976);
and U33478 (N_33478,N_21915,N_20801);
and U33479 (N_33479,N_26022,N_21182);
and U33480 (N_33480,N_29835,N_26946);
and U33481 (N_33481,N_23278,N_20186);
xor U33482 (N_33482,N_27094,N_20017);
nor U33483 (N_33483,N_28898,N_23402);
nor U33484 (N_33484,N_23079,N_25965);
or U33485 (N_33485,N_20691,N_22660);
and U33486 (N_33486,N_29941,N_23373);
nor U33487 (N_33487,N_27329,N_25833);
or U33488 (N_33488,N_25298,N_21183);
or U33489 (N_33489,N_29246,N_29624);
and U33490 (N_33490,N_20347,N_26090);
nor U33491 (N_33491,N_29754,N_25003);
nand U33492 (N_33492,N_26018,N_28559);
or U33493 (N_33493,N_26474,N_23957);
xnor U33494 (N_33494,N_24938,N_27619);
or U33495 (N_33495,N_23883,N_26863);
and U33496 (N_33496,N_22492,N_27163);
or U33497 (N_33497,N_29206,N_28227);
and U33498 (N_33498,N_21587,N_20051);
or U33499 (N_33499,N_24396,N_26310);
nand U33500 (N_33500,N_21407,N_21228);
nor U33501 (N_33501,N_21687,N_24764);
and U33502 (N_33502,N_23443,N_27836);
or U33503 (N_33503,N_21056,N_23685);
and U33504 (N_33504,N_29253,N_28676);
or U33505 (N_33505,N_21987,N_21391);
nand U33506 (N_33506,N_28042,N_26532);
or U33507 (N_33507,N_23380,N_20511);
and U33508 (N_33508,N_24703,N_27709);
nor U33509 (N_33509,N_21812,N_29524);
or U33510 (N_33510,N_20897,N_21105);
and U33511 (N_33511,N_25843,N_28928);
and U33512 (N_33512,N_23806,N_26202);
nand U33513 (N_33513,N_23510,N_23628);
or U33514 (N_33514,N_24389,N_25411);
and U33515 (N_33515,N_28467,N_25306);
xor U33516 (N_33516,N_23427,N_20626);
nand U33517 (N_33517,N_28570,N_22668);
nor U33518 (N_33518,N_21842,N_21210);
and U33519 (N_33519,N_20889,N_22857);
nor U33520 (N_33520,N_27357,N_28764);
or U33521 (N_33521,N_27601,N_26742);
or U33522 (N_33522,N_24351,N_27203);
and U33523 (N_33523,N_26833,N_24683);
nand U33524 (N_33524,N_21782,N_22663);
or U33525 (N_33525,N_20705,N_24908);
or U33526 (N_33526,N_24479,N_21155);
nor U33527 (N_33527,N_27664,N_27488);
and U33528 (N_33528,N_26783,N_20581);
or U33529 (N_33529,N_27623,N_28977);
or U33530 (N_33530,N_27055,N_25084);
and U33531 (N_33531,N_21526,N_24760);
or U33532 (N_33532,N_28094,N_25775);
xnor U33533 (N_33533,N_23865,N_26671);
nor U33534 (N_33534,N_27038,N_26405);
or U33535 (N_33535,N_22873,N_22837);
and U33536 (N_33536,N_21430,N_27696);
nand U33537 (N_33537,N_28840,N_21991);
nor U33538 (N_33538,N_22691,N_28066);
and U33539 (N_33539,N_23256,N_24302);
nand U33540 (N_33540,N_26455,N_23066);
and U33541 (N_33541,N_23989,N_25151);
or U33542 (N_33542,N_22051,N_20746);
nor U33543 (N_33543,N_25307,N_29881);
nor U33544 (N_33544,N_29312,N_22215);
nand U33545 (N_33545,N_29633,N_22194);
and U33546 (N_33546,N_29212,N_28519);
nor U33547 (N_33547,N_22119,N_20019);
and U33548 (N_33548,N_27842,N_20837);
or U33549 (N_33549,N_23398,N_24407);
xnor U33550 (N_33550,N_29579,N_27078);
nor U33551 (N_33551,N_27817,N_22274);
and U33552 (N_33552,N_25521,N_22941);
nand U33553 (N_33553,N_28080,N_22223);
nand U33554 (N_33554,N_29422,N_21339);
nand U33555 (N_33555,N_27688,N_29846);
nor U33556 (N_33556,N_28481,N_21576);
nor U33557 (N_33557,N_22525,N_25674);
nor U33558 (N_33558,N_26327,N_27238);
nor U33559 (N_33559,N_23244,N_20228);
or U33560 (N_33560,N_22338,N_27665);
and U33561 (N_33561,N_23291,N_29089);
and U33562 (N_33562,N_28301,N_23095);
nand U33563 (N_33563,N_24448,N_28825);
xor U33564 (N_33564,N_20063,N_28295);
nand U33565 (N_33565,N_20510,N_24899);
nand U33566 (N_33566,N_20215,N_22477);
xor U33567 (N_33567,N_27827,N_29964);
nor U33568 (N_33568,N_28165,N_20818);
or U33569 (N_33569,N_26138,N_22578);
or U33570 (N_33570,N_24608,N_25891);
nand U33571 (N_33571,N_29351,N_26611);
or U33572 (N_33572,N_20358,N_28852);
nor U33573 (N_33573,N_20477,N_22733);
xnor U33574 (N_33574,N_25077,N_26908);
nor U33575 (N_33575,N_21292,N_29493);
or U33576 (N_33576,N_21974,N_29164);
or U33577 (N_33577,N_22992,N_28344);
nor U33578 (N_33578,N_24223,N_21036);
xnor U33579 (N_33579,N_23771,N_25274);
nand U33580 (N_33580,N_28102,N_24737);
and U33581 (N_33581,N_21829,N_28317);
nor U33582 (N_33582,N_25189,N_22122);
or U33583 (N_33583,N_23463,N_21710);
and U33584 (N_33584,N_20785,N_21286);
nand U33585 (N_33585,N_23195,N_29901);
nand U33586 (N_33586,N_25641,N_28122);
nor U33587 (N_33587,N_26069,N_24783);
nor U33588 (N_33588,N_21760,N_29670);
nor U33589 (N_33589,N_20751,N_28409);
nor U33590 (N_33590,N_23877,N_24332);
and U33591 (N_33591,N_28331,N_29380);
and U33592 (N_33592,N_23541,N_23269);
xnor U33593 (N_33593,N_23328,N_26295);
xnor U33594 (N_33594,N_24464,N_27755);
nand U33595 (N_33595,N_26806,N_28132);
and U33596 (N_33596,N_29588,N_20838);
nand U33597 (N_33597,N_27383,N_23020);
or U33598 (N_33598,N_22939,N_26691);
or U33599 (N_33599,N_23906,N_22711);
or U33600 (N_33600,N_24446,N_28127);
nor U33601 (N_33601,N_27067,N_20995);
xor U33602 (N_33602,N_27427,N_24595);
and U33603 (N_33603,N_26135,N_26043);
nand U33604 (N_33604,N_22709,N_21189);
and U33605 (N_33605,N_29842,N_22821);
nand U33606 (N_33606,N_23540,N_23428);
nor U33607 (N_33607,N_28654,N_26156);
nor U33608 (N_33608,N_26447,N_29310);
xor U33609 (N_33609,N_20823,N_28109);
nand U33610 (N_33610,N_29370,N_22624);
and U33611 (N_33611,N_22662,N_20152);
and U33612 (N_33612,N_28191,N_27683);
or U33613 (N_33613,N_21659,N_23075);
xnor U33614 (N_33614,N_25675,N_25202);
nor U33615 (N_33615,N_24155,N_24465);
or U33616 (N_33616,N_29760,N_24907);
and U33617 (N_33617,N_27475,N_27342);
nor U33618 (N_33618,N_21732,N_22545);
nor U33619 (N_33619,N_26272,N_29974);
or U33620 (N_33620,N_24449,N_27937);
nand U33621 (N_33621,N_22436,N_29903);
and U33622 (N_33622,N_29239,N_26857);
or U33623 (N_33623,N_26220,N_25597);
nor U33624 (N_33624,N_29403,N_29007);
and U33625 (N_33625,N_21207,N_28268);
and U33626 (N_33626,N_29653,N_26674);
and U33627 (N_33627,N_22639,N_21141);
or U33628 (N_33628,N_23023,N_22349);
xnor U33629 (N_33629,N_20420,N_21134);
nand U33630 (N_33630,N_23588,N_24597);
or U33631 (N_33631,N_20381,N_26269);
nor U33632 (N_33632,N_27304,N_28242);
nor U33633 (N_33633,N_21027,N_28553);
and U33634 (N_33634,N_28829,N_20348);
nand U33635 (N_33635,N_22786,N_23770);
xor U33636 (N_33636,N_21279,N_28076);
nand U33637 (N_33637,N_20286,N_20612);
or U33638 (N_33638,N_23166,N_22366);
and U33639 (N_33639,N_23423,N_29991);
and U33640 (N_33640,N_22257,N_27938);
xnor U33641 (N_33641,N_20950,N_29471);
nand U33642 (N_33642,N_22294,N_22262);
nand U33643 (N_33643,N_29232,N_23122);
nor U33644 (N_33644,N_21610,N_25439);
or U33645 (N_33645,N_20576,N_28114);
xor U33646 (N_33646,N_25266,N_24113);
nand U33647 (N_33647,N_26439,N_24394);
and U33648 (N_33648,N_22898,N_28356);
and U33649 (N_33649,N_21030,N_24799);
or U33650 (N_33650,N_21197,N_26609);
nor U33651 (N_33651,N_29216,N_22266);
nand U33652 (N_33652,N_23320,N_24322);
nand U33653 (N_33653,N_22101,N_25682);
and U33654 (N_33654,N_22681,N_25636);
nor U33655 (N_33655,N_21400,N_23225);
or U33656 (N_33656,N_25081,N_26144);
or U33657 (N_33657,N_23899,N_20267);
or U33658 (N_33658,N_23127,N_24832);
and U33659 (N_33659,N_26178,N_22248);
nand U33660 (N_33660,N_27705,N_24475);
and U33661 (N_33661,N_27517,N_22038);
nand U33662 (N_33662,N_24092,N_29419);
or U33663 (N_33663,N_21149,N_20909);
nor U33664 (N_33664,N_25964,N_21741);
nand U33665 (N_33665,N_24026,N_28716);
nand U33666 (N_33666,N_24518,N_29431);
nor U33667 (N_33667,N_29179,N_20577);
xor U33668 (N_33668,N_24724,N_21669);
nor U33669 (N_33669,N_24009,N_24669);
xor U33670 (N_33670,N_21474,N_26936);
nand U33671 (N_33671,N_24882,N_23761);
nand U33672 (N_33672,N_27424,N_20092);
xor U33673 (N_33673,N_24076,N_24450);
nand U33674 (N_33674,N_29857,N_23317);
xnor U33675 (N_33675,N_20093,N_29108);
nand U33676 (N_33676,N_23580,N_22899);
and U33677 (N_33677,N_21804,N_25510);
nor U33678 (N_33678,N_29797,N_29078);
nand U33679 (N_33679,N_20703,N_27420);
or U33680 (N_33680,N_26701,N_21854);
and U33681 (N_33681,N_29014,N_21029);
nand U33682 (N_33682,N_20625,N_24359);
or U33683 (N_33683,N_27185,N_22172);
and U33684 (N_33684,N_28171,N_27351);
and U33685 (N_33685,N_25619,N_26735);
or U33686 (N_33686,N_25662,N_21399);
and U33687 (N_33687,N_26860,N_26612);
or U33688 (N_33688,N_26914,N_25071);
xor U33689 (N_33689,N_27944,N_20980);
xnor U33690 (N_33690,N_27270,N_21242);
xor U33691 (N_33691,N_21237,N_26842);
xor U33692 (N_33692,N_27044,N_27719);
nand U33693 (N_33693,N_22144,N_25280);
nand U33694 (N_33694,N_28588,N_26529);
and U33695 (N_33695,N_20813,N_28434);
and U33696 (N_33696,N_25144,N_26139);
and U33697 (N_33697,N_24329,N_27614);
nand U33698 (N_33698,N_27252,N_27385);
and U33699 (N_33699,N_23639,N_24651);
and U33700 (N_33700,N_29235,N_20718);
nand U33701 (N_33701,N_23702,N_29274);
and U33702 (N_33702,N_24433,N_28810);
nand U33703 (N_33703,N_22757,N_21050);
or U33704 (N_33704,N_26066,N_22649);
nor U33705 (N_33705,N_25565,N_27254);
and U33706 (N_33706,N_22445,N_24145);
and U33707 (N_33707,N_23972,N_24600);
nor U33708 (N_33708,N_27261,N_27898);
nor U33709 (N_33709,N_26670,N_24412);
or U33710 (N_33710,N_27003,N_28621);
nor U33711 (N_33711,N_22945,N_27685);
nand U33712 (N_33712,N_28385,N_27518);
nor U33713 (N_33713,N_24808,N_23956);
nand U33714 (N_33714,N_24005,N_29060);
nand U33715 (N_33715,N_28534,N_21685);
nor U33716 (N_33716,N_20585,N_28880);
or U33717 (N_33717,N_24813,N_29228);
xnor U33718 (N_33718,N_20698,N_27455);
or U33719 (N_33719,N_26085,N_23672);
nor U33720 (N_33720,N_20804,N_23341);
nand U33721 (N_33721,N_21637,N_25451);
nor U33722 (N_33722,N_26078,N_20580);
xnor U33723 (N_33723,N_28763,N_21656);
nor U33724 (N_33724,N_27508,N_25183);
xor U33725 (N_33725,N_26417,N_22413);
nor U33726 (N_33726,N_23911,N_22495);
or U33727 (N_33727,N_21575,N_24773);
and U33728 (N_33728,N_24753,N_23030);
nor U33729 (N_33729,N_29123,N_22412);
or U33730 (N_33730,N_21906,N_21627);
and U33731 (N_33731,N_25617,N_25869);
nor U33732 (N_33732,N_28069,N_29807);
or U33733 (N_33733,N_27922,N_20283);
or U33734 (N_33734,N_26986,N_29892);
nor U33735 (N_33735,N_23696,N_20004);
nor U33736 (N_33736,N_20060,N_20782);
nor U33737 (N_33737,N_29617,N_29932);
and U33738 (N_33738,N_22401,N_25343);
and U33739 (N_33739,N_26282,N_26950);
nor U33740 (N_33740,N_25149,N_29839);
or U33741 (N_33741,N_24087,N_28515);
or U33742 (N_33742,N_28395,N_20061);
nand U33743 (N_33743,N_29328,N_20306);
nand U33744 (N_33744,N_22249,N_23871);
and U33745 (N_33745,N_23932,N_23100);
and U33746 (N_33746,N_24892,N_20068);
and U33747 (N_33747,N_25441,N_23496);
nor U33748 (N_33748,N_21362,N_23288);
xor U33749 (N_33749,N_27041,N_24340);
nor U33750 (N_33750,N_22180,N_28668);
or U33751 (N_33751,N_24142,N_28860);
or U33752 (N_33752,N_22959,N_26889);
nor U33753 (N_33753,N_29059,N_27154);
nand U33754 (N_33754,N_24541,N_26164);
or U33755 (N_33755,N_26118,N_25148);
or U33756 (N_33756,N_25052,N_24995);
nor U33757 (N_33757,N_22217,N_28727);
and U33758 (N_33758,N_26978,N_20084);
nor U33759 (N_33759,N_27173,N_25060);
and U33760 (N_33760,N_21371,N_26113);
and U33761 (N_33761,N_23891,N_26107);
nand U33762 (N_33762,N_26659,N_25533);
nand U33763 (N_33763,N_22402,N_28739);
and U33764 (N_33764,N_21143,N_22535);
and U33765 (N_33765,N_20485,N_21117);
nand U33766 (N_33766,N_26650,N_24503);
nand U33767 (N_33767,N_28823,N_27469);
and U33768 (N_33768,N_26796,N_27822);
and U33769 (N_33769,N_21158,N_20272);
nand U33770 (N_33770,N_28470,N_24150);
nor U33771 (N_33771,N_27546,N_29818);
nor U33772 (N_33772,N_20618,N_28672);
or U33773 (N_33773,N_27023,N_21689);
or U33774 (N_33774,N_21205,N_27177);
and U33775 (N_33775,N_25644,N_29247);
or U33776 (N_33776,N_23052,N_28987);
nand U33777 (N_33777,N_23881,N_23848);
or U33778 (N_33778,N_29296,N_23344);
nor U33779 (N_33779,N_21993,N_27188);
xnor U33780 (N_33780,N_25555,N_23757);
nand U33781 (N_33781,N_22517,N_20905);
and U33782 (N_33782,N_27459,N_22902);
nand U33783 (N_33783,N_27245,N_29485);
nand U33784 (N_33784,N_26319,N_27798);
nor U33785 (N_33785,N_28479,N_26288);
and U33786 (N_33786,N_28465,N_29731);
and U33787 (N_33787,N_28273,N_26314);
nand U33788 (N_33788,N_26781,N_26448);
or U33789 (N_33789,N_27523,N_28002);
nor U33790 (N_33790,N_26921,N_24069);
nor U33791 (N_33791,N_21790,N_26160);
or U33792 (N_33792,N_29597,N_24502);
nand U33793 (N_33793,N_23667,N_21765);
nand U33794 (N_33794,N_28257,N_21004);
or U33795 (N_33795,N_24870,N_21249);
nand U33796 (N_33796,N_20288,N_21508);
nor U33797 (N_33797,N_20715,N_26049);
nor U33798 (N_33798,N_29318,N_23445);
nor U33799 (N_33799,N_27021,N_22056);
xor U33800 (N_33800,N_24182,N_24915);
nand U33801 (N_33801,N_21127,N_21734);
and U33802 (N_33802,N_25342,N_27448);
nor U33803 (N_33803,N_20089,N_21740);
or U33804 (N_33804,N_21060,N_27294);
or U33805 (N_33805,N_24175,N_21212);
nor U33806 (N_33806,N_24358,N_21724);
nand U33807 (N_33807,N_28805,N_24866);
nand U33808 (N_33808,N_20155,N_25895);
and U33809 (N_33809,N_29069,N_27481);
or U33810 (N_33810,N_20643,N_21164);
and U33811 (N_33811,N_27778,N_25542);
nor U33812 (N_33812,N_21274,N_28610);
and U33813 (N_33813,N_23907,N_20290);
or U33814 (N_33814,N_21481,N_26116);
nor U33815 (N_33815,N_24635,N_25402);
and U33816 (N_33816,N_26597,N_28097);
nor U33817 (N_33817,N_26947,N_20144);
nor U33818 (N_33818,N_25598,N_26568);
nand U33819 (N_33819,N_29574,N_22809);
nand U33820 (N_33820,N_26318,N_25217);
nand U33821 (N_33821,N_23048,N_24253);
and U33822 (N_33822,N_24561,N_26279);
nor U33823 (N_33823,N_29551,N_25651);
nand U33824 (N_33824,N_29845,N_26727);
nor U33825 (N_33825,N_29484,N_29199);
nor U33826 (N_33826,N_28204,N_28206);
nand U33827 (N_33827,N_29852,N_27746);
nand U33828 (N_33828,N_25799,N_26147);
or U33829 (N_33829,N_25128,N_20986);
nor U33830 (N_33830,N_28261,N_23845);
and U33831 (N_33831,N_29222,N_26115);
or U33832 (N_33832,N_24632,N_27359);
nor U33833 (N_33833,N_22440,N_29900);
and U33834 (N_33834,N_27868,N_25381);
or U33835 (N_33835,N_26630,N_23994);
or U33836 (N_33836,N_23181,N_27743);
xor U33837 (N_33837,N_21988,N_29178);
nor U33838 (N_33838,N_29137,N_23779);
nand U33839 (N_33839,N_20421,N_29603);
and U33840 (N_33840,N_28329,N_24580);
nand U33841 (N_33841,N_28150,N_27011);
nor U33842 (N_33842,N_28476,N_26723);
nor U33843 (N_33843,N_27736,N_23700);
nand U33844 (N_33844,N_25591,N_27253);
nor U33845 (N_33845,N_28032,N_27332);
nor U33846 (N_33846,N_20653,N_26976);
nor U33847 (N_33847,N_26340,N_23668);
nor U33848 (N_33848,N_28175,N_27289);
nor U33849 (N_33849,N_22252,N_26337);
nor U33850 (N_33850,N_26688,N_25539);
nor U33851 (N_33851,N_25581,N_29793);
nand U33852 (N_33852,N_28159,N_22841);
nand U33853 (N_33853,N_28239,N_23287);
nor U33854 (N_33854,N_22025,N_23376);
and U33855 (N_33855,N_27049,N_20525);
or U33856 (N_33856,N_22629,N_28112);
nor U33857 (N_33857,N_25879,N_20863);
nor U33858 (N_33858,N_29677,N_29536);
or U33859 (N_33859,N_28145,N_27874);
nand U33860 (N_33860,N_26768,N_21830);
and U33861 (N_33861,N_21673,N_24410);
nor U33862 (N_33862,N_21309,N_27820);
or U33863 (N_33863,N_23057,N_27825);
and U33864 (N_33864,N_28541,N_28733);
or U33865 (N_33865,N_20199,N_20120);
and U33866 (N_33866,N_27178,N_24827);
or U33867 (N_33867,N_20606,N_24570);
nand U33868 (N_33868,N_22078,N_25022);
xor U33869 (N_33869,N_24081,N_21472);
and U33870 (N_33870,N_25246,N_24338);
and U33871 (N_33871,N_24445,N_23208);
nand U33872 (N_33872,N_25988,N_26820);
nor U33873 (N_33873,N_21342,N_20278);
and U33874 (N_33874,N_20049,N_24691);
nand U33875 (N_33875,N_21345,N_26411);
nor U33876 (N_33876,N_24493,N_24638);
xnor U33877 (N_33877,N_22414,N_27379);
nor U33878 (N_33878,N_22234,N_29262);
nor U33879 (N_33879,N_28283,N_29584);
xor U33880 (N_33880,N_29621,N_20128);
or U33881 (N_33881,N_27865,N_20891);
nand U33882 (N_33882,N_27161,N_28202);
nor U33883 (N_33883,N_22383,N_29475);
nand U33884 (N_33884,N_27756,N_25671);
nand U33885 (N_33885,N_20293,N_22373);
nand U33886 (N_33886,N_24914,N_28735);
nand U33887 (N_33887,N_26695,N_24272);
nand U33888 (N_33888,N_20328,N_24235);
nand U33889 (N_33889,N_24148,N_24891);
and U33890 (N_33890,N_21209,N_27723);
or U33891 (N_33891,N_29538,N_27325);
and U33892 (N_33892,N_26541,N_26675);
nor U33893 (N_33893,N_22870,N_22597);
or U33894 (N_33894,N_24739,N_20112);
or U33895 (N_33895,N_21884,N_29001);
and U33896 (N_33896,N_22970,N_25605);
nor U33897 (N_33897,N_23447,N_26808);
nor U33898 (N_33898,N_28878,N_29053);
or U33899 (N_33899,N_20575,N_23470);
nor U33900 (N_33900,N_21813,N_25293);
nand U33901 (N_33901,N_24079,N_25781);
and U33902 (N_33902,N_26050,N_26021);
or U33903 (N_33903,N_20617,N_29497);
nor U33904 (N_33904,N_22498,N_29979);
nor U33905 (N_33905,N_22574,N_29221);
nand U33906 (N_33906,N_27754,N_26389);
nor U33907 (N_33907,N_21643,N_26410);
or U33908 (N_33908,N_23262,N_20279);
and U33909 (N_33909,N_26145,N_26774);
or U33910 (N_33910,N_23703,N_20830);
nand U33911 (N_33911,N_20174,N_24554);
nand U33912 (N_33912,N_23687,N_28701);
nand U33913 (N_33913,N_27308,N_27896);
nand U33914 (N_33914,N_23101,N_28229);
nor U33915 (N_33915,N_23070,N_23933);
and U33916 (N_33916,N_28477,N_23698);
and U33917 (N_33917,N_28684,N_20560);
nand U33918 (N_33918,N_27787,N_24224);
xor U33919 (N_33919,N_29833,N_25040);
and U33920 (N_33920,N_25822,N_26913);
or U33921 (N_33921,N_29309,N_20821);
nor U33922 (N_33922,N_28167,N_29739);
xnor U33923 (N_33923,N_21232,N_23361);
nand U33924 (N_33924,N_21674,N_22333);
nand U33925 (N_33925,N_21288,N_22381);
and U33926 (N_33926,N_20769,N_21355);
nand U33927 (N_33927,N_26637,N_27229);
nor U33928 (N_33928,N_26012,N_23162);
nand U33929 (N_33929,N_28157,N_27872);
nor U33930 (N_33930,N_23717,N_21881);
or U33931 (N_33931,N_29113,N_26966);
nor U33932 (N_33932,N_23387,N_27764);
xor U33933 (N_33933,N_25746,N_23138);
or U33934 (N_33934,N_20669,N_23546);
nor U33935 (N_33935,N_29856,N_24519);
and U33936 (N_33936,N_20619,N_20066);
nand U33937 (N_33937,N_25751,N_24192);
nor U33938 (N_33938,N_27086,N_27256);
or U33939 (N_33939,N_26209,N_23358);
nand U33940 (N_33940,N_27873,N_27711);
or U33941 (N_33941,N_21681,N_26212);
or U33942 (N_33942,N_27932,N_29492);
xnor U33943 (N_33943,N_27278,N_25184);
or U33944 (N_33944,N_28148,N_20561);
and U33945 (N_33945,N_28412,N_21236);
nand U33946 (N_33946,N_23316,N_23701);
nor U33947 (N_33947,N_28604,N_20171);
and U33948 (N_33948,N_26201,N_27971);
and U33949 (N_33949,N_27584,N_25688);
and U33950 (N_33950,N_26470,N_25748);
or U33951 (N_33951,N_24804,N_20786);
or U33952 (N_33952,N_24552,N_28607);
or U33953 (N_33953,N_21727,N_28584);
nor U33954 (N_33954,N_28834,N_25992);
nor U33955 (N_33955,N_20209,N_21453);
nand U33956 (N_33956,N_29052,N_22922);
and U33957 (N_33957,N_24080,N_24203);
nand U33958 (N_33958,N_26793,N_28526);
and U33959 (N_33959,N_24129,N_20032);
nand U33960 (N_33960,N_26253,N_20822);
nor U33961 (N_33961,N_22661,N_25129);
nand U33962 (N_33962,N_24021,N_28305);
or U33963 (N_33963,N_25958,N_21276);
and U33964 (N_33964,N_29542,N_20054);
nand U33965 (N_33965,N_28074,N_23226);
and U33966 (N_33966,N_22877,N_25220);
nor U33967 (N_33967,N_27181,N_25714);
or U33968 (N_33968,N_20578,N_27167);
or U33969 (N_33969,N_25715,N_22675);
nor U33970 (N_33970,N_26307,N_27701);
and U33971 (N_33971,N_28070,N_28496);
nor U33972 (N_33972,N_29870,N_21510);
and U33973 (N_33973,N_26859,N_23902);
nor U33974 (N_33974,N_20851,N_23900);
nand U33975 (N_33975,N_28818,N_22780);
or U33976 (N_33976,N_23033,N_28656);
and U33977 (N_33977,N_24806,N_28797);
and U33978 (N_33978,N_23349,N_21218);
or U33979 (N_33979,N_25438,N_27830);
nor U33980 (N_33980,N_26928,N_27180);
and U33981 (N_33981,N_25720,N_26229);
nor U33982 (N_33982,N_29637,N_28423);
nand U33983 (N_33983,N_25136,N_25978);
or U33984 (N_33984,N_25147,N_20994);
nand U33985 (N_33985,N_28264,N_22975);
nor U33986 (N_33986,N_22326,N_20588);
nand U33987 (N_33987,N_25111,N_24054);
or U33988 (N_33988,N_20656,N_23246);
nand U33989 (N_33989,N_27724,N_29396);
xnor U33990 (N_33990,N_21594,N_28049);
nor U33991 (N_33991,N_28466,N_23590);
nor U33992 (N_33992,N_20491,N_21223);
or U33993 (N_33993,N_27201,N_22135);
nand U33994 (N_33994,N_26547,N_26998);
nor U33995 (N_33995,N_26629,N_27072);
nor U33996 (N_33996,N_20825,N_21426);
nand U33997 (N_33997,N_21003,N_20740);
xor U33998 (N_33998,N_24163,N_24501);
or U33999 (N_33999,N_29375,N_24613);
and U34000 (N_34000,N_20006,N_28790);
xor U34001 (N_34001,N_21323,N_26332);
nor U34002 (N_34002,N_25530,N_22811);
nand U34003 (N_34003,N_26933,N_20315);
or U34004 (N_34004,N_22088,N_28418);
and U34005 (N_34005,N_21161,N_24693);
or U34006 (N_34006,N_27132,N_23508);
or U34007 (N_34007,N_23752,N_21199);
nor U34008 (N_34008,N_27784,N_21582);
xnor U34009 (N_34009,N_22672,N_25744);
nand U34010 (N_34010,N_29448,N_23863);
nor U34011 (N_34011,N_22561,N_21666);
xnor U34012 (N_34012,N_27431,N_28176);
nor U34013 (N_34013,N_20263,N_29092);
nand U34014 (N_34014,N_27002,N_28269);
and U34015 (N_34015,N_21454,N_25696);
or U34016 (N_34016,N_22779,N_27190);
and U34017 (N_34017,N_26075,N_21451);
xnor U34018 (N_34018,N_26193,N_22453);
nand U34019 (N_34019,N_23603,N_22491);
xnor U34020 (N_34020,N_29698,N_23498);
nor U34021 (N_34021,N_28469,N_22105);
or U34022 (N_34022,N_26443,N_25687);
or U34023 (N_34023,N_28659,N_26934);
nand U34024 (N_34024,N_20034,N_24222);
nand U34025 (N_34025,N_27881,N_25905);
or U34026 (N_34026,N_28886,N_23613);
or U34027 (N_34027,N_28023,N_27788);
nand U34028 (N_34028,N_26718,N_27557);
nand U34029 (N_34029,N_26938,N_25620);
or U34030 (N_34030,N_27646,N_26326);
nor U34031 (N_34031,N_27525,N_24547);
nand U34032 (N_34032,N_21204,N_27390);
nor U34033 (N_34033,N_21779,N_28757);
nand U34034 (N_34034,N_21487,N_24023);
nand U34035 (N_34035,N_23864,N_28694);
nand U34036 (N_34036,N_22202,N_26578);
and U34037 (N_34037,N_22238,N_29189);
nor U34038 (N_34038,N_27795,N_22827);
xor U34039 (N_34039,N_22354,N_20518);
nor U34040 (N_34040,N_22707,N_25885);
nor U34041 (N_34041,N_26549,N_23975);
or U34042 (N_34042,N_22241,N_26531);
and U34043 (N_34043,N_21930,N_21954);
and U34044 (N_34044,N_26827,N_29152);
or U34045 (N_34045,N_25460,N_20571);
or U34046 (N_34046,N_21518,N_26681);
and U34047 (N_34047,N_24106,N_27695);
nor U34048 (N_34048,N_22526,N_24525);
nor U34049 (N_34049,N_25518,N_27627);
and U34050 (N_34050,N_21496,N_25130);
nand U34051 (N_34051,N_26738,N_22439);
xnor U34052 (N_34052,N_23472,N_22385);
or U34053 (N_34053,N_28100,N_20600);
nand U34054 (N_34054,N_22947,N_23170);
or U34055 (N_34055,N_21752,N_21894);
nor U34056 (N_34056,N_28708,N_28081);
or U34057 (N_34057,N_29514,N_28478);
and U34058 (N_34058,N_23841,N_25957);
or U34059 (N_34059,N_26414,N_26218);
and U34060 (N_34060,N_27704,N_21354);
nor U34061 (N_34061,N_24162,N_29977);
nand U34062 (N_34062,N_20880,N_25660);
nor U34063 (N_34063,N_22867,N_22581);
nor U34064 (N_34064,N_23852,N_26296);
or U34065 (N_34065,N_23738,N_20783);
xor U34066 (N_34066,N_24312,N_24458);
and U34067 (N_34067,N_22693,N_23227);
nor U34068 (N_34068,N_23862,N_20007);
or U34069 (N_34069,N_26460,N_28954);
or U34070 (N_34070,N_25503,N_27581);
xor U34071 (N_34071,N_28393,N_28592);
or U34072 (N_34072,N_25818,N_21556);
and U34073 (N_34073,N_28828,N_22062);
or U34074 (N_34074,N_22805,N_24024);
and U34075 (N_34075,N_28760,N_24072);
or U34076 (N_34076,N_22790,N_28480);
and U34077 (N_34077,N_26822,N_22860);
nand U34078 (N_34078,N_25221,N_24664);
nor U34079 (N_34079,N_22684,N_29981);
or U34080 (N_34080,N_21414,N_21826);
and U34081 (N_34081,N_28215,N_27358);
xnor U34082 (N_34082,N_29805,N_25910);
nor U34083 (N_34083,N_28711,N_20629);
or U34084 (N_34084,N_20379,N_28997);
and U34085 (N_34085,N_27164,N_21043);
nor U34086 (N_34086,N_24831,N_24011);
nand U34087 (N_34087,N_26463,N_28736);
and U34088 (N_34088,N_22893,N_22613);
nand U34089 (N_34089,N_22611,N_26189);
or U34090 (N_34090,N_23308,N_24980);
or U34091 (N_34091,N_24043,N_25479);
nand U34092 (N_34092,N_25918,N_28235);
nand U34093 (N_34093,N_25185,N_22134);
and U34094 (N_34094,N_20748,N_29359);
nand U34095 (N_34095,N_21358,N_29186);
or U34096 (N_34096,N_28737,N_24801);
nor U34097 (N_34097,N_25051,N_28606);
nor U34098 (N_34098,N_26353,N_25616);
nor U34099 (N_34099,N_20461,N_21766);
nor U34100 (N_34100,N_28773,N_25881);
or U34101 (N_34101,N_29980,N_26498);
xnor U34102 (N_34102,N_27947,N_24262);
and U34103 (N_34103,N_29969,N_24588);
or U34104 (N_34104,N_22277,N_27392);
nor U34105 (N_34105,N_29460,N_25417);
nor U34106 (N_34106,N_24127,N_24883);
and U34107 (N_34107,N_24567,N_22066);
and U34108 (N_34108,N_26631,N_26517);
and U34109 (N_34109,N_25755,N_24700);
and U34110 (N_34110,N_23986,N_25421);
or U34111 (N_34111,N_29649,N_22201);
nand U34112 (N_34112,N_29294,N_23809);
and U34113 (N_34113,N_26800,N_22755);
or U34114 (N_34114,N_22372,N_22653);
nor U34115 (N_34115,N_25143,N_29681);
and U34116 (N_34116,N_23815,N_20196);
nor U34117 (N_34117,N_22920,N_25276);
and U34118 (N_34118,N_26956,N_24003);
nand U34119 (N_34119,N_23857,N_28497);
nor U34120 (N_34120,N_29559,N_25496);
nor U34121 (N_34121,N_21965,N_22915);
or U34122 (N_34122,N_21933,N_26899);
nor U34123 (N_34123,N_29000,N_24391);
and U34124 (N_34124,N_26277,N_21593);
and U34125 (N_34125,N_28665,N_20840);
nor U34126 (N_34126,N_27221,N_22888);
xnor U34127 (N_34127,N_25810,N_25976);
or U34128 (N_34128,N_21045,N_28508);
nor U34129 (N_34129,N_22883,N_20788);
and U34130 (N_34130,N_22456,N_29586);
nand U34131 (N_34131,N_23251,N_26354);
or U34132 (N_34132,N_21630,N_28411);
nand U34133 (N_34133,N_27797,N_21692);
or U34134 (N_34134,N_21568,N_23235);
nand U34135 (N_34135,N_24456,N_27069);
and U34136 (N_34136,N_24823,N_20247);
or U34137 (N_34137,N_24636,N_22799);
nor U34138 (N_34138,N_29418,N_28383);
nand U34139 (N_34139,N_25476,N_22114);
xor U34140 (N_34140,N_24418,N_27241);
nor U34141 (N_34141,N_28666,N_22315);
or U34142 (N_34142,N_23642,N_25552);
and U34143 (N_34143,N_26566,N_21825);
nand U34144 (N_34144,N_27323,N_21014);
xor U34145 (N_34145,N_26504,N_29639);
nor U34146 (N_34146,N_26412,N_20681);
nand U34147 (N_34147,N_26605,N_25913);
xor U34148 (N_34148,N_29355,N_27353);
or U34149 (N_34149,N_26106,N_29694);
nor U34150 (N_34150,N_25359,N_28507);
and U34151 (N_34151,N_23378,N_26927);
nor U34152 (N_34152,N_29171,N_23567);
nor U34153 (N_34153,N_26617,N_29875);
or U34154 (N_34154,N_22760,N_26555);
and U34155 (N_34155,N_25215,N_25092);
nor U34156 (N_34156,N_27735,N_26328);
nand U34157 (N_34157,N_24769,N_20330);
nor U34158 (N_34158,N_28658,N_24228);
nand U34159 (N_34159,N_21324,N_29163);
or U34160 (N_34160,N_28724,N_24147);
and U34161 (N_34161,N_28692,N_28931);
nor U34162 (N_34162,N_27096,N_25608);
and U34163 (N_34163,N_29068,N_21074);
or U34164 (N_34164,N_24343,N_26732);
nor U34165 (N_34165,N_23711,N_25519);
and U34166 (N_34166,N_20240,N_25648);
nand U34167 (N_34167,N_28770,N_23520);
and U34168 (N_34168,N_20710,N_26068);
or U34169 (N_34169,N_28725,N_20344);
nand U34170 (N_34170,N_28155,N_21584);
xnor U34171 (N_34171,N_25284,N_25064);
or U34172 (N_34172,N_22365,N_28144);
xnor U34173 (N_34173,N_25433,N_29483);
nand U34174 (N_34174,N_25973,N_26274);
nand U34175 (N_34175,N_20712,N_28919);
and U34176 (N_34176,N_28552,N_26231);
nor U34177 (N_34177,N_24381,N_28460);
xor U34178 (N_34178,N_28567,N_26305);
nand U34179 (N_34179,N_25285,N_25575);
or U34180 (N_34180,N_26762,N_26478);
nor U34181 (N_34181,N_24303,N_26486);
and U34182 (N_34182,N_24881,N_20319);
nor U34183 (N_34183,N_20468,N_24646);
nor U34184 (N_34184,N_21374,N_24656);
nor U34185 (N_34185,N_23679,N_24746);
nand U34186 (N_34186,N_25094,N_25323);
nor U34187 (N_34187,N_27012,N_26939);
or U34188 (N_34188,N_25509,N_27514);
nor U34189 (N_34189,N_23794,N_22910);
or U34190 (N_34190,N_25316,N_21515);
nor U34191 (N_34191,N_27277,N_21623);
or U34192 (N_34192,N_28440,N_21278);
and U34193 (N_34193,N_21388,N_25072);
or U34194 (N_34194,N_23016,N_26880);
and U34195 (N_34195,N_25703,N_22881);
or U34196 (N_34196,N_20069,N_24788);
or U34197 (N_34197,N_29207,N_21293);
nand U34198 (N_34198,N_26618,N_24325);
and U34199 (N_34199,N_24289,N_20697);
and U34200 (N_34200,N_21899,N_22825);
nor U34201 (N_34201,N_28801,N_24984);
nor U34202 (N_34202,N_22616,N_21317);
nor U34203 (N_34203,N_27964,N_29784);
nand U34204 (N_34204,N_25219,N_20025);
nor U34205 (N_34205,N_23749,N_25190);
or U34206 (N_34206,N_22503,N_21529);
nand U34207 (N_34207,N_21377,N_22551);
nand U34208 (N_34208,N_20907,N_25603);
and U34209 (N_34209,N_25007,N_24723);
nand U34210 (N_34210,N_23763,N_20094);
xor U34211 (N_34211,N_24491,N_24385);
or U34212 (N_34212,N_21062,N_29629);
nand U34213 (N_34213,N_27377,N_24083);
nand U34214 (N_34214,N_21121,N_27165);
and U34215 (N_34215,N_22384,N_21565);
or U34216 (N_34216,N_28843,N_24555);
xnor U34217 (N_34217,N_20308,N_28406);
nor U34218 (N_34218,N_20222,N_22466);
and U34219 (N_34219,N_23787,N_20921);
and U34220 (N_34220,N_29085,N_27479);
and U34221 (N_34221,N_20965,N_27341);
xor U34222 (N_34222,N_24034,N_28323);
and U34223 (N_34223,N_21834,N_22914);
nor U34224 (N_34224,N_24405,N_24953);
and U34225 (N_34225,N_22636,N_26039);
and U34226 (N_34226,N_25380,N_27458);
nor U34227 (N_34227,N_24088,N_27246);
nand U34228 (N_34228,N_29682,N_27101);
nand U34229 (N_34229,N_24911,N_29949);
or U34230 (N_34230,N_28266,N_28267);
nor U34231 (N_34231,N_27981,N_21959);
and U34232 (N_34232,N_27655,N_29097);
and U34233 (N_34233,N_28249,N_28979);
nand U34234 (N_34234,N_22996,N_26901);
nand U34235 (N_34235,N_27668,N_26801);
nand U34236 (N_34236,N_24352,N_22839);
xnor U34237 (N_34237,N_24193,N_26268);
and U34238 (N_34238,N_29169,N_24744);
nor U34239 (N_34239,N_20254,N_25989);
xor U34240 (N_34240,N_21176,N_25109);
or U34241 (N_34241,N_28208,N_29423);
and U34242 (N_34242,N_25511,N_29566);
nor U34243 (N_34243,N_22740,N_26311);
xnor U34244 (N_34244,N_28693,N_27439);
and U34245 (N_34245,N_29173,N_28781);
and U34246 (N_34246,N_21037,N_21635);
xor U34247 (N_34247,N_20620,N_27184);
nand U34248 (N_34248,N_25173,N_22874);
nor U34249 (N_34249,N_20683,N_20026);
xnor U34250 (N_34250,N_26551,N_22831);
nand U34251 (N_34251,N_23026,N_27064);
nand U34252 (N_34252,N_24659,N_23778);
nor U34253 (N_34253,N_21463,N_25155);
nor U34254 (N_34254,N_26133,N_25258);
nor U34255 (N_34255,N_22564,N_26580);
nand U34256 (N_34256,N_23489,N_23401);
nand U34257 (N_34257,N_28101,N_26628);
and U34258 (N_34258,N_23136,N_24528);
nor U34259 (N_34259,N_26375,N_23851);
nand U34260 (N_34260,N_26148,N_26142);
and U34261 (N_34261,N_20996,N_24285);
nand U34262 (N_34262,N_25011,N_29925);
or U34263 (N_34263,N_25904,N_27421);
xnor U34264 (N_34264,N_24791,N_20232);
xnor U34265 (N_34265,N_22095,N_26614);
xor U34266 (N_34266,N_24108,N_25713);
xnor U34267 (N_34267,N_25800,N_22659);
and U34268 (N_34268,N_29726,N_28630);
and U34269 (N_34269,N_22444,N_23583);
nand U34270 (N_34270,N_26622,N_23967);
nand U34271 (N_34271,N_25085,N_20091);
xor U34272 (N_34272,N_28556,N_22802);
and U34273 (N_34273,N_26213,N_24283);
nand U34274 (N_34274,N_22118,N_25235);
nand U34275 (N_34275,N_28509,N_26275);
or U34276 (N_34276,N_20857,N_24716);
and U34277 (N_34277,N_20322,N_29590);
and U34278 (N_34278,N_24360,N_27259);
and U34279 (N_34279,N_25567,N_26920);
and U34280 (N_34280,N_28403,N_28593);
nor U34281 (N_34281,N_25456,N_20795);
or U34282 (N_34282,N_27776,N_26926);
nor U34283 (N_34283,N_26588,N_29374);
or U34284 (N_34284,N_26596,N_26054);
or U34285 (N_34285,N_20271,N_21061);
and U34286 (N_34286,N_25614,N_28373);
and U34287 (N_34287,N_20972,N_24179);
or U34288 (N_34288,N_29783,N_29473);
nor U34289 (N_34289,N_24814,N_24123);
nor U34290 (N_34290,N_25240,N_27237);
or U34291 (N_34291,N_25405,N_22800);
or U34292 (N_34292,N_21818,N_20392);
and U34293 (N_34293,N_22982,N_23268);
xnor U34294 (N_34294,N_25640,N_21108);
nand U34295 (N_34295,N_26558,N_21919);
nand U34296 (N_34296,N_25286,N_20592);
nand U34297 (N_34297,N_29031,N_25961);
nor U34298 (N_34298,N_21187,N_27972);
nor U34299 (N_34299,N_26875,N_22965);
xor U34300 (N_34300,N_20799,N_28008);
or U34301 (N_34301,N_29329,N_25120);
or U34302 (N_34302,N_27929,N_29708);
xnor U34303 (N_34303,N_21078,N_28322);
and U34304 (N_34304,N_22471,N_22069);
nand U34305 (N_34305,N_29931,N_23285);
nor U34306 (N_34306,N_22951,N_27634);
or U34307 (N_34307,N_27560,N_21709);
or U34308 (N_34308,N_27955,N_27565);
or U34309 (N_34309,N_27343,N_22647);
nor U34310 (N_34310,N_28747,N_20064);
nand U34311 (N_34311,N_23955,N_28179);
and U34312 (N_34312,N_21132,N_29689);
and U34313 (N_34313,N_21348,N_22882);
and U34314 (N_34314,N_27553,N_23812);
and U34315 (N_34315,N_26120,N_26839);
nand U34316 (N_34316,N_29701,N_27010);
or U34317 (N_34317,N_21751,N_23536);
nor U34318 (N_34318,N_25157,N_25066);
or U34319 (N_34319,N_26181,N_26985);
nor U34320 (N_34320,N_27957,N_27826);
nor U34321 (N_34321,N_22293,N_24300);
or U34322 (N_34322,N_21124,N_28833);
and U34323 (N_34323,N_22108,N_27071);
or U34324 (N_34324,N_22281,N_22300);
and U34325 (N_34325,N_28890,N_28537);
nor U34326 (N_34326,N_25087,N_23720);
and U34327 (N_34327,N_29075,N_24015);
nor U34328 (N_34328,N_27107,N_21559);
nand U34329 (N_34329,N_25955,N_24002);
xor U34330 (N_34330,N_27527,N_27632);
nand U34331 (N_34331,N_23728,N_26061);
and U34332 (N_34332,N_24214,N_21093);
nand U34333 (N_34333,N_25119,N_29960);
and U34334 (N_34334,N_23008,N_26866);
xnor U34335 (N_34335,N_26072,N_26239);
or U34336 (N_34336,N_21597,N_25772);
and U34337 (N_34337,N_27846,N_25897);
or U34338 (N_34338,N_21304,N_23191);
or U34339 (N_34339,N_28514,N_20433);
nor U34340 (N_34340,N_24949,N_27065);
nand U34341 (N_34341,N_24152,N_28623);
or U34342 (N_34342,N_26322,N_21456);
xor U34343 (N_34343,N_23270,N_20827);
or U34344 (N_34344,N_20367,N_20794);
nand U34345 (N_34345,N_27509,N_23924);
and U34346 (N_34346,N_23486,N_27313);
nor U34347 (N_34347,N_27079,N_29762);
nand U34348 (N_34348,N_26997,N_21282);
nor U34349 (N_34349,N_22925,N_25069);
and U34350 (N_34350,N_26721,N_23327);
or U34351 (N_34351,N_26009,N_24936);
xnor U34352 (N_34352,N_21609,N_25639);
and U34353 (N_34353,N_20031,N_25695);
and U34354 (N_34354,N_20742,N_20413);
and U34355 (N_34355,N_29268,N_22481);
nor U34356 (N_34356,N_27512,N_27271);
xnor U34357 (N_34357,N_29369,N_23422);
nor U34358 (N_34358,N_25661,N_20913);
nor U34359 (N_34359,N_20048,N_21853);
and U34360 (N_34360,N_21331,N_24055);
nand U34361 (N_34361,N_28077,N_20282);
nand U34362 (N_34362,N_23886,N_23197);
nand U34363 (N_34363,N_25941,N_24131);
nand U34364 (N_34364,N_24007,N_29176);
and U34365 (N_34365,N_29890,N_21126);
nor U34366 (N_34366,N_23676,N_24511);
and U34367 (N_34367,N_24469,N_23645);
or U34368 (N_34368,N_28474,N_21646);
and U34369 (N_34369,N_22538,N_24124);
and U34370 (N_34370,N_22708,N_24642);
and U34371 (N_34371,N_29368,N_27495);
nor U34372 (N_34372,N_27739,N_24653);
nor U34373 (N_34373,N_23147,N_27659);
nand U34374 (N_34374,N_29303,N_23303);
xor U34375 (N_34375,N_26436,N_20551);
or U34376 (N_34376,N_23228,N_24784);
and U34377 (N_34377,N_21648,N_20753);
nor U34378 (N_34378,N_28033,N_23796);
or U34379 (N_34379,N_26619,N_22036);
nand U34380 (N_34380,N_29401,N_23825);
and U34381 (N_34381,N_23813,N_21742);
or U34382 (N_34382,N_26945,N_20584);
xnor U34383 (N_34383,N_24859,N_23027);
nor U34384 (N_34384,N_20018,N_24426);
and U34385 (N_34385,N_25784,N_29286);
and U34386 (N_34386,N_29067,N_24010);
nor U34387 (N_34387,N_20661,N_29679);
nor U34388 (N_34388,N_25819,N_21791);
nand U34389 (N_34389,N_25573,N_29658);
xor U34390 (N_34390,N_24399,N_21667);
nand U34391 (N_34391,N_21691,N_27428);
nor U34392 (N_34392,N_26520,N_22459);
or U34393 (N_34393,N_27572,N_20530);
nor U34394 (N_34394,N_29776,N_22719);
xor U34395 (N_34395,N_29071,N_22743);
or U34396 (N_34396,N_26511,N_24905);
and U34397 (N_34397,N_28543,N_23534);
or U34398 (N_34398,N_26971,N_24979);
and U34399 (N_34399,N_20074,N_21350);
nor U34400 (N_34400,N_21289,N_22994);
and U34401 (N_34401,N_29747,N_25606);
nor U34402 (N_34402,N_20455,N_23194);
or U34403 (N_34403,N_22566,N_20380);
and U34404 (N_34404,N_26083,N_28027);
xor U34405 (N_34405,N_21103,N_28064);
nand U34406 (N_34406,N_28595,N_29134);
nor U34407 (N_34407,N_22769,N_22127);
nor U34408 (N_34408,N_23372,N_29456);
and U34409 (N_34409,N_29659,N_21438);
nor U34410 (N_34410,N_22627,N_25203);
and U34411 (N_34411,N_29035,N_29706);
or U34412 (N_34412,N_21592,N_24251);
xnor U34413 (N_34413,N_20395,N_20583);
nand U34414 (N_34414,N_24319,N_26343);
nor U34415 (N_34415,N_27477,N_27006);
or U34416 (N_34416,N_28062,N_20476);
nor U34417 (N_34417,N_26014,N_27814);
and U34418 (N_34418,N_21569,N_22371);
or U34419 (N_34419,N_25796,N_29669);
or U34420 (N_34420,N_22764,N_27892);
or U34421 (N_34421,N_23082,N_27346);
xnor U34422 (N_34422,N_23450,N_20418);
or U34423 (N_34423,N_22048,N_27449);
nor U34424 (N_34424,N_29855,N_23302);
xor U34425 (N_34425,N_27833,N_25398);
nand U34426 (N_34426,N_29615,N_25090);
or U34427 (N_34427,N_23110,N_25088);
xor U34428 (N_34428,N_24267,N_26308);
xnor U34429 (N_34429,N_20695,N_22406);
and U34430 (N_34430,N_27473,N_25880);
and U34431 (N_34431,N_27393,N_24280);
and U34432 (N_34432,N_21009,N_26728);
and U34433 (N_34433,N_25971,N_23731);
and U34434 (N_34434,N_29914,N_28090);
nor U34435 (N_34435,N_23096,N_28560);
nor U34436 (N_34436,N_26559,N_24296);
or U34437 (N_34437,N_20948,N_23829);
or U34438 (N_34438,N_23721,N_23579);
or U34439 (N_34439,N_26291,N_28483);
or U34440 (N_34440,N_25112,N_28982);
or U34441 (N_34441,N_24752,N_26306);
nand U34442 (N_34442,N_25795,N_23024);
nand U34443 (N_34443,N_26684,N_26244);
nand U34444 (N_34444,N_21544,N_25981);
or U34445 (N_34445,N_25446,N_28510);
or U34446 (N_34446,N_27160,N_26877);
nand U34447 (N_34447,N_25013,N_20397);
xnor U34448 (N_34448,N_24293,N_28681);
and U34449 (N_34449,N_25558,N_26026);
nand U34450 (N_34450,N_21181,N_20679);
or U34451 (N_34451,N_27073,N_20285);
and U34452 (N_34452,N_22044,N_25929);
or U34453 (N_34453,N_26937,N_21847);
xor U34454 (N_34454,N_23014,N_27578);
or U34455 (N_34455,N_23438,N_26360);
and U34456 (N_34456,N_20630,N_27371);
nor U34457 (N_34457,N_20133,N_27859);
nand U34458 (N_34458,N_23093,N_28601);
nor U34459 (N_34459,N_23333,N_20408);
or U34460 (N_34460,N_22650,N_27376);
nor U34461 (N_34461,N_23418,N_28369);
nand U34462 (N_34462,N_21502,N_24425);
or U34463 (N_34463,N_28500,N_22184);
nand U34464 (N_34464,N_28152,N_20329);
nor U34465 (N_34465,N_21517,N_28691);
nand U34466 (N_34466,N_22425,N_26638);
and U34467 (N_34467,N_21761,N_26157);
or U34468 (N_34468,N_25035,N_25887);
nand U34469 (N_34469,N_27295,N_21283);
nand U34470 (N_34470,N_29346,N_28794);
nor U34471 (N_34471,N_21434,N_29015);
nor U34472 (N_34472,N_21953,N_27629);
and U34473 (N_34473,N_23266,N_27093);
or U34474 (N_34474,N_29550,N_28168);
or U34475 (N_34475,N_21485,N_29254);
and U34476 (N_34476,N_29910,N_22865);
and U34477 (N_34477,N_20998,N_26824);
or U34478 (N_34478,N_27559,N_21693);
or U34479 (N_34479,N_26767,N_23010);
nand U34480 (N_34480,N_24480,N_23245);
nor U34481 (N_34481,N_26521,N_28134);
xor U34482 (N_34482,N_27804,N_25027);
xor U34483 (N_34483,N_27799,N_26344);
xnor U34484 (N_34484,N_27555,N_20862);
nor U34485 (N_34485,N_26524,N_28970);
nor U34486 (N_34486,N_29276,N_27829);
and U34487 (N_34487,N_23415,N_29144);
and U34488 (N_34488,N_23388,N_21952);
nand U34489 (N_34489,N_21890,N_23654);
nand U34490 (N_34490,N_23433,N_29622);
or U34491 (N_34491,N_22174,N_20252);
or U34492 (N_34492,N_21156,N_27850);
xor U34493 (N_34493,N_29605,N_25512);
and U34494 (N_34494,N_26745,N_29155);
and U34495 (N_34495,N_24516,N_23693);
xor U34496 (N_34496,N_24962,N_27996);
or U34497 (N_34497,N_22995,N_26364);
and U34498 (N_34498,N_22729,N_24210);
or U34499 (N_34499,N_21949,N_27622);
and U34500 (N_34500,N_26037,N_21440);
xnor U34501 (N_34501,N_29213,N_23673);
xor U34502 (N_34502,N_27219,N_28232);
nand U34503 (N_34503,N_29512,N_20167);
or U34504 (N_34504,N_25612,N_29929);
nor U34505 (N_34505,N_25002,N_29118);
and U34506 (N_34506,N_29283,N_28141);
xor U34507 (N_34507,N_29790,N_29526);
and U34508 (N_34508,N_29250,N_23306);
and U34509 (N_34509,N_25516,N_28835);
nand U34510 (N_34510,N_23062,N_26171);
and U34511 (N_34511,N_22320,N_23173);
and U34512 (N_34512,N_24388,N_24849);
or U34513 (N_34513,N_22671,N_28915);
or U34514 (N_34514,N_29773,N_26325);
or U34515 (N_34515,N_27537,N_20386);
nand U34516 (N_34516,N_27051,N_28557);
nand U34517 (N_34517,N_26247,N_29349);
nand U34518 (N_34518,N_27480,N_25469);
or U34519 (N_34519,N_23797,N_23788);
nor U34520 (N_34520,N_20713,N_29180);
and U34521 (N_34521,N_29504,N_25419);
and U34522 (N_34522,N_26546,N_27728);
and U34523 (N_34523,N_21079,N_28788);
and U34524 (N_34524,N_22781,N_24640);
nor U34525 (N_34525,N_23115,N_26482);
nor U34526 (N_34526,N_28620,N_27300);
nand U34527 (N_34527,N_25564,N_22107);
nand U34528 (N_34528,N_21024,N_27317);
nand U34529 (N_34529,N_29529,N_22393);
and U34530 (N_34530,N_25448,N_29188);
nand U34531 (N_34531,N_20424,N_23722);
nor U34532 (N_34532,N_27443,N_26885);
nor U34533 (N_34533,N_28012,N_21175);
nand U34534 (N_34534,N_20924,N_20659);
and U34535 (N_34535,N_24782,N_21747);
or U34536 (N_34536,N_27748,N_29861);
or U34537 (N_34537,N_22807,N_27790);
or U34538 (N_34538,N_26792,N_29020);
or U34539 (N_34539,N_21070,N_24727);
or U34540 (N_34540,N_27287,N_24957);
nor U34541 (N_34541,N_22121,N_21694);
and U34542 (N_34542,N_27025,N_22984);
nand U34543 (N_34543,N_27286,N_24860);
and U34544 (N_34544,N_27381,N_26225);
and U34545 (N_34545,N_21521,N_24204);
nand U34546 (N_34546,N_24867,N_29720);
or U34547 (N_34547,N_22843,N_25990);
and U34548 (N_34548,N_20868,N_24919);
and U34549 (N_34549,N_22718,N_21193);
nor U34550 (N_34550,N_24732,N_21248);
nand U34551 (N_34551,N_24586,N_29643);
xor U34552 (N_34552,N_29289,N_28399);
and U34553 (N_34553,N_26753,N_24987);
and U34554 (N_34554,N_25395,N_23996);
nor U34555 (N_34555,N_23200,N_25848);
or U34556 (N_34556,N_27307,N_29751);
or U34557 (N_34557,N_22460,N_24676);
and U34558 (N_34558,N_20893,N_20175);
nand U34559 (N_34559,N_25862,N_24090);
or U34560 (N_34560,N_20930,N_26358);
nand U34561 (N_34561,N_27765,N_29056);
nand U34562 (N_34562,N_24333,N_24311);
nand U34563 (N_34563,N_23368,N_21039);
nand U34564 (N_34564,N_22742,N_27970);
nor U34565 (N_34565,N_22798,N_21683);
xnor U34566 (N_34566,N_22060,N_21858);
xor U34567 (N_34567,N_29667,N_20466);
nand U34568 (N_34568,N_21807,N_20436);
and U34569 (N_34569,N_21996,N_21478);
nor U34570 (N_34570,N_22490,N_29408);
and U34571 (N_34571,N_23764,N_22359);
nand U34572 (N_34572,N_23769,N_23834);
nor U34573 (N_34573,N_21326,N_27483);
xor U34574 (N_34574,N_29759,N_28455);
nor U34575 (N_34575,N_20508,N_27925);
and U34576 (N_34576,N_27899,N_27693);
nor U34577 (N_34577,N_24137,N_23318);
nor U34578 (N_34578,N_25599,N_21998);
nand U34579 (N_34579,N_25506,N_29728);
nand U34580 (N_34580,N_26924,N_24971);
or U34581 (N_34581,N_23575,N_20456);
and U34582 (N_34582,N_26080,N_21449);
and U34583 (N_34583,N_29705,N_21145);
and U34584 (N_34584,N_20310,N_21636);
or U34585 (N_34585,N_27930,N_29699);
or U34586 (N_34586,N_22900,N_25332);
nand U34587 (N_34587,N_27910,N_22619);
and U34588 (N_34588,N_29252,N_21909);
nand U34589 (N_34589,N_29544,N_21413);
or U34590 (N_34590,N_27905,N_28154);
nand U34591 (N_34591,N_27070,N_28709);
xnor U34592 (N_34592,N_28059,N_28240);
xor U34593 (N_34593,N_23038,N_24728);
nor U34594 (N_34594,N_26449,N_27352);
nand U34595 (N_34595,N_23084,N_25021);
and U34596 (N_34596,N_25205,N_24944);
nor U34597 (N_34597,N_26206,N_23371);
and U34598 (N_34598,N_28753,N_24902);
nand U34599 (N_34599,N_21353,N_23077);
nand U34600 (N_34600,N_22149,N_22247);
xor U34601 (N_34601,N_25583,N_21978);
or U34602 (N_34602,N_25104,N_21647);
and U34603 (N_34603,N_27068,N_24893);
or U34604 (N_34604,N_25774,N_21540);
or U34605 (N_34605,N_26283,N_24627);
xnor U34606 (N_34606,N_28670,N_25054);
xor U34607 (N_34607,N_24639,N_27953);
nor U34608 (N_34608,N_27684,N_24705);
nor U34609 (N_34609,N_29717,N_25927);
nor U34610 (N_34610,N_25391,N_27862);
or U34611 (N_34611,N_29710,N_27818);
nor U34612 (N_34612,N_26550,N_28974);
or U34613 (N_34613,N_28071,N_29281);
or U34614 (N_34614,N_20014,N_25723);
nor U34615 (N_34615,N_20467,N_27805);
and U34616 (N_34616,N_26062,N_23963);
nor U34617 (N_34617,N_27205,N_24371);
or U34618 (N_34618,N_23663,N_24620);
xor U34619 (N_34619,N_23058,N_27001);
and U34620 (N_34620,N_22269,N_21922);
or U34621 (N_34621,N_27676,N_20650);
or U34622 (N_34622,N_29240,N_23604);
nor U34623 (N_34623,N_20333,N_26235);
and U34624 (N_34624,N_23683,N_23758);
nor U34625 (N_34625,N_23152,N_25296);
xnor U34626 (N_34626,N_22539,N_29571);
nor U34627 (N_34627,N_21484,N_29540);
or U34628 (N_34628,N_23265,N_26576);
nor U34629 (N_34629,N_28821,N_28427);
or U34630 (N_34630,N_21562,N_24099);
or U34631 (N_34631,N_23293,N_29796);
or U34632 (N_34632,N_23491,N_26329);
or U34633 (N_34633,N_26194,N_27045);
nor U34634 (N_34634,N_23523,N_27520);
nand U34635 (N_34635,N_21318,N_25256);
nor U34636 (N_34636,N_27324,N_22973);
nand U34637 (N_34637,N_20236,N_29338);
and U34638 (N_34638,N_22754,N_25399);
nand U34639 (N_34639,N_21516,N_26500);
nor U34640 (N_34640,N_27708,N_29897);
nor U34641 (N_34641,N_22063,N_28988);
nand U34642 (N_34642,N_25489,N_28287);
nand U34643 (N_34643,N_27890,N_22702);
and U34644 (N_34644,N_27789,N_28935);
or U34645 (N_34645,N_22632,N_21071);
nand U34646 (N_34646,N_24537,N_28963);
xor U34647 (N_34647,N_21112,N_26569);
or U34648 (N_34648,N_26754,N_24947);
xnor U34649 (N_34649,N_23949,N_24633);
and U34650 (N_34650,N_28424,N_25536);
and U34651 (N_34651,N_26779,N_29386);
and U34652 (N_34652,N_24904,N_21224);
nand U34653 (N_34653,N_29585,N_29830);
nand U34654 (N_34654,N_25492,N_23153);
or U34655 (N_34655,N_27861,N_28678);
or U34656 (N_34656,N_25966,N_23511);
and U34657 (N_34657,N_20977,N_24507);
nand U34658 (N_34658,N_26941,N_27029);
or U34659 (N_34659,N_27928,N_28640);
nor U34660 (N_34660,N_29095,N_26747);
or U34661 (N_34661,N_24287,N_29665);
nor U34662 (N_34662,N_27522,N_25824);
nand U34663 (N_34663,N_26260,N_26714);
nand U34664 (N_34664,N_21541,N_24291);
and U34665 (N_34665,N_22505,N_25979);
nor U34666 (N_34666,N_29866,N_23040);
nor U34667 (N_34667,N_24840,N_21470);
nor U34668 (N_34668,N_20962,N_28307);
and U34669 (N_34669,N_29044,N_22980);
nand U34670 (N_34670,N_23537,N_27054);
nand U34671 (N_34671,N_29455,N_21498);
nor U34672 (N_34672,N_20531,N_29606);
nor U34673 (N_34673,N_26444,N_28298);
nand U34674 (N_34674,N_28251,N_28652);
and U34675 (N_34675,N_26536,N_21821);
nor U34676 (N_34676,N_26719,N_22654);
nand U34677 (N_34677,N_23921,N_20663);
nor U34678 (N_34678,N_22540,N_28837);
nand U34679 (N_34679,N_23233,N_27155);
nor U34680 (N_34680,N_23684,N_25543);
xnor U34681 (N_34681,N_24119,N_22751);
nor U34682 (N_34682,N_29026,N_29218);
and U34683 (N_34683,N_21653,N_29547);
nand U34684 (N_34684,N_28535,N_20911);
nor U34685 (N_34685,N_21675,N_20484);
nor U34686 (N_34686,N_26484,N_29711);
xor U34687 (N_34687,N_28330,N_24078);
nor U34688 (N_34688,N_28293,N_29883);
xnor U34689 (N_34689,N_29867,N_22845);
nand U34690 (N_34690,N_26538,N_20398);
nor U34691 (N_34691,N_21911,N_27159);
nand U34692 (N_34692,N_27415,N_21338);
nor U34693 (N_34693,N_25153,N_21387);
nor U34694 (N_34694,N_25711,N_29838);
nand U34695 (N_34695,N_29871,N_23916);
or U34696 (N_34696,N_21243,N_28888);
or U34697 (N_34697,N_26089,N_20944);
or U34698 (N_34698,N_24577,N_25657);
nor U34699 (N_34699,N_27920,N_24886);
or U34700 (N_34700,N_27854,N_21968);
and U34701 (N_34701,N_27660,N_26063);
and U34702 (N_34702,N_25262,N_21490);
nor U34703 (N_34703,N_25991,N_27534);
nor U34704 (N_34704,N_23747,N_24661);
or U34705 (N_34705,N_29320,N_28376);
nor U34706 (N_34706,N_27387,N_28618);
or U34707 (N_34707,N_27362,N_23807);
xnor U34708 (N_34708,N_21940,N_20469);
or U34709 (N_34709,N_26390,N_21013);
and U34710 (N_34710,N_29500,N_20490);
and U34711 (N_34711,N_26648,N_29039);
or U34712 (N_34712,N_29727,N_25786);
and U34713 (N_34713,N_29440,N_24260);
and U34714 (N_34714,N_26183,N_25942);
or U34715 (N_34715,N_20311,N_20475);
or U34716 (N_34716,N_20693,N_25814);
and U34717 (N_34717,N_25029,N_25279);
nor U34718 (N_34718,N_23229,N_28389);
or U34719 (N_34719,N_22697,N_24094);
and U34720 (N_34720,N_26962,N_29517);
and U34721 (N_34721,N_27538,N_21574);
or U34722 (N_34722,N_25665,N_25797);
nand U34723 (N_34723,N_23705,N_20432);
nor U34724 (N_34724,N_20447,N_22442);
and U34725 (N_34725,N_29926,N_21806);
or U34726 (N_34726,N_23798,N_25876);
nand U34727 (N_34727,N_25953,N_26132);
and U34728 (N_34728,N_27585,N_25945);
nor U34729 (N_34729,N_26658,N_26891);
nand U34730 (N_34730,N_28371,N_25046);
or U34731 (N_34731,N_20833,N_25754);
and U34732 (N_34732,N_20873,N_23029);
nor U34733 (N_34733,N_20400,N_21406);
nand U34734 (N_34734,N_20815,N_20058);
or U34735 (N_34735,N_20853,N_22605);
and U34736 (N_34736,N_28791,N_26805);
nand U34737 (N_34737,N_25830,N_21411);
or U34738 (N_34738,N_22423,N_22926);
nand U34739 (N_34739,N_22483,N_29800);
nor U34740 (N_34740,N_28846,N_28813);
or U34741 (N_34741,N_26270,N_27808);
nor U34742 (N_34742,N_24847,N_22879);
and U34743 (N_34743,N_27197,N_20183);
and U34744 (N_34744,N_24006,N_29120);
and U34745 (N_34745,N_20945,N_20415);
nand U34746 (N_34746,N_26543,N_29450);
nor U34747 (N_34747,N_23064,N_25940);
and U34748 (N_34748,N_22167,N_25230);
nand U34749 (N_34749,N_25633,N_27649);
and U34750 (N_34750,N_26246,N_29661);
nand U34751 (N_34751,N_21280,N_28022);
nor U34752 (N_34752,N_24257,N_24574);
and U34753 (N_34753,N_22553,N_24694);
and U34754 (N_34754,N_29196,N_22806);
and U34755 (N_34755,N_21347,N_26528);
or U34756 (N_34756,N_24991,N_27056);
and U34757 (N_34757,N_28671,N_27018);
nand U34758 (N_34758,N_23399,N_25867);
nand U34759 (N_34759,N_28824,N_20338);
nor U34760 (N_34760,N_24434,N_28255);
and U34761 (N_34761,N_29049,N_25718);
and U34762 (N_34762,N_21215,N_22852);
nor U34763 (N_34763,N_27398,N_28945);
nand U34764 (N_34764,N_26303,N_22497);
nor U34765 (N_34765,N_26376,N_28291);
and U34766 (N_34766,N_20978,N_29200);
nor U34767 (N_34767,N_20401,N_28391);
nand U34768 (N_34768,N_29893,N_23530);
and U34769 (N_34769,N_29109,N_24086);
xnor U34770 (N_34770,N_24363,N_24454);
or U34771 (N_34771,N_26372,N_26633);
xor U34772 (N_34772,N_23965,N_24444);
and U34773 (N_34773,N_21185,N_23053);
xor U34774 (N_34774,N_25628,N_23786);
xnor U34775 (N_34775,N_28318,N_24759);
nor U34776 (N_34776,N_24215,N_24544);
or U34777 (N_34777,N_28180,N_24146);
or U34778 (N_34778,N_29360,N_27545);
nor U34779 (N_34779,N_24269,N_28869);
or U34780 (N_34780,N_24504,N_25209);
nor U34781 (N_34781,N_26432,N_27467);
xnor U34782 (N_34782,N_20654,N_24455);
nand U34783 (N_34783,N_26321,N_26897);
nand U34784 (N_34784,N_23234,N_20396);
nor U34785 (N_34785,N_28432,N_29745);
nor U34786 (N_34786,N_23831,N_23898);
and U34787 (N_34787,N_23889,N_25062);
nand U34788 (N_34788,N_27434,N_23021);
and U34789 (N_34789,N_22131,N_21887);
and U34790 (N_34790,N_24234,N_28973);
or U34791 (N_34791,N_22949,N_20865);
nand U34792 (N_34792,N_21986,N_25836);
xnor U34793 (N_34793,N_29811,N_28600);
and U34794 (N_34794,N_25055,N_25326);
or U34795 (N_34795,N_22077,N_29692);
or U34796 (N_34796,N_24529,N_21476);
nor U34797 (N_34797,N_25716,N_24903);
xor U34798 (N_34798,N_25101,N_23736);
and U34799 (N_34799,N_25834,N_20817);
nor U34800 (N_34800,N_25587,N_22579);
or U34801 (N_34801,N_20760,N_26264);
and U34802 (N_34802,N_23931,N_20164);
and U34803 (N_34803,N_27466,N_25780);
and U34804 (N_34804,N_28504,N_25089);
nor U34805 (N_34805,N_29249,N_27590);
nor U34806 (N_34806,N_24064,N_28830);
nand U34807 (N_34807,N_23837,N_23571);
or U34808 (N_34808,N_20153,N_24928);
nor U34809 (N_34809,N_28360,N_21871);
nand U34810 (N_34810,N_28290,N_25224);
nand U34811 (N_34811,N_28140,N_21844);
nor U34812 (N_34812,N_22946,N_28766);
nand U34813 (N_34813,N_21505,N_28245);
xnor U34814 (N_34814,N_24376,N_23185);
nor U34815 (N_34815,N_26663,N_24194);
nor U34816 (N_34816,N_24044,N_22052);
xnor U34817 (N_34817,N_25259,N_22685);
and U34818 (N_34818,N_25804,N_27642);
or U34819 (N_34819,N_21267,N_21266);
and U34820 (N_34820,N_26070,N_27823);
nand U34821 (N_34821,N_27016,N_24828);
and U34822 (N_34822,N_27741,N_27497);
nor U34823 (N_34823,N_23560,N_27179);
or U34824 (N_34824,N_23846,N_24781);
nand U34825 (N_34825,N_25615,N_26893);
and U34826 (N_34826,N_20249,N_25861);
nand U34827 (N_34827,N_25033,N_25632);
or U34828 (N_34828,N_25159,N_25883);
xnor U34829 (N_34829,N_21837,N_21017);
and U34830 (N_34830,N_25346,N_28536);
or U34831 (N_34831,N_22527,N_28511);
nand U34832 (N_34832,N_20902,N_24126);
or U34833 (N_34833,N_22035,N_24151);
and U34834 (N_34834,N_24326,N_27806);
or U34835 (N_34835,N_24367,N_20052);
nand U34836 (N_34836,N_26373,N_29476);
and U34837 (N_34837,N_24199,N_26818);
and U34838 (N_34838,N_29671,N_26233);
nand U34839 (N_34839,N_29515,N_22311);
or U34840 (N_34840,N_29806,N_24670);
nor U34841 (N_34841,N_26255,N_20774);
and U34842 (N_34842,N_25048,N_22152);
and U34843 (N_34843,N_22846,N_24719);
and U34844 (N_34844,N_29452,N_26015);
or U34845 (N_34845,N_22271,N_27118);
and U34846 (N_34846,N_27035,N_23800);
nand U34847 (N_34847,N_22286,N_20658);
or U34848 (N_34848,N_20305,N_25794);
xor U34849 (N_34849,N_27772,N_23958);
or U34850 (N_34850,N_27291,N_24992);
and U34851 (N_34851,N_26413,N_27759);
nand U34852 (N_34852,N_21002,N_29244);
nand U34853 (N_34853,N_25859,N_26769);
and U34854 (N_34854,N_29115,N_26045);
nand U34855 (N_34855,N_23452,N_28992);
or U34856 (N_34856,N_24564,N_21980);
nor U34857 (N_34857,N_27498,N_27887);
nand U34858 (N_34858,N_25500,N_23239);
and U34859 (N_34859,N_21080,N_23620);
and U34860 (N_34860,N_20594,N_24366);
or U34861 (N_34861,N_29714,N_24629);
and U34862 (N_34862,N_22494,N_21701);
or U34863 (N_34863,N_25850,N_29185);
nand U34864 (N_34864,N_25554,N_27149);
nand U34865 (N_34865,N_29704,N_25749);
nor U34866 (N_34866,N_23503,N_28985);
nor U34867 (N_34867,N_20451,N_27236);
and U34868 (N_34868,N_20127,N_21927);
or U34869 (N_34869,N_27906,N_29084);
nand U34870 (N_34870,N_26856,N_29674);
xnor U34871 (N_34871,N_24035,N_22570);
nor U34872 (N_34872,N_23207,N_25878);
nand U34873 (N_34873,N_22594,N_23159);
or U34874 (N_34874,N_26789,N_28884);
xor U34875 (N_34875,N_26245,N_24631);
nand U34876 (N_34876,N_23240,N_20221);
nor U34877 (N_34877,N_25302,N_21950);
or U34878 (N_34878,N_29331,N_23904);
xor U34879 (N_34879,N_27738,N_24978);
nand U34880 (N_34880,N_23072,N_27734);
nand U34881 (N_34881,N_25871,N_27985);
nor U34882 (N_34882,N_22559,N_26383);
nor U34883 (N_34883,N_24958,N_23375);
nor U34884 (N_34884,N_25175,N_27773);
xnor U34885 (N_34885,N_25208,N_22289);
nor U34886 (N_34886,N_20951,N_22084);
or U34887 (N_34887,N_22360,N_28771);
nand U34888 (N_34888,N_21464,N_25757);
nor U34889 (N_34889,N_26415,N_21528);
and U34890 (N_34890,N_21583,N_21462);
and U34891 (N_34891,N_20297,N_21419);
xnor U34892 (N_34892,N_29655,N_27914);
or U34893 (N_34893,N_27474,N_20162);
nor U34894 (N_34894,N_29884,N_22290);
xor U34895 (N_34895,N_21385,N_20422);
and U34896 (N_34896,N_25481,N_24149);
nand U34897 (N_34897,N_21513,N_24114);
nor U34898 (N_34898,N_27214,N_22208);
and U34899 (N_34899,N_23742,N_24022);
and U34900 (N_34900,N_25248,N_22840);
nor U34901 (N_34901,N_21781,N_26667);
and U34902 (N_34902,N_22944,N_27515);
nand U34903 (N_34903,N_20318,N_26594);
or U34904 (N_34904,N_21313,N_22765);
nor U34905 (N_34905,N_24686,N_25828);
nor U34906 (N_34906,N_28224,N_29411);
nand U34907 (N_34907,N_21225,N_27022);
and U34908 (N_34908,N_29607,N_26033);
nand U34909 (N_34909,N_27268,N_24250);
or U34910 (N_34910,N_26126,N_20647);
or U34911 (N_34911,N_23666,N_25832);
and U34912 (N_34912,N_24887,N_25299);
nor U34913 (N_34913,N_29465,N_24754);
and U34914 (N_34914,N_26552,N_21713);
and U34915 (N_34915,N_21275,N_23535);
or U34916 (N_34916,N_23459,N_22562);
nand U34917 (N_34917,N_22145,N_20076);
nor U34918 (N_34918,N_26835,N_24796);
nor U34919 (N_34919,N_28698,N_20628);
or U34920 (N_34920,N_25370,N_23241);
and U34921 (N_34921,N_23482,N_25811);
nor U34922 (N_34922,N_29998,N_23730);
or U34923 (N_34923,N_25154,N_27978);
nand U34924 (N_34924,N_20218,N_27633);
xor U34925 (N_34925,N_24053,N_23120);
or U34926 (N_34926,N_23750,N_29198);
nand U34927 (N_34927,N_24803,N_26904);
nand U34928 (N_34928,N_25537,N_28067);
nand U34929 (N_34929,N_28315,N_25056);
and U34930 (N_34930,N_22560,N_28153);
nand U34931 (N_34931,N_22352,N_25305);
or U34932 (N_34932,N_20161,N_20984);
and U34933 (N_34933,N_29438,N_24973);
nand U34934 (N_34934,N_20341,N_24684);
nor U34935 (N_34935,N_26972,N_25803);
nand U34936 (N_34936,N_20295,N_27394);
nand U34937 (N_34937,N_29935,N_28613);
nor U34938 (N_34938,N_22420,N_24174);
nand U34939 (N_34939,N_22370,N_27679);
nor U34940 (N_34940,N_23502,N_25899);
nand U34941 (N_34941,N_28564,N_24756);
xor U34942 (N_34942,N_23821,N_26428);
nand U34943 (N_34943,N_29752,N_20927);
nor U34944 (N_34944,N_27732,N_26093);
and U34945 (N_34945,N_22652,N_21446);
or U34946 (N_34946,N_27418,N_22357);
and U34947 (N_34947,N_20563,N_28721);
nor U34948 (N_34948,N_27496,N_26999);
nor U34949 (N_34949,N_26351,N_26516);
or U34950 (N_34950,N_20253,N_20359);
nor U34951 (N_34951,N_20337,N_29358);
nor U34952 (N_34952,N_29531,N_28106);
and U34953 (N_34953,N_22462,N_28532);
or U34954 (N_34954,N_23896,N_20983);
nand U34955 (N_34955,N_21246,N_27442);
nor U34956 (N_34956,N_28651,N_27437);
nor U34957 (N_34957,N_25425,N_20482);
or U34958 (N_34958,N_29923,N_25808);
and U34959 (N_34959,N_24361,N_24056);
nor U34960 (N_34960,N_22803,N_22759);
nand U34961 (N_34961,N_23922,N_20529);
and U34962 (N_34962,N_29924,N_22100);
nand U34963 (N_34963,N_26707,N_24689);
nand U34964 (N_34964,N_22667,N_26098);
and U34965 (N_34965,N_26760,N_23878);
or U34966 (N_34966,N_20045,N_20634);
nand U34967 (N_34967,N_22484,N_25197);
nand U34968 (N_34968,N_20534,N_28246);
nor U34969 (N_34969,N_29223,N_27535);
nor U34970 (N_34970,N_24039,N_23993);
nor U34971 (N_34971,N_24531,N_23005);
or U34972 (N_34972,N_24404,N_24557);
or U34973 (N_34973,N_22979,N_29389);
xor U34974 (N_34974,N_26238,N_26840);
xnor U34975 (N_34975,N_21893,N_26236);
or U34976 (N_34976,N_26951,N_23394);
nor U34977 (N_34977,N_28214,N_20259);
xnor U34978 (N_34978,N_21368,N_27367);
and U34979 (N_34979,N_22631,N_21196);
nor U34980 (N_34980,N_26124,N_24990);
nand U34981 (N_34981,N_21758,N_25031);
or U34982 (N_34982,N_22478,N_20727);
nand U34983 (N_34983,N_22302,N_21704);
nand U34984 (N_34984,N_25416,N_24421);
and U34985 (N_34985,N_27786,N_25275);
nor U34986 (N_34986,N_24317,N_24604);
nor U34987 (N_34987,N_22791,N_20716);
or U34988 (N_34988,N_28729,N_20537);
or U34989 (N_34989,N_24277,N_28221);
nor U34990 (N_34990,N_29367,N_22604);
and U34991 (N_34991,N_29427,N_22710);
xor U34992 (N_34992,N_22017,N_20707);
nand U34993 (N_34993,N_24499,N_22683);
or U34994 (N_34994,N_21069,N_27499);
and U34995 (N_34995,N_21421,N_26001);
or U34996 (N_34996,N_28912,N_27710);
nor U34997 (N_34997,N_25379,N_28489);
xnor U34998 (N_34998,N_21077,N_22850);
xnor U34999 (N_34999,N_27960,N_24047);
or U35000 (N_35000,N_20379,N_25700);
xnor U35001 (N_35001,N_20516,N_21211);
nand U35002 (N_35002,N_25488,N_21439);
nand U35003 (N_35003,N_20723,N_28162);
nand U35004 (N_35004,N_21458,N_20614);
and U35005 (N_35005,N_29272,N_21873);
or U35006 (N_35006,N_27875,N_24765);
or U35007 (N_35007,N_25832,N_29319);
or U35008 (N_35008,N_24012,N_22236);
and U35009 (N_35009,N_23079,N_20731);
xor U35010 (N_35010,N_27397,N_25151);
or U35011 (N_35011,N_26327,N_24539);
nor U35012 (N_35012,N_28734,N_26658);
nor U35013 (N_35013,N_27133,N_28542);
and U35014 (N_35014,N_20947,N_21601);
nor U35015 (N_35015,N_29725,N_28329);
nor U35016 (N_35016,N_22197,N_29789);
nor U35017 (N_35017,N_20768,N_21541);
xnor U35018 (N_35018,N_28058,N_21307);
and U35019 (N_35019,N_24694,N_22890);
or U35020 (N_35020,N_26309,N_26055);
and U35021 (N_35021,N_29145,N_23526);
or U35022 (N_35022,N_20424,N_20332);
nor U35023 (N_35023,N_25612,N_22541);
and U35024 (N_35024,N_27555,N_21033);
or U35025 (N_35025,N_22344,N_24679);
or U35026 (N_35026,N_23692,N_21123);
xor U35027 (N_35027,N_29787,N_28433);
and U35028 (N_35028,N_29783,N_20251);
xor U35029 (N_35029,N_22107,N_27781);
and U35030 (N_35030,N_26573,N_23874);
or U35031 (N_35031,N_21399,N_22767);
nor U35032 (N_35032,N_21342,N_27929);
nand U35033 (N_35033,N_22998,N_25263);
or U35034 (N_35034,N_25547,N_23126);
or U35035 (N_35035,N_20080,N_21187);
nor U35036 (N_35036,N_24985,N_22075);
xnor U35037 (N_35037,N_23218,N_29945);
nor U35038 (N_35038,N_20151,N_22297);
and U35039 (N_35039,N_27642,N_22382);
and U35040 (N_35040,N_24314,N_22608);
or U35041 (N_35041,N_28099,N_27880);
nand U35042 (N_35042,N_27973,N_22519);
nand U35043 (N_35043,N_27623,N_29172);
nand U35044 (N_35044,N_26719,N_25697);
nand U35045 (N_35045,N_25406,N_27855);
nor U35046 (N_35046,N_28129,N_27731);
nor U35047 (N_35047,N_24683,N_24856);
and U35048 (N_35048,N_20098,N_27274);
nand U35049 (N_35049,N_24458,N_28963);
and U35050 (N_35050,N_24456,N_28924);
and U35051 (N_35051,N_21573,N_28824);
or U35052 (N_35052,N_26621,N_26533);
nor U35053 (N_35053,N_25206,N_28212);
or U35054 (N_35054,N_28517,N_26350);
nand U35055 (N_35055,N_24004,N_20140);
and U35056 (N_35056,N_24222,N_21615);
nor U35057 (N_35057,N_29338,N_21427);
or U35058 (N_35058,N_20894,N_29362);
and U35059 (N_35059,N_20973,N_25767);
or U35060 (N_35060,N_21013,N_22635);
xnor U35061 (N_35061,N_25051,N_23012);
and U35062 (N_35062,N_26881,N_24759);
nand U35063 (N_35063,N_26593,N_27247);
nor U35064 (N_35064,N_23617,N_27484);
and U35065 (N_35065,N_27908,N_24304);
nor U35066 (N_35066,N_29905,N_20171);
or U35067 (N_35067,N_21615,N_25091);
nor U35068 (N_35068,N_23199,N_26298);
xor U35069 (N_35069,N_21029,N_26663);
or U35070 (N_35070,N_29653,N_21721);
and U35071 (N_35071,N_22304,N_29484);
nand U35072 (N_35072,N_27788,N_22968);
nand U35073 (N_35073,N_29682,N_25844);
or U35074 (N_35074,N_20215,N_28446);
nor U35075 (N_35075,N_21002,N_29982);
and U35076 (N_35076,N_28584,N_26084);
and U35077 (N_35077,N_24141,N_20598);
or U35078 (N_35078,N_24217,N_26230);
and U35079 (N_35079,N_28913,N_24082);
nor U35080 (N_35080,N_24123,N_23938);
nor U35081 (N_35081,N_28707,N_21494);
nor U35082 (N_35082,N_29210,N_24580);
nor U35083 (N_35083,N_20567,N_24768);
or U35084 (N_35084,N_28078,N_22197);
nand U35085 (N_35085,N_23330,N_24598);
nand U35086 (N_35086,N_27052,N_29495);
xor U35087 (N_35087,N_25722,N_27943);
nand U35088 (N_35088,N_22289,N_25237);
and U35089 (N_35089,N_20093,N_26346);
or U35090 (N_35090,N_27088,N_29423);
nor U35091 (N_35091,N_25843,N_24203);
nand U35092 (N_35092,N_24219,N_29882);
nor U35093 (N_35093,N_29521,N_29133);
and U35094 (N_35094,N_23348,N_20596);
or U35095 (N_35095,N_24053,N_26958);
or U35096 (N_35096,N_27290,N_27837);
nand U35097 (N_35097,N_25892,N_21261);
and U35098 (N_35098,N_27569,N_26204);
nand U35099 (N_35099,N_26867,N_28594);
and U35100 (N_35100,N_23928,N_29670);
nor U35101 (N_35101,N_25823,N_27236);
and U35102 (N_35102,N_28186,N_26351);
or U35103 (N_35103,N_24678,N_22915);
nand U35104 (N_35104,N_23331,N_26987);
nor U35105 (N_35105,N_24035,N_23878);
or U35106 (N_35106,N_21993,N_25084);
xor U35107 (N_35107,N_26223,N_27355);
and U35108 (N_35108,N_29599,N_23242);
or U35109 (N_35109,N_26392,N_29615);
and U35110 (N_35110,N_20103,N_24527);
xnor U35111 (N_35111,N_21476,N_27543);
xnor U35112 (N_35112,N_29646,N_22963);
or U35113 (N_35113,N_27066,N_26887);
xor U35114 (N_35114,N_22841,N_20318);
nand U35115 (N_35115,N_27747,N_29158);
xnor U35116 (N_35116,N_20778,N_21684);
or U35117 (N_35117,N_28724,N_20618);
nand U35118 (N_35118,N_24620,N_20594);
xnor U35119 (N_35119,N_22539,N_21333);
or U35120 (N_35120,N_21210,N_24527);
nand U35121 (N_35121,N_26430,N_21764);
nand U35122 (N_35122,N_28467,N_20644);
or U35123 (N_35123,N_24987,N_25224);
or U35124 (N_35124,N_27693,N_21221);
nor U35125 (N_35125,N_22154,N_26227);
and U35126 (N_35126,N_24304,N_22249);
nor U35127 (N_35127,N_27817,N_21899);
and U35128 (N_35128,N_23025,N_28206);
and U35129 (N_35129,N_27882,N_24492);
nand U35130 (N_35130,N_22048,N_22226);
and U35131 (N_35131,N_24987,N_20816);
nand U35132 (N_35132,N_22480,N_29374);
or U35133 (N_35133,N_25872,N_22779);
and U35134 (N_35134,N_21583,N_27453);
and U35135 (N_35135,N_25971,N_29381);
and U35136 (N_35136,N_26254,N_29753);
nand U35137 (N_35137,N_29089,N_23370);
nor U35138 (N_35138,N_28739,N_22271);
and U35139 (N_35139,N_26336,N_29187);
nand U35140 (N_35140,N_23242,N_20358);
nor U35141 (N_35141,N_22641,N_24231);
nor U35142 (N_35142,N_29872,N_27298);
nor U35143 (N_35143,N_20136,N_25827);
nand U35144 (N_35144,N_21237,N_27701);
or U35145 (N_35145,N_23971,N_24966);
nor U35146 (N_35146,N_28105,N_25711);
or U35147 (N_35147,N_28320,N_21214);
nand U35148 (N_35148,N_22526,N_21291);
nor U35149 (N_35149,N_25010,N_22193);
and U35150 (N_35150,N_22905,N_27422);
or U35151 (N_35151,N_26037,N_29055);
or U35152 (N_35152,N_22377,N_21441);
and U35153 (N_35153,N_29760,N_20556);
nor U35154 (N_35154,N_24005,N_26589);
xnor U35155 (N_35155,N_26408,N_27670);
xnor U35156 (N_35156,N_25794,N_21067);
nand U35157 (N_35157,N_28456,N_23421);
and U35158 (N_35158,N_20741,N_27376);
or U35159 (N_35159,N_29268,N_25604);
nor U35160 (N_35160,N_29788,N_22389);
and U35161 (N_35161,N_21935,N_27933);
or U35162 (N_35162,N_25854,N_20543);
and U35163 (N_35163,N_27879,N_21700);
nand U35164 (N_35164,N_20007,N_24187);
or U35165 (N_35165,N_27989,N_24955);
xnor U35166 (N_35166,N_24883,N_20393);
nor U35167 (N_35167,N_20435,N_26825);
nand U35168 (N_35168,N_22109,N_28063);
xnor U35169 (N_35169,N_29793,N_24966);
or U35170 (N_35170,N_21874,N_24840);
or U35171 (N_35171,N_28729,N_20034);
or U35172 (N_35172,N_20284,N_24090);
nor U35173 (N_35173,N_24097,N_20853);
xnor U35174 (N_35174,N_22343,N_21099);
and U35175 (N_35175,N_23720,N_24290);
nand U35176 (N_35176,N_29681,N_23417);
or U35177 (N_35177,N_21152,N_26250);
nor U35178 (N_35178,N_20830,N_20007);
nor U35179 (N_35179,N_21837,N_29753);
xor U35180 (N_35180,N_24276,N_21808);
nor U35181 (N_35181,N_26155,N_26141);
nor U35182 (N_35182,N_20214,N_20215);
and U35183 (N_35183,N_25545,N_29304);
nor U35184 (N_35184,N_24923,N_29521);
nand U35185 (N_35185,N_24702,N_24388);
nand U35186 (N_35186,N_21946,N_22681);
and U35187 (N_35187,N_29056,N_20056);
nand U35188 (N_35188,N_20015,N_26461);
or U35189 (N_35189,N_29902,N_23383);
and U35190 (N_35190,N_28520,N_22060);
nand U35191 (N_35191,N_26563,N_23962);
or U35192 (N_35192,N_26113,N_24178);
nor U35193 (N_35193,N_23133,N_20799);
nand U35194 (N_35194,N_27556,N_28463);
nand U35195 (N_35195,N_25157,N_29170);
or U35196 (N_35196,N_23012,N_29066);
and U35197 (N_35197,N_26316,N_28939);
nand U35198 (N_35198,N_29417,N_27118);
nand U35199 (N_35199,N_23697,N_28211);
nand U35200 (N_35200,N_20166,N_20084);
nand U35201 (N_35201,N_28906,N_20045);
nand U35202 (N_35202,N_25257,N_27506);
xor U35203 (N_35203,N_22450,N_21886);
or U35204 (N_35204,N_24726,N_24300);
xor U35205 (N_35205,N_24723,N_21518);
nor U35206 (N_35206,N_24118,N_24275);
nand U35207 (N_35207,N_26151,N_28070);
and U35208 (N_35208,N_28721,N_25053);
nor U35209 (N_35209,N_20112,N_25180);
nand U35210 (N_35210,N_29109,N_26906);
or U35211 (N_35211,N_21722,N_27400);
nor U35212 (N_35212,N_29726,N_23929);
or U35213 (N_35213,N_25612,N_20562);
and U35214 (N_35214,N_23142,N_20344);
or U35215 (N_35215,N_24515,N_26704);
nor U35216 (N_35216,N_20080,N_29987);
nor U35217 (N_35217,N_20051,N_23694);
nor U35218 (N_35218,N_23233,N_27904);
or U35219 (N_35219,N_29756,N_22134);
or U35220 (N_35220,N_22560,N_25407);
nand U35221 (N_35221,N_24319,N_25988);
xor U35222 (N_35222,N_21143,N_29175);
xnor U35223 (N_35223,N_28119,N_22792);
nand U35224 (N_35224,N_27513,N_22443);
nor U35225 (N_35225,N_29180,N_26919);
and U35226 (N_35226,N_23676,N_29463);
nor U35227 (N_35227,N_29053,N_24101);
nand U35228 (N_35228,N_24880,N_25079);
or U35229 (N_35229,N_26822,N_24390);
nor U35230 (N_35230,N_27663,N_21403);
and U35231 (N_35231,N_21105,N_20523);
nor U35232 (N_35232,N_28220,N_28816);
nand U35233 (N_35233,N_28945,N_26151);
nand U35234 (N_35234,N_28489,N_20764);
nand U35235 (N_35235,N_21897,N_20685);
nand U35236 (N_35236,N_25964,N_22810);
nor U35237 (N_35237,N_28868,N_22901);
xnor U35238 (N_35238,N_21769,N_26590);
nor U35239 (N_35239,N_20269,N_25787);
nor U35240 (N_35240,N_28740,N_27952);
nor U35241 (N_35241,N_20137,N_24462);
nor U35242 (N_35242,N_23993,N_23990);
and U35243 (N_35243,N_21443,N_21704);
and U35244 (N_35244,N_22025,N_25860);
and U35245 (N_35245,N_20951,N_24701);
and U35246 (N_35246,N_21432,N_20515);
xor U35247 (N_35247,N_21212,N_20370);
and U35248 (N_35248,N_27242,N_26421);
nand U35249 (N_35249,N_24635,N_26761);
nor U35250 (N_35250,N_24965,N_22814);
nand U35251 (N_35251,N_24656,N_25312);
or U35252 (N_35252,N_20829,N_22155);
or U35253 (N_35253,N_22900,N_22408);
nand U35254 (N_35254,N_20539,N_20123);
xor U35255 (N_35255,N_21846,N_21654);
nor U35256 (N_35256,N_29364,N_29848);
nor U35257 (N_35257,N_23443,N_27953);
xor U35258 (N_35258,N_26965,N_23931);
and U35259 (N_35259,N_27973,N_28735);
or U35260 (N_35260,N_22500,N_28251);
nand U35261 (N_35261,N_23973,N_24168);
nor U35262 (N_35262,N_22452,N_26671);
and U35263 (N_35263,N_26661,N_29104);
or U35264 (N_35264,N_29675,N_28462);
xor U35265 (N_35265,N_24331,N_22416);
nand U35266 (N_35266,N_24862,N_28797);
and U35267 (N_35267,N_21431,N_21977);
nor U35268 (N_35268,N_26081,N_27634);
and U35269 (N_35269,N_22964,N_23905);
nor U35270 (N_35270,N_20026,N_20758);
nand U35271 (N_35271,N_27466,N_21698);
and U35272 (N_35272,N_20605,N_26329);
nor U35273 (N_35273,N_20586,N_24334);
or U35274 (N_35274,N_20078,N_23252);
or U35275 (N_35275,N_23502,N_23208);
or U35276 (N_35276,N_23065,N_28137);
nand U35277 (N_35277,N_21696,N_24362);
nor U35278 (N_35278,N_22831,N_28038);
and U35279 (N_35279,N_23080,N_28823);
nand U35280 (N_35280,N_27699,N_20002);
and U35281 (N_35281,N_29434,N_29074);
xnor U35282 (N_35282,N_21372,N_21336);
or U35283 (N_35283,N_22665,N_29290);
nand U35284 (N_35284,N_27486,N_24386);
and U35285 (N_35285,N_26487,N_20289);
xnor U35286 (N_35286,N_27641,N_21708);
and U35287 (N_35287,N_24251,N_23445);
and U35288 (N_35288,N_27200,N_28697);
nand U35289 (N_35289,N_24258,N_25127);
xnor U35290 (N_35290,N_21795,N_27146);
and U35291 (N_35291,N_25838,N_27596);
or U35292 (N_35292,N_26729,N_20104);
nor U35293 (N_35293,N_25173,N_27032);
and U35294 (N_35294,N_20148,N_23855);
nor U35295 (N_35295,N_25122,N_22414);
and U35296 (N_35296,N_29896,N_24996);
nor U35297 (N_35297,N_27935,N_22076);
nand U35298 (N_35298,N_23402,N_21581);
or U35299 (N_35299,N_28803,N_29078);
and U35300 (N_35300,N_23274,N_27695);
or U35301 (N_35301,N_22229,N_25273);
xnor U35302 (N_35302,N_26481,N_24413);
nor U35303 (N_35303,N_28908,N_22608);
nand U35304 (N_35304,N_21034,N_24734);
or U35305 (N_35305,N_23194,N_21988);
nor U35306 (N_35306,N_25545,N_29441);
nand U35307 (N_35307,N_20451,N_21090);
and U35308 (N_35308,N_21376,N_24031);
nor U35309 (N_35309,N_22181,N_25389);
xor U35310 (N_35310,N_22856,N_26831);
nand U35311 (N_35311,N_28714,N_26406);
nand U35312 (N_35312,N_24995,N_22157);
nor U35313 (N_35313,N_27213,N_24610);
nand U35314 (N_35314,N_25912,N_21782);
nor U35315 (N_35315,N_29045,N_26766);
or U35316 (N_35316,N_24799,N_25629);
and U35317 (N_35317,N_29515,N_23662);
or U35318 (N_35318,N_22853,N_23754);
xnor U35319 (N_35319,N_23743,N_22480);
xor U35320 (N_35320,N_28842,N_20447);
xor U35321 (N_35321,N_21213,N_24389);
nand U35322 (N_35322,N_22198,N_20940);
nor U35323 (N_35323,N_28539,N_25590);
and U35324 (N_35324,N_26223,N_24970);
nor U35325 (N_35325,N_24787,N_21399);
nand U35326 (N_35326,N_23921,N_28969);
or U35327 (N_35327,N_20622,N_26383);
nand U35328 (N_35328,N_24565,N_29737);
nand U35329 (N_35329,N_27293,N_29561);
nor U35330 (N_35330,N_27230,N_21495);
nand U35331 (N_35331,N_28321,N_24360);
and U35332 (N_35332,N_29281,N_24271);
nand U35333 (N_35333,N_23625,N_27671);
or U35334 (N_35334,N_28299,N_20178);
xnor U35335 (N_35335,N_22833,N_20051);
nand U35336 (N_35336,N_27208,N_26443);
nor U35337 (N_35337,N_27795,N_22443);
nor U35338 (N_35338,N_20818,N_23504);
nand U35339 (N_35339,N_26944,N_20508);
and U35340 (N_35340,N_20085,N_21749);
and U35341 (N_35341,N_24737,N_27321);
nand U35342 (N_35342,N_21258,N_24953);
nand U35343 (N_35343,N_22165,N_25776);
or U35344 (N_35344,N_24533,N_21463);
nor U35345 (N_35345,N_21783,N_23205);
nor U35346 (N_35346,N_26191,N_29359);
nand U35347 (N_35347,N_21849,N_22630);
xor U35348 (N_35348,N_27576,N_20943);
or U35349 (N_35349,N_23197,N_25959);
and U35350 (N_35350,N_20491,N_20742);
and U35351 (N_35351,N_28956,N_21145);
or U35352 (N_35352,N_27283,N_26920);
or U35353 (N_35353,N_22619,N_25931);
nand U35354 (N_35354,N_28079,N_26062);
or U35355 (N_35355,N_26296,N_27209);
nor U35356 (N_35356,N_20379,N_28919);
or U35357 (N_35357,N_27592,N_29160);
nand U35358 (N_35358,N_21781,N_28182);
and U35359 (N_35359,N_26827,N_28320);
or U35360 (N_35360,N_23584,N_20506);
xor U35361 (N_35361,N_21545,N_28814);
nand U35362 (N_35362,N_24569,N_27907);
nand U35363 (N_35363,N_27964,N_24294);
nor U35364 (N_35364,N_24252,N_24875);
nor U35365 (N_35365,N_22529,N_29050);
and U35366 (N_35366,N_25948,N_25682);
nor U35367 (N_35367,N_21759,N_23032);
xnor U35368 (N_35368,N_23327,N_27357);
or U35369 (N_35369,N_29875,N_21388);
nor U35370 (N_35370,N_22457,N_26836);
and U35371 (N_35371,N_29606,N_21928);
or U35372 (N_35372,N_22560,N_26630);
and U35373 (N_35373,N_29351,N_24442);
and U35374 (N_35374,N_20806,N_22125);
and U35375 (N_35375,N_26758,N_23177);
and U35376 (N_35376,N_22264,N_27772);
and U35377 (N_35377,N_22063,N_22467);
or U35378 (N_35378,N_23974,N_29385);
nor U35379 (N_35379,N_29380,N_25298);
and U35380 (N_35380,N_21431,N_22327);
or U35381 (N_35381,N_23553,N_20511);
nor U35382 (N_35382,N_24833,N_27289);
xor U35383 (N_35383,N_28395,N_24463);
nand U35384 (N_35384,N_23790,N_23965);
or U35385 (N_35385,N_29842,N_25858);
nor U35386 (N_35386,N_29773,N_25848);
nand U35387 (N_35387,N_20111,N_20456);
nor U35388 (N_35388,N_25871,N_26127);
nand U35389 (N_35389,N_24740,N_26768);
nand U35390 (N_35390,N_20803,N_24399);
nor U35391 (N_35391,N_23512,N_29146);
nor U35392 (N_35392,N_20012,N_23819);
and U35393 (N_35393,N_20205,N_21112);
and U35394 (N_35394,N_24045,N_29609);
nand U35395 (N_35395,N_29594,N_23034);
nand U35396 (N_35396,N_22130,N_26945);
nand U35397 (N_35397,N_24370,N_23616);
or U35398 (N_35398,N_20503,N_26748);
and U35399 (N_35399,N_21669,N_24100);
xor U35400 (N_35400,N_21774,N_22603);
nand U35401 (N_35401,N_26114,N_26420);
nor U35402 (N_35402,N_29877,N_26684);
nor U35403 (N_35403,N_28107,N_29258);
and U35404 (N_35404,N_28656,N_22554);
nand U35405 (N_35405,N_29360,N_22756);
or U35406 (N_35406,N_28238,N_26121);
nand U35407 (N_35407,N_24899,N_23933);
or U35408 (N_35408,N_29069,N_25172);
xor U35409 (N_35409,N_27301,N_28887);
nand U35410 (N_35410,N_26651,N_20767);
xnor U35411 (N_35411,N_25099,N_22804);
or U35412 (N_35412,N_25586,N_28376);
or U35413 (N_35413,N_28557,N_21066);
or U35414 (N_35414,N_22397,N_24681);
xor U35415 (N_35415,N_28680,N_22976);
nor U35416 (N_35416,N_26669,N_26435);
and U35417 (N_35417,N_20518,N_22262);
nor U35418 (N_35418,N_27221,N_28750);
nor U35419 (N_35419,N_21616,N_27166);
nand U35420 (N_35420,N_23730,N_21492);
nor U35421 (N_35421,N_28936,N_28837);
or U35422 (N_35422,N_23641,N_28588);
xnor U35423 (N_35423,N_28543,N_23689);
and U35424 (N_35424,N_25160,N_28212);
xnor U35425 (N_35425,N_29144,N_26981);
nor U35426 (N_35426,N_28521,N_20003);
or U35427 (N_35427,N_24234,N_26517);
nor U35428 (N_35428,N_25420,N_22229);
nor U35429 (N_35429,N_22377,N_23521);
or U35430 (N_35430,N_21263,N_20498);
nor U35431 (N_35431,N_27972,N_21366);
nand U35432 (N_35432,N_23656,N_21351);
and U35433 (N_35433,N_24112,N_23940);
nor U35434 (N_35434,N_21485,N_28973);
nor U35435 (N_35435,N_25279,N_26985);
or U35436 (N_35436,N_20231,N_21871);
nand U35437 (N_35437,N_20517,N_20385);
nor U35438 (N_35438,N_20837,N_29901);
nand U35439 (N_35439,N_20865,N_25050);
nor U35440 (N_35440,N_27186,N_25642);
nand U35441 (N_35441,N_24990,N_25859);
xor U35442 (N_35442,N_20093,N_20372);
nand U35443 (N_35443,N_20564,N_22118);
nor U35444 (N_35444,N_20558,N_23549);
nor U35445 (N_35445,N_25474,N_24772);
nor U35446 (N_35446,N_22175,N_28810);
nand U35447 (N_35447,N_28983,N_23946);
nand U35448 (N_35448,N_21630,N_28916);
and U35449 (N_35449,N_22087,N_21308);
nand U35450 (N_35450,N_25599,N_25427);
nand U35451 (N_35451,N_27240,N_29526);
nand U35452 (N_35452,N_21462,N_24130);
nand U35453 (N_35453,N_28208,N_21878);
nand U35454 (N_35454,N_20617,N_28138);
nor U35455 (N_35455,N_26440,N_27117);
nand U35456 (N_35456,N_29789,N_28717);
nor U35457 (N_35457,N_27533,N_27545);
or U35458 (N_35458,N_28856,N_27470);
and U35459 (N_35459,N_26912,N_28372);
nand U35460 (N_35460,N_27596,N_29168);
nand U35461 (N_35461,N_25970,N_27226);
or U35462 (N_35462,N_23219,N_27320);
xnor U35463 (N_35463,N_28396,N_20663);
or U35464 (N_35464,N_27916,N_24612);
nor U35465 (N_35465,N_25220,N_24316);
nor U35466 (N_35466,N_25160,N_25722);
nand U35467 (N_35467,N_28923,N_24729);
nor U35468 (N_35468,N_24906,N_26756);
and U35469 (N_35469,N_23184,N_24359);
and U35470 (N_35470,N_23785,N_23371);
nor U35471 (N_35471,N_27921,N_27011);
xnor U35472 (N_35472,N_22429,N_27568);
nand U35473 (N_35473,N_22510,N_26196);
nand U35474 (N_35474,N_22746,N_26691);
nor U35475 (N_35475,N_27892,N_23244);
nand U35476 (N_35476,N_23548,N_27452);
and U35477 (N_35477,N_22989,N_21119);
or U35478 (N_35478,N_28701,N_25886);
and U35479 (N_35479,N_28010,N_29406);
or U35480 (N_35480,N_27462,N_24690);
and U35481 (N_35481,N_28810,N_28404);
nand U35482 (N_35482,N_24578,N_21312);
xnor U35483 (N_35483,N_23180,N_22872);
nand U35484 (N_35484,N_24881,N_26942);
nand U35485 (N_35485,N_24997,N_22231);
nand U35486 (N_35486,N_22726,N_22532);
or U35487 (N_35487,N_20895,N_20962);
or U35488 (N_35488,N_20235,N_24612);
or U35489 (N_35489,N_22126,N_22440);
and U35490 (N_35490,N_22152,N_29587);
nor U35491 (N_35491,N_20826,N_21950);
and U35492 (N_35492,N_27214,N_28020);
nand U35493 (N_35493,N_26170,N_28016);
xnor U35494 (N_35494,N_20956,N_20320);
and U35495 (N_35495,N_20952,N_27127);
nand U35496 (N_35496,N_23343,N_20667);
nand U35497 (N_35497,N_21637,N_23442);
or U35498 (N_35498,N_25763,N_26342);
or U35499 (N_35499,N_21853,N_28666);
nand U35500 (N_35500,N_23341,N_25449);
nand U35501 (N_35501,N_22002,N_21249);
nand U35502 (N_35502,N_23318,N_25735);
nor U35503 (N_35503,N_28311,N_28570);
nand U35504 (N_35504,N_23998,N_24781);
and U35505 (N_35505,N_24656,N_28715);
nand U35506 (N_35506,N_20889,N_25171);
and U35507 (N_35507,N_25051,N_27442);
nor U35508 (N_35508,N_29450,N_25444);
nand U35509 (N_35509,N_23180,N_21337);
nand U35510 (N_35510,N_25492,N_28082);
and U35511 (N_35511,N_24280,N_21491);
or U35512 (N_35512,N_29889,N_27597);
and U35513 (N_35513,N_24196,N_25075);
nand U35514 (N_35514,N_24189,N_20694);
and U35515 (N_35515,N_20334,N_24238);
and U35516 (N_35516,N_26638,N_20810);
and U35517 (N_35517,N_24949,N_28274);
nor U35518 (N_35518,N_25968,N_20202);
nor U35519 (N_35519,N_25234,N_22351);
nor U35520 (N_35520,N_21906,N_25463);
nor U35521 (N_35521,N_29313,N_20866);
and U35522 (N_35522,N_26027,N_24246);
or U35523 (N_35523,N_20164,N_27002);
and U35524 (N_35524,N_23813,N_21722);
and U35525 (N_35525,N_25156,N_20498);
and U35526 (N_35526,N_22917,N_23634);
or U35527 (N_35527,N_21801,N_21033);
nor U35528 (N_35528,N_20546,N_23104);
xnor U35529 (N_35529,N_27769,N_21721);
or U35530 (N_35530,N_29830,N_24601);
xor U35531 (N_35531,N_27424,N_21392);
nand U35532 (N_35532,N_24309,N_26989);
nand U35533 (N_35533,N_25765,N_29667);
or U35534 (N_35534,N_22525,N_25304);
and U35535 (N_35535,N_25587,N_27731);
nor U35536 (N_35536,N_20642,N_23148);
and U35537 (N_35537,N_20642,N_22486);
nor U35538 (N_35538,N_23602,N_29850);
and U35539 (N_35539,N_29533,N_26910);
and U35540 (N_35540,N_24617,N_22580);
nor U35541 (N_35541,N_21853,N_29992);
nand U35542 (N_35542,N_21056,N_26594);
or U35543 (N_35543,N_25761,N_25558);
or U35544 (N_35544,N_28902,N_23836);
nor U35545 (N_35545,N_27925,N_24964);
and U35546 (N_35546,N_22999,N_28414);
and U35547 (N_35547,N_20720,N_24019);
and U35548 (N_35548,N_22181,N_21497);
nor U35549 (N_35549,N_27552,N_23886);
and U35550 (N_35550,N_28219,N_29847);
or U35551 (N_35551,N_21149,N_20718);
nand U35552 (N_35552,N_29926,N_24906);
or U35553 (N_35553,N_23688,N_23950);
nand U35554 (N_35554,N_24330,N_29272);
or U35555 (N_35555,N_28412,N_23727);
nand U35556 (N_35556,N_21503,N_25700);
or U35557 (N_35557,N_22056,N_29963);
or U35558 (N_35558,N_22721,N_25175);
or U35559 (N_35559,N_29255,N_29692);
or U35560 (N_35560,N_26473,N_20738);
or U35561 (N_35561,N_20800,N_20176);
and U35562 (N_35562,N_28405,N_25618);
and U35563 (N_35563,N_25353,N_26451);
and U35564 (N_35564,N_27085,N_23277);
or U35565 (N_35565,N_24897,N_22165);
xor U35566 (N_35566,N_24832,N_28129);
nor U35567 (N_35567,N_29494,N_20209);
nor U35568 (N_35568,N_21008,N_24253);
nand U35569 (N_35569,N_25953,N_29292);
or U35570 (N_35570,N_25598,N_22194);
nor U35571 (N_35571,N_24606,N_21526);
and U35572 (N_35572,N_24597,N_20442);
or U35573 (N_35573,N_24684,N_24233);
nand U35574 (N_35574,N_29578,N_21226);
and U35575 (N_35575,N_26290,N_20992);
and U35576 (N_35576,N_28977,N_22080);
and U35577 (N_35577,N_28490,N_24959);
xnor U35578 (N_35578,N_27922,N_28207);
or U35579 (N_35579,N_24019,N_29986);
nor U35580 (N_35580,N_26602,N_22683);
nor U35581 (N_35581,N_28969,N_26702);
nand U35582 (N_35582,N_28661,N_26222);
nand U35583 (N_35583,N_24456,N_29630);
or U35584 (N_35584,N_24908,N_25282);
or U35585 (N_35585,N_28626,N_26989);
nand U35586 (N_35586,N_28660,N_24857);
or U35587 (N_35587,N_21686,N_23728);
or U35588 (N_35588,N_22360,N_21171);
nor U35589 (N_35589,N_20724,N_23213);
and U35590 (N_35590,N_20406,N_29845);
nand U35591 (N_35591,N_26630,N_21167);
and U35592 (N_35592,N_24470,N_23672);
nor U35593 (N_35593,N_23082,N_25526);
or U35594 (N_35594,N_25386,N_22416);
nor U35595 (N_35595,N_25110,N_20399);
nand U35596 (N_35596,N_27783,N_28683);
nand U35597 (N_35597,N_23792,N_21868);
and U35598 (N_35598,N_27268,N_26963);
or U35599 (N_35599,N_24811,N_26085);
nor U35600 (N_35600,N_23251,N_26385);
nor U35601 (N_35601,N_22417,N_22286);
nand U35602 (N_35602,N_20138,N_21306);
nor U35603 (N_35603,N_28483,N_28524);
or U35604 (N_35604,N_28664,N_24300);
or U35605 (N_35605,N_20848,N_27812);
nor U35606 (N_35606,N_20834,N_26575);
nor U35607 (N_35607,N_21281,N_28111);
and U35608 (N_35608,N_22507,N_24643);
nor U35609 (N_35609,N_29730,N_22373);
nor U35610 (N_35610,N_24670,N_26664);
nand U35611 (N_35611,N_23165,N_28691);
nand U35612 (N_35612,N_26636,N_28760);
nand U35613 (N_35613,N_23513,N_20513);
and U35614 (N_35614,N_28348,N_26567);
and U35615 (N_35615,N_25428,N_23701);
or U35616 (N_35616,N_29405,N_21972);
or U35617 (N_35617,N_25385,N_23991);
nor U35618 (N_35618,N_21589,N_28860);
xor U35619 (N_35619,N_23626,N_29672);
nor U35620 (N_35620,N_21403,N_25894);
nor U35621 (N_35621,N_29223,N_20725);
nor U35622 (N_35622,N_27705,N_21511);
nand U35623 (N_35623,N_25762,N_22257);
nor U35624 (N_35624,N_24900,N_26827);
and U35625 (N_35625,N_25665,N_22212);
or U35626 (N_35626,N_23981,N_29199);
nand U35627 (N_35627,N_22078,N_28231);
nand U35628 (N_35628,N_28999,N_20278);
or U35629 (N_35629,N_26015,N_20329);
and U35630 (N_35630,N_21440,N_21199);
and U35631 (N_35631,N_25758,N_20383);
or U35632 (N_35632,N_23785,N_25465);
and U35633 (N_35633,N_20156,N_21415);
or U35634 (N_35634,N_22380,N_21404);
nand U35635 (N_35635,N_21718,N_22548);
or U35636 (N_35636,N_27892,N_24843);
xor U35637 (N_35637,N_22612,N_22100);
nand U35638 (N_35638,N_28648,N_22795);
or U35639 (N_35639,N_27128,N_27410);
and U35640 (N_35640,N_27174,N_20997);
nand U35641 (N_35641,N_27238,N_25546);
nor U35642 (N_35642,N_26011,N_23518);
nand U35643 (N_35643,N_21517,N_29819);
or U35644 (N_35644,N_27795,N_27395);
nand U35645 (N_35645,N_28273,N_29836);
nor U35646 (N_35646,N_27255,N_29186);
and U35647 (N_35647,N_25311,N_22462);
or U35648 (N_35648,N_22186,N_21951);
nor U35649 (N_35649,N_21264,N_28871);
and U35650 (N_35650,N_24612,N_24350);
and U35651 (N_35651,N_29952,N_26801);
nand U35652 (N_35652,N_22224,N_25549);
xnor U35653 (N_35653,N_21193,N_24040);
and U35654 (N_35654,N_24711,N_28977);
xnor U35655 (N_35655,N_20313,N_27521);
or U35656 (N_35656,N_27403,N_22336);
nor U35657 (N_35657,N_28659,N_25549);
and U35658 (N_35658,N_20166,N_26058);
nand U35659 (N_35659,N_21993,N_21031);
nor U35660 (N_35660,N_28976,N_26311);
nor U35661 (N_35661,N_22430,N_29751);
and U35662 (N_35662,N_29942,N_25641);
nor U35663 (N_35663,N_25952,N_21833);
nor U35664 (N_35664,N_20868,N_29170);
or U35665 (N_35665,N_26209,N_20758);
and U35666 (N_35666,N_25399,N_24604);
nand U35667 (N_35667,N_20276,N_20181);
and U35668 (N_35668,N_22487,N_29098);
nor U35669 (N_35669,N_23070,N_26772);
and U35670 (N_35670,N_29934,N_22079);
nand U35671 (N_35671,N_29562,N_27095);
and U35672 (N_35672,N_24990,N_25811);
or U35673 (N_35673,N_21501,N_29837);
nor U35674 (N_35674,N_24935,N_22985);
and U35675 (N_35675,N_28754,N_22208);
nand U35676 (N_35676,N_29839,N_20813);
or U35677 (N_35677,N_23517,N_22416);
nor U35678 (N_35678,N_28418,N_23246);
or U35679 (N_35679,N_25502,N_29536);
and U35680 (N_35680,N_20825,N_26827);
nand U35681 (N_35681,N_27784,N_22011);
xnor U35682 (N_35682,N_20005,N_22729);
nor U35683 (N_35683,N_21988,N_27516);
nor U35684 (N_35684,N_28169,N_21888);
nor U35685 (N_35685,N_25084,N_23387);
nor U35686 (N_35686,N_22497,N_25922);
nand U35687 (N_35687,N_22889,N_25041);
and U35688 (N_35688,N_23329,N_21492);
nand U35689 (N_35689,N_23789,N_26698);
and U35690 (N_35690,N_28115,N_22806);
or U35691 (N_35691,N_24149,N_23255);
nand U35692 (N_35692,N_25055,N_27952);
nor U35693 (N_35693,N_25886,N_26181);
and U35694 (N_35694,N_25941,N_29688);
nand U35695 (N_35695,N_28589,N_24175);
and U35696 (N_35696,N_20303,N_21077);
xnor U35697 (N_35697,N_24684,N_20830);
and U35698 (N_35698,N_27248,N_20128);
nor U35699 (N_35699,N_20015,N_28528);
or U35700 (N_35700,N_24197,N_25787);
and U35701 (N_35701,N_21597,N_23496);
and U35702 (N_35702,N_28550,N_23063);
nand U35703 (N_35703,N_22796,N_27300);
nand U35704 (N_35704,N_27130,N_21456);
or U35705 (N_35705,N_24176,N_28931);
nand U35706 (N_35706,N_29311,N_20346);
and U35707 (N_35707,N_23872,N_29921);
or U35708 (N_35708,N_21540,N_21885);
or U35709 (N_35709,N_25650,N_21944);
xnor U35710 (N_35710,N_29276,N_21786);
and U35711 (N_35711,N_24578,N_23526);
and U35712 (N_35712,N_20438,N_29583);
nor U35713 (N_35713,N_20264,N_21280);
nand U35714 (N_35714,N_25960,N_27270);
nand U35715 (N_35715,N_25580,N_29329);
and U35716 (N_35716,N_20578,N_27946);
nor U35717 (N_35717,N_29684,N_23858);
xnor U35718 (N_35718,N_27294,N_23312);
xor U35719 (N_35719,N_24091,N_21305);
nand U35720 (N_35720,N_25260,N_21165);
nand U35721 (N_35721,N_25020,N_26825);
nor U35722 (N_35722,N_24199,N_22789);
nand U35723 (N_35723,N_29112,N_25344);
or U35724 (N_35724,N_29919,N_20724);
nor U35725 (N_35725,N_21629,N_27924);
xnor U35726 (N_35726,N_22517,N_21747);
or U35727 (N_35727,N_28438,N_22526);
nand U35728 (N_35728,N_25280,N_25239);
or U35729 (N_35729,N_25487,N_22360);
or U35730 (N_35730,N_24521,N_22782);
nand U35731 (N_35731,N_23621,N_23179);
nand U35732 (N_35732,N_27774,N_24953);
xor U35733 (N_35733,N_22520,N_24366);
nor U35734 (N_35734,N_26151,N_23063);
nor U35735 (N_35735,N_26579,N_20989);
xor U35736 (N_35736,N_20960,N_25892);
or U35737 (N_35737,N_27328,N_28233);
nand U35738 (N_35738,N_20337,N_20523);
and U35739 (N_35739,N_24368,N_24400);
and U35740 (N_35740,N_20477,N_28208);
nand U35741 (N_35741,N_20504,N_21061);
nand U35742 (N_35742,N_24638,N_25498);
or U35743 (N_35743,N_23226,N_24078);
and U35744 (N_35744,N_21472,N_28879);
or U35745 (N_35745,N_29127,N_29913);
nor U35746 (N_35746,N_21795,N_23436);
or U35747 (N_35747,N_23597,N_29575);
or U35748 (N_35748,N_20148,N_27037);
or U35749 (N_35749,N_25832,N_23422);
nand U35750 (N_35750,N_28241,N_20775);
nand U35751 (N_35751,N_25315,N_25632);
nand U35752 (N_35752,N_29551,N_26207);
xnor U35753 (N_35753,N_22095,N_23484);
and U35754 (N_35754,N_23758,N_28474);
nor U35755 (N_35755,N_20054,N_22204);
or U35756 (N_35756,N_25231,N_20478);
nor U35757 (N_35757,N_28318,N_26874);
nand U35758 (N_35758,N_27084,N_25964);
nor U35759 (N_35759,N_29873,N_24046);
or U35760 (N_35760,N_23578,N_26304);
or U35761 (N_35761,N_25619,N_27242);
or U35762 (N_35762,N_23996,N_20773);
nand U35763 (N_35763,N_29353,N_22454);
nor U35764 (N_35764,N_24467,N_20911);
or U35765 (N_35765,N_25661,N_20226);
nor U35766 (N_35766,N_22586,N_22627);
nor U35767 (N_35767,N_25703,N_28076);
nand U35768 (N_35768,N_21095,N_26903);
and U35769 (N_35769,N_29223,N_22992);
and U35770 (N_35770,N_21618,N_27150);
and U35771 (N_35771,N_29880,N_25767);
nand U35772 (N_35772,N_20333,N_29380);
nor U35773 (N_35773,N_29324,N_28839);
nand U35774 (N_35774,N_29010,N_20340);
nand U35775 (N_35775,N_20948,N_26827);
and U35776 (N_35776,N_23416,N_21458);
and U35777 (N_35777,N_24876,N_22763);
xor U35778 (N_35778,N_25958,N_27300);
nor U35779 (N_35779,N_21826,N_26938);
nor U35780 (N_35780,N_22812,N_27644);
nand U35781 (N_35781,N_29402,N_21440);
nor U35782 (N_35782,N_25307,N_20315);
xnor U35783 (N_35783,N_20023,N_27295);
or U35784 (N_35784,N_24574,N_24153);
nor U35785 (N_35785,N_25510,N_20695);
or U35786 (N_35786,N_27877,N_29421);
nor U35787 (N_35787,N_26022,N_27830);
and U35788 (N_35788,N_27663,N_28359);
nor U35789 (N_35789,N_28178,N_24708);
or U35790 (N_35790,N_21278,N_25592);
xor U35791 (N_35791,N_21832,N_21125);
nand U35792 (N_35792,N_25108,N_26167);
and U35793 (N_35793,N_28660,N_26477);
and U35794 (N_35794,N_22366,N_27604);
nor U35795 (N_35795,N_24322,N_29671);
nor U35796 (N_35796,N_26860,N_26878);
nand U35797 (N_35797,N_22807,N_23815);
or U35798 (N_35798,N_22036,N_24695);
or U35799 (N_35799,N_21655,N_22305);
xnor U35800 (N_35800,N_24246,N_28806);
or U35801 (N_35801,N_20954,N_26101);
nand U35802 (N_35802,N_28272,N_21118);
and U35803 (N_35803,N_26143,N_25054);
nor U35804 (N_35804,N_28270,N_25273);
nand U35805 (N_35805,N_27251,N_27454);
and U35806 (N_35806,N_24644,N_24505);
nor U35807 (N_35807,N_24446,N_27012);
nor U35808 (N_35808,N_26852,N_22754);
xor U35809 (N_35809,N_25912,N_20970);
nor U35810 (N_35810,N_22374,N_28792);
and U35811 (N_35811,N_28499,N_27287);
or U35812 (N_35812,N_21276,N_27180);
xor U35813 (N_35813,N_27540,N_25640);
nand U35814 (N_35814,N_21120,N_29002);
nor U35815 (N_35815,N_27334,N_20515);
nor U35816 (N_35816,N_22281,N_29621);
nor U35817 (N_35817,N_23797,N_21146);
and U35818 (N_35818,N_24973,N_24810);
xnor U35819 (N_35819,N_21916,N_27806);
nand U35820 (N_35820,N_20349,N_22371);
nand U35821 (N_35821,N_20744,N_28683);
nor U35822 (N_35822,N_26364,N_21517);
xor U35823 (N_35823,N_25358,N_29418);
nor U35824 (N_35824,N_28548,N_23456);
or U35825 (N_35825,N_27871,N_26840);
nand U35826 (N_35826,N_26435,N_20458);
or U35827 (N_35827,N_22842,N_24278);
nor U35828 (N_35828,N_22083,N_25183);
and U35829 (N_35829,N_21328,N_25060);
xor U35830 (N_35830,N_20568,N_23515);
nand U35831 (N_35831,N_21026,N_20007);
and U35832 (N_35832,N_23414,N_28290);
nand U35833 (N_35833,N_20364,N_24333);
nor U35834 (N_35834,N_26473,N_29853);
nor U35835 (N_35835,N_20901,N_23239);
nor U35836 (N_35836,N_21977,N_22495);
xor U35837 (N_35837,N_29838,N_20308);
and U35838 (N_35838,N_23733,N_28105);
or U35839 (N_35839,N_27406,N_21193);
nor U35840 (N_35840,N_27651,N_28482);
or U35841 (N_35841,N_29003,N_24413);
nand U35842 (N_35842,N_23421,N_29301);
or U35843 (N_35843,N_20132,N_27706);
or U35844 (N_35844,N_22770,N_22200);
and U35845 (N_35845,N_23875,N_22691);
and U35846 (N_35846,N_20673,N_23183);
or U35847 (N_35847,N_26831,N_26430);
or U35848 (N_35848,N_29838,N_24966);
nor U35849 (N_35849,N_22471,N_29454);
nor U35850 (N_35850,N_25890,N_28731);
or U35851 (N_35851,N_20469,N_20905);
nand U35852 (N_35852,N_29618,N_27271);
nor U35853 (N_35853,N_27320,N_22205);
or U35854 (N_35854,N_23894,N_21236);
or U35855 (N_35855,N_20017,N_26219);
and U35856 (N_35856,N_23351,N_23584);
nor U35857 (N_35857,N_27860,N_28476);
or U35858 (N_35858,N_20706,N_21755);
nor U35859 (N_35859,N_22439,N_25697);
and U35860 (N_35860,N_27101,N_21248);
or U35861 (N_35861,N_27651,N_20772);
and U35862 (N_35862,N_21616,N_23697);
and U35863 (N_35863,N_29431,N_21261);
nor U35864 (N_35864,N_25360,N_29750);
nor U35865 (N_35865,N_25872,N_28952);
nand U35866 (N_35866,N_23398,N_29492);
or U35867 (N_35867,N_20688,N_23957);
nand U35868 (N_35868,N_24825,N_21164);
nor U35869 (N_35869,N_26106,N_29344);
and U35870 (N_35870,N_28004,N_21600);
nor U35871 (N_35871,N_21355,N_20613);
nor U35872 (N_35872,N_20532,N_25993);
nand U35873 (N_35873,N_27237,N_25594);
nor U35874 (N_35874,N_29201,N_28090);
and U35875 (N_35875,N_27095,N_28533);
nor U35876 (N_35876,N_27219,N_22684);
nand U35877 (N_35877,N_26893,N_26726);
and U35878 (N_35878,N_25952,N_29212);
or U35879 (N_35879,N_27043,N_26560);
nand U35880 (N_35880,N_21035,N_25271);
nand U35881 (N_35881,N_29494,N_24472);
or U35882 (N_35882,N_26766,N_29853);
nand U35883 (N_35883,N_25981,N_28252);
or U35884 (N_35884,N_25122,N_23181);
nor U35885 (N_35885,N_25168,N_26431);
nor U35886 (N_35886,N_29994,N_29001);
or U35887 (N_35887,N_25747,N_29681);
and U35888 (N_35888,N_27157,N_21303);
or U35889 (N_35889,N_22657,N_22547);
nor U35890 (N_35890,N_28343,N_20700);
nand U35891 (N_35891,N_25821,N_24487);
or U35892 (N_35892,N_28973,N_26505);
nand U35893 (N_35893,N_22634,N_22359);
and U35894 (N_35894,N_23506,N_25515);
xnor U35895 (N_35895,N_22999,N_21868);
nand U35896 (N_35896,N_22525,N_20780);
nand U35897 (N_35897,N_24985,N_23294);
and U35898 (N_35898,N_21841,N_23251);
nand U35899 (N_35899,N_24303,N_25078);
and U35900 (N_35900,N_26911,N_23709);
nand U35901 (N_35901,N_23165,N_22553);
and U35902 (N_35902,N_29793,N_25802);
nand U35903 (N_35903,N_20478,N_22375);
and U35904 (N_35904,N_22143,N_26360);
xor U35905 (N_35905,N_26788,N_26796);
nor U35906 (N_35906,N_25880,N_27932);
nand U35907 (N_35907,N_25740,N_24817);
or U35908 (N_35908,N_22928,N_25014);
nor U35909 (N_35909,N_22869,N_20253);
and U35910 (N_35910,N_25014,N_27243);
nand U35911 (N_35911,N_27391,N_25872);
nor U35912 (N_35912,N_27436,N_25481);
and U35913 (N_35913,N_21549,N_22206);
nand U35914 (N_35914,N_20527,N_29097);
or U35915 (N_35915,N_23233,N_21770);
nor U35916 (N_35916,N_25116,N_27724);
nor U35917 (N_35917,N_23365,N_25353);
xor U35918 (N_35918,N_21816,N_27879);
or U35919 (N_35919,N_25991,N_26873);
nand U35920 (N_35920,N_24390,N_24813);
or U35921 (N_35921,N_29878,N_22233);
and U35922 (N_35922,N_28241,N_20839);
or U35923 (N_35923,N_28261,N_28484);
nor U35924 (N_35924,N_20993,N_27337);
nor U35925 (N_35925,N_25648,N_20147);
nand U35926 (N_35926,N_24823,N_28399);
nor U35927 (N_35927,N_28617,N_22839);
or U35928 (N_35928,N_22424,N_27398);
or U35929 (N_35929,N_28426,N_21261);
or U35930 (N_35930,N_26312,N_25100);
and U35931 (N_35931,N_26227,N_25628);
nor U35932 (N_35932,N_29839,N_25214);
and U35933 (N_35933,N_27399,N_29827);
nor U35934 (N_35934,N_23745,N_21163);
nor U35935 (N_35935,N_20649,N_23669);
or U35936 (N_35936,N_27382,N_29253);
nor U35937 (N_35937,N_26481,N_20761);
nand U35938 (N_35938,N_25862,N_22502);
nor U35939 (N_35939,N_20430,N_28710);
or U35940 (N_35940,N_28146,N_23032);
xor U35941 (N_35941,N_25597,N_29512);
and U35942 (N_35942,N_24331,N_26943);
nand U35943 (N_35943,N_24174,N_23470);
or U35944 (N_35944,N_24838,N_21699);
or U35945 (N_35945,N_22478,N_27965);
nor U35946 (N_35946,N_24775,N_25494);
or U35947 (N_35947,N_26635,N_21884);
nor U35948 (N_35948,N_25784,N_27291);
nand U35949 (N_35949,N_28477,N_27766);
nand U35950 (N_35950,N_24887,N_28722);
nor U35951 (N_35951,N_26164,N_25351);
nand U35952 (N_35952,N_20784,N_26099);
nor U35953 (N_35953,N_20267,N_20226);
or U35954 (N_35954,N_26794,N_27569);
xor U35955 (N_35955,N_20899,N_29991);
and U35956 (N_35956,N_29005,N_29419);
nor U35957 (N_35957,N_24736,N_23821);
nor U35958 (N_35958,N_21985,N_20662);
nand U35959 (N_35959,N_29643,N_26757);
nor U35960 (N_35960,N_29599,N_26398);
nor U35961 (N_35961,N_26777,N_26195);
or U35962 (N_35962,N_23962,N_29425);
and U35963 (N_35963,N_25852,N_26356);
nand U35964 (N_35964,N_21841,N_24215);
and U35965 (N_35965,N_27292,N_26915);
and U35966 (N_35966,N_25626,N_24652);
nand U35967 (N_35967,N_20114,N_21979);
nor U35968 (N_35968,N_27057,N_27655);
nor U35969 (N_35969,N_28484,N_28326);
nor U35970 (N_35970,N_27902,N_28163);
nor U35971 (N_35971,N_27641,N_27981);
nor U35972 (N_35972,N_28346,N_29263);
and U35973 (N_35973,N_23926,N_23610);
nor U35974 (N_35974,N_27326,N_22436);
and U35975 (N_35975,N_26865,N_27417);
and U35976 (N_35976,N_23552,N_29524);
nand U35977 (N_35977,N_29130,N_27072);
or U35978 (N_35978,N_27833,N_22182);
and U35979 (N_35979,N_21479,N_26792);
and U35980 (N_35980,N_28949,N_29876);
or U35981 (N_35981,N_28551,N_28766);
and U35982 (N_35982,N_26534,N_28120);
xor U35983 (N_35983,N_28821,N_29499);
nor U35984 (N_35984,N_23947,N_29241);
xnor U35985 (N_35985,N_29666,N_26047);
or U35986 (N_35986,N_23406,N_25641);
or U35987 (N_35987,N_22355,N_29771);
nand U35988 (N_35988,N_28824,N_28030);
nor U35989 (N_35989,N_27619,N_26048);
xnor U35990 (N_35990,N_25102,N_26212);
or U35991 (N_35991,N_28884,N_26577);
nand U35992 (N_35992,N_26942,N_23169);
or U35993 (N_35993,N_26863,N_28604);
nand U35994 (N_35994,N_21714,N_24306);
or U35995 (N_35995,N_22843,N_21571);
or U35996 (N_35996,N_27488,N_26230);
nor U35997 (N_35997,N_21403,N_26360);
nand U35998 (N_35998,N_27518,N_28933);
and U35999 (N_35999,N_24306,N_28051);
nand U36000 (N_36000,N_21106,N_26602);
nor U36001 (N_36001,N_26953,N_26962);
nor U36002 (N_36002,N_26574,N_27345);
nand U36003 (N_36003,N_29613,N_22630);
or U36004 (N_36004,N_21253,N_27421);
xnor U36005 (N_36005,N_25614,N_24661);
nor U36006 (N_36006,N_20446,N_29238);
or U36007 (N_36007,N_23184,N_25967);
nand U36008 (N_36008,N_26372,N_27057);
nor U36009 (N_36009,N_21412,N_24263);
nor U36010 (N_36010,N_29796,N_20442);
or U36011 (N_36011,N_23991,N_29439);
nand U36012 (N_36012,N_26424,N_28601);
and U36013 (N_36013,N_29701,N_26247);
nand U36014 (N_36014,N_26107,N_20031);
or U36015 (N_36015,N_23653,N_25615);
nand U36016 (N_36016,N_29656,N_22874);
or U36017 (N_36017,N_22172,N_20787);
or U36018 (N_36018,N_25993,N_27144);
and U36019 (N_36019,N_29927,N_20242);
xnor U36020 (N_36020,N_26472,N_26498);
xor U36021 (N_36021,N_28866,N_25644);
xor U36022 (N_36022,N_21457,N_22340);
and U36023 (N_36023,N_22875,N_25153);
or U36024 (N_36024,N_20342,N_20079);
nor U36025 (N_36025,N_27125,N_22704);
and U36026 (N_36026,N_24647,N_22426);
nor U36027 (N_36027,N_27523,N_28469);
or U36028 (N_36028,N_22950,N_20159);
nor U36029 (N_36029,N_20912,N_20998);
xor U36030 (N_36030,N_27428,N_23279);
or U36031 (N_36031,N_29847,N_20872);
or U36032 (N_36032,N_21397,N_28287);
and U36033 (N_36033,N_22272,N_23029);
or U36034 (N_36034,N_22991,N_20374);
and U36035 (N_36035,N_24654,N_22215);
xor U36036 (N_36036,N_22504,N_26268);
nor U36037 (N_36037,N_23257,N_27914);
or U36038 (N_36038,N_23132,N_28439);
nand U36039 (N_36039,N_20954,N_26426);
nor U36040 (N_36040,N_29473,N_21958);
nand U36041 (N_36041,N_28713,N_26962);
nor U36042 (N_36042,N_20697,N_27615);
and U36043 (N_36043,N_20303,N_21414);
or U36044 (N_36044,N_23469,N_20248);
nor U36045 (N_36045,N_23765,N_28758);
and U36046 (N_36046,N_27210,N_21028);
or U36047 (N_36047,N_21804,N_22271);
or U36048 (N_36048,N_23227,N_22324);
xnor U36049 (N_36049,N_21856,N_23469);
and U36050 (N_36050,N_26434,N_21148);
or U36051 (N_36051,N_28779,N_25101);
and U36052 (N_36052,N_27536,N_21715);
or U36053 (N_36053,N_28021,N_22620);
nor U36054 (N_36054,N_21661,N_20672);
or U36055 (N_36055,N_23205,N_23960);
nand U36056 (N_36056,N_25597,N_25377);
nor U36057 (N_36057,N_24987,N_21845);
xnor U36058 (N_36058,N_27624,N_28859);
nand U36059 (N_36059,N_25142,N_22265);
and U36060 (N_36060,N_23359,N_23757);
or U36061 (N_36061,N_27507,N_21957);
nand U36062 (N_36062,N_23900,N_24795);
or U36063 (N_36063,N_29091,N_24173);
or U36064 (N_36064,N_25819,N_26004);
nor U36065 (N_36065,N_25096,N_29963);
or U36066 (N_36066,N_25926,N_23807);
and U36067 (N_36067,N_24960,N_27419);
nand U36068 (N_36068,N_29725,N_23872);
nand U36069 (N_36069,N_25645,N_29942);
nand U36070 (N_36070,N_28553,N_27037);
or U36071 (N_36071,N_20196,N_27123);
and U36072 (N_36072,N_23710,N_22626);
xnor U36073 (N_36073,N_23092,N_26528);
nand U36074 (N_36074,N_29114,N_23398);
xor U36075 (N_36075,N_23436,N_22911);
xnor U36076 (N_36076,N_27651,N_24133);
and U36077 (N_36077,N_23231,N_29258);
and U36078 (N_36078,N_20042,N_22985);
nand U36079 (N_36079,N_28322,N_21067);
nor U36080 (N_36080,N_22498,N_28753);
and U36081 (N_36081,N_20325,N_23420);
xnor U36082 (N_36082,N_22499,N_22475);
and U36083 (N_36083,N_23059,N_27578);
nor U36084 (N_36084,N_26900,N_25176);
nor U36085 (N_36085,N_26371,N_27552);
or U36086 (N_36086,N_27360,N_20132);
and U36087 (N_36087,N_22973,N_23404);
or U36088 (N_36088,N_28147,N_22835);
or U36089 (N_36089,N_28507,N_21476);
nand U36090 (N_36090,N_23224,N_24323);
nand U36091 (N_36091,N_23692,N_25725);
nor U36092 (N_36092,N_25336,N_26362);
and U36093 (N_36093,N_21988,N_26637);
and U36094 (N_36094,N_24023,N_27304);
and U36095 (N_36095,N_23014,N_27717);
nand U36096 (N_36096,N_26023,N_25009);
or U36097 (N_36097,N_25879,N_23868);
nor U36098 (N_36098,N_21371,N_28678);
nor U36099 (N_36099,N_29779,N_27513);
nor U36100 (N_36100,N_24639,N_21429);
or U36101 (N_36101,N_20683,N_27413);
nand U36102 (N_36102,N_24684,N_24304);
nand U36103 (N_36103,N_23888,N_24752);
xnor U36104 (N_36104,N_22209,N_22117);
xnor U36105 (N_36105,N_23205,N_20360);
nand U36106 (N_36106,N_29504,N_21611);
nor U36107 (N_36107,N_25610,N_27646);
nand U36108 (N_36108,N_21273,N_20048);
and U36109 (N_36109,N_24810,N_25238);
nand U36110 (N_36110,N_24508,N_20963);
or U36111 (N_36111,N_24508,N_25222);
nor U36112 (N_36112,N_21708,N_21191);
nor U36113 (N_36113,N_20694,N_23798);
nand U36114 (N_36114,N_29259,N_22825);
nor U36115 (N_36115,N_26793,N_29060);
nor U36116 (N_36116,N_20576,N_20152);
and U36117 (N_36117,N_22855,N_28552);
or U36118 (N_36118,N_20766,N_27945);
nor U36119 (N_36119,N_21799,N_25093);
nand U36120 (N_36120,N_29778,N_29285);
nor U36121 (N_36121,N_27186,N_24942);
or U36122 (N_36122,N_29206,N_29478);
xnor U36123 (N_36123,N_20870,N_20350);
nor U36124 (N_36124,N_28225,N_28363);
or U36125 (N_36125,N_27002,N_27848);
nor U36126 (N_36126,N_27811,N_23289);
and U36127 (N_36127,N_26802,N_21118);
or U36128 (N_36128,N_24312,N_29329);
and U36129 (N_36129,N_28876,N_29387);
nor U36130 (N_36130,N_25927,N_24831);
nand U36131 (N_36131,N_20142,N_29098);
and U36132 (N_36132,N_25932,N_22326);
nor U36133 (N_36133,N_29347,N_26599);
nor U36134 (N_36134,N_25940,N_26695);
or U36135 (N_36135,N_29217,N_20622);
and U36136 (N_36136,N_21932,N_22178);
nand U36137 (N_36137,N_22592,N_29096);
xnor U36138 (N_36138,N_22614,N_27656);
nor U36139 (N_36139,N_28434,N_25153);
and U36140 (N_36140,N_24626,N_26635);
or U36141 (N_36141,N_23646,N_26420);
nand U36142 (N_36142,N_27486,N_21232);
and U36143 (N_36143,N_20757,N_23722);
or U36144 (N_36144,N_27232,N_21476);
and U36145 (N_36145,N_24507,N_26578);
nand U36146 (N_36146,N_21361,N_25827);
nand U36147 (N_36147,N_24820,N_23692);
xnor U36148 (N_36148,N_26912,N_28682);
nand U36149 (N_36149,N_29484,N_28658);
nor U36150 (N_36150,N_27491,N_21637);
and U36151 (N_36151,N_22525,N_24661);
nand U36152 (N_36152,N_26537,N_26430);
and U36153 (N_36153,N_27171,N_24522);
xor U36154 (N_36154,N_27577,N_20075);
or U36155 (N_36155,N_24569,N_27187);
and U36156 (N_36156,N_26339,N_26679);
xor U36157 (N_36157,N_23808,N_24265);
or U36158 (N_36158,N_20233,N_25317);
nand U36159 (N_36159,N_27835,N_29170);
xor U36160 (N_36160,N_21027,N_26783);
nand U36161 (N_36161,N_29241,N_22993);
or U36162 (N_36162,N_27993,N_28023);
nand U36163 (N_36163,N_21581,N_22196);
nor U36164 (N_36164,N_21863,N_21710);
or U36165 (N_36165,N_23869,N_22375);
and U36166 (N_36166,N_25671,N_26722);
nand U36167 (N_36167,N_22557,N_27646);
or U36168 (N_36168,N_27543,N_26637);
or U36169 (N_36169,N_24034,N_21789);
or U36170 (N_36170,N_28834,N_20423);
xnor U36171 (N_36171,N_22218,N_27348);
or U36172 (N_36172,N_28553,N_20005);
and U36173 (N_36173,N_24395,N_24558);
nor U36174 (N_36174,N_23651,N_28485);
or U36175 (N_36175,N_26519,N_26337);
or U36176 (N_36176,N_29955,N_27301);
or U36177 (N_36177,N_26008,N_25248);
nor U36178 (N_36178,N_25571,N_21134);
nand U36179 (N_36179,N_27738,N_26972);
or U36180 (N_36180,N_25307,N_26705);
nor U36181 (N_36181,N_21895,N_27309);
or U36182 (N_36182,N_21526,N_21433);
and U36183 (N_36183,N_22422,N_27313);
nand U36184 (N_36184,N_21954,N_28836);
nor U36185 (N_36185,N_22447,N_29170);
or U36186 (N_36186,N_22186,N_20525);
or U36187 (N_36187,N_23542,N_22257);
or U36188 (N_36188,N_21895,N_27214);
or U36189 (N_36189,N_26673,N_22052);
nor U36190 (N_36190,N_21175,N_23770);
or U36191 (N_36191,N_21914,N_25436);
or U36192 (N_36192,N_26622,N_27246);
and U36193 (N_36193,N_23781,N_23207);
nor U36194 (N_36194,N_22056,N_29669);
nand U36195 (N_36195,N_25048,N_27953);
or U36196 (N_36196,N_28880,N_25206);
nand U36197 (N_36197,N_20249,N_27151);
nor U36198 (N_36198,N_28134,N_28105);
or U36199 (N_36199,N_27204,N_27304);
nand U36200 (N_36200,N_22287,N_28465);
nand U36201 (N_36201,N_25734,N_24016);
and U36202 (N_36202,N_22569,N_29952);
and U36203 (N_36203,N_21487,N_26606);
nand U36204 (N_36204,N_28142,N_20426);
and U36205 (N_36205,N_25235,N_27688);
xor U36206 (N_36206,N_20260,N_26659);
xnor U36207 (N_36207,N_26279,N_24386);
or U36208 (N_36208,N_29893,N_26141);
nand U36209 (N_36209,N_20682,N_28623);
nand U36210 (N_36210,N_29884,N_24771);
nor U36211 (N_36211,N_27933,N_20280);
and U36212 (N_36212,N_28106,N_20176);
nor U36213 (N_36213,N_22123,N_21144);
nand U36214 (N_36214,N_27064,N_28709);
nor U36215 (N_36215,N_28480,N_25939);
nor U36216 (N_36216,N_27486,N_29815);
and U36217 (N_36217,N_24428,N_21090);
nand U36218 (N_36218,N_28885,N_22859);
nor U36219 (N_36219,N_29909,N_29463);
and U36220 (N_36220,N_29403,N_20378);
xnor U36221 (N_36221,N_28842,N_23899);
nor U36222 (N_36222,N_28249,N_26122);
and U36223 (N_36223,N_25601,N_21812);
nor U36224 (N_36224,N_25086,N_21650);
xor U36225 (N_36225,N_21152,N_21086);
nor U36226 (N_36226,N_28101,N_27119);
and U36227 (N_36227,N_29303,N_23037);
or U36228 (N_36228,N_22888,N_29408);
nor U36229 (N_36229,N_25009,N_28306);
nor U36230 (N_36230,N_26465,N_29314);
nor U36231 (N_36231,N_27175,N_29930);
or U36232 (N_36232,N_29640,N_29345);
or U36233 (N_36233,N_28210,N_22230);
nor U36234 (N_36234,N_29469,N_27813);
or U36235 (N_36235,N_27276,N_23959);
and U36236 (N_36236,N_20611,N_20363);
nor U36237 (N_36237,N_20904,N_23193);
and U36238 (N_36238,N_22801,N_28593);
nand U36239 (N_36239,N_25498,N_29774);
nand U36240 (N_36240,N_27260,N_22600);
or U36241 (N_36241,N_23823,N_22745);
nand U36242 (N_36242,N_21025,N_22990);
nor U36243 (N_36243,N_28927,N_26819);
xnor U36244 (N_36244,N_24958,N_29953);
and U36245 (N_36245,N_28113,N_27724);
nor U36246 (N_36246,N_25376,N_24573);
nor U36247 (N_36247,N_23441,N_24151);
or U36248 (N_36248,N_26816,N_28515);
nand U36249 (N_36249,N_26041,N_25741);
nand U36250 (N_36250,N_26673,N_24030);
nand U36251 (N_36251,N_22021,N_27937);
or U36252 (N_36252,N_20024,N_28974);
and U36253 (N_36253,N_20061,N_21331);
nor U36254 (N_36254,N_23453,N_21981);
or U36255 (N_36255,N_28003,N_23785);
and U36256 (N_36256,N_27653,N_25072);
or U36257 (N_36257,N_29201,N_25219);
and U36258 (N_36258,N_26181,N_26947);
nand U36259 (N_36259,N_27488,N_28398);
or U36260 (N_36260,N_25264,N_20750);
and U36261 (N_36261,N_23663,N_29799);
nand U36262 (N_36262,N_22824,N_27830);
nand U36263 (N_36263,N_25577,N_27480);
or U36264 (N_36264,N_26700,N_28714);
or U36265 (N_36265,N_27896,N_21968);
and U36266 (N_36266,N_28527,N_25741);
nor U36267 (N_36267,N_21813,N_22720);
and U36268 (N_36268,N_26567,N_23370);
or U36269 (N_36269,N_25478,N_20982);
nand U36270 (N_36270,N_25023,N_29270);
nand U36271 (N_36271,N_28635,N_22504);
nand U36272 (N_36272,N_28582,N_24756);
nor U36273 (N_36273,N_29117,N_21103);
and U36274 (N_36274,N_29390,N_20389);
and U36275 (N_36275,N_21876,N_23952);
or U36276 (N_36276,N_25273,N_24505);
nand U36277 (N_36277,N_25209,N_27258);
or U36278 (N_36278,N_21555,N_27303);
and U36279 (N_36279,N_24675,N_23902);
nor U36280 (N_36280,N_23208,N_29515);
and U36281 (N_36281,N_27596,N_24742);
and U36282 (N_36282,N_21897,N_21914);
or U36283 (N_36283,N_22781,N_28621);
nor U36284 (N_36284,N_22198,N_28155);
nor U36285 (N_36285,N_25383,N_29903);
nand U36286 (N_36286,N_29687,N_28358);
nor U36287 (N_36287,N_25001,N_26018);
and U36288 (N_36288,N_23590,N_25397);
nand U36289 (N_36289,N_25321,N_28720);
and U36290 (N_36290,N_20167,N_22254);
nand U36291 (N_36291,N_20482,N_23843);
xnor U36292 (N_36292,N_29270,N_23948);
and U36293 (N_36293,N_22127,N_25299);
xor U36294 (N_36294,N_22132,N_28281);
or U36295 (N_36295,N_23478,N_28099);
and U36296 (N_36296,N_28839,N_21756);
and U36297 (N_36297,N_23455,N_20791);
and U36298 (N_36298,N_27561,N_25507);
nor U36299 (N_36299,N_28228,N_23450);
nor U36300 (N_36300,N_24867,N_22328);
nor U36301 (N_36301,N_24526,N_27794);
nor U36302 (N_36302,N_23379,N_26187);
nand U36303 (N_36303,N_20224,N_24012);
or U36304 (N_36304,N_21654,N_25247);
nand U36305 (N_36305,N_23339,N_24940);
or U36306 (N_36306,N_28224,N_21541);
and U36307 (N_36307,N_26760,N_28459);
nor U36308 (N_36308,N_20772,N_28233);
nand U36309 (N_36309,N_28483,N_25742);
nor U36310 (N_36310,N_28187,N_26026);
and U36311 (N_36311,N_22349,N_26793);
and U36312 (N_36312,N_26382,N_21744);
and U36313 (N_36313,N_26932,N_26742);
nor U36314 (N_36314,N_21032,N_24096);
or U36315 (N_36315,N_26779,N_28836);
xor U36316 (N_36316,N_22697,N_22155);
nor U36317 (N_36317,N_28679,N_24552);
nor U36318 (N_36318,N_25390,N_24459);
or U36319 (N_36319,N_24657,N_28121);
or U36320 (N_36320,N_24073,N_29835);
or U36321 (N_36321,N_22853,N_22826);
and U36322 (N_36322,N_26721,N_28414);
nor U36323 (N_36323,N_20924,N_25345);
nand U36324 (N_36324,N_25159,N_23948);
nand U36325 (N_36325,N_20561,N_24210);
nand U36326 (N_36326,N_22308,N_26749);
or U36327 (N_36327,N_22748,N_21781);
xor U36328 (N_36328,N_25255,N_22152);
nand U36329 (N_36329,N_25838,N_22862);
xnor U36330 (N_36330,N_27534,N_26582);
xor U36331 (N_36331,N_21740,N_27097);
xor U36332 (N_36332,N_27010,N_25956);
and U36333 (N_36333,N_29984,N_23513);
nand U36334 (N_36334,N_23254,N_23485);
nor U36335 (N_36335,N_21100,N_27880);
nor U36336 (N_36336,N_20230,N_23470);
or U36337 (N_36337,N_24166,N_23301);
nand U36338 (N_36338,N_23359,N_24652);
nand U36339 (N_36339,N_28085,N_22758);
nand U36340 (N_36340,N_24405,N_29035);
nand U36341 (N_36341,N_24618,N_24870);
and U36342 (N_36342,N_28511,N_26514);
and U36343 (N_36343,N_22465,N_29137);
nand U36344 (N_36344,N_23359,N_28755);
and U36345 (N_36345,N_29272,N_25837);
xnor U36346 (N_36346,N_28778,N_24023);
and U36347 (N_36347,N_20282,N_20841);
or U36348 (N_36348,N_21968,N_29947);
and U36349 (N_36349,N_28240,N_28191);
xnor U36350 (N_36350,N_24400,N_20049);
nor U36351 (N_36351,N_24131,N_25156);
nor U36352 (N_36352,N_24127,N_29766);
or U36353 (N_36353,N_28442,N_23505);
and U36354 (N_36354,N_22306,N_28592);
nand U36355 (N_36355,N_20233,N_24390);
and U36356 (N_36356,N_28396,N_23438);
nor U36357 (N_36357,N_27502,N_28158);
and U36358 (N_36358,N_29157,N_21918);
and U36359 (N_36359,N_25743,N_22188);
nand U36360 (N_36360,N_28326,N_25397);
and U36361 (N_36361,N_21699,N_29195);
nor U36362 (N_36362,N_24230,N_23752);
or U36363 (N_36363,N_29946,N_28385);
and U36364 (N_36364,N_28800,N_23873);
nor U36365 (N_36365,N_25249,N_21167);
nand U36366 (N_36366,N_20185,N_20673);
or U36367 (N_36367,N_21491,N_20018);
nor U36368 (N_36368,N_26340,N_21830);
and U36369 (N_36369,N_28782,N_28780);
or U36370 (N_36370,N_29163,N_26569);
and U36371 (N_36371,N_22679,N_22739);
and U36372 (N_36372,N_22719,N_25554);
nor U36373 (N_36373,N_23755,N_24031);
nor U36374 (N_36374,N_21368,N_24731);
nand U36375 (N_36375,N_25154,N_21070);
and U36376 (N_36376,N_23006,N_25997);
nand U36377 (N_36377,N_21801,N_24068);
nor U36378 (N_36378,N_26670,N_25107);
and U36379 (N_36379,N_29303,N_24129);
xor U36380 (N_36380,N_26984,N_21210);
nor U36381 (N_36381,N_22001,N_28207);
or U36382 (N_36382,N_27536,N_22948);
nand U36383 (N_36383,N_26574,N_29042);
and U36384 (N_36384,N_25604,N_24772);
or U36385 (N_36385,N_27324,N_26806);
or U36386 (N_36386,N_26172,N_27432);
nor U36387 (N_36387,N_23258,N_25295);
nand U36388 (N_36388,N_27649,N_22255);
and U36389 (N_36389,N_27108,N_29405);
or U36390 (N_36390,N_26365,N_24161);
nand U36391 (N_36391,N_28287,N_24452);
or U36392 (N_36392,N_24558,N_26958);
nand U36393 (N_36393,N_25083,N_23149);
xor U36394 (N_36394,N_26549,N_28308);
xor U36395 (N_36395,N_20697,N_20049);
or U36396 (N_36396,N_26491,N_23461);
or U36397 (N_36397,N_22788,N_23805);
nor U36398 (N_36398,N_22992,N_22604);
or U36399 (N_36399,N_27127,N_28909);
nor U36400 (N_36400,N_25785,N_22653);
or U36401 (N_36401,N_27482,N_27374);
nor U36402 (N_36402,N_21097,N_23514);
nand U36403 (N_36403,N_24768,N_23103);
nand U36404 (N_36404,N_26597,N_23870);
xor U36405 (N_36405,N_20864,N_26943);
nand U36406 (N_36406,N_24482,N_21055);
nor U36407 (N_36407,N_20196,N_26168);
nor U36408 (N_36408,N_22212,N_22954);
nand U36409 (N_36409,N_23391,N_22152);
xnor U36410 (N_36410,N_26059,N_25863);
nor U36411 (N_36411,N_25275,N_28591);
nand U36412 (N_36412,N_26904,N_24004);
and U36413 (N_36413,N_27571,N_23337);
xnor U36414 (N_36414,N_20563,N_24794);
and U36415 (N_36415,N_29977,N_29413);
and U36416 (N_36416,N_25167,N_26677);
or U36417 (N_36417,N_20342,N_26754);
nor U36418 (N_36418,N_26181,N_22016);
or U36419 (N_36419,N_23459,N_20323);
and U36420 (N_36420,N_29225,N_24923);
nor U36421 (N_36421,N_27373,N_29931);
nor U36422 (N_36422,N_26984,N_24509);
nor U36423 (N_36423,N_26588,N_22956);
nor U36424 (N_36424,N_25072,N_20524);
and U36425 (N_36425,N_24794,N_25823);
and U36426 (N_36426,N_26665,N_29349);
nor U36427 (N_36427,N_25247,N_20549);
xor U36428 (N_36428,N_28782,N_23560);
nand U36429 (N_36429,N_29357,N_28581);
or U36430 (N_36430,N_22486,N_25444);
nand U36431 (N_36431,N_22961,N_22172);
xnor U36432 (N_36432,N_24991,N_23119);
nor U36433 (N_36433,N_28715,N_25383);
xnor U36434 (N_36434,N_23090,N_22536);
or U36435 (N_36435,N_25559,N_24625);
nand U36436 (N_36436,N_20468,N_23191);
and U36437 (N_36437,N_23617,N_20056);
or U36438 (N_36438,N_24401,N_21672);
nand U36439 (N_36439,N_28167,N_20628);
nand U36440 (N_36440,N_22196,N_20007);
nor U36441 (N_36441,N_20586,N_23559);
nor U36442 (N_36442,N_20020,N_21308);
xor U36443 (N_36443,N_28336,N_24385);
nand U36444 (N_36444,N_25176,N_27191);
and U36445 (N_36445,N_22428,N_20436);
nor U36446 (N_36446,N_21079,N_22743);
and U36447 (N_36447,N_22395,N_23321);
or U36448 (N_36448,N_20833,N_22016);
xor U36449 (N_36449,N_27617,N_21015);
or U36450 (N_36450,N_28335,N_26066);
nand U36451 (N_36451,N_25841,N_23391);
nor U36452 (N_36452,N_29106,N_27269);
nor U36453 (N_36453,N_20752,N_26837);
nor U36454 (N_36454,N_24597,N_21754);
nor U36455 (N_36455,N_24651,N_29134);
nand U36456 (N_36456,N_23117,N_29587);
nor U36457 (N_36457,N_26591,N_28410);
nor U36458 (N_36458,N_20079,N_26212);
and U36459 (N_36459,N_20531,N_20044);
nand U36460 (N_36460,N_27764,N_21930);
nand U36461 (N_36461,N_29625,N_24790);
and U36462 (N_36462,N_22870,N_20038);
or U36463 (N_36463,N_26251,N_22921);
xor U36464 (N_36464,N_29031,N_29975);
or U36465 (N_36465,N_28468,N_21202);
and U36466 (N_36466,N_24031,N_21413);
nor U36467 (N_36467,N_26011,N_28315);
xnor U36468 (N_36468,N_22044,N_24300);
or U36469 (N_36469,N_28817,N_21283);
and U36470 (N_36470,N_28372,N_28997);
and U36471 (N_36471,N_26998,N_24107);
nand U36472 (N_36472,N_20439,N_28022);
or U36473 (N_36473,N_22074,N_25205);
xor U36474 (N_36474,N_20323,N_29585);
nand U36475 (N_36475,N_25928,N_22720);
or U36476 (N_36476,N_20450,N_23125);
nor U36477 (N_36477,N_23386,N_28955);
or U36478 (N_36478,N_27266,N_26648);
nor U36479 (N_36479,N_28133,N_22164);
and U36480 (N_36480,N_22308,N_25523);
xor U36481 (N_36481,N_26403,N_21687);
nand U36482 (N_36482,N_26781,N_21591);
nor U36483 (N_36483,N_28876,N_20762);
nor U36484 (N_36484,N_25573,N_27278);
nor U36485 (N_36485,N_29069,N_27588);
nand U36486 (N_36486,N_24522,N_25348);
or U36487 (N_36487,N_28389,N_20712);
nand U36488 (N_36488,N_21312,N_24259);
nor U36489 (N_36489,N_21897,N_21184);
and U36490 (N_36490,N_24995,N_23670);
and U36491 (N_36491,N_28445,N_23977);
xor U36492 (N_36492,N_26537,N_25690);
nor U36493 (N_36493,N_22456,N_26159);
and U36494 (N_36494,N_21165,N_23169);
and U36495 (N_36495,N_22100,N_29572);
and U36496 (N_36496,N_27310,N_27791);
and U36497 (N_36497,N_21543,N_27078);
or U36498 (N_36498,N_23841,N_20425);
nor U36499 (N_36499,N_20874,N_26034);
nand U36500 (N_36500,N_22646,N_25726);
and U36501 (N_36501,N_26232,N_21603);
xnor U36502 (N_36502,N_26768,N_24562);
nand U36503 (N_36503,N_28134,N_27214);
and U36504 (N_36504,N_25821,N_21147);
nand U36505 (N_36505,N_23855,N_24856);
and U36506 (N_36506,N_29422,N_24020);
nor U36507 (N_36507,N_27162,N_25898);
and U36508 (N_36508,N_22291,N_28284);
and U36509 (N_36509,N_20696,N_23054);
nand U36510 (N_36510,N_25991,N_26916);
and U36511 (N_36511,N_29467,N_29685);
or U36512 (N_36512,N_29236,N_24055);
or U36513 (N_36513,N_27119,N_27601);
and U36514 (N_36514,N_29864,N_28854);
xnor U36515 (N_36515,N_25405,N_22593);
or U36516 (N_36516,N_23756,N_24649);
or U36517 (N_36517,N_29410,N_26225);
or U36518 (N_36518,N_24720,N_28065);
or U36519 (N_36519,N_26874,N_25676);
nor U36520 (N_36520,N_27541,N_27544);
nor U36521 (N_36521,N_26568,N_24483);
and U36522 (N_36522,N_25913,N_23293);
nand U36523 (N_36523,N_26380,N_25551);
nor U36524 (N_36524,N_23352,N_22533);
and U36525 (N_36525,N_27675,N_28936);
and U36526 (N_36526,N_26291,N_23682);
nor U36527 (N_36527,N_22709,N_29545);
or U36528 (N_36528,N_22285,N_28818);
nor U36529 (N_36529,N_21598,N_20440);
or U36530 (N_36530,N_26236,N_28611);
nor U36531 (N_36531,N_20904,N_29017);
nand U36532 (N_36532,N_22399,N_29647);
and U36533 (N_36533,N_23784,N_25091);
nand U36534 (N_36534,N_26012,N_24790);
nor U36535 (N_36535,N_24044,N_27814);
or U36536 (N_36536,N_29521,N_28777);
and U36537 (N_36537,N_22338,N_22743);
and U36538 (N_36538,N_27351,N_20421);
nand U36539 (N_36539,N_23767,N_29831);
and U36540 (N_36540,N_20642,N_29797);
and U36541 (N_36541,N_25848,N_22903);
nor U36542 (N_36542,N_27895,N_26514);
nand U36543 (N_36543,N_24101,N_24023);
and U36544 (N_36544,N_21544,N_20493);
nor U36545 (N_36545,N_23863,N_20122);
nand U36546 (N_36546,N_22464,N_20883);
or U36547 (N_36547,N_20824,N_20275);
or U36548 (N_36548,N_23594,N_23661);
nand U36549 (N_36549,N_23833,N_20589);
nand U36550 (N_36550,N_29235,N_22448);
and U36551 (N_36551,N_26462,N_21825);
and U36552 (N_36552,N_27776,N_22416);
nand U36553 (N_36553,N_24117,N_23179);
nand U36554 (N_36554,N_25127,N_23878);
or U36555 (N_36555,N_22217,N_26498);
nor U36556 (N_36556,N_24237,N_27844);
nand U36557 (N_36557,N_23863,N_27588);
and U36558 (N_36558,N_21109,N_25397);
and U36559 (N_36559,N_22012,N_27521);
nor U36560 (N_36560,N_21337,N_23175);
or U36561 (N_36561,N_22956,N_24945);
and U36562 (N_36562,N_27100,N_24575);
nand U36563 (N_36563,N_28859,N_27254);
nand U36564 (N_36564,N_28322,N_28819);
and U36565 (N_36565,N_20050,N_26132);
nor U36566 (N_36566,N_25204,N_23228);
nor U36567 (N_36567,N_21958,N_24041);
or U36568 (N_36568,N_20366,N_21319);
nand U36569 (N_36569,N_22196,N_27547);
or U36570 (N_36570,N_21683,N_25780);
or U36571 (N_36571,N_28166,N_25230);
or U36572 (N_36572,N_20813,N_27168);
nor U36573 (N_36573,N_28579,N_25964);
or U36574 (N_36574,N_23150,N_22715);
and U36575 (N_36575,N_22677,N_22537);
or U36576 (N_36576,N_22906,N_25544);
nor U36577 (N_36577,N_25554,N_20188);
and U36578 (N_36578,N_28795,N_25994);
or U36579 (N_36579,N_27247,N_23617);
nor U36580 (N_36580,N_23734,N_23231);
xor U36581 (N_36581,N_28647,N_24128);
nand U36582 (N_36582,N_26713,N_27524);
nand U36583 (N_36583,N_29342,N_23517);
or U36584 (N_36584,N_23612,N_23457);
nand U36585 (N_36585,N_23412,N_29351);
or U36586 (N_36586,N_20439,N_21251);
nor U36587 (N_36587,N_24553,N_27838);
nand U36588 (N_36588,N_25184,N_26010);
and U36589 (N_36589,N_24042,N_23360);
nor U36590 (N_36590,N_21730,N_24054);
nor U36591 (N_36591,N_25532,N_27523);
nor U36592 (N_36592,N_24462,N_24534);
nand U36593 (N_36593,N_23452,N_24699);
or U36594 (N_36594,N_21553,N_23247);
xor U36595 (N_36595,N_29925,N_25277);
nor U36596 (N_36596,N_26161,N_29670);
or U36597 (N_36597,N_25804,N_24483);
nor U36598 (N_36598,N_27643,N_21882);
and U36599 (N_36599,N_29526,N_28558);
nand U36600 (N_36600,N_23566,N_25500);
nand U36601 (N_36601,N_27181,N_23767);
or U36602 (N_36602,N_22608,N_28290);
nor U36603 (N_36603,N_27170,N_20636);
and U36604 (N_36604,N_22591,N_24914);
nand U36605 (N_36605,N_21952,N_20453);
nor U36606 (N_36606,N_21354,N_24426);
xor U36607 (N_36607,N_20214,N_27019);
or U36608 (N_36608,N_27126,N_29014);
and U36609 (N_36609,N_26131,N_29525);
nand U36610 (N_36610,N_26129,N_27825);
nand U36611 (N_36611,N_24272,N_23838);
nand U36612 (N_36612,N_24953,N_27822);
and U36613 (N_36613,N_28784,N_29420);
or U36614 (N_36614,N_27796,N_23668);
or U36615 (N_36615,N_28060,N_26838);
nor U36616 (N_36616,N_23465,N_24570);
nand U36617 (N_36617,N_28541,N_26117);
nor U36618 (N_36618,N_26466,N_29659);
nor U36619 (N_36619,N_22570,N_23737);
xor U36620 (N_36620,N_29679,N_22748);
nand U36621 (N_36621,N_26320,N_23447);
nor U36622 (N_36622,N_22363,N_24639);
nand U36623 (N_36623,N_22757,N_28635);
nor U36624 (N_36624,N_26294,N_29226);
nand U36625 (N_36625,N_24487,N_22396);
and U36626 (N_36626,N_23858,N_23672);
nand U36627 (N_36627,N_24040,N_20096);
or U36628 (N_36628,N_21439,N_25732);
nand U36629 (N_36629,N_26188,N_29469);
nand U36630 (N_36630,N_29397,N_23717);
or U36631 (N_36631,N_27088,N_26183);
nand U36632 (N_36632,N_23366,N_20660);
and U36633 (N_36633,N_20193,N_28583);
or U36634 (N_36634,N_25304,N_24888);
or U36635 (N_36635,N_22869,N_25898);
or U36636 (N_36636,N_23185,N_25282);
xor U36637 (N_36637,N_22941,N_25290);
xnor U36638 (N_36638,N_28124,N_22426);
xnor U36639 (N_36639,N_25358,N_21233);
nand U36640 (N_36640,N_29109,N_23255);
and U36641 (N_36641,N_26601,N_28161);
xor U36642 (N_36642,N_21660,N_24905);
xor U36643 (N_36643,N_26285,N_24838);
and U36644 (N_36644,N_28130,N_26423);
nor U36645 (N_36645,N_29130,N_23850);
nand U36646 (N_36646,N_26022,N_25275);
and U36647 (N_36647,N_21777,N_26478);
and U36648 (N_36648,N_24313,N_23279);
nor U36649 (N_36649,N_23490,N_21635);
nor U36650 (N_36650,N_26225,N_22229);
nand U36651 (N_36651,N_26217,N_25707);
nor U36652 (N_36652,N_26614,N_20893);
and U36653 (N_36653,N_21731,N_23023);
nor U36654 (N_36654,N_27899,N_24159);
xor U36655 (N_36655,N_29713,N_28695);
nor U36656 (N_36656,N_29417,N_23864);
and U36657 (N_36657,N_29620,N_26777);
xnor U36658 (N_36658,N_25130,N_20035);
nor U36659 (N_36659,N_21166,N_27456);
and U36660 (N_36660,N_28108,N_21551);
nor U36661 (N_36661,N_23051,N_20138);
or U36662 (N_36662,N_26348,N_20647);
nor U36663 (N_36663,N_21044,N_23776);
nand U36664 (N_36664,N_21762,N_26209);
or U36665 (N_36665,N_25801,N_22158);
nor U36666 (N_36666,N_20118,N_21917);
or U36667 (N_36667,N_20498,N_20999);
or U36668 (N_36668,N_25200,N_29632);
nand U36669 (N_36669,N_24732,N_26550);
nand U36670 (N_36670,N_21272,N_28582);
or U36671 (N_36671,N_24829,N_29219);
nand U36672 (N_36672,N_28201,N_28697);
nand U36673 (N_36673,N_23415,N_21480);
and U36674 (N_36674,N_26899,N_22001);
nor U36675 (N_36675,N_28833,N_26420);
and U36676 (N_36676,N_25421,N_25635);
and U36677 (N_36677,N_24856,N_28291);
or U36678 (N_36678,N_26911,N_22374);
nand U36679 (N_36679,N_25695,N_24429);
xnor U36680 (N_36680,N_29782,N_24540);
and U36681 (N_36681,N_22041,N_24619);
nor U36682 (N_36682,N_21419,N_23434);
and U36683 (N_36683,N_26812,N_27183);
and U36684 (N_36684,N_27811,N_20487);
nor U36685 (N_36685,N_26473,N_23504);
and U36686 (N_36686,N_25107,N_29883);
or U36687 (N_36687,N_28451,N_21872);
nand U36688 (N_36688,N_29169,N_20209);
nor U36689 (N_36689,N_20293,N_24435);
nand U36690 (N_36690,N_28471,N_23303);
nand U36691 (N_36691,N_28164,N_22822);
nor U36692 (N_36692,N_27023,N_24045);
nand U36693 (N_36693,N_22996,N_28104);
nand U36694 (N_36694,N_24437,N_24441);
or U36695 (N_36695,N_21199,N_25554);
and U36696 (N_36696,N_29247,N_28445);
nand U36697 (N_36697,N_26071,N_24552);
or U36698 (N_36698,N_24561,N_22512);
and U36699 (N_36699,N_29540,N_21483);
nor U36700 (N_36700,N_28468,N_22357);
xnor U36701 (N_36701,N_29130,N_26795);
or U36702 (N_36702,N_20654,N_27059);
nand U36703 (N_36703,N_27842,N_25215);
nand U36704 (N_36704,N_26454,N_27260);
xor U36705 (N_36705,N_23254,N_24644);
and U36706 (N_36706,N_21124,N_26889);
or U36707 (N_36707,N_24687,N_27316);
nor U36708 (N_36708,N_25427,N_24143);
nor U36709 (N_36709,N_20206,N_26363);
or U36710 (N_36710,N_25745,N_27632);
nor U36711 (N_36711,N_20568,N_25058);
nand U36712 (N_36712,N_28807,N_27477);
and U36713 (N_36713,N_22791,N_27467);
or U36714 (N_36714,N_26421,N_25944);
or U36715 (N_36715,N_26818,N_25243);
xor U36716 (N_36716,N_21657,N_25061);
xnor U36717 (N_36717,N_22087,N_26199);
or U36718 (N_36718,N_23289,N_24235);
xnor U36719 (N_36719,N_20738,N_28906);
nor U36720 (N_36720,N_22310,N_24860);
or U36721 (N_36721,N_23109,N_26784);
or U36722 (N_36722,N_29561,N_22942);
or U36723 (N_36723,N_26894,N_24019);
nor U36724 (N_36724,N_23280,N_21181);
nand U36725 (N_36725,N_25099,N_23030);
nand U36726 (N_36726,N_20782,N_28952);
and U36727 (N_36727,N_23652,N_21957);
or U36728 (N_36728,N_20006,N_24409);
nand U36729 (N_36729,N_25037,N_20380);
or U36730 (N_36730,N_22790,N_23468);
or U36731 (N_36731,N_23665,N_24985);
and U36732 (N_36732,N_22775,N_28305);
or U36733 (N_36733,N_24381,N_22238);
or U36734 (N_36734,N_28203,N_27400);
nand U36735 (N_36735,N_20639,N_22896);
nor U36736 (N_36736,N_27288,N_28032);
and U36737 (N_36737,N_22276,N_28968);
xnor U36738 (N_36738,N_29642,N_22880);
or U36739 (N_36739,N_26540,N_20774);
and U36740 (N_36740,N_25832,N_25948);
and U36741 (N_36741,N_27571,N_29789);
nand U36742 (N_36742,N_20078,N_26952);
nor U36743 (N_36743,N_22922,N_23882);
nor U36744 (N_36744,N_24713,N_24116);
or U36745 (N_36745,N_23129,N_28625);
xor U36746 (N_36746,N_21804,N_20873);
nand U36747 (N_36747,N_27015,N_26687);
nor U36748 (N_36748,N_28357,N_27071);
nor U36749 (N_36749,N_21785,N_22084);
nor U36750 (N_36750,N_25065,N_27394);
xor U36751 (N_36751,N_20268,N_21645);
or U36752 (N_36752,N_29144,N_25998);
nand U36753 (N_36753,N_22201,N_26271);
and U36754 (N_36754,N_21398,N_20940);
nand U36755 (N_36755,N_24673,N_24772);
nand U36756 (N_36756,N_20912,N_28610);
and U36757 (N_36757,N_22284,N_23349);
and U36758 (N_36758,N_20322,N_21776);
or U36759 (N_36759,N_24626,N_20814);
nand U36760 (N_36760,N_29957,N_20868);
or U36761 (N_36761,N_21245,N_26337);
and U36762 (N_36762,N_25843,N_29484);
and U36763 (N_36763,N_29824,N_28982);
xnor U36764 (N_36764,N_24869,N_21847);
xor U36765 (N_36765,N_29625,N_28083);
nor U36766 (N_36766,N_23831,N_23884);
nand U36767 (N_36767,N_20205,N_20933);
nand U36768 (N_36768,N_25566,N_28189);
and U36769 (N_36769,N_24886,N_29820);
nand U36770 (N_36770,N_29415,N_25545);
nand U36771 (N_36771,N_21807,N_20115);
nand U36772 (N_36772,N_22029,N_22378);
nor U36773 (N_36773,N_29075,N_24914);
nand U36774 (N_36774,N_23880,N_29326);
and U36775 (N_36775,N_25640,N_20328);
xnor U36776 (N_36776,N_20627,N_22987);
or U36777 (N_36777,N_25222,N_23050);
nand U36778 (N_36778,N_28081,N_21077);
nand U36779 (N_36779,N_20934,N_21748);
nand U36780 (N_36780,N_21194,N_21721);
nor U36781 (N_36781,N_26429,N_24934);
nand U36782 (N_36782,N_22607,N_22289);
and U36783 (N_36783,N_22641,N_25891);
nor U36784 (N_36784,N_24339,N_21019);
nor U36785 (N_36785,N_21981,N_26006);
nor U36786 (N_36786,N_26384,N_22838);
or U36787 (N_36787,N_21009,N_27786);
nand U36788 (N_36788,N_27299,N_22589);
and U36789 (N_36789,N_26295,N_26270);
xor U36790 (N_36790,N_27355,N_24818);
or U36791 (N_36791,N_21638,N_23512);
or U36792 (N_36792,N_21626,N_20087);
and U36793 (N_36793,N_28963,N_27254);
nand U36794 (N_36794,N_21038,N_26862);
nand U36795 (N_36795,N_21558,N_27084);
and U36796 (N_36796,N_21031,N_27793);
and U36797 (N_36797,N_21402,N_20520);
nor U36798 (N_36798,N_26519,N_24928);
nor U36799 (N_36799,N_20688,N_27875);
nor U36800 (N_36800,N_29340,N_20286);
or U36801 (N_36801,N_26053,N_22523);
xor U36802 (N_36802,N_23047,N_22095);
nor U36803 (N_36803,N_25041,N_23706);
nor U36804 (N_36804,N_26075,N_21040);
nor U36805 (N_36805,N_23392,N_20885);
xnor U36806 (N_36806,N_20767,N_27442);
nand U36807 (N_36807,N_27630,N_25501);
nand U36808 (N_36808,N_20066,N_28367);
or U36809 (N_36809,N_22224,N_22936);
and U36810 (N_36810,N_23761,N_25060);
or U36811 (N_36811,N_21053,N_29605);
nand U36812 (N_36812,N_28392,N_24607);
or U36813 (N_36813,N_24105,N_24158);
nor U36814 (N_36814,N_25871,N_23185);
nor U36815 (N_36815,N_29036,N_29284);
nand U36816 (N_36816,N_26705,N_23921);
or U36817 (N_36817,N_26084,N_21584);
xnor U36818 (N_36818,N_20705,N_25285);
and U36819 (N_36819,N_27638,N_22362);
nor U36820 (N_36820,N_21287,N_23930);
nand U36821 (N_36821,N_22965,N_24710);
or U36822 (N_36822,N_28619,N_29952);
and U36823 (N_36823,N_20485,N_24867);
and U36824 (N_36824,N_26676,N_23690);
nand U36825 (N_36825,N_20994,N_23901);
and U36826 (N_36826,N_27155,N_27241);
and U36827 (N_36827,N_29322,N_25203);
xnor U36828 (N_36828,N_27522,N_26265);
or U36829 (N_36829,N_29366,N_20110);
and U36830 (N_36830,N_24864,N_21082);
nor U36831 (N_36831,N_23375,N_24082);
nand U36832 (N_36832,N_20848,N_26542);
and U36833 (N_36833,N_20331,N_29181);
or U36834 (N_36834,N_22847,N_27147);
nand U36835 (N_36835,N_23008,N_23986);
nor U36836 (N_36836,N_24187,N_24480);
or U36837 (N_36837,N_26094,N_20929);
nand U36838 (N_36838,N_26065,N_21159);
nand U36839 (N_36839,N_26337,N_25258);
nor U36840 (N_36840,N_22405,N_23419);
and U36841 (N_36841,N_28735,N_26160);
or U36842 (N_36842,N_20608,N_24723);
nand U36843 (N_36843,N_22624,N_24396);
or U36844 (N_36844,N_21761,N_22743);
or U36845 (N_36845,N_29219,N_22282);
and U36846 (N_36846,N_26181,N_21369);
xnor U36847 (N_36847,N_20282,N_24685);
or U36848 (N_36848,N_29814,N_21595);
and U36849 (N_36849,N_24612,N_20947);
or U36850 (N_36850,N_24803,N_24876);
and U36851 (N_36851,N_23051,N_20746);
xor U36852 (N_36852,N_26405,N_25614);
and U36853 (N_36853,N_24108,N_21768);
nor U36854 (N_36854,N_22809,N_22465);
nand U36855 (N_36855,N_22635,N_23565);
or U36856 (N_36856,N_27413,N_23374);
and U36857 (N_36857,N_22788,N_23156);
or U36858 (N_36858,N_27014,N_25061);
nand U36859 (N_36859,N_21273,N_22100);
or U36860 (N_36860,N_27393,N_21529);
or U36861 (N_36861,N_21195,N_28267);
nor U36862 (N_36862,N_23541,N_20892);
and U36863 (N_36863,N_23287,N_28041);
nor U36864 (N_36864,N_28150,N_24303);
or U36865 (N_36865,N_23024,N_26834);
nor U36866 (N_36866,N_25156,N_28610);
nand U36867 (N_36867,N_23505,N_24475);
or U36868 (N_36868,N_25811,N_24175);
nand U36869 (N_36869,N_26443,N_27868);
nor U36870 (N_36870,N_21808,N_28596);
nor U36871 (N_36871,N_20956,N_22308);
nand U36872 (N_36872,N_26665,N_27112);
or U36873 (N_36873,N_21418,N_24706);
nand U36874 (N_36874,N_25345,N_29678);
and U36875 (N_36875,N_26377,N_26877);
nor U36876 (N_36876,N_29447,N_23127);
or U36877 (N_36877,N_21852,N_20105);
or U36878 (N_36878,N_26883,N_26783);
and U36879 (N_36879,N_26441,N_23338);
and U36880 (N_36880,N_29537,N_28313);
and U36881 (N_36881,N_26427,N_22207);
xnor U36882 (N_36882,N_22888,N_28413);
and U36883 (N_36883,N_25402,N_24997);
xor U36884 (N_36884,N_21705,N_21386);
and U36885 (N_36885,N_21278,N_25901);
nor U36886 (N_36886,N_20789,N_26876);
xor U36887 (N_36887,N_22269,N_24680);
or U36888 (N_36888,N_22810,N_21609);
nand U36889 (N_36889,N_22156,N_26991);
or U36890 (N_36890,N_28050,N_20184);
nand U36891 (N_36891,N_22903,N_27508);
or U36892 (N_36892,N_22668,N_27691);
nor U36893 (N_36893,N_25447,N_26479);
nand U36894 (N_36894,N_26252,N_25820);
or U36895 (N_36895,N_27289,N_26154);
nor U36896 (N_36896,N_28858,N_28173);
xnor U36897 (N_36897,N_21728,N_20826);
nor U36898 (N_36898,N_24587,N_27129);
or U36899 (N_36899,N_28649,N_21816);
or U36900 (N_36900,N_22824,N_27737);
nand U36901 (N_36901,N_26607,N_26707);
nor U36902 (N_36902,N_28501,N_25875);
or U36903 (N_36903,N_29709,N_21357);
nand U36904 (N_36904,N_20104,N_20612);
nor U36905 (N_36905,N_20019,N_23252);
or U36906 (N_36906,N_23097,N_20299);
and U36907 (N_36907,N_29375,N_26829);
nand U36908 (N_36908,N_29654,N_23495);
nor U36909 (N_36909,N_23568,N_24796);
nor U36910 (N_36910,N_27571,N_29092);
nor U36911 (N_36911,N_26791,N_22337);
and U36912 (N_36912,N_26918,N_25412);
or U36913 (N_36913,N_27383,N_29677);
and U36914 (N_36914,N_23329,N_28889);
nand U36915 (N_36915,N_27414,N_29189);
nand U36916 (N_36916,N_20159,N_25673);
or U36917 (N_36917,N_22576,N_29492);
nand U36918 (N_36918,N_27661,N_20872);
nand U36919 (N_36919,N_22316,N_29383);
or U36920 (N_36920,N_22362,N_29597);
nor U36921 (N_36921,N_29618,N_26607);
or U36922 (N_36922,N_24160,N_21739);
nand U36923 (N_36923,N_26767,N_23093);
or U36924 (N_36924,N_28060,N_24037);
nor U36925 (N_36925,N_28411,N_28837);
nor U36926 (N_36926,N_29361,N_22226);
nand U36927 (N_36927,N_29176,N_23343);
nand U36928 (N_36928,N_26764,N_28245);
nor U36929 (N_36929,N_21546,N_22165);
nor U36930 (N_36930,N_28614,N_26066);
or U36931 (N_36931,N_25418,N_25681);
or U36932 (N_36932,N_26649,N_28569);
nor U36933 (N_36933,N_21935,N_20384);
or U36934 (N_36934,N_21809,N_27920);
and U36935 (N_36935,N_23922,N_24557);
and U36936 (N_36936,N_23814,N_28976);
nand U36937 (N_36937,N_28100,N_29690);
or U36938 (N_36938,N_24695,N_21341);
nand U36939 (N_36939,N_20501,N_27596);
and U36940 (N_36940,N_29887,N_28613);
or U36941 (N_36941,N_28709,N_22613);
or U36942 (N_36942,N_25308,N_26185);
nor U36943 (N_36943,N_21531,N_21898);
and U36944 (N_36944,N_29349,N_26005);
nand U36945 (N_36945,N_20092,N_21012);
and U36946 (N_36946,N_28032,N_22278);
or U36947 (N_36947,N_29384,N_21435);
or U36948 (N_36948,N_28801,N_22561);
and U36949 (N_36949,N_22919,N_28719);
xnor U36950 (N_36950,N_25563,N_21216);
nand U36951 (N_36951,N_23238,N_28045);
and U36952 (N_36952,N_28972,N_23149);
nand U36953 (N_36953,N_25091,N_29477);
and U36954 (N_36954,N_22467,N_28681);
nand U36955 (N_36955,N_20150,N_24999);
or U36956 (N_36956,N_25432,N_26524);
xor U36957 (N_36957,N_23347,N_28743);
nor U36958 (N_36958,N_20082,N_24706);
nor U36959 (N_36959,N_25030,N_20154);
or U36960 (N_36960,N_25883,N_29032);
and U36961 (N_36961,N_24691,N_24403);
and U36962 (N_36962,N_21263,N_28323);
nor U36963 (N_36963,N_29486,N_27281);
xor U36964 (N_36964,N_24846,N_29902);
and U36965 (N_36965,N_20219,N_26701);
and U36966 (N_36966,N_26454,N_22521);
nor U36967 (N_36967,N_29258,N_27635);
nor U36968 (N_36968,N_25333,N_24290);
xor U36969 (N_36969,N_26476,N_27272);
or U36970 (N_36970,N_26776,N_27578);
nor U36971 (N_36971,N_28928,N_20282);
and U36972 (N_36972,N_26954,N_24077);
or U36973 (N_36973,N_28887,N_24406);
xor U36974 (N_36974,N_25522,N_24260);
xor U36975 (N_36975,N_29907,N_29492);
nor U36976 (N_36976,N_20997,N_28509);
xor U36977 (N_36977,N_28338,N_29024);
xnor U36978 (N_36978,N_21008,N_26138);
nor U36979 (N_36979,N_27707,N_21805);
or U36980 (N_36980,N_25211,N_23276);
or U36981 (N_36981,N_21224,N_28427);
nand U36982 (N_36982,N_20809,N_28108);
and U36983 (N_36983,N_20241,N_21700);
and U36984 (N_36984,N_25854,N_25097);
and U36985 (N_36985,N_24742,N_25063);
nand U36986 (N_36986,N_21052,N_24068);
nand U36987 (N_36987,N_23600,N_26767);
xor U36988 (N_36988,N_21983,N_28042);
and U36989 (N_36989,N_21917,N_20812);
and U36990 (N_36990,N_28379,N_26977);
nand U36991 (N_36991,N_22399,N_25146);
and U36992 (N_36992,N_21606,N_23594);
or U36993 (N_36993,N_28440,N_22020);
xnor U36994 (N_36994,N_26647,N_25991);
and U36995 (N_36995,N_23623,N_28986);
nor U36996 (N_36996,N_26791,N_23050);
nand U36997 (N_36997,N_29639,N_22355);
xor U36998 (N_36998,N_26122,N_21636);
or U36999 (N_36999,N_29276,N_21194);
xnor U37000 (N_37000,N_20442,N_22647);
nand U37001 (N_37001,N_25331,N_23283);
or U37002 (N_37002,N_28169,N_28516);
or U37003 (N_37003,N_28954,N_26050);
nor U37004 (N_37004,N_27244,N_28543);
nor U37005 (N_37005,N_29026,N_21691);
nor U37006 (N_37006,N_23564,N_23835);
and U37007 (N_37007,N_27122,N_20474);
nand U37008 (N_37008,N_21924,N_26067);
and U37009 (N_37009,N_29519,N_21855);
or U37010 (N_37010,N_27104,N_22649);
nand U37011 (N_37011,N_24873,N_22659);
nor U37012 (N_37012,N_25878,N_22023);
nor U37013 (N_37013,N_22335,N_27014);
or U37014 (N_37014,N_24773,N_24215);
nand U37015 (N_37015,N_20649,N_22773);
nor U37016 (N_37016,N_23968,N_22037);
nand U37017 (N_37017,N_29990,N_27113);
nand U37018 (N_37018,N_22164,N_29844);
or U37019 (N_37019,N_29776,N_25963);
xnor U37020 (N_37020,N_27949,N_20546);
nand U37021 (N_37021,N_23787,N_25059);
and U37022 (N_37022,N_21595,N_21839);
nor U37023 (N_37023,N_21530,N_27803);
and U37024 (N_37024,N_23272,N_20994);
and U37025 (N_37025,N_24971,N_22793);
nand U37026 (N_37026,N_24150,N_26712);
or U37027 (N_37027,N_24232,N_24399);
nand U37028 (N_37028,N_22218,N_21005);
nor U37029 (N_37029,N_24165,N_26883);
and U37030 (N_37030,N_28531,N_25386);
and U37031 (N_37031,N_27441,N_29423);
and U37032 (N_37032,N_28744,N_22791);
nand U37033 (N_37033,N_21785,N_25687);
and U37034 (N_37034,N_25301,N_23325);
nor U37035 (N_37035,N_24212,N_25287);
nor U37036 (N_37036,N_27537,N_25001);
nand U37037 (N_37037,N_27428,N_22948);
and U37038 (N_37038,N_29769,N_24332);
nor U37039 (N_37039,N_20307,N_21782);
xnor U37040 (N_37040,N_27508,N_21099);
nand U37041 (N_37041,N_23856,N_20431);
nand U37042 (N_37042,N_25053,N_20173);
xnor U37043 (N_37043,N_22563,N_27150);
or U37044 (N_37044,N_21157,N_21933);
nor U37045 (N_37045,N_28539,N_27573);
nand U37046 (N_37046,N_21244,N_23450);
and U37047 (N_37047,N_29187,N_25601);
nor U37048 (N_37048,N_23102,N_27044);
nand U37049 (N_37049,N_28443,N_27912);
nand U37050 (N_37050,N_29493,N_24965);
xnor U37051 (N_37051,N_22361,N_22516);
nor U37052 (N_37052,N_28758,N_29039);
nor U37053 (N_37053,N_25166,N_28062);
nor U37054 (N_37054,N_20195,N_23913);
or U37055 (N_37055,N_27108,N_27280);
or U37056 (N_37056,N_22645,N_24643);
and U37057 (N_37057,N_23730,N_21119);
xnor U37058 (N_37058,N_24444,N_21435);
and U37059 (N_37059,N_28050,N_21279);
or U37060 (N_37060,N_20515,N_22628);
nor U37061 (N_37061,N_22676,N_23924);
nor U37062 (N_37062,N_20714,N_29024);
and U37063 (N_37063,N_20246,N_25872);
nand U37064 (N_37064,N_22472,N_23382);
xor U37065 (N_37065,N_20446,N_28468);
or U37066 (N_37066,N_23218,N_21914);
xor U37067 (N_37067,N_20399,N_21928);
nor U37068 (N_37068,N_21378,N_26417);
and U37069 (N_37069,N_20859,N_28844);
nand U37070 (N_37070,N_21738,N_25148);
xnor U37071 (N_37071,N_20889,N_20414);
and U37072 (N_37072,N_21654,N_29719);
nand U37073 (N_37073,N_20738,N_20532);
or U37074 (N_37074,N_26230,N_22517);
and U37075 (N_37075,N_28970,N_25856);
xor U37076 (N_37076,N_25631,N_28445);
nand U37077 (N_37077,N_25554,N_28560);
nor U37078 (N_37078,N_20433,N_27537);
nor U37079 (N_37079,N_20982,N_27581);
or U37080 (N_37080,N_23916,N_20315);
or U37081 (N_37081,N_23389,N_29847);
nor U37082 (N_37082,N_25559,N_21980);
nand U37083 (N_37083,N_21237,N_24397);
and U37084 (N_37084,N_22596,N_27845);
and U37085 (N_37085,N_25191,N_28442);
and U37086 (N_37086,N_24822,N_26534);
nor U37087 (N_37087,N_27731,N_26887);
nand U37088 (N_37088,N_21998,N_26696);
xor U37089 (N_37089,N_29040,N_20533);
nand U37090 (N_37090,N_21068,N_24824);
nor U37091 (N_37091,N_24795,N_24013);
nor U37092 (N_37092,N_27313,N_24215);
and U37093 (N_37093,N_23998,N_25594);
nand U37094 (N_37094,N_22189,N_23089);
nor U37095 (N_37095,N_24801,N_26796);
nand U37096 (N_37096,N_21450,N_26468);
nand U37097 (N_37097,N_26970,N_28908);
xnor U37098 (N_37098,N_25380,N_22172);
and U37099 (N_37099,N_26079,N_29958);
or U37100 (N_37100,N_29604,N_24610);
xor U37101 (N_37101,N_22817,N_29466);
xnor U37102 (N_37102,N_24334,N_20015);
and U37103 (N_37103,N_23385,N_20401);
and U37104 (N_37104,N_26777,N_23498);
nor U37105 (N_37105,N_26484,N_27211);
nand U37106 (N_37106,N_20496,N_26912);
nor U37107 (N_37107,N_29153,N_25760);
and U37108 (N_37108,N_26396,N_28035);
or U37109 (N_37109,N_28108,N_29962);
nand U37110 (N_37110,N_21236,N_26811);
and U37111 (N_37111,N_24834,N_22388);
or U37112 (N_37112,N_27010,N_29955);
and U37113 (N_37113,N_27150,N_25284);
nand U37114 (N_37114,N_28339,N_21849);
nor U37115 (N_37115,N_25479,N_26718);
nand U37116 (N_37116,N_29165,N_23610);
and U37117 (N_37117,N_23508,N_23222);
or U37118 (N_37118,N_22393,N_29756);
nand U37119 (N_37119,N_26506,N_25731);
and U37120 (N_37120,N_28320,N_21048);
nor U37121 (N_37121,N_22005,N_26361);
and U37122 (N_37122,N_28306,N_27350);
nand U37123 (N_37123,N_24885,N_20088);
nand U37124 (N_37124,N_20797,N_29910);
nand U37125 (N_37125,N_21604,N_28137);
nand U37126 (N_37126,N_24697,N_20182);
or U37127 (N_37127,N_21711,N_25688);
nor U37128 (N_37128,N_20298,N_23928);
nand U37129 (N_37129,N_25392,N_22060);
or U37130 (N_37130,N_26437,N_23483);
nor U37131 (N_37131,N_21319,N_21227);
and U37132 (N_37132,N_21891,N_28167);
nand U37133 (N_37133,N_26117,N_29689);
or U37134 (N_37134,N_23763,N_29582);
nor U37135 (N_37135,N_28110,N_23764);
or U37136 (N_37136,N_25025,N_25164);
or U37137 (N_37137,N_21542,N_28032);
nand U37138 (N_37138,N_27207,N_27652);
nor U37139 (N_37139,N_24881,N_26883);
nor U37140 (N_37140,N_22300,N_25292);
nor U37141 (N_37141,N_26570,N_28834);
nor U37142 (N_37142,N_22179,N_21822);
nor U37143 (N_37143,N_23572,N_24308);
nand U37144 (N_37144,N_20020,N_21563);
nor U37145 (N_37145,N_28423,N_29183);
nand U37146 (N_37146,N_28326,N_28884);
or U37147 (N_37147,N_26511,N_28036);
and U37148 (N_37148,N_25700,N_23347);
nor U37149 (N_37149,N_26587,N_24831);
nor U37150 (N_37150,N_20216,N_24369);
nand U37151 (N_37151,N_26654,N_21447);
or U37152 (N_37152,N_24061,N_22165);
and U37153 (N_37153,N_25102,N_22069);
or U37154 (N_37154,N_24473,N_25222);
xor U37155 (N_37155,N_25913,N_26594);
or U37156 (N_37156,N_23783,N_27072);
nor U37157 (N_37157,N_26299,N_25051);
or U37158 (N_37158,N_28947,N_21569);
nor U37159 (N_37159,N_29524,N_29132);
or U37160 (N_37160,N_23831,N_29569);
nor U37161 (N_37161,N_28391,N_26830);
nand U37162 (N_37162,N_26171,N_29587);
and U37163 (N_37163,N_23753,N_29568);
and U37164 (N_37164,N_23479,N_28444);
or U37165 (N_37165,N_21457,N_23015);
nor U37166 (N_37166,N_22419,N_23398);
or U37167 (N_37167,N_21041,N_23058);
or U37168 (N_37168,N_23781,N_29961);
nor U37169 (N_37169,N_25902,N_26489);
and U37170 (N_37170,N_29716,N_21485);
nor U37171 (N_37171,N_24143,N_27246);
and U37172 (N_37172,N_23147,N_21431);
nor U37173 (N_37173,N_21489,N_28745);
and U37174 (N_37174,N_26285,N_20269);
and U37175 (N_37175,N_29515,N_22062);
and U37176 (N_37176,N_27562,N_20208);
xor U37177 (N_37177,N_22114,N_20314);
xnor U37178 (N_37178,N_28337,N_23967);
and U37179 (N_37179,N_23504,N_27768);
or U37180 (N_37180,N_25125,N_23387);
or U37181 (N_37181,N_25395,N_23134);
nand U37182 (N_37182,N_27831,N_22254);
nand U37183 (N_37183,N_24951,N_23749);
or U37184 (N_37184,N_25993,N_23683);
and U37185 (N_37185,N_25194,N_29993);
or U37186 (N_37186,N_22170,N_29520);
nand U37187 (N_37187,N_21000,N_21312);
or U37188 (N_37188,N_29470,N_23506);
or U37189 (N_37189,N_21289,N_20096);
or U37190 (N_37190,N_27306,N_25855);
and U37191 (N_37191,N_24772,N_27582);
or U37192 (N_37192,N_29746,N_23665);
nand U37193 (N_37193,N_26540,N_28238);
nand U37194 (N_37194,N_20874,N_23883);
nor U37195 (N_37195,N_20368,N_21872);
and U37196 (N_37196,N_20787,N_20655);
or U37197 (N_37197,N_25587,N_27000);
and U37198 (N_37198,N_29293,N_28359);
nand U37199 (N_37199,N_28470,N_25609);
and U37200 (N_37200,N_20935,N_27557);
nor U37201 (N_37201,N_28230,N_29773);
xor U37202 (N_37202,N_29956,N_29949);
xor U37203 (N_37203,N_27466,N_25933);
nand U37204 (N_37204,N_22670,N_29830);
and U37205 (N_37205,N_29712,N_21292);
nor U37206 (N_37206,N_29274,N_28751);
xnor U37207 (N_37207,N_21572,N_21161);
or U37208 (N_37208,N_20502,N_23853);
nand U37209 (N_37209,N_21234,N_28186);
nand U37210 (N_37210,N_20757,N_20096);
and U37211 (N_37211,N_29219,N_24892);
nor U37212 (N_37212,N_26286,N_25156);
nor U37213 (N_37213,N_26053,N_28677);
and U37214 (N_37214,N_29677,N_29567);
xnor U37215 (N_37215,N_24934,N_28460);
nand U37216 (N_37216,N_29469,N_21790);
and U37217 (N_37217,N_23372,N_22219);
and U37218 (N_37218,N_20519,N_27302);
xnor U37219 (N_37219,N_23764,N_25507);
and U37220 (N_37220,N_29855,N_20280);
and U37221 (N_37221,N_24852,N_28042);
nand U37222 (N_37222,N_21923,N_23334);
nand U37223 (N_37223,N_23996,N_21393);
nand U37224 (N_37224,N_20192,N_25293);
nand U37225 (N_37225,N_23616,N_29952);
nor U37226 (N_37226,N_23387,N_24713);
nor U37227 (N_37227,N_29138,N_28222);
and U37228 (N_37228,N_26844,N_23779);
or U37229 (N_37229,N_29356,N_25577);
nand U37230 (N_37230,N_27218,N_23130);
or U37231 (N_37231,N_29587,N_27278);
or U37232 (N_37232,N_27342,N_27783);
or U37233 (N_37233,N_21619,N_25735);
nand U37234 (N_37234,N_21336,N_27449);
and U37235 (N_37235,N_27512,N_25929);
nor U37236 (N_37236,N_24902,N_23258);
nor U37237 (N_37237,N_22016,N_22747);
and U37238 (N_37238,N_23312,N_26351);
and U37239 (N_37239,N_27291,N_21482);
or U37240 (N_37240,N_29158,N_22423);
xor U37241 (N_37241,N_22149,N_26644);
or U37242 (N_37242,N_20645,N_24762);
xnor U37243 (N_37243,N_29682,N_22393);
xnor U37244 (N_37244,N_28363,N_25115);
or U37245 (N_37245,N_28176,N_28793);
nand U37246 (N_37246,N_22674,N_20819);
and U37247 (N_37247,N_20177,N_29438);
xnor U37248 (N_37248,N_25118,N_22883);
or U37249 (N_37249,N_24386,N_22461);
nand U37250 (N_37250,N_29420,N_21307);
and U37251 (N_37251,N_26608,N_29745);
nand U37252 (N_37252,N_24274,N_20861);
and U37253 (N_37253,N_26390,N_22801);
nand U37254 (N_37254,N_28674,N_21355);
nand U37255 (N_37255,N_21459,N_20087);
nand U37256 (N_37256,N_23856,N_22090);
or U37257 (N_37257,N_20861,N_20834);
nor U37258 (N_37258,N_26048,N_29986);
nand U37259 (N_37259,N_27861,N_27605);
nor U37260 (N_37260,N_25146,N_28385);
nand U37261 (N_37261,N_20119,N_20436);
and U37262 (N_37262,N_21391,N_23024);
and U37263 (N_37263,N_20377,N_20577);
nor U37264 (N_37264,N_29650,N_20753);
nand U37265 (N_37265,N_23621,N_20035);
or U37266 (N_37266,N_24110,N_29268);
and U37267 (N_37267,N_25244,N_22184);
and U37268 (N_37268,N_24571,N_21737);
nand U37269 (N_37269,N_21900,N_21459);
or U37270 (N_37270,N_20671,N_22080);
or U37271 (N_37271,N_23200,N_26638);
nand U37272 (N_37272,N_23613,N_22555);
nand U37273 (N_37273,N_24754,N_24822);
or U37274 (N_37274,N_25998,N_20339);
and U37275 (N_37275,N_26274,N_21268);
nand U37276 (N_37276,N_21533,N_28604);
nand U37277 (N_37277,N_23326,N_28298);
nor U37278 (N_37278,N_26536,N_25890);
nand U37279 (N_37279,N_26898,N_24416);
xnor U37280 (N_37280,N_29194,N_20749);
nand U37281 (N_37281,N_23597,N_26211);
xnor U37282 (N_37282,N_29302,N_21535);
nand U37283 (N_37283,N_24187,N_23661);
nor U37284 (N_37284,N_20105,N_23415);
nand U37285 (N_37285,N_29423,N_27513);
nand U37286 (N_37286,N_22194,N_29352);
nor U37287 (N_37287,N_21549,N_24058);
or U37288 (N_37288,N_28083,N_25615);
nor U37289 (N_37289,N_25944,N_23019);
or U37290 (N_37290,N_28217,N_28247);
nor U37291 (N_37291,N_20373,N_24466);
xor U37292 (N_37292,N_23082,N_29734);
or U37293 (N_37293,N_21708,N_20126);
nor U37294 (N_37294,N_28463,N_27394);
nand U37295 (N_37295,N_27425,N_23735);
xor U37296 (N_37296,N_29948,N_26223);
nand U37297 (N_37297,N_24155,N_21835);
nor U37298 (N_37298,N_24691,N_28270);
xor U37299 (N_37299,N_28251,N_26667);
nor U37300 (N_37300,N_24628,N_25756);
nor U37301 (N_37301,N_24433,N_20194);
nor U37302 (N_37302,N_22326,N_26337);
and U37303 (N_37303,N_23697,N_21909);
or U37304 (N_37304,N_22479,N_22796);
or U37305 (N_37305,N_20534,N_25966);
nor U37306 (N_37306,N_26432,N_22220);
nand U37307 (N_37307,N_22926,N_22703);
or U37308 (N_37308,N_23493,N_26732);
nand U37309 (N_37309,N_20085,N_21548);
or U37310 (N_37310,N_21293,N_27558);
nor U37311 (N_37311,N_26916,N_29063);
or U37312 (N_37312,N_23276,N_20570);
nor U37313 (N_37313,N_25811,N_26536);
and U37314 (N_37314,N_22758,N_28413);
or U37315 (N_37315,N_22026,N_25619);
nand U37316 (N_37316,N_20098,N_24395);
xor U37317 (N_37317,N_29407,N_25892);
xor U37318 (N_37318,N_24843,N_27937);
or U37319 (N_37319,N_26827,N_23955);
nor U37320 (N_37320,N_22196,N_21724);
nor U37321 (N_37321,N_21725,N_29248);
xnor U37322 (N_37322,N_23286,N_28721);
nand U37323 (N_37323,N_24647,N_25748);
xnor U37324 (N_37324,N_26107,N_28854);
xnor U37325 (N_37325,N_29431,N_23185);
nor U37326 (N_37326,N_27345,N_22318);
and U37327 (N_37327,N_26784,N_20067);
nor U37328 (N_37328,N_24423,N_26262);
and U37329 (N_37329,N_27780,N_20121);
or U37330 (N_37330,N_29917,N_29100);
xor U37331 (N_37331,N_21851,N_28028);
nor U37332 (N_37332,N_21020,N_28394);
or U37333 (N_37333,N_21564,N_25517);
and U37334 (N_37334,N_24781,N_25282);
or U37335 (N_37335,N_29839,N_21996);
xnor U37336 (N_37336,N_20449,N_23511);
or U37337 (N_37337,N_29930,N_25322);
nor U37338 (N_37338,N_23826,N_29951);
or U37339 (N_37339,N_24916,N_23877);
and U37340 (N_37340,N_22423,N_26567);
or U37341 (N_37341,N_23921,N_22820);
or U37342 (N_37342,N_20856,N_27815);
and U37343 (N_37343,N_20845,N_26537);
and U37344 (N_37344,N_21294,N_28165);
nor U37345 (N_37345,N_24202,N_21261);
and U37346 (N_37346,N_24039,N_26288);
and U37347 (N_37347,N_29689,N_29003);
nor U37348 (N_37348,N_22623,N_21814);
or U37349 (N_37349,N_26940,N_26021);
nand U37350 (N_37350,N_25213,N_27218);
or U37351 (N_37351,N_28680,N_24853);
or U37352 (N_37352,N_23590,N_21652);
or U37353 (N_37353,N_29142,N_22104);
and U37354 (N_37354,N_27344,N_20270);
nand U37355 (N_37355,N_24499,N_20171);
nor U37356 (N_37356,N_20320,N_23017);
or U37357 (N_37357,N_21090,N_29741);
or U37358 (N_37358,N_28634,N_21189);
and U37359 (N_37359,N_21222,N_27402);
or U37360 (N_37360,N_25384,N_27826);
or U37361 (N_37361,N_28414,N_23196);
nor U37362 (N_37362,N_26135,N_28520);
or U37363 (N_37363,N_24583,N_26936);
and U37364 (N_37364,N_21901,N_24447);
and U37365 (N_37365,N_21145,N_26136);
nor U37366 (N_37366,N_25224,N_20419);
nor U37367 (N_37367,N_29055,N_26826);
nand U37368 (N_37368,N_23744,N_28033);
and U37369 (N_37369,N_22886,N_22957);
nor U37370 (N_37370,N_29108,N_29962);
or U37371 (N_37371,N_26802,N_20375);
nand U37372 (N_37372,N_24150,N_23401);
nand U37373 (N_37373,N_21677,N_20279);
or U37374 (N_37374,N_24790,N_21924);
and U37375 (N_37375,N_22582,N_22403);
nor U37376 (N_37376,N_29399,N_29782);
nand U37377 (N_37377,N_25145,N_21200);
and U37378 (N_37378,N_21871,N_21127);
and U37379 (N_37379,N_27694,N_21797);
or U37380 (N_37380,N_21289,N_26590);
nand U37381 (N_37381,N_25169,N_22432);
or U37382 (N_37382,N_25020,N_29363);
and U37383 (N_37383,N_27133,N_26609);
or U37384 (N_37384,N_22228,N_29986);
nand U37385 (N_37385,N_22178,N_29923);
or U37386 (N_37386,N_27463,N_20944);
nor U37387 (N_37387,N_26988,N_27946);
nand U37388 (N_37388,N_26881,N_28339);
nand U37389 (N_37389,N_28008,N_20797);
or U37390 (N_37390,N_27476,N_29531);
and U37391 (N_37391,N_22271,N_26914);
nor U37392 (N_37392,N_27395,N_25661);
nor U37393 (N_37393,N_20368,N_29035);
nand U37394 (N_37394,N_22600,N_26877);
xor U37395 (N_37395,N_26411,N_24708);
and U37396 (N_37396,N_22199,N_21328);
and U37397 (N_37397,N_20886,N_24575);
xnor U37398 (N_37398,N_23833,N_29478);
and U37399 (N_37399,N_29339,N_22096);
xnor U37400 (N_37400,N_21161,N_24559);
nand U37401 (N_37401,N_21247,N_25050);
nor U37402 (N_37402,N_20461,N_25933);
nor U37403 (N_37403,N_23888,N_23549);
or U37404 (N_37404,N_20024,N_27675);
xnor U37405 (N_37405,N_21409,N_29059);
or U37406 (N_37406,N_29009,N_25524);
and U37407 (N_37407,N_21306,N_22663);
nand U37408 (N_37408,N_20180,N_21928);
nor U37409 (N_37409,N_20361,N_27474);
or U37410 (N_37410,N_21497,N_25914);
nor U37411 (N_37411,N_29778,N_29467);
nand U37412 (N_37412,N_22004,N_23107);
nand U37413 (N_37413,N_26124,N_23233);
or U37414 (N_37414,N_24927,N_22044);
or U37415 (N_37415,N_20561,N_22857);
nand U37416 (N_37416,N_27257,N_29502);
nor U37417 (N_37417,N_28430,N_25068);
and U37418 (N_37418,N_24217,N_26001);
or U37419 (N_37419,N_21146,N_21856);
or U37420 (N_37420,N_29338,N_27876);
and U37421 (N_37421,N_24029,N_22716);
nand U37422 (N_37422,N_25819,N_21351);
nand U37423 (N_37423,N_22847,N_20457);
nor U37424 (N_37424,N_26458,N_23786);
and U37425 (N_37425,N_25361,N_29456);
nand U37426 (N_37426,N_28354,N_20093);
nor U37427 (N_37427,N_28494,N_25178);
and U37428 (N_37428,N_21939,N_25964);
nor U37429 (N_37429,N_27662,N_23186);
xnor U37430 (N_37430,N_20334,N_24556);
or U37431 (N_37431,N_27030,N_26122);
nand U37432 (N_37432,N_23956,N_25335);
or U37433 (N_37433,N_20435,N_21294);
or U37434 (N_37434,N_27410,N_21342);
and U37435 (N_37435,N_22487,N_26175);
or U37436 (N_37436,N_27263,N_22668);
nand U37437 (N_37437,N_28544,N_27040);
nor U37438 (N_37438,N_22164,N_29701);
or U37439 (N_37439,N_25453,N_27461);
nand U37440 (N_37440,N_22496,N_27231);
nand U37441 (N_37441,N_25147,N_23214);
xor U37442 (N_37442,N_24631,N_21662);
nor U37443 (N_37443,N_23096,N_26023);
nand U37444 (N_37444,N_22652,N_26512);
or U37445 (N_37445,N_26591,N_22867);
nor U37446 (N_37446,N_28933,N_27512);
nand U37447 (N_37447,N_29544,N_28221);
xnor U37448 (N_37448,N_21404,N_22765);
xor U37449 (N_37449,N_24027,N_23494);
nand U37450 (N_37450,N_29156,N_27402);
nand U37451 (N_37451,N_21233,N_23489);
nand U37452 (N_37452,N_26642,N_24371);
or U37453 (N_37453,N_23566,N_20796);
nor U37454 (N_37454,N_24780,N_27234);
or U37455 (N_37455,N_21292,N_28745);
or U37456 (N_37456,N_21843,N_27032);
nor U37457 (N_37457,N_21215,N_26868);
xnor U37458 (N_37458,N_20203,N_29377);
xnor U37459 (N_37459,N_20899,N_20244);
or U37460 (N_37460,N_24543,N_25781);
or U37461 (N_37461,N_27749,N_28341);
or U37462 (N_37462,N_23488,N_20390);
or U37463 (N_37463,N_21432,N_27816);
nor U37464 (N_37464,N_21309,N_24177);
nor U37465 (N_37465,N_29911,N_23135);
nand U37466 (N_37466,N_21170,N_26492);
and U37467 (N_37467,N_28669,N_20961);
and U37468 (N_37468,N_25779,N_29581);
and U37469 (N_37469,N_29460,N_21119);
and U37470 (N_37470,N_29314,N_28490);
or U37471 (N_37471,N_23864,N_29414);
or U37472 (N_37472,N_27858,N_29603);
and U37473 (N_37473,N_27269,N_23843);
or U37474 (N_37474,N_25021,N_21474);
nand U37475 (N_37475,N_24523,N_24542);
nor U37476 (N_37476,N_22487,N_27328);
nand U37477 (N_37477,N_20028,N_20638);
nor U37478 (N_37478,N_24220,N_28125);
or U37479 (N_37479,N_25447,N_25065);
or U37480 (N_37480,N_21985,N_26320);
and U37481 (N_37481,N_28514,N_20810);
and U37482 (N_37482,N_21703,N_28093);
nand U37483 (N_37483,N_26084,N_26346);
nand U37484 (N_37484,N_27051,N_21382);
xnor U37485 (N_37485,N_28562,N_28450);
or U37486 (N_37486,N_27906,N_28406);
and U37487 (N_37487,N_27630,N_23677);
xnor U37488 (N_37488,N_29033,N_20370);
nand U37489 (N_37489,N_26124,N_24079);
and U37490 (N_37490,N_28127,N_26782);
and U37491 (N_37491,N_22288,N_23532);
nand U37492 (N_37492,N_28685,N_26430);
nand U37493 (N_37493,N_22824,N_22153);
or U37494 (N_37494,N_26182,N_24101);
and U37495 (N_37495,N_23245,N_27400);
nor U37496 (N_37496,N_28552,N_21045);
and U37497 (N_37497,N_26652,N_24695);
nand U37498 (N_37498,N_23622,N_24663);
or U37499 (N_37499,N_26935,N_21592);
nor U37500 (N_37500,N_25552,N_27452);
or U37501 (N_37501,N_25425,N_24362);
or U37502 (N_37502,N_29035,N_20802);
xnor U37503 (N_37503,N_26107,N_23204);
xor U37504 (N_37504,N_29023,N_28922);
nand U37505 (N_37505,N_20674,N_25812);
and U37506 (N_37506,N_27140,N_25143);
nand U37507 (N_37507,N_20212,N_27176);
nand U37508 (N_37508,N_23519,N_25575);
or U37509 (N_37509,N_21804,N_29445);
or U37510 (N_37510,N_22773,N_26208);
and U37511 (N_37511,N_26426,N_20293);
and U37512 (N_37512,N_22850,N_25482);
and U37513 (N_37513,N_26468,N_25120);
or U37514 (N_37514,N_24364,N_26286);
nand U37515 (N_37515,N_28828,N_27588);
and U37516 (N_37516,N_26666,N_26148);
or U37517 (N_37517,N_28111,N_28493);
nand U37518 (N_37518,N_21509,N_25969);
and U37519 (N_37519,N_23088,N_28011);
xnor U37520 (N_37520,N_27444,N_21413);
nand U37521 (N_37521,N_24758,N_28346);
nor U37522 (N_37522,N_28869,N_21354);
nand U37523 (N_37523,N_25770,N_28126);
or U37524 (N_37524,N_20722,N_20399);
and U37525 (N_37525,N_29722,N_23742);
nand U37526 (N_37526,N_23872,N_21926);
nand U37527 (N_37527,N_28680,N_28209);
nand U37528 (N_37528,N_24570,N_28437);
and U37529 (N_37529,N_27879,N_21182);
xnor U37530 (N_37530,N_22727,N_26945);
or U37531 (N_37531,N_25841,N_28604);
or U37532 (N_37532,N_22188,N_23925);
nor U37533 (N_37533,N_27301,N_20253);
or U37534 (N_37534,N_25253,N_28561);
nor U37535 (N_37535,N_27964,N_29589);
and U37536 (N_37536,N_28837,N_28919);
nand U37537 (N_37537,N_20857,N_29693);
nor U37538 (N_37538,N_20096,N_28296);
and U37539 (N_37539,N_27702,N_26881);
and U37540 (N_37540,N_28313,N_21862);
nand U37541 (N_37541,N_25806,N_22000);
nor U37542 (N_37542,N_28709,N_24287);
nor U37543 (N_37543,N_26280,N_27028);
nand U37544 (N_37544,N_26374,N_24985);
nand U37545 (N_37545,N_24875,N_23417);
nand U37546 (N_37546,N_29942,N_22272);
nand U37547 (N_37547,N_26790,N_28654);
and U37548 (N_37548,N_25339,N_28434);
nand U37549 (N_37549,N_25157,N_27992);
or U37550 (N_37550,N_26882,N_22828);
and U37551 (N_37551,N_21190,N_25780);
and U37552 (N_37552,N_28786,N_29919);
nand U37553 (N_37553,N_25545,N_20466);
and U37554 (N_37554,N_23103,N_22824);
nor U37555 (N_37555,N_27009,N_24593);
and U37556 (N_37556,N_20815,N_24795);
or U37557 (N_37557,N_22217,N_24090);
and U37558 (N_37558,N_24273,N_20265);
nor U37559 (N_37559,N_28515,N_21769);
or U37560 (N_37560,N_27902,N_20689);
xnor U37561 (N_37561,N_24330,N_20919);
xnor U37562 (N_37562,N_29413,N_28433);
and U37563 (N_37563,N_20271,N_24194);
xnor U37564 (N_37564,N_20053,N_28768);
and U37565 (N_37565,N_27941,N_27310);
nand U37566 (N_37566,N_27183,N_22155);
and U37567 (N_37567,N_24372,N_27037);
nand U37568 (N_37568,N_21486,N_29677);
xor U37569 (N_37569,N_29481,N_22591);
xor U37570 (N_37570,N_20395,N_20786);
xnor U37571 (N_37571,N_24808,N_27222);
xnor U37572 (N_37572,N_24166,N_28620);
or U37573 (N_37573,N_22647,N_25394);
nand U37574 (N_37574,N_27942,N_24497);
or U37575 (N_37575,N_26062,N_29784);
nor U37576 (N_37576,N_27504,N_29194);
nand U37577 (N_37577,N_21500,N_27403);
nand U37578 (N_37578,N_20959,N_26486);
or U37579 (N_37579,N_28841,N_27238);
nand U37580 (N_37580,N_25284,N_26064);
nor U37581 (N_37581,N_20892,N_22107);
and U37582 (N_37582,N_23746,N_24774);
and U37583 (N_37583,N_26146,N_28680);
and U37584 (N_37584,N_27205,N_24693);
and U37585 (N_37585,N_22590,N_25809);
nor U37586 (N_37586,N_22733,N_20479);
nor U37587 (N_37587,N_27892,N_28199);
or U37588 (N_37588,N_28722,N_23576);
or U37589 (N_37589,N_23906,N_20370);
and U37590 (N_37590,N_29048,N_26170);
nand U37591 (N_37591,N_26994,N_25269);
nand U37592 (N_37592,N_23141,N_22386);
or U37593 (N_37593,N_23503,N_20161);
xor U37594 (N_37594,N_22253,N_25572);
nor U37595 (N_37595,N_27595,N_25235);
and U37596 (N_37596,N_27922,N_23355);
and U37597 (N_37597,N_29594,N_21439);
nor U37598 (N_37598,N_20932,N_24821);
nand U37599 (N_37599,N_20981,N_27029);
nor U37600 (N_37600,N_21788,N_21882);
or U37601 (N_37601,N_21118,N_29415);
and U37602 (N_37602,N_25733,N_22887);
xnor U37603 (N_37603,N_29691,N_25924);
nand U37604 (N_37604,N_27259,N_26278);
and U37605 (N_37605,N_23556,N_22474);
and U37606 (N_37606,N_26185,N_20679);
and U37607 (N_37607,N_23273,N_23857);
or U37608 (N_37608,N_20675,N_27836);
nand U37609 (N_37609,N_29564,N_27911);
xnor U37610 (N_37610,N_21498,N_26157);
or U37611 (N_37611,N_25317,N_21719);
nor U37612 (N_37612,N_21092,N_28672);
and U37613 (N_37613,N_28368,N_20821);
or U37614 (N_37614,N_29654,N_21337);
xor U37615 (N_37615,N_27206,N_24309);
or U37616 (N_37616,N_20045,N_22739);
and U37617 (N_37617,N_23764,N_26258);
nand U37618 (N_37618,N_26903,N_25163);
nor U37619 (N_37619,N_26663,N_26575);
nand U37620 (N_37620,N_20834,N_29970);
and U37621 (N_37621,N_23089,N_25096);
nand U37622 (N_37622,N_23761,N_27626);
nor U37623 (N_37623,N_24232,N_20036);
xnor U37624 (N_37624,N_23879,N_25748);
nor U37625 (N_37625,N_21389,N_21136);
nor U37626 (N_37626,N_28622,N_27829);
or U37627 (N_37627,N_26793,N_20163);
or U37628 (N_37628,N_28596,N_25849);
or U37629 (N_37629,N_28409,N_24701);
and U37630 (N_37630,N_23372,N_24822);
and U37631 (N_37631,N_24781,N_26952);
or U37632 (N_37632,N_22043,N_23696);
nor U37633 (N_37633,N_26027,N_27178);
xor U37634 (N_37634,N_28912,N_20887);
and U37635 (N_37635,N_29207,N_21488);
and U37636 (N_37636,N_22882,N_24411);
or U37637 (N_37637,N_20961,N_28472);
nor U37638 (N_37638,N_24738,N_27199);
or U37639 (N_37639,N_20926,N_24027);
nor U37640 (N_37640,N_29839,N_27050);
nand U37641 (N_37641,N_27788,N_26670);
and U37642 (N_37642,N_29400,N_20372);
and U37643 (N_37643,N_28595,N_27171);
nand U37644 (N_37644,N_23636,N_25159);
and U37645 (N_37645,N_27532,N_27082);
and U37646 (N_37646,N_29046,N_22840);
xor U37647 (N_37647,N_20734,N_25092);
nor U37648 (N_37648,N_23023,N_29872);
nor U37649 (N_37649,N_27612,N_20050);
nand U37650 (N_37650,N_26969,N_21959);
nand U37651 (N_37651,N_27333,N_25990);
xor U37652 (N_37652,N_21632,N_23573);
nand U37653 (N_37653,N_28847,N_28598);
nand U37654 (N_37654,N_27065,N_22614);
xor U37655 (N_37655,N_20709,N_27182);
xnor U37656 (N_37656,N_29834,N_24431);
and U37657 (N_37657,N_25353,N_22363);
nor U37658 (N_37658,N_22186,N_20668);
and U37659 (N_37659,N_28327,N_21932);
nor U37660 (N_37660,N_28490,N_26577);
nand U37661 (N_37661,N_27344,N_20733);
or U37662 (N_37662,N_22392,N_20718);
nor U37663 (N_37663,N_26918,N_28215);
nor U37664 (N_37664,N_29532,N_27341);
and U37665 (N_37665,N_23370,N_22815);
or U37666 (N_37666,N_26977,N_25351);
nor U37667 (N_37667,N_28643,N_22178);
xnor U37668 (N_37668,N_28396,N_29737);
or U37669 (N_37669,N_24429,N_23627);
nor U37670 (N_37670,N_29873,N_24919);
or U37671 (N_37671,N_28845,N_29521);
nand U37672 (N_37672,N_24394,N_28515);
nand U37673 (N_37673,N_24965,N_22607);
nor U37674 (N_37674,N_21369,N_28527);
and U37675 (N_37675,N_28086,N_25792);
nand U37676 (N_37676,N_27093,N_24641);
xnor U37677 (N_37677,N_21638,N_27237);
nor U37678 (N_37678,N_23870,N_25658);
xnor U37679 (N_37679,N_24755,N_29851);
nand U37680 (N_37680,N_20980,N_21116);
or U37681 (N_37681,N_22995,N_21334);
or U37682 (N_37682,N_28110,N_28229);
and U37683 (N_37683,N_22213,N_26048);
and U37684 (N_37684,N_23815,N_25912);
nor U37685 (N_37685,N_27766,N_23714);
and U37686 (N_37686,N_25823,N_29125);
or U37687 (N_37687,N_23397,N_22781);
nand U37688 (N_37688,N_25592,N_21845);
nand U37689 (N_37689,N_22160,N_21678);
nand U37690 (N_37690,N_29139,N_20224);
and U37691 (N_37691,N_26896,N_26294);
nand U37692 (N_37692,N_26307,N_25867);
xnor U37693 (N_37693,N_26441,N_27836);
xor U37694 (N_37694,N_28438,N_20806);
and U37695 (N_37695,N_25191,N_22289);
and U37696 (N_37696,N_29028,N_23459);
nand U37697 (N_37697,N_22659,N_24023);
and U37698 (N_37698,N_23133,N_25350);
nand U37699 (N_37699,N_26871,N_23494);
and U37700 (N_37700,N_25038,N_20257);
or U37701 (N_37701,N_27702,N_27071);
nor U37702 (N_37702,N_20927,N_21361);
nor U37703 (N_37703,N_26331,N_27242);
and U37704 (N_37704,N_21290,N_22278);
nand U37705 (N_37705,N_26366,N_28749);
or U37706 (N_37706,N_29287,N_20883);
xnor U37707 (N_37707,N_23777,N_26353);
and U37708 (N_37708,N_27196,N_28667);
nand U37709 (N_37709,N_21913,N_27747);
and U37710 (N_37710,N_25238,N_28155);
xor U37711 (N_37711,N_28089,N_28172);
nand U37712 (N_37712,N_26741,N_26798);
nand U37713 (N_37713,N_22458,N_25700);
or U37714 (N_37714,N_29050,N_20949);
nand U37715 (N_37715,N_20118,N_23635);
nand U37716 (N_37716,N_23913,N_27418);
or U37717 (N_37717,N_26568,N_24554);
and U37718 (N_37718,N_22650,N_23922);
or U37719 (N_37719,N_22840,N_25545);
nand U37720 (N_37720,N_28652,N_28326);
nor U37721 (N_37721,N_20601,N_24402);
xnor U37722 (N_37722,N_28330,N_21618);
or U37723 (N_37723,N_27648,N_28760);
and U37724 (N_37724,N_26985,N_22602);
and U37725 (N_37725,N_23634,N_27514);
nor U37726 (N_37726,N_29615,N_25416);
xor U37727 (N_37727,N_28835,N_20716);
nor U37728 (N_37728,N_27483,N_21446);
nand U37729 (N_37729,N_29668,N_23687);
nor U37730 (N_37730,N_22169,N_22243);
and U37731 (N_37731,N_26333,N_28085);
nor U37732 (N_37732,N_20641,N_26833);
xnor U37733 (N_37733,N_25403,N_21081);
nor U37734 (N_37734,N_22021,N_24410);
and U37735 (N_37735,N_28556,N_26267);
nand U37736 (N_37736,N_23984,N_28942);
nand U37737 (N_37737,N_20004,N_20515);
nand U37738 (N_37738,N_22268,N_23487);
or U37739 (N_37739,N_27535,N_25987);
nor U37740 (N_37740,N_21213,N_29787);
or U37741 (N_37741,N_21161,N_25976);
and U37742 (N_37742,N_28645,N_26817);
nand U37743 (N_37743,N_27386,N_28488);
or U37744 (N_37744,N_22603,N_29160);
nand U37745 (N_37745,N_28505,N_27244);
nand U37746 (N_37746,N_23627,N_23848);
nand U37747 (N_37747,N_26325,N_23657);
and U37748 (N_37748,N_20554,N_22077);
nor U37749 (N_37749,N_28190,N_26633);
and U37750 (N_37750,N_21772,N_29255);
or U37751 (N_37751,N_27366,N_20570);
and U37752 (N_37752,N_29361,N_25854);
or U37753 (N_37753,N_29229,N_27825);
nand U37754 (N_37754,N_26850,N_28703);
nand U37755 (N_37755,N_22810,N_24048);
nand U37756 (N_37756,N_28263,N_29010);
or U37757 (N_37757,N_20180,N_26783);
and U37758 (N_37758,N_27197,N_21771);
and U37759 (N_37759,N_27765,N_28170);
or U37760 (N_37760,N_26545,N_29830);
nor U37761 (N_37761,N_25756,N_24034);
or U37762 (N_37762,N_26528,N_23613);
and U37763 (N_37763,N_26218,N_24221);
xnor U37764 (N_37764,N_24021,N_29900);
nand U37765 (N_37765,N_22424,N_24143);
or U37766 (N_37766,N_22812,N_22252);
or U37767 (N_37767,N_27334,N_27400);
and U37768 (N_37768,N_21144,N_26298);
xnor U37769 (N_37769,N_22178,N_21458);
xnor U37770 (N_37770,N_24090,N_23438);
nor U37771 (N_37771,N_28009,N_24944);
or U37772 (N_37772,N_28056,N_29970);
nor U37773 (N_37773,N_27669,N_23495);
and U37774 (N_37774,N_24736,N_21230);
nand U37775 (N_37775,N_24271,N_20595);
or U37776 (N_37776,N_24462,N_23548);
or U37777 (N_37777,N_24027,N_28433);
xor U37778 (N_37778,N_26958,N_25050);
or U37779 (N_37779,N_29325,N_25410);
nand U37780 (N_37780,N_29817,N_29296);
or U37781 (N_37781,N_26261,N_24640);
nand U37782 (N_37782,N_26479,N_24408);
nor U37783 (N_37783,N_25348,N_24671);
nand U37784 (N_37784,N_26475,N_29226);
and U37785 (N_37785,N_29983,N_21274);
and U37786 (N_37786,N_20961,N_21804);
nand U37787 (N_37787,N_20659,N_29230);
nand U37788 (N_37788,N_22134,N_29563);
nand U37789 (N_37789,N_26673,N_29314);
or U37790 (N_37790,N_24205,N_25477);
and U37791 (N_37791,N_29672,N_25569);
or U37792 (N_37792,N_27755,N_28341);
nor U37793 (N_37793,N_25569,N_27414);
or U37794 (N_37794,N_21305,N_22656);
or U37795 (N_37795,N_24056,N_29101);
and U37796 (N_37796,N_28649,N_24767);
nor U37797 (N_37797,N_23892,N_28883);
or U37798 (N_37798,N_26977,N_29452);
or U37799 (N_37799,N_21737,N_24828);
nand U37800 (N_37800,N_20502,N_25449);
or U37801 (N_37801,N_28872,N_21723);
and U37802 (N_37802,N_20372,N_20681);
nand U37803 (N_37803,N_23770,N_21461);
or U37804 (N_37804,N_23192,N_26968);
nor U37805 (N_37805,N_23696,N_20858);
xor U37806 (N_37806,N_26388,N_25594);
and U37807 (N_37807,N_24426,N_24820);
nand U37808 (N_37808,N_24400,N_20888);
nor U37809 (N_37809,N_23550,N_22732);
nand U37810 (N_37810,N_20104,N_21442);
nor U37811 (N_37811,N_26799,N_27673);
and U37812 (N_37812,N_29021,N_20696);
xor U37813 (N_37813,N_29027,N_20837);
nor U37814 (N_37814,N_25361,N_24705);
nor U37815 (N_37815,N_27599,N_27250);
nor U37816 (N_37816,N_20546,N_27916);
nor U37817 (N_37817,N_23822,N_24587);
or U37818 (N_37818,N_29684,N_25552);
nor U37819 (N_37819,N_20844,N_22437);
nand U37820 (N_37820,N_20662,N_28518);
nor U37821 (N_37821,N_24448,N_26450);
or U37822 (N_37822,N_21833,N_22430);
and U37823 (N_37823,N_26597,N_21230);
nor U37824 (N_37824,N_26756,N_23817);
xnor U37825 (N_37825,N_27566,N_26970);
nor U37826 (N_37826,N_20315,N_29085);
or U37827 (N_37827,N_23363,N_25051);
nand U37828 (N_37828,N_26009,N_23709);
nor U37829 (N_37829,N_21368,N_20880);
xor U37830 (N_37830,N_28773,N_24767);
and U37831 (N_37831,N_20892,N_23208);
or U37832 (N_37832,N_26769,N_28889);
or U37833 (N_37833,N_25885,N_21412);
nor U37834 (N_37834,N_27171,N_22127);
nor U37835 (N_37835,N_24652,N_20275);
or U37836 (N_37836,N_21649,N_29367);
or U37837 (N_37837,N_20889,N_24167);
and U37838 (N_37838,N_28384,N_22472);
xnor U37839 (N_37839,N_29220,N_27576);
nand U37840 (N_37840,N_25922,N_21427);
nand U37841 (N_37841,N_29113,N_26398);
nand U37842 (N_37842,N_29214,N_21761);
or U37843 (N_37843,N_25425,N_28778);
or U37844 (N_37844,N_22797,N_27912);
nor U37845 (N_37845,N_25797,N_28799);
nand U37846 (N_37846,N_27910,N_27449);
and U37847 (N_37847,N_20098,N_28020);
and U37848 (N_37848,N_25183,N_20061);
nor U37849 (N_37849,N_29921,N_28705);
xor U37850 (N_37850,N_23469,N_27775);
and U37851 (N_37851,N_27924,N_24363);
or U37852 (N_37852,N_26135,N_20714);
nor U37853 (N_37853,N_21169,N_25039);
and U37854 (N_37854,N_24425,N_22075);
and U37855 (N_37855,N_28595,N_27858);
nor U37856 (N_37856,N_22637,N_27562);
and U37857 (N_37857,N_25624,N_27576);
nor U37858 (N_37858,N_24784,N_21347);
and U37859 (N_37859,N_20788,N_25865);
nor U37860 (N_37860,N_26959,N_28714);
and U37861 (N_37861,N_20878,N_24779);
and U37862 (N_37862,N_22045,N_23075);
and U37863 (N_37863,N_23581,N_26161);
nor U37864 (N_37864,N_24504,N_27178);
nand U37865 (N_37865,N_27292,N_20323);
xnor U37866 (N_37866,N_29102,N_27191);
nor U37867 (N_37867,N_20794,N_28190);
or U37868 (N_37868,N_26192,N_20192);
nor U37869 (N_37869,N_24986,N_20755);
nand U37870 (N_37870,N_21008,N_21103);
xor U37871 (N_37871,N_26378,N_24165);
and U37872 (N_37872,N_28509,N_20822);
nand U37873 (N_37873,N_28450,N_23058);
and U37874 (N_37874,N_20342,N_24098);
or U37875 (N_37875,N_27829,N_20587);
nor U37876 (N_37876,N_21062,N_24604);
and U37877 (N_37877,N_25627,N_25141);
or U37878 (N_37878,N_28885,N_28501);
or U37879 (N_37879,N_22689,N_27480);
nor U37880 (N_37880,N_26515,N_28127);
nand U37881 (N_37881,N_27893,N_28072);
nor U37882 (N_37882,N_29576,N_26487);
and U37883 (N_37883,N_28508,N_24235);
nor U37884 (N_37884,N_23116,N_24307);
xor U37885 (N_37885,N_25805,N_26612);
nand U37886 (N_37886,N_20790,N_23730);
or U37887 (N_37887,N_22187,N_22181);
nand U37888 (N_37888,N_26240,N_28066);
nand U37889 (N_37889,N_24918,N_20198);
nand U37890 (N_37890,N_22197,N_22101);
and U37891 (N_37891,N_23473,N_22115);
and U37892 (N_37892,N_20235,N_28718);
xor U37893 (N_37893,N_20161,N_29138);
or U37894 (N_37894,N_29981,N_23601);
nor U37895 (N_37895,N_25565,N_23809);
nand U37896 (N_37896,N_26318,N_24704);
xor U37897 (N_37897,N_29632,N_21171);
nand U37898 (N_37898,N_26900,N_24252);
nor U37899 (N_37899,N_24867,N_23773);
nor U37900 (N_37900,N_26900,N_22035);
or U37901 (N_37901,N_29086,N_20563);
and U37902 (N_37902,N_28620,N_27291);
and U37903 (N_37903,N_27351,N_21730);
xnor U37904 (N_37904,N_24127,N_28953);
or U37905 (N_37905,N_23307,N_23716);
and U37906 (N_37906,N_21411,N_23532);
and U37907 (N_37907,N_22133,N_28215);
nand U37908 (N_37908,N_28646,N_23104);
and U37909 (N_37909,N_22889,N_21477);
or U37910 (N_37910,N_24281,N_20994);
nand U37911 (N_37911,N_26911,N_28504);
and U37912 (N_37912,N_23882,N_28771);
nor U37913 (N_37913,N_20789,N_27821);
nand U37914 (N_37914,N_29177,N_24854);
nor U37915 (N_37915,N_21837,N_21983);
xnor U37916 (N_37916,N_25325,N_20404);
and U37917 (N_37917,N_22791,N_28381);
nor U37918 (N_37918,N_28119,N_20362);
or U37919 (N_37919,N_21805,N_27803);
nand U37920 (N_37920,N_25739,N_24029);
or U37921 (N_37921,N_22344,N_28634);
nor U37922 (N_37922,N_20410,N_23245);
nand U37923 (N_37923,N_21781,N_29831);
and U37924 (N_37924,N_23893,N_28126);
xor U37925 (N_37925,N_23706,N_25923);
or U37926 (N_37926,N_24753,N_22274);
or U37927 (N_37927,N_28357,N_20296);
xnor U37928 (N_37928,N_25098,N_27495);
nand U37929 (N_37929,N_26813,N_20072);
or U37930 (N_37930,N_27247,N_25316);
xnor U37931 (N_37931,N_26529,N_27302);
or U37932 (N_37932,N_20773,N_25819);
xnor U37933 (N_37933,N_20539,N_24567);
and U37934 (N_37934,N_26372,N_22027);
and U37935 (N_37935,N_25097,N_21716);
and U37936 (N_37936,N_20665,N_24305);
nand U37937 (N_37937,N_24017,N_22893);
and U37938 (N_37938,N_24608,N_28661);
and U37939 (N_37939,N_22446,N_25156);
nand U37940 (N_37940,N_21899,N_28038);
nand U37941 (N_37941,N_28817,N_21379);
and U37942 (N_37942,N_21389,N_28482);
or U37943 (N_37943,N_29509,N_28853);
or U37944 (N_37944,N_27186,N_21725);
and U37945 (N_37945,N_27980,N_28026);
or U37946 (N_37946,N_26982,N_25726);
and U37947 (N_37947,N_21163,N_28545);
or U37948 (N_37948,N_26954,N_26753);
and U37949 (N_37949,N_28179,N_22118);
nand U37950 (N_37950,N_24199,N_24364);
nor U37951 (N_37951,N_29946,N_21005);
or U37952 (N_37952,N_26233,N_21675);
nor U37953 (N_37953,N_24010,N_28991);
nor U37954 (N_37954,N_25694,N_21763);
and U37955 (N_37955,N_21021,N_27823);
nand U37956 (N_37956,N_23637,N_26773);
and U37957 (N_37957,N_27494,N_24256);
and U37958 (N_37958,N_24599,N_29477);
or U37959 (N_37959,N_22865,N_20917);
or U37960 (N_37960,N_23472,N_26209);
and U37961 (N_37961,N_26049,N_29964);
xnor U37962 (N_37962,N_24793,N_28457);
or U37963 (N_37963,N_29100,N_26682);
nor U37964 (N_37964,N_27227,N_29237);
or U37965 (N_37965,N_26959,N_29258);
or U37966 (N_37966,N_21650,N_26044);
nor U37967 (N_37967,N_22267,N_28536);
nor U37968 (N_37968,N_24653,N_26069);
nand U37969 (N_37969,N_21185,N_21872);
nor U37970 (N_37970,N_23642,N_27191);
nand U37971 (N_37971,N_23007,N_20747);
nor U37972 (N_37972,N_29314,N_23889);
or U37973 (N_37973,N_26047,N_27792);
nand U37974 (N_37974,N_24325,N_26219);
nor U37975 (N_37975,N_25035,N_20188);
or U37976 (N_37976,N_25755,N_21875);
or U37977 (N_37977,N_20398,N_21043);
xnor U37978 (N_37978,N_21771,N_25875);
nand U37979 (N_37979,N_25428,N_24142);
and U37980 (N_37980,N_22016,N_29609);
nor U37981 (N_37981,N_28501,N_20699);
xor U37982 (N_37982,N_21779,N_24606);
xnor U37983 (N_37983,N_27900,N_25983);
nand U37984 (N_37984,N_21871,N_23134);
or U37985 (N_37985,N_28708,N_25066);
nand U37986 (N_37986,N_21813,N_25482);
and U37987 (N_37987,N_25647,N_24257);
and U37988 (N_37988,N_20817,N_25497);
and U37989 (N_37989,N_26511,N_24293);
and U37990 (N_37990,N_21789,N_24194);
xnor U37991 (N_37991,N_22138,N_23139);
and U37992 (N_37992,N_24243,N_20197);
nand U37993 (N_37993,N_22152,N_29895);
or U37994 (N_37994,N_27834,N_20784);
nor U37995 (N_37995,N_29927,N_25500);
and U37996 (N_37996,N_22437,N_23137);
xnor U37997 (N_37997,N_27490,N_23896);
and U37998 (N_37998,N_21004,N_24633);
or U37999 (N_37999,N_26207,N_20982);
or U38000 (N_38000,N_24679,N_20316);
or U38001 (N_38001,N_20837,N_20801);
nand U38002 (N_38002,N_25804,N_24119);
or U38003 (N_38003,N_23975,N_26170);
and U38004 (N_38004,N_24478,N_27178);
nand U38005 (N_38005,N_20394,N_23748);
nand U38006 (N_38006,N_20511,N_25589);
or U38007 (N_38007,N_23137,N_25143);
or U38008 (N_38008,N_24591,N_26147);
xor U38009 (N_38009,N_28712,N_29310);
or U38010 (N_38010,N_23497,N_27564);
xnor U38011 (N_38011,N_27302,N_24585);
or U38012 (N_38012,N_27111,N_20933);
or U38013 (N_38013,N_29802,N_23809);
or U38014 (N_38014,N_22933,N_27589);
or U38015 (N_38015,N_29871,N_29808);
nand U38016 (N_38016,N_25965,N_25198);
xor U38017 (N_38017,N_28381,N_24066);
or U38018 (N_38018,N_24128,N_23604);
or U38019 (N_38019,N_24368,N_25495);
nand U38020 (N_38020,N_24596,N_20956);
nand U38021 (N_38021,N_29208,N_26868);
nor U38022 (N_38022,N_26653,N_28180);
or U38023 (N_38023,N_28078,N_21434);
or U38024 (N_38024,N_22636,N_21472);
nand U38025 (N_38025,N_21599,N_21272);
and U38026 (N_38026,N_26639,N_22557);
xor U38027 (N_38027,N_21790,N_21275);
and U38028 (N_38028,N_25074,N_26784);
nand U38029 (N_38029,N_28303,N_21265);
and U38030 (N_38030,N_20155,N_27218);
nand U38031 (N_38031,N_20902,N_27366);
or U38032 (N_38032,N_20843,N_25965);
xnor U38033 (N_38033,N_27856,N_25374);
nor U38034 (N_38034,N_26728,N_20936);
nor U38035 (N_38035,N_27062,N_26240);
nand U38036 (N_38036,N_26213,N_23994);
nor U38037 (N_38037,N_22988,N_27575);
nand U38038 (N_38038,N_29038,N_27653);
and U38039 (N_38039,N_20776,N_23173);
nor U38040 (N_38040,N_22030,N_28641);
or U38041 (N_38041,N_22645,N_27157);
and U38042 (N_38042,N_23108,N_21180);
nor U38043 (N_38043,N_21341,N_28683);
or U38044 (N_38044,N_29747,N_23622);
nand U38045 (N_38045,N_21460,N_29655);
and U38046 (N_38046,N_21284,N_24662);
and U38047 (N_38047,N_20982,N_26298);
or U38048 (N_38048,N_22403,N_26983);
nor U38049 (N_38049,N_29660,N_27198);
nand U38050 (N_38050,N_26660,N_23004);
or U38051 (N_38051,N_28489,N_26327);
xnor U38052 (N_38052,N_24742,N_21597);
nand U38053 (N_38053,N_27205,N_24368);
nand U38054 (N_38054,N_29038,N_25492);
and U38055 (N_38055,N_21305,N_21521);
and U38056 (N_38056,N_29227,N_24956);
or U38057 (N_38057,N_29675,N_23073);
and U38058 (N_38058,N_26422,N_27820);
nand U38059 (N_38059,N_24949,N_23138);
or U38060 (N_38060,N_25001,N_26232);
nand U38061 (N_38061,N_28523,N_22905);
and U38062 (N_38062,N_22841,N_23731);
nand U38063 (N_38063,N_29279,N_20212);
or U38064 (N_38064,N_20197,N_28994);
xor U38065 (N_38065,N_29155,N_29284);
or U38066 (N_38066,N_24225,N_24105);
nor U38067 (N_38067,N_22417,N_21911);
and U38068 (N_38068,N_20985,N_26936);
nor U38069 (N_38069,N_21775,N_26671);
xor U38070 (N_38070,N_24843,N_20860);
or U38071 (N_38071,N_24285,N_21965);
nor U38072 (N_38072,N_21183,N_20486);
or U38073 (N_38073,N_23327,N_24374);
or U38074 (N_38074,N_28636,N_24314);
or U38075 (N_38075,N_23472,N_26469);
and U38076 (N_38076,N_26309,N_26836);
and U38077 (N_38077,N_21864,N_28884);
nor U38078 (N_38078,N_25022,N_28527);
xnor U38079 (N_38079,N_20870,N_28935);
or U38080 (N_38080,N_24432,N_28834);
and U38081 (N_38081,N_22367,N_22582);
nand U38082 (N_38082,N_28197,N_27474);
nand U38083 (N_38083,N_21018,N_27156);
nand U38084 (N_38084,N_28530,N_20462);
nand U38085 (N_38085,N_24984,N_29875);
nor U38086 (N_38086,N_26240,N_21759);
and U38087 (N_38087,N_21888,N_23967);
nand U38088 (N_38088,N_28986,N_25862);
or U38089 (N_38089,N_28638,N_25293);
or U38090 (N_38090,N_28022,N_27088);
or U38091 (N_38091,N_20690,N_25810);
nor U38092 (N_38092,N_25862,N_21142);
and U38093 (N_38093,N_26256,N_26381);
or U38094 (N_38094,N_25396,N_23092);
and U38095 (N_38095,N_20180,N_22682);
and U38096 (N_38096,N_29534,N_29046);
nor U38097 (N_38097,N_27549,N_22674);
nand U38098 (N_38098,N_22120,N_24047);
nor U38099 (N_38099,N_22500,N_22526);
nand U38100 (N_38100,N_24093,N_29429);
nand U38101 (N_38101,N_28083,N_27963);
xor U38102 (N_38102,N_20123,N_29981);
or U38103 (N_38103,N_20043,N_20098);
and U38104 (N_38104,N_25803,N_22983);
xor U38105 (N_38105,N_23567,N_29945);
or U38106 (N_38106,N_21893,N_29385);
and U38107 (N_38107,N_25784,N_21239);
nor U38108 (N_38108,N_25703,N_28088);
and U38109 (N_38109,N_26442,N_22385);
and U38110 (N_38110,N_23217,N_24964);
and U38111 (N_38111,N_21615,N_25168);
and U38112 (N_38112,N_20683,N_28829);
xnor U38113 (N_38113,N_22150,N_20956);
or U38114 (N_38114,N_28710,N_23973);
nand U38115 (N_38115,N_28193,N_23157);
nand U38116 (N_38116,N_28783,N_22530);
xor U38117 (N_38117,N_28321,N_21325);
or U38118 (N_38118,N_20268,N_29327);
and U38119 (N_38119,N_25927,N_21862);
nor U38120 (N_38120,N_24010,N_22548);
nand U38121 (N_38121,N_20335,N_23659);
or U38122 (N_38122,N_24106,N_26508);
nor U38123 (N_38123,N_25985,N_26121);
and U38124 (N_38124,N_29900,N_23362);
and U38125 (N_38125,N_23331,N_26777);
nand U38126 (N_38126,N_27614,N_25078);
nand U38127 (N_38127,N_22147,N_27410);
and U38128 (N_38128,N_21417,N_24977);
nand U38129 (N_38129,N_27394,N_29018);
and U38130 (N_38130,N_23367,N_23511);
or U38131 (N_38131,N_29108,N_22218);
nor U38132 (N_38132,N_23885,N_25676);
and U38133 (N_38133,N_24373,N_22684);
nor U38134 (N_38134,N_21438,N_23387);
nand U38135 (N_38135,N_25550,N_25750);
nand U38136 (N_38136,N_26705,N_27075);
and U38137 (N_38137,N_22549,N_25568);
and U38138 (N_38138,N_26715,N_29679);
and U38139 (N_38139,N_26821,N_28218);
nor U38140 (N_38140,N_24889,N_22108);
nor U38141 (N_38141,N_28780,N_21268);
and U38142 (N_38142,N_25435,N_25592);
nand U38143 (N_38143,N_21757,N_26039);
nor U38144 (N_38144,N_27308,N_26325);
and U38145 (N_38145,N_28972,N_27424);
or U38146 (N_38146,N_28736,N_24789);
nand U38147 (N_38147,N_22652,N_21494);
nor U38148 (N_38148,N_22455,N_27489);
nand U38149 (N_38149,N_22777,N_29544);
nand U38150 (N_38150,N_29578,N_27476);
and U38151 (N_38151,N_26450,N_24434);
nand U38152 (N_38152,N_25387,N_20282);
nor U38153 (N_38153,N_23059,N_29999);
nor U38154 (N_38154,N_21578,N_27265);
or U38155 (N_38155,N_29159,N_24508);
and U38156 (N_38156,N_21520,N_22548);
and U38157 (N_38157,N_26363,N_27300);
nor U38158 (N_38158,N_28283,N_20123);
and U38159 (N_38159,N_20998,N_29208);
nand U38160 (N_38160,N_25953,N_20230);
and U38161 (N_38161,N_24786,N_23574);
nand U38162 (N_38162,N_24812,N_20241);
nand U38163 (N_38163,N_27821,N_26015);
and U38164 (N_38164,N_28501,N_21669);
nor U38165 (N_38165,N_22558,N_28315);
and U38166 (N_38166,N_28137,N_21988);
and U38167 (N_38167,N_20275,N_29439);
or U38168 (N_38168,N_25294,N_25275);
xor U38169 (N_38169,N_24351,N_22533);
nor U38170 (N_38170,N_23218,N_25381);
xnor U38171 (N_38171,N_21076,N_20333);
and U38172 (N_38172,N_27671,N_26669);
or U38173 (N_38173,N_29895,N_22758);
nor U38174 (N_38174,N_23900,N_24827);
xor U38175 (N_38175,N_27453,N_27363);
and U38176 (N_38176,N_26869,N_23365);
or U38177 (N_38177,N_23905,N_28416);
and U38178 (N_38178,N_20503,N_25007);
nor U38179 (N_38179,N_28005,N_25848);
or U38180 (N_38180,N_23022,N_24773);
nand U38181 (N_38181,N_24473,N_22534);
nor U38182 (N_38182,N_29680,N_23225);
or U38183 (N_38183,N_23228,N_24030);
and U38184 (N_38184,N_20171,N_23479);
nor U38185 (N_38185,N_29566,N_21414);
nor U38186 (N_38186,N_24780,N_24861);
and U38187 (N_38187,N_23833,N_20670);
nand U38188 (N_38188,N_25785,N_24210);
nor U38189 (N_38189,N_20804,N_29426);
and U38190 (N_38190,N_21976,N_25569);
and U38191 (N_38191,N_27288,N_26886);
nor U38192 (N_38192,N_21769,N_26639);
nor U38193 (N_38193,N_25637,N_22865);
or U38194 (N_38194,N_22280,N_25264);
and U38195 (N_38195,N_27386,N_21821);
nor U38196 (N_38196,N_20504,N_29640);
or U38197 (N_38197,N_21998,N_22108);
and U38198 (N_38198,N_27018,N_25243);
and U38199 (N_38199,N_24368,N_21089);
nand U38200 (N_38200,N_28615,N_26858);
and U38201 (N_38201,N_26003,N_29328);
or U38202 (N_38202,N_22578,N_27897);
nand U38203 (N_38203,N_25910,N_22744);
xnor U38204 (N_38204,N_27872,N_21993);
or U38205 (N_38205,N_28026,N_24695);
nor U38206 (N_38206,N_27172,N_25462);
or U38207 (N_38207,N_27670,N_24114);
nand U38208 (N_38208,N_25994,N_23690);
nand U38209 (N_38209,N_25990,N_27789);
nand U38210 (N_38210,N_27333,N_26345);
nand U38211 (N_38211,N_22717,N_28889);
xnor U38212 (N_38212,N_28150,N_24657);
or U38213 (N_38213,N_23296,N_25799);
or U38214 (N_38214,N_28397,N_27499);
nand U38215 (N_38215,N_26620,N_29147);
and U38216 (N_38216,N_21509,N_27355);
xnor U38217 (N_38217,N_20507,N_25417);
nand U38218 (N_38218,N_29772,N_26395);
and U38219 (N_38219,N_27996,N_29274);
and U38220 (N_38220,N_24769,N_20082);
and U38221 (N_38221,N_27896,N_20562);
nor U38222 (N_38222,N_28996,N_28362);
and U38223 (N_38223,N_29743,N_28134);
nand U38224 (N_38224,N_26419,N_26930);
or U38225 (N_38225,N_26915,N_27428);
and U38226 (N_38226,N_24050,N_25562);
or U38227 (N_38227,N_24355,N_29085);
nor U38228 (N_38228,N_26927,N_27912);
or U38229 (N_38229,N_27409,N_20278);
nand U38230 (N_38230,N_29764,N_23048);
nand U38231 (N_38231,N_26012,N_26257);
nor U38232 (N_38232,N_23315,N_21559);
or U38233 (N_38233,N_21093,N_20269);
nand U38234 (N_38234,N_29841,N_26365);
nor U38235 (N_38235,N_22694,N_20049);
nor U38236 (N_38236,N_20064,N_27962);
nand U38237 (N_38237,N_20851,N_24347);
nand U38238 (N_38238,N_22889,N_21383);
or U38239 (N_38239,N_21549,N_25232);
or U38240 (N_38240,N_22462,N_25564);
nand U38241 (N_38241,N_24039,N_24061);
nand U38242 (N_38242,N_25039,N_29059);
and U38243 (N_38243,N_23249,N_25542);
and U38244 (N_38244,N_29904,N_22679);
nand U38245 (N_38245,N_26179,N_28272);
nor U38246 (N_38246,N_23098,N_26835);
xor U38247 (N_38247,N_28809,N_21789);
or U38248 (N_38248,N_29941,N_26883);
and U38249 (N_38249,N_26860,N_24774);
and U38250 (N_38250,N_25638,N_21158);
nand U38251 (N_38251,N_20203,N_20820);
or U38252 (N_38252,N_20496,N_27924);
nor U38253 (N_38253,N_26811,N_23349);
or U38254 (N_38254,N_23649,N_26419);
xnor U38255 (N_38255,N_22307,N_29250);
xor U38256 (N_38256,N_23588,N_29425);
nand U38257 (N_38257,N_22502,N_21041);
nor U38258 (N_38258,N_21081,N_26937);
and U38259 (N_38259,N_20005,N_29643);
nor U38260 (N_38260,N_23227,N_29803);
nand U38261 (N_38261,N_23023,N_20887);
and U38262 (N_38262,N_28059,N_28351);
xnor U38263 (N_38263,N_28777,N_22009);
nand U38264 (N_38264,N_28665,N_20732);
xor U38265 (N_38265,N_23017,N_27228);
and U38266 (N_38266,N_28064,N_20289);
or U38267 (N_38267,N_28820,N_20056);
nand U38268 (N_38268,N_26363,N_27202);
nor U38269 (N_38269,N_20932,N_27383);
nor U38270 (N_38270,N_21145,N_25502);
nor U38271 (N_38271,N_29098,N_21482);
nand U38272 (N_38272,N_28859,N_27944);
and U38273 (N_38273,N_23398,N_22531);
and U38274 (N_38274,N_25020,N_28776);
nor U38275 (N_38275,N_27883,N_28091);
or U38276 (N_38276,N_21051,N_28686);
or U38277 (N_38277,N_20822,N_28474);
nor U38278 (N_38278,N_29595,N_25710);
or U38279 (N_38279,N_23671,N_27282);
and U38280 (N_38280,N_26702,N_29975);
nor U38281 (N_38281,N_22703,N_23627);
or U38282 (N_38282,N_23478,N_20101);
and U38283 (N_38283,N_21779,N_21898);
or U38284 (N_38284,N_28030,N_20556);
nor U38285 (N_38285,N_29677,N_27181);
nand U38286 (N_38286,N_26519,N_22342);
nand U38287 (N_38287,N_26065,N_21313);
nand U38288 (N_38288,N_29804,N_25239);
xor U38289 (N_38289,N_21550,N_27442);
nand U38290 (N_38290,N_27111,N_22461);
and U38291 (N_38291,N_23171,N_21257);
or U38292 (N_38292,N_27317,N_24403);
and U38293 (N_38293,N_26278,N_29987);
or U38294 (N_38294,N_23591,N_20002);
and U38295 (N_38295,N_27468,N_24369);
or U38296 (N_38296,N_29790,N_27735);
and U38297 (N_38297,N_21204,N_21912);
or U38298 (N_38298,N_26125,N_23141);
nor U38299 (N_38299,N_24721,N_24172);
xnor U38300 (N_38300,N_21586,N_20605);
nor U38301 (N_38301,N_22432,N_27530);
nor U38302 (N_38302,N_22372,N_28627);
nand U38303 (N_38303,N_22035,N_25762);
or U38304 (N_38304,N_23286,N_23024);
xnor U38305 (N_38305,N_24238,N_28818);
nand U38306 (N_38306,N_22336,N_25988);
and U38307 (N_38307,N_20422,N_21534);
nor U38308 (N_38308,N_26649,N_24685);
or U38309 (N_38309,N_23833,N_24889);
nor U38310 (N_38310,N_26522,N_23007);
nand U38311 (N_38311,N_29480,N_29633);
and U38312 (N_38312,N_29519,N_24479);
and U38313 (N_38313,N_27084,N_27778);
nand U38314 (N_38314,N_24132,N_27583);
nor U38315 (N_38315,N_21675,N_29041);
and U38316 (N_38316,N_21113,N_25072);
nand U38317 (N_38317,N_27009,N_28226);
nand U38318 (N_38318,N_21081,N_20625);
nand U38319 (N_38319,N_25186,N_24846);
xnor U38320 (N_38320,N_21984,N_22818);
or U38321 (N_38321,N_28615,N_21890);
nor U38322 (N_38322,N_23679,N_22412);
or U38323 (N_38323,N_20563,N_22866);
nor U38324 (N_38324,N_24927,N_25406);
xnor U38325 (N_38325,N_22604,N_24257);
and U38326 (N_38326,N_23584,N_27917);
nand U38327 (N_38327,N_26091,N_26108);
or U38328 (N_38328,N_20388,N_24084);
and U38329 (N_38329,N_22769,N_29816);
nand U38330 (N_38330,N_29382,N_28933);
nor U38331 (N_38331,N_29760,N_21816);
and U38332 (N_38332,N_26661,N_23584);
and U38333 (N_38333,N_29384,N_25469);
xnor U38334 (N_38334,N_29341,N_21021);
or U38335 (N_38335,N_24148,N_21490);
nor U38336 (N_38336,N_20995,N_23038);
and U38337 (N_38337,N_22722,N_25478);
nand U38338 (N_38338,N_23293,N_29051);
nand U38339 (N_38339,N_22494,N_28609);
or U38340 (N_38340,N_27043,N_26172);
or U38341 (N_38341,N_24672,N_29622);
nor U38342 (N_38342,N_27545,N_25327);
or U38343 (N_38343,N_22944,N_24799);
or U38344 (N_38344,N_22828,N_26172);
or U38345 (N_38345,N_20394,N_23570);
or U38346 (N_38346,N_21393,N_24769);
nor U38347 (N_38347,N_22594,N_26996);
and U38348 (N_38348,N_28642,N_29272);
or U38349 (N_38349,N_22609,N_27320);
xnor U38350 (N_38350,N_23223,N_26825);
or U38351 (N_38351,N_20577,N_22732);
nor U38352 (N_38352,N_27686,N_24581);
nand U38353 (N_38353,N_27426,N_27074);
nand U38354 (N_38354,N_24169,N_27620);
or U38355 (N_38355,N_24087,N_28151);
nor U38356 (N_38356,N_25993,N_26852);
or U38357 (N_38357,N_24907,N_20497);
or U38358 (N_38358,N_26235,N_25483);
nand U38359 (N_38359,N_25925,N_25785);
and U38360 (N_38360,N_22939,N_22955);
or U38361 (N_38361,N_23671,N_21031);
or U38362 (N_38362,N_27939,N_28086);
nor U38363 (N_38363,N_28264,N_24113);
or U38364 (N_38364,N_20904,N_27318);
xor U38365 (N_38365,N_28721,N_23586);
nor U38366 (N_38366,N_23316,N_29243);
or U38367 (N_38367,N_24437,N_26711);
xnor U38368 (N_38368,N_25934,N_24810);
nor U38369 (N_38369,N_22785,N_28664);
and U38370 (N_38370,N_23562,N_27447);
or U38371 (N_38371,N_25547,N_23221);
and U38372 (N_38372,N_29746,N_25321);
or U38373 (N_38373,N_27831,N_28707);
nor U38374 (N_38374,N_26790,N_22042);
nand U38375 (N_38375,N_27984,N_24055);
and U38376 (N_38376,N_24505,N_24076);
or U38377 (N_38377,N_23704,N_29927);
or U38378 (N_38378,N_27595,N_20113);
nor U38379 (N_38379,N_22909,N_25388);
xnor U38380 (N_38380,N_25372,N_21197);
and U38381 (N_38381,N_23000,N_23148);
or U38382 (N_38382,N_23832,N_29808);
nand U38383 (N_38383,N_29868,N_27913);
and U38384 (N_38384,N_29246,N_29393);
nor U38385 (N_38385,N_25234,N_25969);
or U38386 (N_38386,N_24668,N_29108);
nand U38387 (N_38387,N_25092,N_27936);
and U38388 (N_38388,N_27886,N_20528);
nor U38389 (N_38389,N_25162,N_27495);
and U38390 (N_38390,N_21322,N_27975);
nor U38391 (N_38391,N_29073,N_28642);
or U38392 (N_38392,N_20237,N_27437);
nand U38393 (N_38393,N_21995,N_26854);
nand U38394 (N_38394,N_27678,N_23827);
nor U38395 (N_38395,N_29593,N_24761);
or U38396 (N_38396,N_26254,N_24803);
or U38397 (N_38397,N_21174,N_22995);
xor U38398 (N_38398,N_25491,N_22603);
and U38399 (N_38399,N_24405,N_21439);
and U38400 (N_38400,N_26712,N_28415);
or U38401 (N_38401,N_25652,N_21385);
nand U38402 (N_38402,N_26496,N_27422);
xor U38403 (N_38403,N_23648,N_24833);
nor U38404 (N_38404,N_27984,N_23952);
or U38405 (N_38405,N_20334,N_23947);
and U38406 (N_38406,N_27614,N_28452);
nand U38407 (N_38407,N_27380,N_29100);
and U38408 (N_38408,N_25510,N_25466);
nor U38409 (N_38409,N_24649,N_27022);
xor U38410 (N_38410,N_22670,N_20303);
and U38411 (N_38411,N_26371,N_22257);
nand U38412 (N_38412,N_27412,N_25850);
and U38413 (N_38413,N_27186,N_24571);
or U38414 (N_38414,N_29203,N_27723);
and U38415 (N_38415,N_24599,N_25434);
and U38416 (N_38416,N_26081,N_23915);
or U38417 (N_38417,N_27705,N_27566);
or U38418 (N_38418,N_23232,N_23889);
or U38419 (N_38419,N_20587,N_22836);
and U38420 (N_38420,N_25219,N_27654);
or U38421 (N_38421,N_27812,N_20492);
xor U38422 (N_38422,N_23824,N_25916);
xnor U38423 (N_38423,N_20543,N_28047);
and U38424 (N_38424,N_25877,N_27324);
xnor U38425 (N_38425,N_24103,N_23983);
and U38426 (N_38426,N_20823,N_25328);
nand U38427 (N_38427,N_24820,N_20805);
and U38428 (N_38428,N_22082,N_21103);
or U38429 (N_38429,N_26668,N_25001);
xor U38430 (N_38430,N_23041,N_22565);
nand U38431 (N_38431,N_26875,N_28850);
nand U38432 (N_38432,N_24019,N_22017);
or U38433 (N_38433,N_27652,N_24790);
and U38434 (N_38434,N_21751,N_25528);
nand U38435 (N_38435,N_23219,N_22368);
nor U38436 (N_38436,N_21878,N_29904);
or U38437 (N_38437,N_21097,N_26612);
nor U38438 (N_38438,N_20179,N_26517);
nor U38439 (N_38439,N_26808,N_22414);
nor U38440 (N_38440,N_27201,N_23963);
and U38441 (N_38441,N_25860,N_29865);
nand U38442 (N_38442,N_25434,N_24689);
xnor U38443 (N_38443,N_20753,N_27362);
or U38444 (N_38444,N_27920,N_21545);
xnor U38445 (N_38445,N_21248,N_23796);
and U38446 (N_38446,N_20227,N_23569);
nor U38447 (N_38447,N_28741,N_24816);
or U38448 (N_38448,N_26693,N_27273);
and U38449 (N_38449,N_25564,N_21196);
nor U38450 (N_38450,N_26185,N_21629);
nor U38451 (N_38451,N_29424,N_27113);
nand U38452 (N_38452,N_23676,N_25085);
nand U38453 (N_38453,N_26772,N_25463);
nand U38454 (N_38454,N_29042,N_25636);
nand U38455 (N_38455,N_26070,N_23899);
or U38456 (N_38456,N_25403,N_20755);
and U38457 (N_38457,N_21913,N_28781);
nand U38458 (N_38458,N_27775,N_20645);
nand U38459 (N_38459,N_28224,N_26582);
and U38460 (N_38460,N_27651,N_29374);
nor U38461 (N_38461,N_29252,N_28032);
or U38462 (N_38462,N_28059,N_26862);
nand U38463 (N_38463,N_26703,N_23690);
nor U38464 (N_38464,N_23956,N_29811);
xor U38465 (N_38465,N_27986,N_27282);
nand U38466 (N_38466,N_28998,N_28314);
nand U38467 (N_38467,N_20802,N_29722);
nand U38468 (N_38468,N_20572,N_20200);
or U38469 (N_38469,N_29123,N_23505);
or U38470 (N_38470,N_29098,N_28705);
nand U38471 (N_38471,N_24772,N_22026);
or U38472 (N_38472,N_27090,N_25069);
nor U38473 (N_38473,N_29627,N_23360);
and U38474 (N_38474,N_20683,N_29824);
nand U38475 (N_38475,N_29661,N_20027);
or U38476 (N_38476,N_26029,N_20764);
nor U38477 (N_38477,N_23336,N_29339);
nor U38478 (N_38478,N_20667,N_29515);
or U38479 (N_38479,N_29983,N_25651);
nor U38480 (N_38480,N_24372,N_22894);
and U38481 (N_38481,N_25007,N_21127);
or U38482 (N_38482,N_29535,N_20268);
nor U38483 (N_38483,N_27619,N_28298);
nor U38484 (N_38484,N_29901,N_24443);
nor U38485 (N_38485,N_25944,N_20497);
and U38486 (N_38486,N_20896,N_29160);
or U38487 (N_38487,N_29314,N_26240);
nand U38488 (N_38488,N_21218,N_20133);
nand U38489 (N_38489,N_28546,N_25528);
nand U38490 (N_38490,N_27661,N_24260);
nand U38491 (N_38491,N_20736,N_29233);
xor U38492 (N_38492,N_23881,N_27873);
nand U38493 (N_38493,N_25999,N_22164);
or U38494 (N_38494,N_20349,N_25536);
and U38495 (N_38495,N_22302,N_23910);
xor U38496 (N_38496,N_24644,N_26207);
xnor U38497 (N_38497,N_25371,N_29002);
nand U38498 (N_38498,N_20001,N_21941);
nor U38499 (N_38499,N_25520,N_23268);
nor U38500 (N_38500,N_22210,N_20519);
nand U38501 (N_38501,N_28175,N_28942);
nand U38502 (N_38502,N_29057,N_29343);
nor U38503 (N_38503,N_21071,N_21255);
or U38504 (N_38504,N_25971,N_28628);
nor U38505 (N_38505,N_29578,N_24690);
and U38506 (N_38506,N_20358,N_20153);
xnor U38507 (N_38507,N_21100,N_21370);
or U38508 (N_38508,N_21460,N_20137);
or U38509 (N_38509,N_20388,N_26566);
nor U38510 (N_38510,N_26044,N_28987);
or U38511 (N_38511,N_23060,N_29208);
and U38512 (N_38512,N_23752,N_28523);
xnor U38513 (N_38513,N_21378,N_27869);
nand U38514 (N_38514,N_28247,N_29273);
and U38515 (N_38515,N_23431,N_22483);
nand U38516 (N_38516,N_22283,N_27407);
nand U38517 (N_38517,N_28551,N_29965);
nand U38518 (N_38518,N_29648,N_28230);
xor U38519 (N_38519,N_27994,N_21860);
xnor U38520 (N_38520,N_26192,N_22630);
and U38521 (N_38521,N_20719,N_25496);
or U38522 (N_38522,N_21798,N_27972);
or U38523 (N_38523,N_22334,N_27383);
and U38524 (N_38524,N_27626,N_26104);
or U38525 (N_38525,N_23023,N_25886);
nand U38526 (N_38526,N_25056,N_23010);
xnor U38527 (N_38527,N_27496,N_27543);
or U38528 (N_38528,N_24789,N_26863);
and U38529 (N_38529,N_28854,N_22959);
and U38530 (N_38530,N_23728,N_22481);
or U38531 (N_38531,N_20501,N_29505);
xor U38532 (N_38532,N_25622,N_20271);
or U38533 (N_38533,N_27770,N_20290);
nand U38534 (N_38534,N_28154,N_29487);
and U38535 (N_38535,N_20177,N_22194);
nor U38536 (N_38536,N_26885,N_29934);
nand U38537 (N_38537,N_20856,N_24420);
xor U38538 (N_38538,N_24135,N_29512);
or U38539 (N_38539,N_20118,N_22817);
or U38540 (N_38540,N_24495,N_24444);
or U38541 (N_38541,N_23099,N_24829);
xnor U38542 (N_38542,N_28915,N_27391);
xnor U38543 (N_38543,N_21846,N_27289);
or U38544 (N_38544,N_25549,N_20053);
nor U38545 (N_38545,N_29633,N_21512);
or U38546 (N_38546,N_21293,N_26042);
or U38547 (N_38547,N_27955,N_21620);
nor U38548 (N_38548,N_24489,N_28175);
nor U38549 (N_38549,N_20452,N_29064);
nand U38550 (N_38550,N_20599,N_25671);
and U38551 (N_38551,N_26691,N_25501);
nor U38552 (N_38552,N_29908,N_23790);
or U38553 (N_38553,N_26916,N_22036);
or U38554 (N_38554,N_27095,N_22111);
or U38555 (N_38555,N_20050,N_29480);
or U38556 (N_38556,N_26506,N_23194);
or U38557 (N_38557,N_20690,N_23459);
nand U38558 (N_38558,N_20684,N_23997);
and U38559 (N_38559,N_25090,N_29929);
xor U38560 (N_38560,N_25464,N_27633);
nor U38561 (N_38561,N_24889,N_21450);
xnor U38562 (N_38562,N_20812,N_23452);
or U38563 (N_38563,N_29786,N_27972);
nand U38564 (N_38564,N_28394,N_25872);
nand U38565 (N_38565,N_24795,N_24251);
or U38566 (N_38566,N_29363,N_27964);
nor U38567 (N_38567,N_26749,N_29819);
nor U38568 (N_38568,N_29685,N_25120);
or U38569 (N_38569,N_26912,N_29866);
nand U38570 (N_38570,N_23976,N_24638);
and U38571 (N_38571,N_25884,N_27830);
nand U38572 (N_38572,N_26263,N_27841);
nor U38573 (N_38573,N_25784,N_21704);
nor U38574 (N_38574,N_20463,N_28411);
and U38575 (N_38575,N_25630,N_24818);
xor U38576 (N_38576,N_27408,N_29330);
nor U38577 (N_38577,N_25456,N_24784);
nor U38578 (N_38578,N_20455,N_22301);
nand U38579 (N_38579,N_21157,N_25815);
nand U38580 (N_38580,N_21256,N_22164);
and U38581 (N_38581,N_25260,N_26410);
nor U38582 (N_38582,N_22730,N_28278);
and U38583 (N_38583,N_24121,N_24390);
nor U38584 (N_38584,N_24221,N_21608);
nor U38585 (N_38585,N_24167,N_20888);
nand U38586 (N_38586,N_23354,N_22756);
and U38587 (N_38587,N_27774,N_22383);
nand U38588 (N_38588,N_23804,N_24176);
nand U38589 (N_38589,N_20478,N_22959);
nand U38590 (N_38590,N_27243,N_23425);
nor U38591 (N_38591,N_24756,N_21682);
nand U38592 (N_38592,N_25090,N_24536);
or U38593 (N_38593,N_27672,N_26766);
nor U38594 (N_38594,N_20641,N_28481);
or U38595 (N_38595,N_28557,N_29263);
and U38596 (N_38596,N_28743,N_21574);
and U38597 (N_38597,N_24357,N_24860);
nand U38598 (N_38598,N_23217,N_29987);
nand U38599 (N_38599,N_22703,N_28784);
nand U38600 (N_38600,N_22851,N_27556);
nand U38601 (N_38601,N_23300,N_24288);
xnor U38602 (N_38602,N_27418,N_26655);
and U38603 (N_38603,N_27351,N_22394);
nand U38604 (N_38604,N_22533,N_28704);
nor U38605 (N_38605,N_21834,N_29976);
xor U38606 (N_38606,N_20464,N_28377);
nor U38607 (N_38607,N_28958,N_22497);
and U38608 (N_38608,N_27129,N_27978);
or U38609 (N_38609,N_29034,N_24305);
nand U38610 (N_38610,N_21778,N_20976);
nor U38611 (N_38611,N_23674,N_29116);
xnor U38612 (N_38612,N_29752,N_27272);
or U38613 (N_38613,N_26057,N_27176);
nor U38614 (N_38614,N_28702,N_21404);
nor U38615 (N_38615,N_29454,N_28251);
and U38616 (N_38616,N_25943,N_22412);
nand U38617 (N_38617,N_26259,N_24880);
and U38618 (N_38618,N_24666,N_20322);
nand U38619 (N_38619,N_20145,N_25466);
nor U38620 (N_38620,N_22104,N_21369);
and U38621 (N_38621,N_28238,N_28171);
and U38622 (N_38622,N_24463,N_20062);
and U38623 (N_38623,N_29777,N_22905);
nand U38624 (N_38624,N_22216,N_29580);
nor U38625 (N_38625,N_24116,N_22701);
xor U38626 (N_38626,N_26190,N_25721);
nor U38627 (N_38627,N_21267,N_20588);
nand U38628 (N_38628,N_20297,N_22375);
and U38629 (N_38629,N_22549,N_20650);
xnor U38630 (N_38630,N_24399,N_20573);
xor U38631 (N_38631,N_24298,N_25070);
and U38632 (N_38632,N_26357,N_27399);
nand U38633 (N_38633,N_28829,N_21433);
or U38634 (N_38634,N_21876,N_21455);
nor U38635 (N_38635,N_23124,N_22864);
nand U38636 (N_38636,N_26896,N_24175);
nor U38637 (N_38637,N_24587,N_28402);
nand U38638 (N_38638,N_29589,N_24574);
nor U38639 (N_38639,N_26474,N_23777);
nand U38640 (N_38640,N_26074,N_25755);
and U38641 (N_38641,N_20058,N_22876);
or U38642 (N_38642,N_22566,N_29933);
nand U38643 (N_38643,N_28848,N_27295);
and U38644 (N_38644,N_26903,N_28683);
nor U38645 (N_38645,N_22976,N_25487);
xor U38646 (N_38646,N_25647,N_25692);
nor U38647 (N_38647,N_23444,N_27306);
and U38648 (N_38648,N_24582,N_20104);
or U38649 (N_38649,N_20087,N_29116);
nor U38650 (N_38650,N_24742,N_29951);
nand U38651 (N_38651,N_22485,N_24289);
nor U38652 (N_38652,N_20404,N_26616);
nand U38653 (N_38653,N_27060,N_27762);
nor U38654 (N_38654,N_20585,N_21594);
nor U38655 (N_38655,N_24604,N_26883);
nor U38656 (N_38656,N_21176,N_22364);
xnor U38657 (N_38657,N_20841,N_28500);
and U38658 (N_38658,N_28354,N_20982);
or U38659 (N_38659,N_29949,N_28328);
nand U38660 (N_38660,N_24840,N_29258);
nor U38661 (N_38661,N_27422,N_26568);
nor U38662 (N_38662,N_23046,N_22903);
xor U38663 (N_38663,N_29293,N_25850);
nor U38664 (N_38664,N_21580,N_28252);
or U38665 (N_38665,N_21350,N_20903);
nand U38666 (N_38666,N_25304,N_23455);
nor U38667 (N_38667,N_25879,N_27493);
and U38668 (N_38668,N_21123,N_23953);
nor U38669 (N_38669,N_20193,N_25493);
nor U38670 (N_38670,N_21814,N_28811);
or U38671 (N_38671,N_29632,N_28316);
nand U38672 (N_38672,N_26745,N_25949);
nor U38673 (N_38673,N_26529,N_26212);
or U38674 (N_38674,N_25956,N_21042);
nand U38675 (N_38675,N_26011,N_26470);
nand U38676 (N_38676,N_21075,N_25803);
nor U38677 (N_38677,N_21136,N_20510);
nand U38678 (N_38678,N_26553,N_25278);
and U38679 (N_38679,N_22790,N_21741);
nand U38680 (N_38680,N_25564,N_29612);
or U38681 (N_38681,N_22634,N_23909);
or U38682 (N_38682,N_21310,N_28153);
and U38683 (N_38683,N_22159,N_26564);
or U38684 (N_38684,N_20731,N_27924);
or U38685 (N_38685,N_20394,N_22785);
xor U38686 (N_38686,N_21056,N_20774);
nand U38687 (N_38687,N_24164,N_26134);
and U38688 (N_38688,N_29425,N_24338);
and U38689 (N_38689,N_22707,N_24741);
nand U38690 (N_38690,N_20802,N_25028);
or U38691 (N_38691,N_23341,N_26975);
or U38692 (N_38692,N_25673,N_21536);
nand U38693 (N_38693,N_22962,N_28211);
nand U38694 (N_38694,N_24756,N_25632);
or U38695 (N_38695,N_24660,N_24288);
and U38696 (N_38696,N_26433,N_23096);
and U38697 (N_38697,N_29169,N_22921);
nor U38698 (N_38698,N_26032,N_28911);
nor U38699 (N_38699,N_20525,N_24991);
nor U38700 (N_38700,N_24229,N_28495);
nor U38701 (N_38701,N_29926,N_25755);
and U38702 (N_38702,N_26759,N_23154);
nand U38703 (N_38703,N_27393,N_27108);
or U38704 (N_38704,N_24849,N_20099);
nor U38705 (N_38705,N_23624,N_28908);
or U38706 (N_38706,N_23886,N_25833);
and U38707 (N_38707,N_29505,N_26956);
nor U38708 (N_38708,N_28819,N_20352);
nor U38709 (N_38709,N_21870,N_26073);
and U38710 (N_38710,N_21905,N_24034);
and U38711 (N_38711,N_26677,N_21992);
and U38712 (N_38712,N_21351,N_23682);
nor U38713 (N_38713,N_29327,N_28559);
and U38714 (N_38714,N_27890,N_25950);
and U38715 (N_38715,N_28484,N_23473);
or U38716 (N_38716,N_29140,N_28103);
or U38717 (N_38717,N_22255,N_27734);
nand U38718 (N_38718,N_29765,N_23822);
nor U38719 (N_38719,N_20004,N_24917);
and U38720 (N_38720,N_25726,N_27768);
or U38721 (N_38721,N_24609,N_29415);
xnor U38722 (N_38722,N_27987,N_29623);
nor U38723 (N_38723,N_24442,N_23330);
xor U38724 (N_38724,N_23337,N_26120);
and U38725 (N_38725,N_23476,N_22259);
nor U38726 (N_38726,N_21066,N_20208);
nor U38727 (N_38727,N_25902,N_22563);
nor U38728 (N_38728,N_26761,N_28277);
nor U38729 (N_38729,N_29728,N_23082);
nor U38730 (N_38730,N_27179,N_27266);
xor U38731 (N_38731,N_21836,N_25301);
and U38732 (N_38732,N_23627,N_26518);
and U38733 (N_38733,N_29930,N_27111);
xnor U38734 (N_38734,N_29890,N_22575);
nand U38735 (N_38735,N_28682,N_28374);
nor U38736 (N_38736,N_20014,N_29281);
xor U38737 (N_38737,N_26596,N_20239);
nand U38738 (N_38738,N_29412,N_25687);
and U38739 (N_38739,N_25244,N_22965);
or U38740 (N_38740,N_25795,N_20280);
and U38741 (N_38741,N_26240,N_20997);
nand U38742 (N_38742,N_25079,N_22374);
nand U38743 (N_38743,N_22771,N_23696);
and U38744 (N_38744,N_26456,N_26943);
xnor U38745 (N_38745,N_27625,N_23006);
nand U38746 (N_38746,N_23998,N_27105);
and U38747 (N_38747,N_29473,N_29239);
nand U38748 (N_38748,N_24126,N_24390);
nand U38749 (N_38749,N_25282,N_21756);
or U38750 (N_38750,N_27972,N_24980);
and U38751 (N_38751,N_21840,N_28369);
nor U38752 (N_38752,N_27995,N_22236);
xnor U38753 (N_38753,N_28582,N_24072);
or U38754 (N_38754,N_24019,N_24871);
or U38755 (N_38755,N_22007,N_20175);
nand U38756 (N_38756,N_24556,N_20461);
nor U38757 (N_38757,N_21644,N_27336);
nor U38758 (N_38758,N_21123,N_29492);
nor U38759 (N_38759,N_23871,N_23739);
or U38760 (N_38760,N_26135,N_29692);
or U38761 (N_38761,N_26467,N_22744);
and U38762 (N_38762,N_27616,N_23596);
nor U38763 (N_38763,N_21197,N_21413);
nor U38764 (N_38764,N_21216,N_24351);
nor U38765 (N_38765,N_26178,N_23746);
nor U38766 (N_38766,N_21592,N_29761);
and U38767 (N_38767,N_28650,N_26916);
or U38768 (N_38768,N_24211,N_27292);
xnor U38769 (N_38769,N_29487,N_24721);
nor U38770 (N_38770,N_24480,N_21304);
and U38771 (N_38771,N_24170,N_28860);
nand U38772 (N_38772,N_25211,N_24703);
or U38773 (N_38773,N_27242,N_25671);
nand U38774 (N_38774,N_29960,N_29528);
xnor U38775 (N_38775,N_24702,N_28882);
and U38776 (N_38776,N_28299,N_21837);
xor U38777 (N_38777,N_23387,N_24961);
and U38778 (N_38778,N_20506,N_25037);
or U38779 (N_38779,N_25558,N_26441);
nor U38780 (N_38780,N_26362,N_20514);
nand U38781 (N_38781,N_26320,N_22676);
and U38782 (N_38782,N_29976,N_25133);
nor U38783 (N_38783,N_24324,N_29361);
nand U38784 (N_38784,N_22367,N_25545);
nor U38785 (N_38785,N_20303,N_28943);
or U38786 (N_38786,N_26974,N_24387);
nand U38787 (N_38787,N_27847,N_22070);
and U38788 (N_38788,N_20916,N_25381);
nor U38789 (N_38789,N_24151,N_28265);
nor U38790 (N_38790,N_28845,N_21706);
xnor U38791 (N_38791,N_21978,N_25666);
and U38792 (N_38792,N_25895,N_29666);
nor U38793 (N_38793,N_26451,N_26677);
or U38794 (N_38794,N_29520,N_23701);
or U38795 (N_38795,N_22563,N_21884);
xnor U38796 (N_38796,N_29498,N_26471);
nand U38797 (N_38797,N_24185,N_28812);
nand U38798 (N_38798,N_28741,N_22912);
nand U38799 (N_38799,N_21640,N_26541);
or U38800 (N_38800,N_22181,N_25579);
nand U38801 (N_38801,N_25987,N_27790);
or U38802 (N_38802,N_24929,N_29356);
and U38803 (N_38803,N_25664,N_29834);
nand U38804 (N_38804,N_27232,N_29638);
xor U38805 (N_38805,N_22500,N_24189);
nor U38806 (N_38806,N_21036,N_24699);
or U38807 (N_38807,N_21747,N_29135);
or U38808 (N_38808,N_24821,N_23212);
nor U38809 (N_38809,N_24145,N_26831);
nor U38810 (N_38810,N_23415,N_28446);
and U38811 (N_38811,N_28555,N_29233);
and U38812 (N_38812,N_24726,N_25945);
nand U38813 (N_38813,N_26471,N_29517);
nand U38814 (N_38814,N_24278,N_20762);
and U38815 (N_38815,N_26929,N_24967);
xnor U38816 (N_38816,N_22469,N_25378);
and U38817 (N_38817,N_22958,N_20809);
and U38818 (N_38818,N_25172,N_22979);
and U38819 (N_38819,N_22998,N_27521);
nand U38820 (N_38820,N_24805,N_27768);
or U38821 (N_38821,N_22584,N_22647);
and U38822 (N_38822,N_25476,N_27606);
nand U38823 (N_38823,N_22019,N_21473);
nand U38824 (N_38824,N_20126,N_27189);
and U38825 (N_38825,N_27942,N_20306);
xnor U38826 (N_38826,N_22056,N_27123);
and U38827 (N_38827,N_22275,N_29486);
nor U38828 (N_38828,N_29471,N_29411);
and U38829 (N_38829,N_21175,N_21162);
and U38830 (N_38830,N_29425,N_28976);
xnor U38831 (N_38831,N_20502,N_29538);
xnor U38832 (N_38832,N_24553,N_27976);
or U38833 (N_38833,N_22931,N_24740);
nor U38834 (N_38834,N_29979,N_23621);
or U38835 (N_38835,N_20110,N_20683);
or U38836 (N_38836,N_25873,N_20529);
nand U38837 (N_38837,N_24363,N_29318);
and U38838 (N_38838,N_21472,N_23532);
xor U38839 (N_38839,N_26668,N_21130);
nand U38840 (N_38840,N_27182,N_29325);
nor U38841 (N_38841,N_23900,N_20294);
nor U38842 (N_38842,N_22980,N_24437);
or U38843 (N_38843,N_21576,N_24847);
and U38844 (N_38844,N_26486,N_28478);
nor U38845 (N_38845,N_20061,N_28425);
or U38846 (N_38846,N_25422,N_27765);
or U38847 (N_38847,N_20343,N_26512);
nand U38848 (N_38848,N_25838,N_24284);
and U38849 (N_38849,N_20231,N_20258);
xnor U38850 (N_38850,N_29918,N_29364);
and U38851 (N_38851,N_25734,N_21519);
nor U38852 (N_38852,N_21643,N_20723);
nand U38853 (N_38853,N_23388,N_22836);
nor U38854 (N_38854,N_20007,N_20119);
nor U38855 (N_38855,N_24120,N_20279);
nor U38856 (N_38856,N_24492,N_20656);
and U38857 (N_38857,N_23796,N_21578);
and U38858 (N_38858,N_21041,N_26512);
and U38859 (N_38859,N_25311,N_28588);
nor U38860 (N_38860,N_26266,N_21819);
or U38861 (N_38861,N_26830,N_26754);
nor U38862 (N_38862,N_25955,N_20447);
nand U38863 (N_38863,N_28455,N_29093);
nor U38864 (N_38864,N_23976,N_22294);
xor U38865 (N_38865,N_22946,N_27675);
or U38866 (N_38866,N_24537,N_28549);
and U38867 (N_38867,N_28000,N_22471);
nor U38868 (N_38868,N_28631,N_27225);
nor U38869 (N_38869,N_22507,N_23076);
nand U38870 (N_38870,N_20571,N_24033);
and U38871 (N_38871,N_25118,N_28173);
xor U38872 (N_38872,N_29733,N_28621);
xnor U38873 (N_38873,N_25857,N_28099);
nor U38874 (N_38874,N_25917,N_25273);
and U38875 (N_38875,N_22900,N_28994);
and U38876 (N_38876,N_28359,N_22899);
and U38877 (N_38877,N_28350,N_26358);
nand U38878 (N_38878,N_20178,N_21674);
nand U38879 (N_38879,N_29487,N_26640);
nor U38880 (N_38880,N_24736,N_26985);
nor U38881 (N_38881,N_29408,N_22655);
and U38882 (N_38882,N_22850,N_25378);
or U38883 (N_38883,N_20058,N_27318);
or U38884 (N_38884,N_23073,N_29264);
or U38885 (N_38885,N_20283,N_28114);
and U38886 (N_38886,N_24171,N_27035);
or U38887 (N_38887,N_25163,N_22453);
and U38888 (N_38888,N_27118,N_27049);
and U38889 (N_38889,N_25371,N_26011);
nor U38890 (N_38890,N_24187,N_23458);
or U38891 (N_38891,N_21454,N_29243);
nand U38892 (N_38892,N_27323,N_23314);
xnor U38893 (N_38893,N_20973,N_20502);
nor U38894 (N_38894,N_29462,N_21493);
xor U38895 (N_38895,N_29196,N_29158);
and U38896 (N_38896,N_28540,N_22648);
or U38897 (N_38897,N_27980,N_20216);
or U38898 (N_38898,N_20644,N_24774);
and U38899 (N_38899,N_20016,N_28623);
nor U38900 (N_38900,N_20031,N_20522);
xnor U38901 (N_38901,N_27765,N_20531);
xor U38902 (N_38902,N_20552,N_24129);
nor U38903 (N_38903,N_27585,N_25389);
xor U38904 (N_38904,N_25399,N_29458);
and U38905 (N_38905,N_24925,N_27405);
xor U38906 (N_38906,N_20813,N_25399);
xnor U38907 (N_38907,N_25215,N_28515);
nand U38908 (N_38908,N_22700,N_27884);
or U38909 (N_38909,N_25171,N_21402);
nand U38910 (N_38910,N_20436,N_25925);
xor U38911 (N_38911,N_21984,N_23638);
nand U38912 (N_38912,N_20561,N_21544);
nand U38913 (N_38913,N_29640,N_23814);
nand U38914 (N_38914,N_23439,N_25919);
or U38915 (N_38915,N_20600,N_27513);
and U38916 (N_38916,N_24505,N_24397);
nor U38917 (N_38917,N_29705,N_27795);
nor U38918 (N_38918,N_24375,N_22301);
nor U38919 (N_38919,N_28479,N_23222);
and U38920 (N_38920,N_25916,N_26977);
and U38921 (N_38921,N_21413,N_22943);
or U38922 (N_38922,N_27674,N_21256);
and U38923 (N_38923,N_22607,N_29791);
or U38924 (N_38924,N_21396,N_28147);
or U38925 (N_38925,N_23558,N_22253);
nor U38926 (N_38926,N_24967,N_29452);
nand U38927 (N_38927,N_22700,N_27486);
or U38928 (N_38928,N_27547,N_23309);
and U38929 (N_38929,N_26076,N_25435);
or U38930 (N_38930,N_25060,N_25869);
nor U38931 (N_38931,N_21700,N_23275);
and U38932 (N_38932,N_27210,N_29249);
or U38933 (N_38933,N_29925,N_22254);
nand U38934 (N_38934,N_29917,N_24387);
nand U38935 (N_38935,N_21731,N_26872);
and U38936 (N_38936,N_25651,N_24560);
nand U38937 (N_38937,N_20972,N_23495);
and U38938 (N_38938,N_27208,N_21660);
nand U38939 (N_38939,N_25538,N_27464);
nor U38940 (N_38940,N_21973,N_28028);
and U38941 (N_38941,N_28226,N_23418);
nor U38942 (N_38942,N_28695,N_26593);
nand U38943 (N_38943,N_26685,N_20987);
nor U38944 (N_38944,N_24917,N_29042);
xor U38945 (N_38945,N_23672,N_23969);
nor U38946 (N_38946,N_21428,N_20952);
nand U38947 (N_38947,N_25215,N_20978);
nand U38948 (N_38948,N_22945,N_26261);
or U38949 (N_38949,N_24955,N_20590);
nand U38950 (N_38950,N_22928,N_25653);
and U38951 (N_38951,N_28778,N_26496);
xor U38952 (N_38952,N_28894,N_25422);
or U38953 (N_38953,N_21801,N_26863);
and U38954 (N_38954,N_29647,N_21024);
nand U38955 (N_38955,N_29283,N_20350);
and U38956 (N_38956,N_22678,N_29779);
xnor U38957 (N_38957,N_27632,N_27084);
xnor U38958 (N_38958,N_26140,N_29185);
or U38959 (N_38959,N_21500,N_20637);
nand U38960 (N_38960,N_20811,N_27152);
nand U38961 (N_38961,N_22568,N_27278);
nand U38962 (N_38962,N_26496,N_29435);
nor U38963 (N_38963,N_29020,N_20925);
nand U38964 (N_38964,N_23620,N_23948);
or U38965 (N_38965,N_24174,N_26780);
and U38966 (N_38966,N_25410,N_27412);
or U38967 (N_38967,N_25086,N_28813);
xnor U38968 (N_38968,N_27920,N_24739);
or U38969 (N_38969,N_27706,N_29904);
nand U38970 (N_38970,N_29276,N_28054);
nand U38971 (N_38971,N_28827,N_27412);
nand U38972 (N_38972,N_23858,N_28150);
and U38973 (N_38973,N_28401,N_24340);
or U38974 (N_38974,N_27651,N_27921);
and U38975 (N_38975,N_21177,N_29582);
and U38976 (N_38976,N_21179,N_24578);
nor U38977 (N_38977,N_29421,N_28518);
or U38978 (N_38978,N_29052,N_28149);
nor U38979 (N_38979,N_20181,N_21308);
nand U38980 (N_38980,N_24436,N_29719);
nor U38981 (N_38981,N_26749,N_22403);
xor U38982 (N_38982,N_20227,N_21926);
or U38983 (N_38983,N_29936,N_24978);
or U38984 (N_38984,N_26581,N_28353);
xor U38985 (N_38985,N_25778,N_23457);
or U38986 (N_38986,N_21044,N_21908);
nand U38987 (N_38987,N_23531,N_26537);
nor U38988 (N_38988,N_22371,N_26362);
nand U38989 (N_38989,N_25033,N_24489);
nor U38990 (N_38990,N_29910,N_29034);
xnor U38991 (N_38991,N_20843,N_23613);
nor U38992 (N_38992,N_23758,N_26214);
and U38993 (N_38993,N_27887,N_21339);
and U38994 (N_38994,N_27877,N_29294);
or U38995 (N_38995,N_27027,N_29620);
or U38996 (N_38996,N_26752,N_22220);
nand U38997 (N_38997,N_21585,N_25695);
or U38998 (N_38998,N_23393,N_25823);
or U38999 (N_38999,N_22455,N_22870);
nand U39000 (N_39000,N_27992,N_21600);
xor U39001 (N_39001,N_22489,N_29790);
or U39002 (N_39002,N_20076,N_24549);
or U39003 (N_39003,N_29566,N_20501);
xnor U39004 (N_39004,N_26501,N_22571);
nand U39005 (N_39005,N_26079,N_24461);
and U39006 (N_39006,N_26774,N_23113);
nand U39007 (N_39007,N_29264,N_25827);
nand U39008 (N_39008,N_23934,N_21610);
nand U39009 (N_39009,N_26673,N_24811);
xnor U39010 (N_39010,N_27825,N_25311);
nand U39011 (N_39011,N_28852,N_26342);
nor U39012 (N_39012,N_28596,N_22114);
or U39013 (N_39013,N_20671,N_23352);
nor U39014 (N_39014,N_28594,N_23535);
nor U39015 (N_39015,N_28722,N_25279);
or U39016 (N_39016,N_20473,N_25583);
or U39017 (N_39017,N_26493,N_26492);
or U39018 (N_39018,N_27696,N_26303);
nand U39019 (N_39019,N_25591,N_23637);
or U39020 (N_39020,N_26025,N_28594);
nand U39021 (N_39021,N_22127,N_22882);
xor U39022 (N_39022,N_29393,N_25926);
nand U39023 (N_39023,N_28202,N_25210);
xnor U39024 (N_39024,N_23954,N_26709);
and U39025 (N_39025,N_25896,N_24332);
nand U39026 (N_39026,N_22135,N_22702);
and U39027 (N_39027,N_22312,N_28879);
or U39028 (N_39028,N_25315,N_22993);
xnor U39029 (N_39029,N_22610,N_27250);
or U39030 (N_39030,N_28720,N_28495);
nand U39031 (N_39031,N_22148,N_20241);
or U39032 (N_39032,N_21001,N_29097);
and U39033 (N_39033,N_23260,N_23019);
or U39034 (N_39034,N_27052,N_23999);
or U39035 (N_39035,N_25083,N_27468);
nand U39036 (N_39036,N_25846,N_21092);
or U39037 (N_39037,N_28461,N_27319);
or U39038 (N_39038,N_20300,N_22159);
or U39039 (N_39039,N_26510,N_27249);
and U39040 (N_39040,N_24041,N_25542);
nor U39041 (N_39041,N_23230,N_29768);
and U39042 (N_39042,N_21615,N_24899);
or U39043 (N_39043,N_20639,N_24169);
nand U39044 (N_39044,N_29142,N_29998);
or U39045 (N_39045,N_20320,N_20809);
xnor U39046 (N_39046,N_21172,N_23795);
and U39047 (N_39047,N_27627,N_23319);
nand U39048 (N_39048,N_29129,N_24549);
nand U39049 (N_39049,N_27781,N_28697);
or U39050 (N_39050,N_20088,N_20676);
or U39051 (N_39051,N_22396,N_29873);
and U39052 (N_39052,N_23517,N_24123);
and U39053 (N_39053,N_28394,N_29601);
xnor U39054 (N_39054,N_27739,N_24428);
and U39055 (N_39055,N_27313,N_27119);
xor U39056 (N_39056,N_25350,N_29990);
and U39057 (N_39057,N_29226,N_23268);
xor U39058 (N_39058,N_21589,N_28287);
or U39059 (N_39059,N_23889,N_26854);
nand U39060 (N_39060,N_22270,N_24997);
xnor U39061 (N_39061,N_26776,N_21400);
and U39062 (N_39062,N_25921,N_25696);
nor U39063 (N_39063,N_25138,N_23364);
or U39064 (N_39064,N_21509,N_26448);
nor U39065 (N_39065,N_21475,N_20216);
nand U39066 (N_39066,N_21715,N_25957);
xor U39067 (N_39067,N_29462,N_25815);
nor U39068 (N_39068,N_22962,N_29100);
or U39069 (N_39069,N_26787,N_21734);
and U39070 (N_39070,N_25494,N_29515);
or U39071 (N_39071,N_23236,N_22069);
and U39072 (N_39072,N_29424,N_25774);
nor U39073 (N_39073,N_24830,N_24212);
nor U39074 (N_39074,N_25082,N_28795);
or U39075 (N_39075,N_24050,N_24983);
and U39076 (N_39076,N_25192,N_25669);
nand U39077 (N_39077,N_20464,N_22967);
or U39078 (N_39078,N_23088,N_24511);
or U39079 (N_39079,N_23202,N_23568);
or U39080 (N_39080,N_20114,N_23256);
xnor U39081 (N_39081,N_24735,N_26751);
xnor U39082 (N_39082,N_26551,N_25774);
and U39083 (N_39083,N_29183,N_27580);
nor U39084 (N_39084,N_28378,N_26289);
nand U39085 (N_39085,N_24275,N_21613);
and U39086 (N_39086,N_27116,N_28179);
or U39087 (N_39087,N_26883,N_23874);
and U39088 (N_39088,N_29179,N_27128);
nor U39089 (N_39089,N_24763,N_20964);
and U39090 (N_39090,N_20905,N_29038);
nand U39091 (N_39091,N_21469,N_24024);
or U39092 (N_39092,N_22156,N_20534);
nand U39093 (N_39093,N_23273,N_25294);
and U39094 (N_39094,N_29435,N_24434);
nand U39095 (N_39095,N_21382,N_21372);
or U39096 (N_39096,N_22101,N_29532);
or U39097 (N_39097,N_22931,N_25082);
and U39098 (N_39098,N_29460,N_28708);
nor U39099 (N_39099,N_28493,N_25279);
and U39100 (N_39100,N_20362,N_24683);
or U39101 (N_39101,N_25873,N_25311);
nand U39102 (N_39102,N_21773,N_27539);
and U39103 (N_39103,N_22491,N_22201);
or U39104 (N_39104,N_24388,N_26210);
xor U39105 (N_39105,N_23232,N_24257);
or U39106 (N_39106,N_21683,N_20130);
nor U39107 (N_39107,N_25881,N_28410);
and U39108 (N_39108,N_21226,N_24898);
nor U39109 (N_39109,N_20996,N_27716);
or U39110 (N_39110,N_20457,N_25038);
or U39111 (N_39111,N_28019,N_25550);
nand U39112 (N_39112,N_25003,N_23380);
nor U39113 (N_39113,N_23374,N_21894);
nand U39114 (N_39114,N_26313,N_21170);
or U39115 (N_39115,N_22139,N_26756);
nand U39116 (N_39116,N_29135,N_23928);
or U39117 (N_39117,N_28462,N_26600);
and U39118 (N_39118,N_20966,N_20112);
and U39119 (N_39119,N_25507,N_20923);
nor U39120 (N_39120,N_21250,N_27245);
nand U39121 (N_39121,N_28550,N_28453);
nand U39122 (N_39122,N_25466,N_28242);
nor U39123 (N_39123,N_24101,N_21406);
or U39124 (N_39124,N_27668,N_23244);
nor U39125 (N_39125,N_23210,N_22758);
or U39126 (N_39126,N_25637,N_24231);
or U39127 (N_39127,N_22676,N_28029);
nand U39128 (N_39128,N_27176,N_21928);
nor U39129 (N_39129,N_29196,N_20138);
or U39130 (N_39130,N_22210,N_27123);
or U39131 (N_39131,N_20800,N_26798);
nor U39132 (N_39132,N_26109,N_28600);
or U39133 (N_39133,N_24173,N_27179);
xnor U39134 (N_39134,N_22345,N_28136);
xor U39135 (N_39135,N_25119,N_20664);
and U39136 (N_39136,N_21103,N_21947);
and U39137 (N_39137,N_23785,N_28583);
or U39138 (N_39138,N_22593,N_21249);
nor U39139 (N_39139,N_26915,N_23206);
nand U39140 (N_39140,N_28861,N_20321);
nor U39141 (N_39141,N_29700,N_29685);
nor U39142 (N_39142,N_28837,N_25582);
or U39143 (N_39143,N_27556,N_29486);
nand U39144 (N_39144,N_28139,N_29410);
nand U39145 (N_39145,N_22020,N_21910);
or U39146 (N_39146,N_28235,N_22223);
or U39147 (N_39147,N_25854,N_22721);
and U39148 (N_39148,N_24909,N_26415);
and U39149 (N_39149,N_28349,N_29287);
nand U39150 (N_39150,N_21848,N_24723);
and U39151 (N_39151,N_28468,N_24257);
and U39152 (N_39152,N_23157,N_20949);
nor U39153 (N_39153,N_29885,N_21626);
or U39154 (N_39154,N_22085,N_24311);
and U39155 (N_39155,N_23722,N_28387);
xnor U39156 (N_39156,N_23057,N_23299);
nor U39157 (N_39157,N_20192,N_25287);
nor U39158 (N_39158,N_20989,N_21037);
nor U39159 (N_39159,N_29014,N_24340);
and U39160 (N_39160,N_22739,N_23126);
nand U39161 (N_39161,N_20209,N_25996);
nand U39162 (N_39162,N_28287,N_20972);
nor U39163 (N_39163,N_21876,N_23014);
and U39164 (N_39164,N_26071,N_22634);
nor U39165 (N_39165,N_25632,N_22989);
nor U39166 (N_39166,N_29496,N_25908);
xor U39167 (N_39167,N_25182,N_20907);
or U39168 (N_39168,N_23610,N_22117);
or U39169 (N_39169,N_27385,N_29318);
nor U39170 (N_39170,N_21199,N_20322);
xor U39171 (N_39171,N_27849,N_21945);
or U39172 (N_39172,N_29378,N_21305);
nand U39173 (N_39173,N_24142,N_25477);
nor U39174 (N_39174,N_20989,N_24674);
nor U39175 (N_39175,N_29691,N_24208);
or U39176 (N_39176,N_21960,N_25432);
nand U39177 (N_39177,N_28645,N_20027);
nand U39178 (N_39178,N_29697,N_22623);
and U39179 (N_39179,N_29051,N_22448);
nor U39180 (N_39180,N_23874,N_21122);
nor U39181 (N_39181,N_25255,N_21097);
or U39182 (N_39182,N_24442,N_20996);
nand U39183 (N_39183,N_20407,N_24674);
and U39184 (N_39184,N_26420,N_27055);
nand U39185 (N_39185,N_24181,N_26889);
nor U39186 (N_39186,N_22871,N_25720);
and U39187 (N_39187,N_28501,N_20739);
or U39188 (N_39188,N_23317,N_28056);
nor U39189 (N_39189,N_22635,N_25974);
or U39190 (N_39190,N_28325,N_28336);
nor U39191 (N_39191,N_26297,N_25739);
or U39192 (N_39192,N_22974,N_21079);
nor U39193 (N_39193,N_28471,N_21151);
nor U39194 (N_39194,N_27076,N_20777);
and U39195 (N_39195,N_23348,N_24698);
and U39196 (N_39196,N_22803,N_27869);
nor U39197 (N_39197,N_23724,N_21727);
and U39198 (N_39198,N_28570,N_26451);
nor U39199 (N_39199,N_26087,N_21613);
nand U39200 (N_39200,N_26245,N_28682);
nand U39201 (N_39201,N_26505,N_20371);
or U39202 (N_39202,N_21253,N_22472);
nand U39203 (N_39203,N_21666,N_26504);
nand U39204 (N_39204,N_27508,N_22403);
or U39205 (N_39205,N_20772,N_26358);
and U39206 (N_39206,N_28205,N_24638);
or U39207 (N_39207,N_25460,N_20407);
nor U39208 (N_39208,N_29770,N_25898);
nor U39209 (N_39209,N_24955,N_23779);
nand U39210 (N_39210,N_26069,N_24442);
nand U39211 (N_39211,N_20100,N_20345);
nand U39212 (N_39212,N_25300,N_23288);
or U39213 (N_39213,N_28371,N_22462);
nand U39214 (N_39214,N_27175,N_28009);
or U39215 (N_39215,N_23342,N_23225);
nand U39216 (N_39216,N_27407,N_23452);
xor U39217 (N_39217,N_23008,N_28807);
and U39218 (N_39218,N_23124,N_23370);
nor U39219 (N_39219,N_20960,N_20429);
nor U39220 (N_39220,N_29228,N_25149);
and U39221 (N_39221,N_26913,N_28186);
and U39222 (N_39222,N_24194,N_28883);
nand U39223 (N_39223,N_22307,N_22376);
nand U39224 (N_39224,N_22003,N_21654);
nand U39225 (N_39225,N_20712,N_23442);
nand U39226 (N_39226,N_20308,N_21873);
nand U39227 (N_39227,N_27931,N_28321);
or U39228 (N_39228,N_25803,N_21503);
or U39229 (N_39229,N_24911,N_22335);
and U39230 (N_39230,N_29756,N_25392);
nor U39231 (N_39231,N_27855,N_22478);
nand U39232 (N_39232,N_26040,N_23357);
or U39233 (N_39233,N_24609,N_26960);
nor U39234 (N_39234,N_23453,N_28019);
nand U39235 (N_39235,N_27259,N_27447);
or U39236 (N_39236,N_22859,N_21738);
nand U39237 (N_39237,N_21164,N_29678);
nor U39238 (N_39238,N_29136,N_23034);
nand U39239 (N_39239,N_20521,N_26933);
or U39240 (N_39240,N_26726,N_24448);
or U39241 (N_39241,N_27489,N_29186);
and U39242 (N_39242,N_26021,N_24795);
or U39243 (N_39243,N_21176,N_28403);
and U39244 (N_39244,N_21096,N_27603);
nand U39245 (N_39245,N_21382,N_20132);
and U39246 (N_39246,N_27114,N_20008);
nand U39247 (N_39247,N_26953,N_21332);
and U39248 (N_39248,N_28343,N_29557);
and U39249 (N_39249,N_23338,N_22995);
or U39250 (N_39250,N_23257,N_25157);
nand U39251 (N_39251,N_29933,N_28076);
and U39252 (N_39252,N_24364,N_24553);
or U39253 (N_39253,N_21627,N_24200);
or U39254 (N_39254,N_21788,N_22848);
nand U39255 (N_39255,N_27900,N_27855);
or U39256 (N_39256,N_26649,N_28107);
nor U39257 (N_39257,N_20384,N_28402);
nor U39258 (N_39258,N_27871,N_26837);
nand U39259 (N_39259,N_21711,N_22724);
or U39260 (N_39260,N_25365,N_22210);
or U39261 (N_39261,N_21276,N_23108);
and U39262 (N_39262,N_23909,N_27204);
and U39263 (N_39263,N_21921,N_27675);
nor U39264 (N_39264,N_21660,N_27072);
nor U39265 (N_39265,N_27025,N_26349);
nand U39266 (N_39266,N_25327,N_23417);
or U39267 (N_39267,N_24132,N_23228);
nand U39268 (N_39268,N_28812,N_23378);
nor U39269 (N_39269,N_23961,N_26990);
and U39270 (N_39270,N_28990,N_29962);
nand U39271 (N_39271,N_25532,N_20782);
and U39272 (N_39272,N_29947,N_29203);
nor U39273 (N_39273,N_24231,N_25486);
nand U39274 (N_39274,N_23717,N_28180);
nor U39275 (N_39275,N_20390,N_23567);
and U39276 (N_39276,N_22840,N_21022);
nor U39277 (N_39277,N_21969,N_21447);
nor U39278 (N_39278,N_23210,N_21894);
nand U39279 (N_39279,N_27429,N_23471);
xor U39280 (N_39280,N_24635,N_21696);
xor U39281 (N_39281,N_27735,N_24482);
nor U39282 (N_39282,N_23406,N_26286);
and U39283 (N_39283,N_29204,N_28613);
or U39284 (N_39284,N_28923,N_27845);
nor U39285 (N_39285,N_21160,N_24088);
and U39286 (N_39286,N_20492,N_25160);
and U39287 (N_39287,N_24476,N_28771);
nand U39288 (N_39288,N_23591,N_23377);
and U39289 (N_39289,N_28281,N_27539);
or U39290 (N_39290,N_20870,N_21000);
nor U39291 (N_39291,N_23176,N_20283);
nor U39292 (N_39292,N_26956,N_23799);
and U39293 (N_39293,N_26658,N_22263);
or U39294 (N_39294,N_26700,N_29023);
or U39295 (N_39295,N_26584,N_24019);
or U39296 (N_39296,N_28654,N_22077);
nor U39297 (N_39297,N_28219,N_21389);
or U39298 (N_39298,N_21809,N_27079);
or U39299 (N_39299,N_23077,N_20156);
xnor U39300 (N_39300,N_25884,N_24352);
and U39301 (N_39301,N_24763,N_25557);
nor U39302 (N_39302,N_24458,N_20065);
nand U39303 (N_39303,N_20232,N_29315);
nor U39304 (N_39304,N_21047,N_23905);
nand U39305 (N_39305,N_22076,N_26110);
nand U39306 (N_39306,N_21133,N_22514);
and U39307 (N_39307,N_23129,N_24456);
nand U39308 (N_39308,N_27270,N_23685);
and U39309 (N_39309,N_27891,N_26741);
or U39310 (N_39310,N_26746,N_28816);
nor U39311 (N_39311,N_28755,N_25160);
and U39312 (N_39312,N_21913,N_23537);
nand U39313 (N_39313,N_22477,N_27709);
or U39314 (N_39314,N_26687,N_23550);
nand U39315 (N_39315,N_21556,N_23380);
or U39316 (N_39316,N_28864,N_28396);
nand U39317 (N_39317,N_20036,N_22111);
and U39318 (N_39318,N_22906,N_21749);
nand U39319 (N_39319,N_29164,N_29839);
nand U39320 (N_39320,N_25904,N_20141);
or U39321 (N_39321,N_22527,N_22332);
or U39322 (N_39322,N_22962,N_22364);
nor U39323 (N_39323,N_27738,N_29781);
or U39324 (N_39324,N_23002,N_25095);
or U39325 (N_39325,N_28375,N_29607);
nand U39326 (N_39326,N_29039,N_28828);
nand U39327 (N_39327,N_22891,N_23526);
and U39328 (N_39328,N_29589,N_28475);
and U39329 (N_39329,N_23429,N_25722);
nor U39330 (N_39330,N_22040,N_28281);
or U39331 (N_39331,N_29196,N_27642);
nand U39332 (N_39332,N_23621,N_26264);
or U39333 (N_39333,N_20083,N_20694);
nor U39334 (N_39334,N_21498,N_26011);
nor U39335 (N_39335,N_27610,N_28729);
and U39336 (N_39336,N_28696,N_20355);
nor U39337 (N_39337,N_25705,N_29543);
and U39338 (N_39338,N_25330,N_22174);
xor U39339 (N_39339,N_27067,N_20713);
nor U39340 (N_39340,N_27553,N_29336);
nor U39341 (N_39341,N_27866,N_24191);
and U39342 (N_39342,N_20367,N_27591);
nor U39343 (N_39343,N_28662,N_27442);
xor U39344 (N_39344,N_26848,N_25699);
nand U39345 (N_39345,N_26189,N_24044);
nand U39346 (N_39346,N_20665,N_29158);
or U39347 (N_39347,N_27782,N_27615);
xnor U39348 (N_39348,N_28081,N_29178);
nor U39349 (N_39349,N_28947,N_21015);
xnor U39350 (N_39350,N_28928,N_28895);
nor U39351 (N_39351,N_24986,N_20733);
and U39352 (N_39352,N_25684,N_20832);
and U39353 (N_39353,N_29110,N_26583);
nor U39354 (N_39354,N_25736,N_28981);
nand U39355 (N_39355,N_20123,N_25822);
or U39356 (N_39356,N_25754,N_24958);
or U39357 (N_39357,N_29032,N_21185);
and U39358 (N_39358,N_22088,N_27327);
and U39359 (N_39359,N_25461,N_25810);
nor U39360 (N_39360,N_22859,N_28334);
nor U39361 (N_39361,N_23236,N_22752);
nor U39362 (N_39362,N_29716,N_21668);
and U39363 (N_39363,N_20266,N_28625);
nand U39364 (N_39364,N_27213,N_20024);
nand U39365 (N_39365,N_29911,N_23810);
or U39366 (N_39366,N_26157,N_23786);
xor U39367 (N_39367,N_25742,N_29918);
nand U39368 (N_39368,N_24379,N_22173);
nor U39369 (N_39369,N_21609,N_22252);
or U39370 (N_39370,N_21735,N_29865);
or U39371 (N_39371,N_28366,N_27044);
nor U39372 (N_39372,N_21814,N_24141);
nand U39373 (N_39373,N_20899,N_28710);
nor U39374 (N_39374,N_27568,N_27473);
nand U39375 (N_39375,N_27769,N_22578);
and U39376 (N_39376,N_23208,N_23983);
nand U39377 (N_39377,N_29122,N_29735);
nand U39378 (N_39378,N_20458,N_27380);
nand U39379 (N_39379,N_28755,N_25494);
nor U39380 (N_39380,N_27494,N_28326);
or U39381 (N_39381,N_25987,N_29859);
nor U39382 (N_39382,N_25462,N_24696);
xor U39383 (N_39383,N_24552,N_24108);
nor U39384 (N_39384,N_27117,N_23123);
or U39385 (N_39385,N_24781,N_24297);
nor U39386 (N_39386,N_28997,N_20311);
nand U39387 (N_39387,N_26041,N_28952);
and U39388 (N_39388,N_23515,N_25601);
xor U39389 (N_39389,N_25468,N_23205);
nor U39390 (N_39390,N_28380,N_25630);
nand U39391 (N_39391,N_23609,N_24550);
and U39392 (N_39392,N_22118,N_23372);
nor U39393 (N_39393,N_26752,N_21512);
or U39394 (N_39394,N_20030,N_29762);
nand U39395 (N_39395,N_26567,N_26513);
nand U39396 (N_39396,N_28686,N_28946);
nor U39397 (N_39397,N_24309,N_21127);
nor U39398 (N_39398,N_25960,N_22447);
and U39399 (N_39399,N_26558,N_23392);
or U39400 (N_39400,N_29926,N_20394);
or U39401 (N_39401,N_25030,N_24061);
or U39402 (N_39402,N_28420,N_23202);
and U39403 (N_39403,N_25346,N_26867);
and U39404 (N_39404,N_29043,N_20960);
nand U39405 (N_39405,N_21279,N_22317);
nor U39406 (N_39406,N_27602,N_21380);
or U39407 (N_39407,N_22011,N_21455);
or U39408 (N_39408,N_23864,N_20165);
and U39409 (N_39409,N_21829,N_22681);
nand U39410 (N_39410,N_29446,N_29281);
nor U39411 (N_39411,N_21482,N_28815);
nand U39412 (N_39412,N_24101,N_29992);
and U39413 (N_39413,N_27563,N_22451);
and U39414 (N_39414,N_22167,N_20155);
nand U39415 (N_39415,N_28233,N_25136);
nor U39416 (N_39416,N_28186,N_28944);
and U39417 (N_39417,N_29995,N_21026);
or U39418 (N_39418,N_22398,N_28340);
nand U39419 (N_39419,N_21317,N_23062);
or U39420 (N_39420,N_27589,N_24927);
and U39421 (N_39421,N_27983,N_22882);
and U39422 (N_39422,N_25314,N_28172);
and U39423 (N_39423,N_26485,N_24479);
nor U39424 (N_39424,N_29908,N_20428);
and U39425 (N_39425,N_21663,N_22710);
or U39426 (N_39426,N_26937,N_27475);
or U39427 (N_39427,N_28990,N_23821);
xnor U39428 (N_39428,N_26210,N_22218);
or U39429 (N_39429,N_27152,N_22896);
or U39430 (N_39430,N_25612,N_21268);
nor U39431 (N_39431,N_23505,N_29866);
nand U39432 (N_39432,N_27775,N_27220);
and U39433 (N_39433,N_27911,N_23981);
nor U39434 (N_39434,N_26146,N_26549);
or U39435 (N_39435,N_29347,N_29926);
nand U39436 (N_39436,N_28982,N_26516);
nand U39437 (N_39437,N_29608,N_24059);
and U39438 (N_39438,N_23151,N_20078);
nand U39439 (N_39439,N_26369,N_24264);
or U39440 (N_39440,N_29530,N_24024);
nand U39441 (N_39441,N_20774,N_28263);
nand U39442 (N_39442,N_20548,N_22270);
nor U39443 (N_39443,N_25215,N_26522);
and U39444 (N_39444,N_23566,N_29504);
and U39445 (N_39445,N_26551,N_26750);
nor U39446 (N_39446,N_24671,N_24711);
nand U39447 (N_39447,N_25012,N_22842);
nor U39448 (N_39448,N_24345,N_21983);
nand U39449 (N_39449,N_27652,N_22277);
nor U39450 (N_39450,N_24429,N_25260);
or U39451 (N_39451,N_24613,N_25332);
or U39452 (N_39452,N_25059,N_24432);
nand U39453 (N_39453,N_23023,N_27512);
or U39454 (N_39454,N_27393,N_28561);
or U39455 (N_39455,N_20245,N_21089);
nor U39456 (N_39456,N_29720,N_23862);
nand U39457 (N_39457,N_26620,N_27225);
and U39458 (N_39458,N_28457,N_25370);
nand U39459 (N_39459,N_28257,N_28300);
nand U39460 (N_39460,N_27261,N_23426);
xnor U39461 (N_39461,N_24620,N_26533);
and U39462 (N_39462,N_24992,N_27149);
or U39463 (N_39463,N_23027,N_20573);
and U39464 (N_39464,N_22156,N_23471);
nor U39465 (N_39465,N_26186,N_24908);
xor U39466 (N_39466,N_29141,N_29673);
and U39467 (N_39467,N_26991,N_28367);
nand U39468 (N_39468,N_29745,N_22235);
or U39469 (N_39469,N_23991,N_23776);
or U39470 (N_39470,N_24526,N_20437);
and U39471 (N_39471,N_21850,N_29641);
and U39472 (N_39472,N_27873,N_28403);
nand U39473 (N_39473,N_23643,N_26239);
or U39474 (N_39474,N_29477,N_21290);
xor U39475 (N_39475,N_27979,N_27967);
and U39476 (N_39476,N_27706,N_26265);
nor U39477 (N_39477,N_21953,N_27279);
and U39478 (N_39478,N_28753,N_24038);
and U39479 (N_39479,N_28070,N_29933);
nor U39480 (N_39480,N_24820,N_21870);
and U39481 (N_39481,N_23838,N_22855);
or U39482 (N_39482,N_27535,N_29639);
and U39483 (N_39483,N_23271,N_29813);
nor U39484 (N_39484,N_24852,N_21439);
nand U39485 (N_39485,N_28503,N_27987);
nand U39486 (N_39486,N_23577,N_24356);
or U39487 (N_39487,N_23338,N_27261);
or U39488 (N_39488,N_22235,N_26338);
and U39489 (N_39489,N_20315,N_28449);
nand U39490 (N_39490,N_24756,N_26904);
and U39491 (N_39491,N_24361,N_27660);
nand U39492 (N_39492,N_26849,N_29430);
and U39493 (N_39493,N_28662,N_24675);
nand U39494 (N_39494,N_20608,N_25400);
or U39495 (N_39495,N_26741,N_21230);
nor U39496 (N_39496,N_27797,N_25091);
nor U39497 (N_39497,N_29221,N_26684);
xor U39498 (N_39498,N_29252,N_20081);
and U39499 (N_39499,N_25702,N_27761);
and U39500 (N_39500,N_25697,N_26095);
and U39501 (N_39501,N_28342,N_21328);
and U39502 (N_39502,N_25770,N_22586);
and U39503 (N_39503,N_22987,N_23451);
or U39504 (N_39504,N_22077,N_23686);
nand U39505 (N_39505,N_23576,N_21873);
or U39506 (N_39506,N_26808,N_26284);
or U39507 (N_39507,N_20095,N_21811);
nand U39508 (N_39508,N_23599,N_24374);
or U39509 (N_39509,N_21412,N_24638);
nor U39510 (N_39510,N_24249,N_29610);
nand U39511 (N_39511,N_28580,N_20167);
or U39512 (N_39512,N_25262,N_26050);
xnor U39513 (N_39513,N_27487,N_26351);
or U39514 (N_39514,N_29436,N_27766);
or U39515 (N_39515,N_21509,N_21544);
or U39516 (N_39516,N_26613,N_28094);
or U39517 (N_39517,N_27505,N_28215);
or U39518 (N_39518,N_27286,N_21571);
nand U39519 (N_39519,N_21585,N_20073);
and U39520 (N_39520,N_29787,N_23937);
nand U39521 (N_39521,N_20361,N_22558);
nand U39522 (N_39522,N_24852,N_26575);
nand U39523 (N_39523,N_24586,N_22848);
or U39524 (N_39524,N_23089,N_24554);
or U39525 (N_39525,N_24316,N_25323);
nand U39526 (N_39526,N_26769,N_25613);
and U39527 (N_39527,N_26546,N_28656);
nor U39528 (N_39528,N_24221,N_28985);
or U39529 (N_39529,N_21752,N_20848);
or U39530 (N_39530,N_25838,N_21016);
nor U39531 (N_39531,N_25848,N_25914);
or U39532 (N_39532,N_28544,N_28320);
nand U39533 (N_39533,N_26059,N_28246);
nand U39534 (N_39534,N_21469,N_24562);
or U39535 (N_39535,N_26352,N_28211);
nor U39536 (N_39536,N_24193,N_23446);
or U39537 (N_39537,N_24450,N_27778);
or U39538 (N_39538,N_28957,N_21199);
or U39539 (N_39539,N_22211,N_22732);
nor U39540 (N_39540,N_27669,N_23293);
and U39541 (N_39541,N_22690,N_28139);
or U39542 (N_39542,N_28678,N_20169);
and U39543 (N_39543,N_21780,N_27674);
or U39544 (N_39544,N_24377,N_24829);
nor U39545 (N_39545,N_24622,N_28681);
nand U39546 (N_39546,N_21736,N_25861);
and U39547 (N_39547,N_27901,N_28879);
and U39548 (N_39548,N_27709,N_26518);
or U39549 (N_39549,N_21513,N_22133);
nor U39550 (N_39550,N_22251,N_24341);
nand U39551 (N_39551,N_20160,N_29337);
and U39552 (N_39552,N_25422,N_20491);
or U39553 (N_39553,N_22042,N_26464);
or U39554 (N_39554,N_24780,N_26621);
and U39555 (N_39555,N_20540,N_24850);
and U39556 (N_39556,N_28814,N_21502);
and U39557 (N_39557,N_29047,N_20608);
nand U39558 (N_39558,N_21441,N_23825);
nor U39559 (N_39559,N_29038,N_27364);
xor U39560 (N_39560,N_21079,N_28918);
or U39561 (N_39561,N_24777,N_21688);
and U39562 (N_39562,N_24969,N_28422);
and U39563 (N_39563,N_26842,N_20301);
nor U39564 (N_39564,N_23133,N_26514);
nand U39565 (N_39565,N_27937,N_23541);
or U39566 (N_39566,N_23153,N_20779);
or U39567 (N_39567,N_20529,N_29969);
nand U39568 (N_39568,N_20292,N_22087);
nand U39569 (N_39569,N_27998,N_25187);
or U39570 (N_39570,N_23920,N_26657);
or U39571 (N_39571,N_24130,N_21865);
or U39572 (N_39572,N_27819,N_24617);
and U39573 (N_39573,N_27954,N_24339);
or U39574 (N_39574,N_21362,N_25276);
nor U39575 (N_39575,N_28705,N_24104);
nor U39576 (N_39576,N_22108,N_24841);
or U39577 (N_39577,N_29793,N_26651);
xnor U39578 (N_39578,N_21677,N_29266);
nor U39579 (N_39579,N_22074,N_23725);
or U39580 (N_39580,N_28089,N_25235);
or U39581 (N_39581,N_22474,N_27732);
and U39582 (N_39582,N_24433,N_23341);
xnor U39583 (N_39583,N_20965,N_20912);
and U39584 (N_39584,N_27693,N_23104);
and U39585 (N_39585,N_25306,N_25757);
nand U39586 (N_39586,N_21024,N_26241);
nor U39587 (N_39587,N_20456,N_21085);
and U39588 (N_39588,N_20389,N_25141);
or U39589 (N_39589,N_22214,N_25511);
xnor U39590 (N_39590,N_28246,N_21212);
and U39591 (N_39591,N_23877,N_29189);
and U39592 (N_39592,N_26336,N_28064);
and U39593 (N_39593,N_20535,N_28836);
nand U39594 (N_39594,N_20263,N_25052);
and U39595 (N_39595,N_21770,N_23106);
nand U39596 (N_39596,N_27415,N_27820);
and U39597 (N_39597,N_21342,N_20335);
and U39598 (N_39598,N_22438,N_21122);
or U39599 (N_39599,N_24902,N_23075);
or U39600 (N_39600,N_22172,N_28793);
nand U39601 (N_39601,N_27533,N_20432);
nor U39602 (N_39602,N_26379,N_20600);
nor U39603 (N_39603,N_21666,N_24285);
or U39604 (N_39604,N_27334,N_25404);
nor U39605 (N_39605,N_27425,N_23536);
or U39606 (N_39606,N_24121,N_29024);
and U39607 (N_39607,N_27429,N_26034);
or U39608 (N_39608,N_22873,N_28385);
nor U39609 (N_39609,N_27971,N_28007);
or U39610 (N_39610,N_24989,N_25840);
and U39611 (N_39611,N_21301,N_20960);
nor U39612 (N_39612,N_20664,N_27765);
nand U39613 (N_39613,N_23458,N_29395);
or U39614 (N_39614,N_27617,N_23924);
nand U39615 (N_39615,N_29805,N_27157);
nand U39616 (N_39616,N_26595,N_23013);
or U39617 (N_39617,N_25561,N_29329);
or U39618 (N_39618,N_22926,N_24559);
xnor U39619 (N_39619,N_25769,N_25040);
or U39620 (N_39620,N_20369,N_21324);
and U39621 (N_39621,N_23512,N_29105);
and U39622 (N_39622,N_23076,N_22237);
and U39623 (N_39623,N_23376,N_23316);
xnor U39624 (N_39624,N_29246,N_20131);
nand U39625 (N_39625,N_25980,N_26746);
and U39626 (N_39626,N_28098,N_28927);
or U39627 (N_39627,N_29123,N_29507);
and U39628 (N_39628,N_21617,N_21575);
or U39629 (N_39629,N_25701,N_27268);
and U39630 (N_39630,N_27486,N_29971);
and U39631 (N_39631,N_24263,N_20229);
nor U39632 (N_39632,N_29536,N_27348);
or U39633 (N_39633,N_23791,N_26025);
xnor U39634 (N_39634,N_26206,N_27723);
or U39635 (N_39635,N_28973,N_26959);
nor U39636 (N_39636,N_23709,N_24143);
or U39637 (N_39637,N_29831,N_25372);
or U39638 (N_39638,N_20640,N_20533);
nor U39639 (N_39639,N_22645,N_21528);
and U39640 (N_39640,N_28751,N_21862);
or U39641 (N_39641,N_29286,N_23530);
nor U39642 (N_39642,N_25196,N_20314);
nand U39643 (N_39643,N_21661,N_20663);
or U39644 (N_39644,N_21868,N_26380);
nand U39645 (N_39645,N_25307,N_21399);
nand U39646 (N_39646,N_22609,N_22955);
xnor U39647 (N_39647,N_22035,N_22087);
or U39648 (N_39648,N_22106,N_29472);
nand U39649 (N_39649,N_26220,N_23090);
or U39650 (N_39650,N_21894,N_23217);
nor U39651 (N_39651,N_20116,N_25859);
nor U39652 (N_39652,N_22508,N_24696);
nor U39653 (N_39653,N_22047,N_23299);
nand U39654 (N_39654,N_20878,N_27869);
nor U39655 (N_39655,N_29773,N_20434);
nor U39656 (N_39656,N_27810,N_25955);
xnor U39657 (N_39657,N_21687,N_24267);
nor U39658 (N_39658,N_26712,N_22170);
or U39659 (N_39659,N_20734,N_24314);
nand U39660 (N_39660,N_24107,N_24900);
xnor U39661 (N_39661,N_23710,N_24929);
nor U39662 (N_39662,N_29266,N_22859);
nand U39663 (N_39663,N_29778,N_27925);
xnor U39664 (N_39664,N_28860,N_21575);
and U39665 (N_39665,N_26388,N_23850);
or U39666 (N_39666,N_27309,N_23051);
and U39667 (N_39667,N_29402,N_24348);
nand U39668 (N_39668,N_20613,N_27004);
xnor U39669 (N_39669,N_21124,N_28998);
xor U39670 (N_39670,N_26591,N_22752);
xnor U39671 (N_39671,N_24232,N_20781);
or U39672 (N_39672,N_23743,N_26844);
xnor U39673 (N_39673,N_23677,N_24788);
xnor U39674 (N_39674,N_24942,N_20697);
nand U39675 (N_39675,N_29124,N_27811);
nand U39676 (N_39676,N_28467,N_20688);
or U39677 (N_39677,N_27992,N_29186);
and U39678 (N_39678,N_23846,N_20531);
xor U39679 (N_39679,N_27013,N_28621);
nor U39680 (N_39680,N_28073,N_23937);
or U39681 (N_39681,N_28798,N_25254);
nand U39682 (N_39682,N_25518,N_22985);
nor U39683 (N_39683,N_26482,N_28278);
and U39684 (N_39684,N_24105,N_29901);
nand U39685 (N_39685,N_28488,N_20223);
or U39686 (N_39686,N_27052,N_25470);
and U39687 (N_39687,N_20340,N_25878);
nor U39688 (N_39688,N_21151,N_26050);
and U39689 (N_39689,N_26676,N_23998);
or U39690 (N_39690,N_26877,N_26768);
nor U39691 (N_39691,N_21389,N_26980);
nor U39692 (N_39692,N_27013,N_27876);
xnor U39693 (N_39693,N_25667,N_24459);
nor U39694 (N_39694,N_24840,N_25556);
and U39695 (N_39695,N_23917,N_29658);
or U39696 (N_39696,N_26239,N_20863);
nand U39697 (N_39697,N_27234,N_23612);
and U39698 (N_39698,N_22808,N_22853);
nand U39699 (N_39699,N_27421,N_24561);
and U39700 (N_39700,N_29195,N_28539);
nand U39701 (N_39701,N_25047,N_23691);
and U39702 (N_39702,N_22062,N_29987);
or U39703 (N_39703,N_22253,N_24168);
xnor U39704 (N_39704,N_28076,N_20971);
xor U39705 (N_39705,N_25051,N_24680);
or U39706 (N_39706,N_26936,N_20775);
or U39707 (N_39707,N_29304,N_29668);
or U39708 (N_39708,N_21702,N_22305);
or U39709 (N_39709,N_22970,N_22934);
and U39710 (N_39710,N_21569,N_24191);
nand U39711 (N_39711,N_22179,N_20847);
and U39712 (N_39712,N_25666,N_24815);
nand U39713 (N_39713,N_21323,N_27723);
nor U39714 (N_39714,N_28721,N_29652);
nand U39715 (N_39715,N_22156,N_29141);
nor U39716 (N_39716,N_26835,N_23311);
nand U39717 (N_39717,N_22551,N_24772);
or U39718 (N_39718,N_27102,N_24194);
nand U39719 (N_39719,N_21368,N_26096);
or U39720 (N_39720,N_23789,N_24660);
and U39721 (N_39721,N_29071,N_25983);
nor U39722 (N_39722,N_29403,N_23211);
and U39723 (N_39723,N_27373,N_23603);
nand U39724 (N_39724,N_23148,N_24013);
and U39725 (N_39725,N_20567,N_25151);
nand U39726 (N_39726,N_26440,N_27350);
nor U39727 (N_39727,N_24724,N_20779);
or U39728 (N_39728,N_26859,N_23281);
nand U39729 (N_39729,N_28796,N_28102);
and U39730 (N_39730,N_24423,N_28447);
xnor U39731 (N_39731,N_25766,N_21144);
xor U39732 (N_39732,N_22094,N_27266);
nor U39733 (N_39733,N_27411,N_26978);
and U39734 (N_39734,N_22651,N_21238);
nand U39735 (N_39735,N_29147,N_29620);
nor U39736 (N_39736,N_20097,N_26632);
and U39737 (N_39737,N_27490,N_25963);
and U39738 (N_39738,N_29928,N_20615);
and U39739 (N_39739,N_20789,N_23864);
and U39740 (N_39740,N_20848,N_21451);
nand U39741 (N_39741,N_22505,N_29952);
nor U39742 (N_39742,N_22901,N_23144);
nand U39743 (N_39743,N_25396,N_28197);
nand U39744 (N_39744,N_27755,N_23889);
or U39745 (N_39745,N_27657,N_28166);
nand U39746 (N_39746,N_21608,N_24782);
and U39747 (N_39747,N_28756,N_20054);
or U39748 (N_39748,N_23484,N_24847);
xor U39749 (N_39749,N_21709,N_27206);
and U39750 (N_39750,N_20530,N_25247);
nand U39751 (N_39751,N_21071,N_25942);
nor U39752 (N_39752,N_28330,N_27236);
nand U39753 (N_39753,N_20724,N_20698);
or U39754 (N_39754,N_27249,N_23533);
nor U39755 (N_39755,N_22910,N_28669);
or U39756 (N_39756,N_28776,N_29755);
and U39757 (N_39757,N_28926,N_20095);
nor U39758 (N_39758,N_28819,N_28665);
nand U39759 (N_39759,N_28701,N_27344);
xnor U39760 (N_39760,N_29401,N_29067);
nand U39761 (N_39761,N_24112,N_24161);
nand U39762 (N_39762,N_25550,N_27519);
nand U39763 (N_39763,N_24420,N_22901);
nor U39764 (N_39764,N_26839,N_26981);
nand U39765 (N_39765,N_28482,N_23479);
nand U39766 (N_39766,N_26485,N_21369);
and U39767 (N_39767,N_22208,N_20166);
nor U39768 (N_39768,N_25498,N_21316);
nor U39769 (N_39769,N_26721,N_27704);
xnor U39770 (N_39770,N_29978,N_22356);
nand U39771 (N_39771,N_21459,N_24026);
or U39772 (N_39772,N_24398,N_27920);
or U39773 (N_39773,N_23206,N_21276);
and U39774 (N_39774,N_26813,N_26933);
xnor U39775 (N_39775,N_25777,N_27931);
or U39776 (N_39776,N_22479,N_22820);
and U39777 (N_39777,N_21115,N_20157);
nor U39778 (N_39778,N_23473,N_28318);
nand U39779 (N_39779,N_27355,N_22173);
nor U39780 (N_39780,N_25322,N_26672);
xor U39781 (N_39781,N_26233,N_28457);
or U39782 (N_39782,N_22451,N_21214);
or U39783 (N_39783,N_20265,N_27032);
and U39784 (N_39784,N_23357,N_24271);
and U39785 (N_39785,N_22583,N_28535);
or U39786 (N_39786,N_22868,N_20552);
nand U39787 (N_39787,N_28311,N_28507);
and U39788 (N_39788,N_27551,N_24763);
nor U39789 (N_39789,N_23852,N_26379);
and U39790 (N_39790,N_28437,N_24580);
nand U39791 (N_39791,N_20447,N_26906);
or U39792 (N_39792,N_29152,N_23063);
or U39793 (N_39793,N_29363,N_22894);
nor U39794 (N_39794,N_28944,N_21542);
or U39795 (N_39795,N_29161,N_25138);
nand U39796 (N_39796,N_26653,N_23691);
nor U39797 (N_39797,N_20980,N_22794);
nand U39798 (N_39798,N_20358,N_29647);
nand U39799 (N_39799,N_25016,N_26267);
and U39800 (N_39800,N_26989,N_27510);
nor U39801 (N_39801,N_21201,N_27160);
and U39802 (N_39802,N_28360,N_20408);
or U39803 (N_39803,N_23701,N_26682);
or U39804 (N_39804,N_29969,N_23797);
nor U39805 (N_39805,N_22506,N_22976);
xnor U39806 (N_39806,N_22231,N_23844);
or U39807 (N_39807,N_23819,N_28276);
nor U39808 (N_39808,N_29433,N_23899);
nand U39809 (N_39809,N_25202,N_27257);
nand U39810 (N_39810,N_25602,N_28345);
nor U39811 (N_39811,N_28945,N_27120);
and U39812 (N_39812,N_22123,N_25232);
and U39813 (N_39813,N_20202,N_20065);
or U39814 (N_39814,N_25950,N_29060);
nor U39815 (N_39815,N_27182,N_21719);
nand U39816 (N_39816,N_26652,N_23454);
and U39817 (N_39817,N_25008,N_29925);
and U39818 (N_39818,N_26722,N_24196);
or U39819 (N_39819,N_25010,N_25548);
nand U39820 (N_39820,N_20275,N_26143);
nand U39821 (N_39821,N_26061,N_27054);
or U39822 (N_39822,N_22318,N_22369);
xnor U39823 (N_39823,N_29910,N_23852);
nor U39824 (N_39824,N_27879,N_22773);
or U39825 (N_39825,N_27551,N_22417);
and U39826 (N_39826,N_23746,N_27744);
xor U39827 (N_39827,N_27274,N_28573);
nor U39828 (N_39828,N_21230,N_20596);
and U39829 (N_39829,N_22597,N_28692);
and U39830 (N_39830,N_28231,N_25670);
or U39831 (N_39831,N_24150,N_24483);
nand U39832 (N_39832,N_22488,N_25404);
nand U39833 (N_39833,N_26383,N_23471);
and U39834 (N_39834,N_26407,N_25203);
nand U39835 (N_39835,N_28664,N_21381);
xor U39836 (N_39836,N_27012,N_21499);
and U39837 (N_39837,N_27610,N_24645);
nor U39838 (N_39838,N_29687,N_22588);
nand U39839 (N_39839,N_22355,N_20387);
nor U39840 (N_39840,N_23838,N_23161);
xor U39841 (N_39841,N_22010,N_27105);
nand U39842 (N_39842,N_23699,N_27792);
nor U39843 (N_39843,N_27326,N_20169);
nand U39844 (N_39844,N_22156,N_21248);
and U39845 (N_39845,N_20087,N_22847);
nor U39846 (N_39846,N_27899,N_22349);
nor U39847 (N_39847,N_22210,N_21022);
nand U39848 (N_39848,N_21746,N_26199);
nand U39849 (N_39849,N_29566,N_23907);
or U39850 (N_39850,N_25091,N_28412);
or U39851 (N_39851,N_23014,N_25937);
and U39852 (N_39852,N_22131,N_29972);
nor U39853 (N_39853,N_22064,N_21884);
nand U39854 (N_39854,N_27120,N_24205);
and U39855 (N_39855,N_23386,N_20316);
or U39856 (N_39856,N_20040,N_21274);
or U39857 (N_39857,N_27326,N_24352);
xnor U39858 (N_39858,N_27403,N_27205);
nor U39859 (N_39859,N_27607,N_29235);
or U39860 (N_39860,N_24283,N_21269);
or U39861 (N_39861,N_29340,N_25485);
or U39862 (N_39862,N_27606,N_29991);
nand U39863 (N_39863,N_21206,N_20855);
nor U39864 (N_39864,N_22902,N_21661);
and U39865 (N_39865,N_29931,N_20532);
nor U39866 (N_39866,N_25537,N_24514);
or U39867 (N_39867,N_27233,N_24204);
xnor U39868 (N_39868,N_20722,N_20940);
nor U39869 (N_39869,N_25428,N_29098);
nand U39870 (N_39870,N_29480,N_27518);
nand U39871 (N_39871,N_20444,N_21063);
nor U39872 (N_39872,N_21041,N_21465);
or U39873 (N_39873,N_29523,N_26345);
or U39874 (N_39874,N_29565,N_26101);
nand U39875 (N_39875,N_23649,N_29644);
nand U39876 (N_39876,N_24710,N_24040);
and U39877 (N_39877,N_20741,N_28671);
nor U39878 (N_39878,N_21898,N_28701);
and U39879 (N_39879,N_29421,N_26968);
xor U39880 (N_39880,N_27796,N_25175);
and U39881 (N_39881,N_23800,N_26752);
xnor U39882 (N_39882,N_25093,N_25512);
and U39883 (N_39883,N_29223,N_27483);
and U39884 (N_39884,N_29592,N_25062);
nor U39885 (N_39885,N_20097,N_22342);
or U39886 (N_39886,N_28788,N_23285);
nor U39887 (N_39887,N_21380,N_23996);
or U39888 (N_39888,N_21670,N_28073);
nor U39889 (N_39889,N_24094,N_22926);
and U39890 (N_39890,N_28522,N_28217);
xor U39891 (N_39891,N_27783,N_23416);
or U39892 (N_39892,N_25987,N_27687);
and U39893 (N_39893,N_27830,N_22628);
and U39894 (N_39894,N_26948,N_21895);
nand U39895 (N_39895,N_20160,N_25436);
nand U39896 (N_39896,N_26490,N_20733);
or U39897 (N_39897,N_25590,N_24982);
and U39898 (N_39898,N_20550,N_21845);
and U39899 (N_39899,N_28628,N_23231);
nor U39900 (N_39900,N_26203,N_22199);
or U39901 (N_39901,N_20159,N_21175);
or U39902 (N_39902,N_26070,N_20775);
nand U39903 (N_39903,N_24875,N_28790);
nor U39904 (N_39904,N_28999,N_27653);
and U39905 (N_39905,N_29747,N_28515);
and U39906 (N_39906,N_27227,N_20378);
and U39907 (N_39907,N_29257,N_26514);
nand U39908 (N_39908,N_26232,N_23355);
nand U39909 (N_39909,N_26215,N_25420);
and U39910 (N_39910,N_24621,N_28221);
or U39911 (N_39911,N_27110,N_20206);
nand U39912 (N_39912,N_27105,N_23405);
or U39913 (N_39913,N_28778,N_26084);
and U39914 (N_39914,N_29380,N_26579);
nand U39915 (N_39915,N_27540,N_28546);
nand U39916 (N_39916,N_26079,N_23780);
and U39917 (N_39917,N_25414,N_20862);
xor U39918 (N_39918,N_20583,N_24932);
nand U39919 (N_39919,N_23330,N_26987);
nor U39920 (N_39920,N_28046,N_24135);
or U39921 (N_39921,N_28890,N_23103);
xnor U39922 (N_39922,N_21357,N_26875);
nand U39923 (N_39923,N_21990,N_22915);
nor U39924 (N_39924,N_25289,N_28132);
and U39925 (N_39925,N_26879,N_27664);
nand U39926 (N_39926,N_29463,N_26411);
nor U39927 (N_39927,N_29775,N_28271);
or U39928 (N_39928,N_23885,N_23113);
and U39929 (N_39929,N_20645,N_20155);
nand U39930 (N_39930,N_22574,N_25451);
and U39931 (N_39931,N_23704,N_25511);
or U39932 (N_39932,N_24963,N_22226);
and U39933 (N_39933,N_25065,N_27952);
xnor U39934 (N_39934,N_20393,N_27252);
or U39935 (N_39935,N_29273,N_23754);
nor U39936 (N_39936,N_25882,N_20180);
or U39937 (N_39937,N_23355,N_25177);
nor U39938 (N_39938,N_29212,N_21308);
or U39939 (N_39939,N_23267,N_22643);
nor U39940 (N_39940,N_20314,N_25580);
and U39941 (N_39941,N_22064,N_24763);
nor U39942 (N_39942,N_25269,N_21111);
nand U39943 (N_39943,N_27442,N_27453);
and U39944 (N_39944,N_24003,N_21324);
or U39945 (N_39945,N_20830,N_29192);
nor U39946 (N_39946,N_26805,N_23426);
nor U39947 (N_39947,N_22996,N_25700);
and U39948 (N_39948,N_29963,N_26904);
or U39949 (N_39949,N_22694,N_20998);
or U39950 (N_39950,N_27826,N_28727);
and U39951 (N_39951,N_21050,N_20029);
and U39952 (N_39952,N_25868,N_25609);
and U39953 (N_39953,N_26783,N_24528);
and U39954 (N_39954,N_20793,N_23045);
nor U39955 (N_39955,N_21057,N_28822);
nand U39956 (N_39956,N_26644,N_22941);
or U39957 (N_39957,N_22570,N_26680);
nor U39958 (N_39958,N_27338,N_24993);
and U39959 (N_39959,N_28370,N_25012);
nor U39960 (N_39960,N_24207,N_20209);
and U39961 (N_39961,N_20878,N_27517);
or U39962 (N_39962,N_29440,N_24620);
or U39963 (N_39963,N_25011,N_25188);
or U39964 (N_39964,N_20015,N_27356);
and U39965 (N_39965,N_27122,N_27336);
or U39966 (N_39966,N_29239,N_26344);
and U39967 (N_39967,N_20425,N_20546);
and U39968 (N_39968,N_25460,N_22509);
nand U39969 (N_39969,N_25013,N_23127);
nand U39970 (N_39970,N_20203,N_27543);
and U39971 (N_39971,N_23520,N_21043);
and U39972 (N_39972,N_21716,N_28615);
xor U39973 (N_39973,N_23273,N_21600);
or U39974 (N_39974,N_28688,N_29194);
and U39975 (N_39975,N_27620,N_20211);
nor U39976 (N_39976,N_21751,N_24973);
and U39977 (N_39977,N_21650,N_26451);
nand U39978 (N_39978,N_26602,N_27413);
nor U39979 (N_39979,N_26585,N_22873);
and U39980 (N_39980,N_29860,N_25524);
or U39981 (N_39981,N_24260,N_20769);
or U39982 (N_39982,N_28403,N_24383);
and U39983 (N_39983,N_20441,N_21840);
and U39984 (N_39984,N_27676,N_20235);
and U39985 (N_39985,N_21783,N_25512);
nor U39986 (N_39986,N_24242,N_22626);
nor U39987 (N_39987,N_22301,N_22877);
and U39988 (N_39988,N_28208,N_29068);
xor U39989 (N_39989,N_24985,N_21856);
or U39990 (N_39990,N_27165,N_23227);
or U39991 (N_39991,N_26309,N_21002);
xnor U39992 (N_39992,N_26944,N_26825);
nand U39993 (N_39993,N_28749,N_24922);
and U39994 (N_39994,N_21076,N_20765);
or U39995 (N_39995,N_24119,N_27082);
xnor U39996 (N_39996,N_27988,N_29473);
or U39997 (N_39997,N_24048,N_27736);
nand U39998 (N_39998,N_27257,N_29634);
and U39999 (N_39999,N_23405,N_22717);
and U40000 (N_40000,N_39267,N_38303);
or U40001 (N_40001,N_30679,N_37368);
nor U40002 (N_40002,N_37921,N_37924);
and U40003 (N_40003,N_32699,N_35509);
nand U40004 (N_40004,N_32194,N_35243);
nor U40005 (N_40005,N_34135,N_33383);
xnor U40006 (N_40006,N_32628,N_38276);
nor U40007 (N_40007,N_38043,N_33297);
or U40008 (N_40008,N_31592,N_34603);
nor U40009 (N_40009,N_32635,N_36200);
and U40010 (N_40010,N_30757,N_34666);
nor U40011 (N_40011,N_30887,N_39732);
nor U40012 (N_40012,N_31596,N_35705);
nor U40013 (N_40013,N_37615,N_38518);
and U40014 (N_40014,N_39708,N_38740);
and U40015 (N_40015,N_34590,N_35681);
and U40016 (N_40016,N_39776,N_36327);
and U40017 (N_40017,N_38090,N_31409);
nand U40018 (N_40018,N_37735,N_33667);
nor U40019 (N_40019,N_33930,N_33006);
and U40020 (N_40020,N_39991,N_31452);
nor U40021 (N_40021,N_38466,N_35129);
and U40022 (N_40022,N_39538,N_39699);
or U40023 (N_40023,N_39152,N_34083);
nor U40024 (N_40024,N_33105,N_35311);
xnor U40025 (N_40025,N_37261,N_31263);
or U40026 (N_40026,N_31634,N_30405);
nand U40027 (N_40027,N_33863,N_35900);
nor U40028 (N_40028,N_32557,N_36594);
and U40029 (N_40029,N_32659,N_30023);
or U40030 (N_40030,N_38501,N_36446);
or U40031 (N_40031,N_37610,N_32221);
nand U40032 (N_40032,N_35207,N_39832);
or U40033 (N_40033,N_38441,N_30375);
nand U40034 (N_40034,N_30704,N_30613);
and U40035 (N_40035,N_35343,N_30616);
and U40036 (N_40036,N_36007,N_36840);
or U40037 (N_40037,N_37360,N_32377);
or U40038 (N_40038,N_35807,N_37148);
or U40039 (N_40039,N_30753,N_36253);
xnor U40040 (N_40040,N_32772,N_30296);
nand U40041 (N_40041,N_35692,N_33306);
and U40042 (N_40042,N_33528,N_37556);
or U40043 (N_40043,N_37432,N_31973);
and U40044 (N_40044,N_36247,N_35322);
nand U40045 (N_40045,N_33823,N_34341);
nand U40046 (N_40046,N_35654,N_34589);
xnor U40047 (N_40047,N_37363,N_39506);
nor U40048 (N_40048,N_39995,N_35893);
or U40049 (N_40049,N_34195,N_32288);
nand U40050 (N_40050,N_34880,N_33399);
nor U40051 (N_40051,N_30149,N_35615);
nand U40052 (N_40052,N_38702,N_32418);
nand U40053 (N_40053,N_30147,N_38000);
nor U40054 (N_40054,N_31123,N_35298);
and U40055 (N_40055,N_32296,N_34786);
nor U40056 (N_40056,N_39333,N_33213);
and U40057 (N_40057,N_33599,N_30448);
or U40058 (N_40058,N_31725,N_34322);
nor U40059 (N_40059,N_37025,N_37003);
nand U40060 (N_40060,N_33073,N_35437);
and U40061 (N_40061,N_32530,N_39956);
nand U40062 (N_40062,N_32059,N_39783);
nand U40063 (N_40063,N_33608,N_35915);
nor U40064 (N_40064,N_34310,N_33908);
and U40065 (N_40065,N_38834,N_39357);
and U40066 (N_40066,N_36503,N_32770);
or U40067 (N_40067,N_31354,N_30304);
and U40068 (N_40068,N_39246,N_39702);
or U40069 (N_40069,N_31867,N_34556);
nand U40070 (N_40070,N_35271,N_34464);
xnor U40071 (N_40071,N_30131,N_37062);
and U40072 (N_40072,N_36097,N_34718);
and U40073 (N_40073,N_36784,N_30633);
and U40074 (N_40074,N_31662,N_38705);
and U40075 (N_40075,N_36801,N_36514);
nor U40076 (N_40076,N_34405,N_37970);
nor U40077 (N_40077,N_34392,N_37066);
and U40078 (N_40078,N_31307,N_32731);
and U40079 (N_40079,N_33158,N_38822);
or U40080 (N_40080,N_32141,N_33226);
nand U40081 (N_40081,N_38263,N_35055);
or U40082 (N_40082,N_31115,N_32780);
xnor U40083 (N_40083,N_34487,N_30766);
and U40084 (N_40084,N_36796,N_35548);
nor U40085 (N_40085,N_38726,N_30860);
nor U40086 (N_40086,N_30854,N_34584);
or U40087 (N_40087,N_32959,N_37930);
or U40088 (N_40088,N_30465,N_33428);
and U40089 (N_40089,N_39265,N_39053);
nand U40090 (N_40090,N_35411,N_35710);
or U40091 (N_40091,N_33392,N_33502);
or U40092 (N_40092,N_30064,N_38475);
and U40093 (N_40093,N_33047,N_30276);
nor U40094 (N_40094,N_31543,N_38869);
nand U40095 (N_40095,N_38437,N_32613);
nor U40096 (N_40096,N_33311,N_36480);
nand U40097 (N_40097,N_36323,N_30552);
nor U40098 (N_40098,N_38841,N_33115);
nor U40099 (N_40099,N_34363,N_31157);
and U40100 (N_40100,N_31727,N_38152);
nand U40101 (N_40101,N_32816,N_38250);
or U40102 (N_40102,N_31081,N_34335);
or U40103 (N_40103,N_33779,N_31532);
nor U40104 (N_40104,N_34501,N_38863);
nand U40105 (N_40105,N_32153,N_38577);
nand U40106 (N_40106,N_36414,N_30282);
nand U40107 (N_40107,N_32186,N_38891);
or U40108 (N_40108,N_38407,N_34023);
and U40109 (N_40109,N_38102,N_36006);
nand U40110 (N_40110,N_30966,N_37012);
nand U40111 (N_40111,N_33648,N_39735);
nand U40112 (N_40112,N_33294,N_31387);
and U40113 (N_40113,N_38362,N_34126);
nand U40114 (N_40114,N_36482,N_33475);
and U40115 (N_40115,N_37466,N_31346);
or U40116 (N_40116,N_38420,N_36451);
or U40117 (N_40117,N_36072,N_37652);
xnor U40118 (N_40118,N_37591,N_33664);
nor U40119 (N_40119,N_39034,N_31892);
or U40120 (N_40120,N_36215,N_30072);
or U40121 (N_40121,N_36279,N_33893);
and U40122 (N_40122,N_37902,N_32159);
and U40123 (N_40123,N_36959,N_31051);
nand U40124 (N_40124,N_36056,N_34780);
nor U40125 (N_40125,N_32592,N_37719);
xor U40126 (N_40126,N_30603,N_32002);
or U40127 (N_40127,N_35353,N_32478);
nand U40128 (N_40128,N_34554,N_31395);
nand U40129 (N_40129,N_35952,N_33053);
and U40130 (N_40130,N_37553,N_30581);
and U40131 (N_40131,N_38288,N_36459);
nor U40132 (N_40132,N_35483,N_35042);
nor U40133 (N_40133,N_31693,N_30577);
and U40134 (N_40134,N_35659,N_36165);
nor U40135 (N_40135,N_31002,N_38225);
xor U40136 (N_40136,N_31842,N_30436);
nand U40137 (N_40137,N_30476,N_39639);
nand U40138 (N_40138,N_33194,N_32054);
nor U40139 (N_40139,N_38129,N_30223);
xor U40140 (N_40140,N_36483,N_37771);
and U40141 (N_40141,N_37871,N_34003);
and U40142 (N_40142,N_35494,N_33822);
and U40143 (N_40143,N_36589,N_35410);
and U40144 (N_40144,N_33285,N_37082);
or U40145 (N_40145,N_38548,N_34885);
and U40146 (N_40146,N_39280,N_37969);
or U40147 (N_40147,N_35318,N_38190);
or U40148 (N_40148,N_39349,N_38473);
and U40149 (N_40149,N_32974,N_35975);
nor U40150 (N_40150,N_31249,N_37545);
nand U40151 (N_40151,N_34388,N_36568);
xnor U40152 (N_40152,N_31447,N_35961);
nand U40153 (N_40153,N_31760,N_32853);
nor U40154 (N_40154,N_36660,N_30882);
or U40155 (N_40155,N_37341,N_30014);
nor U40156 (N_40156,N_32585,N_39046);
or U40157 (N_40157,N_32163,N_33040);
nand U40158 (N_40158,N_38742,N_38949);
or U40159 (N_40159,N_36089,N_30817);
or U40160 (N_40160,N_35285,N_31764);
nor U40161 (N_40161,N_36887,N_37822);
nor U40162 (N_40162,N_39204,N_37660);
nor U40163 (N_40163,N_39017,N_36272);
nand U40164 (N_40164,N_34707,N_35673);
nor U40165 (N_40165,N_35663,N_34670);
nand U40166 (N_40166,N_31968,N_32705);
or U40167 (N_40167,N_35054,N_32474);
nand U40168 (N_40168,N_32740,N_35753);
xor U40169 (N_40169,N_39108,N_37035);
nor U40170 (N_40170,N_34991,N_39450);
or U40171 (N_40171,N_38097,N_34695);
nor U40172 (N_40172,N_31880,N_32073);
or U40173 (N_40173,N_33868,N_36046);
and U40174 (N_40174,N_37205,N_36750);
xor U40175 (N_40175,N_35779,N_36655);
or U40176 (N_40176,N_35881,N_39717);
or U40177 (N_40177,N_33741,N_31528);
and U40178 (N_40178,N_37536,N_32229);
nor U40179 (N_40179,N_36286,N_36449);
xnor U40180 (N_40180,N_31981,N_37589);
nor U40181 (N_40181,N_36017,N_30019);
nor U40182 (N_40182,N_37163,N_36021);
nand U40183 (N_40183,N_38093,N_31568);
or U40184 (N_40184,N_33258,N_38789);
and U40185 (N_40185,N_34594,N_37884);
and U40186 (N_40186,N_37827,N_34898);
or U40187 (N_40187,N_30517,N_35036);
or U40188 (N_40188,N_33722,N_33296);
and U40189 (N_40189,N_31321,N_37953);
and U40190 (N_40190,N_33074,N_35527);
nand U40191 (N_40191,N_32090,N_32022);
nand U40192 (N_40192,N_36118,N_35022);
and U40193 (N_40193,N_36318,N_38648);
and U40194 (N_40194,N_33852,N_30009);
and U40195 (N_40195,N_38353,N_35469);
nand U40196 (N_40196,N_37980,N_34399);
or U40197 (N_40197,N_32038,N_32996);
nor U40198 (N_40198,N_34605,N_36032);
and U40199 (N_40199,N_36038,N_34920);
nor U40200 (N_40200,N_37241,N_39888);
nor U40201 (N_40201,N_30449,N_33869);
or U40202 (N_40202,N_38487,N_39883);
and U40203 (N_40203,N_31237,N_30203);
or U40204 (N_40204,N_30337,N_35909);
nand U40205 (N_40205,N_37699,N_37484);
or U40206 (N_40206,N_34987,N_36742);
and U40207 (N_40207,N_35872,N_36546);
nor U40208 (N_40208,N_37430,N_38823);
nor U40209 (N_40209,N_37317,N_31812);
nor U40210 (N_40210,N_39295,N_35273);
nand U40211 (N_40211,N_31449,N_30016);
nand U40212 (N_40212,N_30050,N_33338);
or U40213 (N_40213,N_34642,N_39033);
nor U40214 (N_40214,N_37567,N_34496);
or U40215 (N_40215,N_38065,N_39595);
nor U40216 (N_40216,N_34519,N_30780);
nor U40217 (N_40217,N_37764,N_30361);
and U40218 (N_40218,N_37635,N_36229);
nor U40219 (N_40219,N_32923,N_35544);
nand U40220 (N_40220,N_32497,N_31530);
and U40221 (N_40221,N_34230,N_36837);
or U40222 (N_40222,N_34832,N_37096);
xor U40223 (N_40223,N_39879,N_37626);
or U40224 (N_40224,N_39426,N_35372);
and U40225 (N_40225,N_36189,N_34444);
nor U40226 (N_40226,N_37785,N_31691);
nand U40227 (N_40227,N_35995,N_34610);
nor U40228 (N_40228,N_30240,N_34451);
or U40229 (N_40229,N_31475,N_37369);
nor U40230 (N_40230,N_39941,N_35334);
xor U40231 (N_40231,N_38240,N_30784);
nand U40232 (N_40232,N_32366,N_32978);
nor U40233 (N_40233,N_35922,N_32994);
or U40234 (N_40234,N_32105,N_35073);
nor U40235 (N_40235,N_36878,N_35308);
nor U40236 (N_40236,N_35015,N_31770);
nand U40237 (N_40237,N_35519,N_38213);
and U40238 (N_40238,N_34583,N_33402);
nand U40239 (N_40239,N_31878,N_31772);
or U40240 (N_40240,N_34409,N_37632);
nor U40241 (N_40241,N_31443,N_35350);
or U40242 (N_40242,N_35759,N_39010);
and U40243 (N_40243,N_39600,N_36799);
nand U40244 (N_40244,N_36930,N_38981);
xnor U40245 (N_40245,N_39039,N_33321);
nor U40246 (N_40246,N_35623,N_35943);
or U40247 (N_40247,N_31006,N_32815);
and U40248 (N_40248,N_35084,N_35229);
or U40249 (N_40249,N_30848,N_32445);
nand U40250 (N_40250,N_34785,N_37490);
nand U40251 (N_40251,N_32878,N_38652);
nor U40252 (N_40252,N_38242,N_33916);
nor U40253 (N_40253,N_38578,N_35404);
nand U40254 (N_40254,N_32476,N_38616);
and U40255 (N_40255,N_36102,N_33231);
or U40256 (N_40256,N_30807,N_37837);
xnor U40257 (N_40257,N_37940,N_37200);
and U40258 (N_40258,N_37858,N_37910);
nor U40259 (N_40259,N_37122,N_35014);
xnor U40260 (N_40260,N_39323,N_36310);
nor U40261 (N_40261,N_31291,N_39686);
xor U40262 (N_40262,N_30176,N_35780);
nor U40263 (N_40263,N_32103,N_36425);
and U40264 (N_40264,N_32297,N_36979);
nand U40265 (N_40265,N_34120,N_38366);
or U40266 (N_40266,N_30238,N_32428);
and U40267 (N_40267,N_33957,N_36988);
nand U40268 (N_40268,N_38428,N_30635);
nor U40269 (N_40269,N_39096,N_30665);
nor U40270 (N_40270,N_38507,N_31987);
xnor U40271 (N_40271,N_32256,N_31955);
nand U40272 (N_40272,N_32488,N_33791);
and U40273 (N_40273,N_32304,N_35282);
nor U40274 (N_40274,N_32126,N_35647);
and U40275 (N_40275,N_32202,N_34917);
or U40276 (N_40276,N_33694,N_31881);
nor U40277 (N_40277,N_30832,N_33339);
nand U40278 (N_40278,N_32847,N_39528);
nand U40279 (N_40279,N_30742,N_37105);
nor U40280 (N_40280,N_38044,N_31649);
or U40281 (N_40281,N_38772,N_38748);
and U40282 (N_40282,N_33892,N_39143);
or U40283 (N_40283,N_38530,N_33501);
or U40284 (N_40284,N_37332,N_32665);
nand U40285 (N_40285,N_33715,N_38576);
or U40286 (N_40286,N_37019,N_37600);
nand U40287 (N_40287,N_36539,N_37880);
nand U40288 (N_40288,N_30835,N_31431);
or U40289 (N_40289,N_33026,N_31534);
nor U40290 (N_40290,N_31914,N_33538);
nand U40291 (N_40291,N_33699,N_38892);
xnor U40292 (N_40292,N_38820,N_32837);
nand U40293 (N_40293,N_30070,N_32465);
nand U40294 (N_40294,N_37027,N_35933);
nor U40295 (N_40295,N_30795,N_38955);
nor U40296 (N_40296,N_34402,N_35508);
or U40297 (N_40297,N_37541,N_34735);
xor U40298 (N_40298,N_34370,N_31654);
nand U40299 (N_40299,N_38650,N_37008);
nor U40300 (N_40300,N_38858,N_31539);
or U40301 (N_40301,N_31236,N_30094);
xnor U40302 (N_40302,N_38006,N_37869);
and U40303 (N_40303,N_31303,N_32786);
nand U40304 (N_40304,N_30508,N_36154);
nand U40305 (N_40305,N_33028,N_33515);
nor U40306 (N_40306,N_36800,N_39156);
and U40307 (N_40307,N_34152,N_37853);
and U40308 (N_40308,N_35296,N_34173);
and U40309 (N_40309,N_39861,N_32005);
or U40310 (N_40310,N_35850,N_38266);
xnor U40311 (N_40311,N_30877,N_36468);
nor U40312 (N_40312,N_37784,N_36682);
nor U40313 (N_40313,N_36732,N_38503);
nand U40314 (N_40314,N_30320,N_35037);
and U40315 (N_40315,N_33736,N_37401);
and U40316 (N_40316,N_31069,N_39396);
nor U40317 (N_40317,N_35139,N_35599);
or U40318 (N_40318,N_33577,N_34582);
nand U40319 (N_40319,N_37744,N_37267);
nand U40320 (N_40320,N_32564,N_33163);
and U40321 (N_40321,N_30153,N_38515);
xnor U40322 (N_40322,N_35109,N_38312);
and U40323 (N_40323,N_33628,N_30002);
nor U40324 (N_40324,N_33064,N_33448);
and U40325 (N_40325,N_39677,N_32627);
nand U40326 (N_40326,N_30255,N_39020);
or U40327 (N_40327,N_38598,N_38332);
nand U40328 (N_40328,N_32515,N_39574);
or U40329 (N_40329,N_31692,N_33887);
nand U40330 (N_40330,N_34941,N_36782);
xor U40331 (N_40331,N_30912,N_31416);
nor U40332 (N_40332,N_33041,N_33286);
nand U40333 (N_40333,N_39530,N_31477);
and U40334 (N_40334,N_35454,N_38930);
or U40335 (N_40335,N_39649,N_39689);
or U40336 (N_40336,N_30226,N_32892);
and U40337 (N_40337,N_31509,N_31716);
xnor U40338 (N_40338,N_30696,N_37471);
nand U40339 (N_40339,N_36115,N_34804);
xor U40340 (N_40340,N_31800,N_33171);
nand U40341 (N_40341,N_35091,N_38080);
or U40342 (N_40342,N_36168,N_32451);
nand U40343 (N_40343,N_38424,N_36158);
nor U40344 (N_40344,N_32872,N_35957);
and U40345 (N_40345,N_36845,N_33956);
nand U40346 (N_40346,N_39721,N_38711);
xnor U40347 (N_40347,N_36130,N_30080);
or U40348 (N_40348,N_31983,N_30682);
or U40349 (N_40349,N_38232,N_38377);
xor U40350 (N_40350,N_37239,N_38386);
nand U40351 (N_40351,N_38825,N_36283);
and U40352 (N_40352,N_33910,N_30587);
xor U40353 (N_40353,N_39692,N_37925);
nand U40354 (N_40354,N_35168,N_34954);
nor U40355 (N_40355,N_31919,N_35789);
nor U40356 (N_40356,N_35457,N_30157);
xnor U40357 (N_40357,N_31333,N_37964);
xor U40358 (N_40358,N_37621,N_32968);
or U40359 (N_40359,N_38181,N_36411);
nand U40360 (N_40360,N_38510,N_36358);
nor U40361 (N_40361,N_32121,N_33506);
nor U40362 (N_40362,N_35189,N_34441);
nor U40363 (N_40363,N_36735,N_37537);
xnor U40364 (N_40364,N_39014,N_32679);
nand U40365 (N_40365,N_31086,N_37642);
or U40366 (N_40366,N_35179,N_33003);
nand U40367 (N_40367,N_36345,N_35682);
or U40368 (N_40368,N_33732,N_32236);
nor U40369 (N_40369,N_33111,N_37936);
nand U40370 (N_40370,N_30847,N_33136);
nand U40371 (N_40371,N_36760,N_33637);
xnor U40372 (N_40372,N_34883,N_33295);
and U40373 (N_40373,N_31524,N_39245);
xnor U40374 (N_40374,N_34478,N_33821);
nor U40375 (N_40375,N_38078,N_36462);
nand U40376 (N_40376,N_39091,N_36051);
nand U40377 (N_40377,N_34193,N_32006);
nand U40378 (N_40378,N_35305,N_30516);
nor U40379 (N_40379,N_33187,N_32417);
and U40380 (N_40380,N_34044,N_39392);
nand U40381 (N_40381,N_30253,N_38538);
xor U40382 (N_40382,N_38958,N_34979);
nand U40383 (N_40383,N_33190,N_30749);
and U40384 (N_40384,N_31124,N_39196);
nand U40385 (N_40385,N_32057,N_35863);
nor U40386 (N_40386,N_35734,N_38990);
xor U40387 (N_40387,N_33875,N_39160);
nand U40388 (N_40388,N_35421,N_39367);
or U40389 (N_40389,N_30724,N_32191);
nor U40390 (N_40390,N_39035,N_32388);
nand U40391 (N_40391,N_36481,N_36396);
nand U40392 (N_40392,N_31635,N_39957);
nand U40393 (N_40393,N_37742,N_35792);
nand U40394 (N_40394,N_39442,N_36769);
xor U40395 (N_40395,N_34475,N_36520);
nand U40396 (N_40396,N_39688,N_31762);
nand U40397 (N_40397,N_39777,N_37480);
nor U40398 (N_40398,N_39161,N_39958);
or U40399 (N_40399,N_36094,N_30555);
nor U40400 (N_40400,N_35571,N_37102);
nand U40401 (N_40401,N_30055,N_30840);
nor U40402 (N_40402,N_39533,N_35012);
or U40403 (N_40403,N_34181,N_38984);
and U40404 (N_40404,N_30089,N_38026);
or U40405 (N_40405,N_30411,N_39235);
nand U40406 (N_40406,N_36075,N_35423);
or U40407 (N_40407,N_31154,N_37636);
and U40408 (N_40408,N_31996,N_32633);
and U40409 (N_40409,N_37527,N_31771);
or U40410 (N_40410,N_30129,N_36378);
nand U40411 (N_40411,N_39909,N_34524);
nor U40412 (N_40412,N_31756,N_37667);
and U40413 (N_40413,N_39572,N_31313);
and U40414 (N_40414,N_33658,N_38189);
nand U40415 (N_40415,N_39347,N_31611);
or U40416 (N_40416,N_31527,N_32719);
or U40417 (N_40417,N_31480,N_37438);
and U40418 (N_40418,N_32177,N_39980);
xnor U40419 (N_40419,N_32622,N_37656);
or U40420 (N_40420,N_36246,N_36371);
and U40421 (N_40421,N_34090,N_37631);
or U40422 (N_40422,N_30105,N_31967);
nand U40423 (N_40423,N_30799,N_33920);
nor U40424 (N_40424,N_38954,N_31434);
nand U40425 (N_40425,N_35278,N_39446);
nand U40426 (N_40426,N_38290,N_31407);
nor U40427 (N_40427,N_35602,N_32611);
nor U40428 (N_40428,N_34282,N_32479);
nand U40429 (N_40429,N_37232,N_38910);
and U40430 (N_40430,N_39753,N_34354);
nor U40431 (N_40431,N_32263,N_39230);
nor U40432 (N_40432,N_34779,N_37961);
and U40433 (N_40433,N_34537,N_39172);
nand U40434 (N_40434,N_34355,N_31011);
xnor U40435 (N_40435,N_30185,N_31595);
xor U40436 (N_40436,N_39065,N_32132);
nand U40437 (N_40437,N_30108,N_32449);
nand U40438 (N_40438,N_39374,N_34535);
nor U40439 (N_40439,N_39343,N_30617);
nor U40440 (N_40440,N_35707,N_34473);
nor U40441 (N_40441,N_37175,N_36931);
or U40442 (N_40442,N_35335,N_30843);
nor U40443 (N_40443,N_33627,N_33873);
nor U40444 (N_40444,N_31863,N_30861);
and U40445 (N_40445,N_34286,N_32089);
and U40446 (N_40446,N_35316,N_32753);
and U40447 (N_40447,N_38034,N_33324);
nand U40448 (N_40448,N_34243,N_36302);
nand U40449 (N_40449,N_32317,N_39487);
nand U40450 (N_40450,N_32537,N_31792);
or U40451 (N_40451,N_39191,N_31697);
xnor U40452 (N_40452,N_32039,N_33967);
or U40453 (N_40453,N_34709,N_31245);
or U40454 (N_40454,N_33420,N_32300);
and U40455 (N_40455,N_32950,N_35879);
or U40456 (N_40456,N_34332,N_30627);
and U40457 (N_40457,N_34940,N_36472);
nor U40458 (N_40458,N_37913,N_38111);
nand U40459 (N_40459,N_38490,N_36675);
nor U40460 (N_40460,N_34965,N_32997);
or U40461 (N_40461,N_39545,N_38294);
and U40462 (N_40462,N_32732,N_33576);
nand U40463 (N_40463,N_31751,N_35176);
and U40464 (N_40464,N_34776,N_37138);
nand U40465 (N_40465,N_33993,N_30953);
nand U40466 (N_40466,N_37286,N_33874);
nor U40467 (N_40467,N_31413,N_39497);
nor U40468 (N_40468,N_30473,N_39681);
nand U40469 (N_40469,N_32657,N_35808);
and U40470 (N_40470,N_39599,N_38516);
and U40471 (N_40471,N_36549,N_30003);
nand U40472 (N_40472,N_37551,N_32410);
or U40473 (N_40473,N_34404,N_30015);
nor U40474 (N_40474,N_30041,N_31938);
or U40475 (N_40475,N_38371,N_37045);
and U40476 (N_40476,N_32711,N_32251);
and U40477 (N_40477,N_38761,N_35644);
nand U40478 (N_40478,N_35913,N_35198);
and U40479 (N_40479,N_39264,N_34613);
nand U40480 (N_40480,N_37220,N_33499);
xnor U40481 (N_40481,N_37130,N_37752);
nor U40482 (N_40482,N_34942,N_32315);
and U40483 (N_40483,N_36139,N_30352);
nor U40484 (N_40484,N_38231,N_33561);
or U40485 (N_40485,N_30327,N_36152);
and U40486 (N_40486,N_39582,N_31023);
nand U40487 (N_40487,N_38704,N_31060);
nor U40488 (N_40488,N_36180,N_36771);
or U40489 (N_40489,N_38145,N_37979);
nand U40490 (N_40490,N_38649,N_37834);
and U40491 (N_40491,N_38547,N_30731);
nor U40492 (N_40492,N_38131,N_39175);
and U40493 (N_40493,N_33175,N_34704);
nor U40494 (N_40494,N_30038,N_34039);
nand U40495 (N_40495,N_30434,N_37741);
nor U40496 (N_40496,N_33900,N_33408);
or U40497 (N_40497,N_35435,N_36122);
or U40498 (N_40498,N_30355,N_37039);
nand U40499 (N_40499,N_36521,N_35034);
nor U40500 (N_40500,N_34591,N_31496);
nand U40501 (N_40501,N_32310,N_38574);
or U40502 (N_40502,N_37740,N_39561);
xnor U40503 (N_40503,N_33899,N_34936);
and U40504 (N_40504,N_36453,N_35228);
xor U40505 (N_40505,N_38791,N_37451);
nand U40506 (N_40506,N_30717,N_39840);
nor U40507 (N_40507,N_38096,N_33256);
and U40508 (N_40508,N_31225,N_33191);
nand U40509 (N_40509,N_33122,N_36002);
or U40510 (N_40510,N_35203,N_39872);
or U40511 (N_40511,N_32278,N_35880);
nand U40512 (N_40512,N_32211,N_32795);
and U40513 (N_40513,N_33586,N_33375);
and U40514 (N_40514,N_37057,N_37352);
and U40515 (N_40515,N_31639,N_36248);
and U40516 (N_40516,N_34053,N_35937);
and U40517 (N_40517,N_33990,N_34374);
nand U40518 (N_40518,N_35754,N_38457);
or U40519 (N_40519,N_35063,N_39388);
or U40520 (N_40520,N_38928,N_31365);
nor U40521 (N_40521,N_39019,N_32130);
nor U40522 (N_40522,N_31441,N_33534);
or U40523 (N_40523,N_37738,N_39402);
or U40524 (N_40524,N_33197,N_32827);
nor U40525 (N_40525,N_31493,N_39276);
or U40526 (N_40526,N_37185,N_30576);
nand U40527 (N_40527,N_39354,N_33298);
and U40528 (N_40528,N_30984,N_38104);
nor U40529 (N_40529,N_32675,N_33139);
or U40530 (N_40530,N_31037,N_36213);
and U40531 (N_40531,N_38223,N_30641);
nor U40532 (N_40532,N_34679,N_39710);
or U40533 (N_40533,N_32380,N_38683);
xor U40534 (N_40534,N_35810,N_39130);
and U40535 (N_40535,N_30263,N_33354);
or U40536 (N_40536,N_39327,N_36496);
and U40537 (N_40537,N_33313,N_36785);
or U40538 (N_40538,N_33300,N_39871);
or U40539 (N_40539,N_33498,N_33353);
or U40540 (N_40540,N_38315,N_34961);
or U40541 (N_40541,N_34612,N_39332);
nand U40542 (N_40542,N_30634,N_35344);
xnor U40543 (N_40543,N_35101,N_39762);
or U40544 (N_40544,N_32291,N_33720);
nor U40545 (N_40545,N_33391,N_34254);
nor U40546 (N_40546,N_30900,N_37813);
nor U40547 (N_40547,N_32914,N_34650);
or U40548 (N_40548,N_32678,N_36294);
nand U40549 (N_40549,N_30325,N_34606);
nor U40550 (N_40550,N_39071,N_38157);
and U40551 (N_40551,N_36625,N_31554);
or U40552 (N_40552,N_32562,N_34510);
nand U40553 (N_40553,N_38585,N_32215);
nand U40554 (N_40554,N_38209,N_34909);
nor U40555 (N_40555,N_35104,N_33477);
xor U40556 (N_40556,N_37302,N_37065);
and U40557 (N_40557,N_39643,N_36633);
xor U40558 (N_40558,N_35152,N_38019);
nand U40559 (N_40559,N_32626,N_33834);
or U40560 (N_40560,N_32246,N_36599);
nor U40561 (N_40561,N_35314,N_30338);
or U40562 (N_40562,N_32342,N_35712);
xor U40563 (N_40563,N_38691,N_34418);
nor U40564 (N_40564,N_37613,N_37762);
nand U40565 (N_40565,N_37005,N_38861);
or U40566 (N_40566,N_34675,N_31678);
nor U40567 (N_40567,N_32116,N_30640);
and U40568 (N_40568,N_32835,N_37355);
or U40569 (N_40569,N_33316,N_37174);
nor U40570 (N_40570,N_38663,N_33148);
and U40571 (N_40571,N_37743,N_39464);
and U40572 (N_40572,N_35584,N_37210);
or U40573 (N_40573,N_30721,N_36049);
nor U40574 (N_40574,N_31617,N_37119);
nand U40575 (N_40575,N_32559,N_39424);
xor U40576 (N_40576,N_35652,N_36553);
nand U40577 (N_40577,N_38037,N_37881);
xor U40578 (N_40578,N_34134,N_37625);
and U40579 (N_40579,N_35489,N_35375);
or U40580 (N_40580,N_33570,N_34852);
or U40581 (N_40581,N_30424,N_32239);
nor U40582 (N_40582,N_36196,N_30888);
or U40583 (N_40583,N_33415,N_35052);
xor U40584 (N_40584,N_31076,N_33160);
and U40585 (N_40585,N_33442,N_36967);
nand U40586 (N_40586,N_33302,N_35523);
nand U40587 (N_40587,N_31427,N_36707);
and U40588 (N_40588,N_31273,N_30996);
or U40589 (N_40589,N_37439,N_35757);
nor U40590 (N_40590,N_38206,N_35230);
or U40591 (N_40591,N_35488,N_35235);
nand U40592 (N_40592,N_39546,N_38450);
or U40593 (N_40593,N_33048,N_36540);
or U40594 (N_40594,N_33325,N_35517);
nand U40595 (N_40595,N_38281,N_33343);
nand U40596 (N_40596,N_38793,N_35566);
nor U40597 (N_40597,N_31306,N_32069);
nor U40598 (N_40598,N_39036,N_31949);
nand U40599 (N_40599,N_31979,N_36157);
or U40600 (N_40600,N_30745,N_39429);
and U40601 (N_40601,N_32962,N_37245);
and U40602 (N_40602,N_37386,N_33283);
nand U40603 (N_40603,N_38074,N_34611);
or U40604 (N_40604,N_37755,N_38582);
and U40605 (N_40605,N_34862,N_37149);
xor U40606 (N_40606,N_35722,N_36418);
and U40607 (N_40607,N_30422,N_37051);
or U40608 (N_40608,N_30609,N_35569);
and U40609 (N_40609,N_38939,N_30227);
xnor U40610 (N_40610,N_30880,N_38766);
xnor U40611 (N_40611,N_37595,N_33978);
and U40612 (N_40612,N_39860,N_33937);
and U40613 (N_40613,N_33985,N_33202);
nor U40614 (N_40614,N_38745,N_31557);
nor U40615 (N_40615,N_32469,N_36174);
xor U40616 (N_40616,N_34869,N_31053);
xnor U40617 (N_40617,N_38234,N_38708);
and U40618 (N_40618,N_39734,N_38381);
nor U40619 (N_40619,N_37971,N_36647);
nor U40620 (N_40620,N_39996,N_31308);
nor U40621 (N_40621,N_33676,N_35332);
and U40622 (N_40622,N_33457,N_34902);
and U40623 (N_40623,N_31140,N_30787);
nor U40624 (N_40624,N_36960,N_34746);
and U40625 (N_40625,N_32325,N_35007);
and U40626 (N_40626,N_30591,N_35743);
xnor U40627 (N_40627,N_32097,N_30018);
and U40628 (N_40628,N_33252,N_30740);
nand U40629 (N_40629,N_34689,N_36701);
and U40630 (N_40630,N_34261,N_30993);
and U40631 (N_40631,N_39365,N_33866);
and U40632 (N_40632,N_35397,N_35408);
or U40633 (N_40633,N_35876,N_30174);
nor U40634 (N_40634,N_35126,N_39166);
or U40635 (N_40635,N_38376,N_36330);
xor U40636 (N_40636,N_32716,N_38040);
nand U40637 (N_40637,N_37833,N_33407);
nand U40638 (N_40638,N_31796,N_35174);
nor U40639 (N_40639,N_30087,N_32983);
or U40640 (N_40640,N_36001,N_30259);
nor U40641 (N_40641,N_38166,N_39012);
or U40642 (N_40642,N_34312,N_37357);
or U40643 (N_40643,N_34235,N_36117);
xnor U40644 (N_40644,N_32843,N_32900);
nor U40645 (N_40645,N_38725,N_30841);
or U40646 (N_40646,N_38757,N_30462);
nor U40647 (N_40647,N_34856,N_39408);
or U40648 (N_40648,N_31934,N_34963);
nor U40649 (N_40649,N_31254,N_31201);
nor U40650 (N_40650,N_36686,N_36605);
nor U40651 (N_40651,N_33059,N_38794);
or U40652 (N_40652,N_32661,N_37448);
and U40653 (N_40653,N_38900,N_31018);
or U40654 (N_40654,N_30769,N_30229);
nand U40655 (N_40655,N_36515,N_39287);
and U40656 (N_40656,N_31262,N_34360);
and U40657 (N_40657,N_36216,N_34375);
nand U40658 (N_40658,N_36252,N_39744);
or U40659 (N_40659,N_30090,N_32701);
and U40660 (N_40660,N_39437,N_34622);
nor U40661 (N_40661,N_39461,N_39570);
nand U40662 (N_40662,N_38716,N_32283);
nand U40663 (N_40663,N_39218,N_36195);
nand U40664 (N_40664,N_36563,N_31674);
nor U40665 (N_40665,N_32461,N_39373);
nand U40666 (N_40666,N_31778,N_38644);
nand U40667 (N_40667,N_36717,N_34696);
and U40668 (N_40668,N_34084,N_31104);
nand U40669 (N_40669,N_36194,N_35570);
nor U40670 (N_40670,N_33565,N_38968);
nor U40671 (N_40671,N_38321,N_34391);
nand U40672 (N_40672,N_30022,N_36754);
or U40673 (N_40673,N_36419,N_36569);
nand U40674 (N_40674,N_36486,N_39905);
nand U40675 (N_40675,N_37144,N_33574);
or U40676 (N_40676,N_38836,N_34813);
or U40677 (N_40677,N_37830,N_31813);
nor U40678 (N_40678,N_31984,N_33649);
nor U40679 (N_40679,N_31373,N_31468);
and U40680 (N_40680,N_34687,N_30669);
xnor U40681 (N_40681,N_33696,N_39038);
and U40682 (N_40682,N_34291,N_30853);
and U40683 (N_40683,N_33456,N_39814);
or U40684 (N_40684,N_37824,N_38454);
and U40685 (N_40685,N_35409,N_31562);
and U40686 (N_40686,N_35865,N_37593);
nand U40687 (N_40687,N_31767,N_35358);
nand U40688 (N_40688,N_35528,N_34732);
xnor U40689 (N_40689,N_30901,N_38947);
nor U40690 (N_40690,N_33812,N_37578);
and U40691 (N_40691,N_32981,N_36678);
and U40692 (N_40692,N_39986,N_37932);
nand U40693 (N_40693,N_33562,N_34128);
xnor U40694 (N_40694,N_30150,N_36178);
or U40695 (N_40695,N_36787,N_33646);
or U40696 (N_40696,N_39656,N_39551);
or U40697 (N_40697,N_36217,N_37086);
nor U40698 (N_40698,N_38293,N_39760);
nand U40699 (N_40699,N_37729,N_30389);
nand U40700 (N_40700,N_36582,N_30393);
nand U40701 (N_40701,N_30313,N_37330);
and U40702 (N_40702,N_36374,N_30260);
xnor U40703 (N_40703,N_37696,N_39748);
nand U40704 (N_40704,N_35732,N_36913);
nand U40705 (N_40705,N_39640,N_36705);
nand U40706 (N_40706,N_31171,N_32395);
nor U40707 (N_40707,N_39819,N_37101);
and U40708 (N_40708,N_38323,N_39824);
nor U40709 (N_40709,N_38647,N_30756);
nor U40710 (N_40710,N_37224,N_36973);
and U40711 (N_40711,N_37552,N_32112);
nor U40712 (N_40712,N_33524,N_30979);
nand U40713 (N_40713,N_33011,N_31864);
nor U40714 (N_40714,N_32225,N_39363);
and U40715 (N_40715,N_33884,N_36571);
nand U40716 (N_40716,N_33367,N_33384);
nor U40717 (N_40717,N_39766,N_32205);
nor U40718 (N_40718,N_38079,N_37554);
nor U40719 (N_40719,N_33345,N_35163);
and U40720 (N_40720,N_36505,N_30565);
nor U40721 (N_40721,N_33530,N_35035);
and U40722 (N_40722,N_38729,N_39737);
and U40723 (N_40723,N_33424,N_38115);
nor U40724 (N_40724,N_37404,N_33591);
nor U40725 (N_40725,N_33103,N_32343);
or U40726 (N_40726,N_33083,N_37178);
or U40727 (N_40727,N_32148,N_30865);
and U40728 (N_40728,N_33847,N_32187);
and U40729 (N_40729,N_35160,N_32118);
or U40730 (N_40730,N_33429,N_34321);
nand U40731 (N_40731,N_30805,N_35043);
nand U40732 (N_40732,N_33487,N_37162);
and U40733 (N_40733,N_35325,N_37844);
nor U40734 (N_40734,N_34888,N_33926);
and U40735 (N_40735,N_33037,N_30036);
nand U40736 (N_40736,N_36810,N_33953);
and U40737 (N_40737,N_32819,N_34030);
and U40738 (N_40738,N_30469,N_31470);
and U40739 (N_40739,N_33626,N_35921);
nand U40740 (N_40740,N_34249,N_39110);
nand U40741 (N_40741,N_38395,N_31935);
nand U40742 (N_40742,N_32360,N_36382);
xnor U40743 (N_40743,N_33092,N_30432);
or U40744 (N_40744,N_37897,N_32432);
nor U40745 (N_40745,N_39848,N_30708);
or U40746 (N_40746,N_31451,N_30189);
or U40747 (N_40747,N_35095,N_35582);
or U40748 (N_40748,N_38368,N_31886);
nand U40749 (N_40749,N_36644,N_38670);
or U40750 (N_40750,N_33971,N_39521);
or U40751 (N_40751,N_34016,N_38608);
xnor U40752 (N_40752,N_34726,N_33211);
and U40753 (N_40753,N_33760,N_31839);
or U40754 (N_40754,N_38489,N_35854);
and U40755 (N_40755,N_34579,N_34148);
and U40756 (N_40756,N_33513,N_35525);
nand U40757 (N_40757,N_31694,N_30045);
or U40758 (N_40758,N_30876,N_32344);
nor U40759 (N_40759,N_33643,N_39478);
and U40760 (N_40760,N_31675,N_37733);
and U40761 (N_40761,N_34320,N_32690);
nor U40762 (N_40762,N_31334,N_34753);
nor U40763 (N_40763,N_38542,N_32178);
or U40764 (N_40764,N_36651,N_36809);
nand U40765 (N_40765,N_30933,N_37221);
xnor U40766 (N_40766,N_35279,N_35442);
or U40767 (N_40767,N_31500,N_37395);
and U40768 (N_40768,N_30410,N_39992);
and U40769 (N_40769,N_32875,N_32970);
and U40770 (N_40770,N_38777,N_33949);
and U40771 (N_40771,N_33793,N_34616);
and U40772 (N_40772,N_35875,N_37508);
or U40773 (N_40773,N_34356,N_35708);
or U40774 (N_40774,N_34769,N_34867);
or U40775 (N_40775,N_38655,N_36222);
and U40776 (N_40776,N_39716,N_37171);
or U40777 (N_40777,N_38831,N_39647);
or U40778 (N_40778,N_33802,N_31194);
nor U40779 (N_40779,N_34114,N_37006);
and U40780 (N_40780,N_39340,N_35297);
or U40781 (N_40781,N_32901,N_36205);
or U40782 (N_40782,N_38673,N_36506);
and U40783 (N_40783,N_39050,N_34298);
and U40784 (N_40784,N_30830,N_31329);
xnor U40785 (N_40785,N_34210,N_30358);
nor U40786 (N_40786,N_34734,N_31486);
xnor U40787 (N_40787,N_37305,N_35672);
and U40788 (N_40788,N_30533,N_37805);
and U40789 (N_40789,N_35604,N_34624);
nand U40790 (N_40790,N_32355,N_36048);
xor U40791 (N_40791,N_30596,N_38087);
or U40792 (N_40792,N_35930,N_39344);
nand U40793 (N_40793,N_36727,N_31116);
nand U40794 (N_40794,N_33009,N_34870);
nor U40795 (N_40795,N_37004,N_38137);
nor U40796 (N_40796,N_36938,N_37633);
nand U40797 (N_40797,N_32742,N_36649);
and U40798 (N_40798,N_36580,N_37974);
xnor U40799 (N_40799,N_30166,N_35979);
or U40800 (N_40800,N_36548,N_30505);
nand U40801 (N_40801,N_32572,N_39510);
and U40802 (N_40802,N_37889,N_33669);
nor U40803 (N_40803,N_39209,N_30879);
and U40804 (N_40804,N_34446,N_30791);
xnor U40805 (N_40805,N_31640,N_39061);
or U40806 (N_40806,N_38357,N_31275);
nor U40807 (N_40807,N_39138,N_34454);
nand U40808 (N_40808,N_36356,N_36781);
nand U40809 (N_40809,N_33238,N_35799);
nand U40810 (N_40810,N_31754,N_32327);
nand U40811 (N_40811,N_36729,N_31749);
or U40812 (N_40812,N_37887,N_30541);
nor U40813 (N_40813,N_32939,N_32382);
nand U40814 (N_40814,N_31335,N_32767);
nand U40815 (N_40815,N_35533,N_36499);
and U40816 (N_40816,N_31971,N_38699);
nand U40817 (N_40817,N_32424,N_34764);
and U40818 (N_40818,N_31369,N_36295);
nand U40819 (N_40819,N_33170,N_33598);
nor U40820 (N_40820,N_36383,N_37040);
and U40821 (N_40821,N_39654,N_37321);
nand U40822 (N_40822,N_38541,N_37503);
nand U40823 (N_40823,N_35147,N_39469);
nor U40824 (N_40824,N_37765,N_39697);
or U40825 (N_40825,N_38069,N_36074);
nand U40826 (N_40826,N_39281,N_31908);
or U40827 (N_40827,N_36368,N_38522);
or U40828 (N_40828,N_31482,N_39578);
nor U40829 (N_40829,N_31047,N_33889);
and U40830 (N_40830,N_31420,N_32810);
nor U40831 (N_40831,N_33436,N_30069);
or U40832 (N_40832,N_39989,N_36036);
or U40833 (N_40833,N_30453,N_34766);
nor U40834 (N_40834,N_30573,N_33262);
nor U40835 (N_40835,N_36024,N_31710);
nor U40836 (N_40836,N_39794,N_32932);
nor U40837 (N_40837,N_34096,N_39389);
and U40838 (N_40838,N_37264,N_33394);
nor U40839 (N_40839,N_38902,N_34819);
nand U40840 (N_40840,N_37001,N_36170);
and U40841 (N_40841,N_31830,N_34770);
or U40842 (N_40842,N_32852,N_37054);
nor U40843 (N_40843,N_33072,N_30197);
nand U40844 (N_40844,N_38088,N_32727);
nand U40845 (N_40845,N_36066,N_32881);
or U40846 (N_40846,N_37426,N_39701);
and U40847 (N_40847,N_33199,N_35088);
nor U40848 (N_40848,N_36209,N_34179);
xor U40849 (N_40849,N_33473,N_39935);
nor U40850 (N_40850,N_32227,N_30027);
nor U40851 (N_40851,N_36714,N_37611);
xor U40852 (N_40852,N_39738,N_33804);
and U40853 (N_40853,N_39678,N_36053);
and U40854 (N_40854,N_35346,N_37661);
xor U40855 (N_40855,N_38324,N_34199);
nor U40856 (N_40856,N_31219,N_39049);
and U40857 (N_40857,N_31364,N_34643);
nand U40858 (N_40858,N_37020,N_39803);
and U40859 (N_40859,N_30188,N_30899);
xor U40860 (N_40860,N_39543,N_39316);
or U40861 (N_40861,N_32653,N_33309);
nand U40862 (N_40862,N_32528,N_36688);
and U40863 (N_40863,N_30081,N_39718);
nand U40864 (N_40864,N_38847,N_39214);
nor U40865 (N_40865,N_36889,N_36558);
xnor U40866 (N_40866,N_36316,N_31853);
nand U40867 (N_40867,N_31894,N_31466);
or U40868 (N_40868,N_31454,N_32838);
nand U40869 (N_40869,N_32352,N_36946);
nor U40870 (N_40870,N_39844,N_39409);
and U40871 (N_40871,N_38809,N_37643);
nor U40872 (N_40872,N_37710,N_33989);
and U40873 (N_40873,N_38373,N_39567);
nand U40874 (N_40874,N_30217,N_32535);
or U40875 (N_40875,N_30233,N_32928);
nand U40876 (N_40876,N_32989,N_34079);
nand U40877 (N_40877,N_38511,N_33143);
nand U40878 (N_40878,N_31309,N_36912);
or U40879 (N_40879,N_30109,N_30892);
nor U40880 (N_40880,N_31553,N_38798);
nor U40881 (N_40881,N_35502,N_36029);
nor U40882 (N_40882,N_39252,N_38036);
nor U40883 (N_40883,N_31964,N_33395);
and U40884 (N_40884,N_33098,N_34943);
nor U40885 (N_40885,N_31746,N_31859);
nand U40886 (N_40886,N_33902,N_34380);
nand U40887 (N_40887,N_36942,N_35529);
nor U40888 (N_40888,N_35790,N_37962);
or U40889 (N_40889,N_39770,N_36901);
and U40890 (N_40890,N_37896,N_30857);
nor U40891 (N_40891,N_35060,N_31631);
nand U40892 (N_40892,N_30074,N_33445);
xor U40893 (N_40893,N_37294,N_36076);
nor U40894 (N_40894,N_38812,N_36551);
and U40895 (N_40895,N_34914,N_36221);
nor U40896 (N_40896,N_39043,N_38369);
nor U40897 (N_40897,N_33263,N_36757);
or U40898 (N_40898,N_38611,N_37124);
nor U40899 (N_40899,N_35420,N_35837);
xor U40900 (N_40900,N_30726,N_31538);
xnor U40901 (N_40901,N_36037,N_36597);
xnor U40902 (N_40902,N_34115,N_39669);
nor U40903 (N_40903,N_34705,N_31074);
or U40904 (N_40904,N_37419,N_37867);
or U40905 (N_40905,N_36448,N_35620);
nand U40906 (N_40906,N_38316,N_36654);
nor U40907 (N_40907,N_39809,N_32268);
or U40908 (N_40908,N_34669,N_31923);
and U40909 (N_40909,N_32745,N_32253);
nor U40910 (N_40910,N_39443,N_30778);
and U40911 (N_40911,N_35622,N_33124);
xnor U40912 (N_40912,N_31436,N_31223);
nand U40913 (N_40913,N_30154,N_39151);
nand U40914 (N_40914,N_31721,N_31755);
nor U40915 (N_40915,N_33130,N_30605);
or U40916 (N_40916,N_37411,N_38438);
nor U40917 (N_40917,N_31844,N_30796);
and U40918 (N_40918,N_39625,N_35270);
and U40919 (N_40919,N_33447,N_38835);
or U40920 (N_40920,N_30232,N_39356);
or U40921 (N_40921,N_30883,N_32400);
or U40922 (N_40922,N_34692,N_38221);
nand U40923 (N_40923,N_37976,N_33329);
or U40924 (N_40924,N_32385,N_34433);
nand U40925 (N_40925,N_35833,N_33337);
nor U40926 (N_40926,N_33214,N_32230);
nor U40927 (N_40927,N_35986,N_36573);
nor U40928 (N_40928,N_30909,N_34797);
and U40929 (N_40929,N_33068,N_39165);
nor U40930 (N_40930,N_35561,N_35626);
nand U40931 (N_40931,N_31247,N_32652);
and U40932 (N_40932,N_31614,N_35157);
nor U40933 (N_40933,N_33243,N_37088);
and U40934 (N_40934,N_36559,N_34659);
or U40935 (N_40935,N_32691,N_31479);
nor U40936 (N_40936,N_36343,N_33460);
and U40937 (N_40937,N_34546,N_30928);
and U40938 (N_40938,N_32561,N_33636);
nand U40939 (N_40939,N_30507,N_39666);
and U40940 (N_40940,N_36214,N_33723);
and U40941 (N_40941,N_38273,N_38313);
xnor U40942 (N_40942,N_30652,N_31874);
and U40943 (N_40943,N_38054,N_34369);
or U40944 (N_40944,N_34364,N_36460);
or U40945 (N_40945,N_35996,N_36284);
nor U40946 (N_40946,N_38612,N_31686);
or U40947 (N_40947,N_39622,N_36377);
and U40948 (N_40948,N_33520,N_39971);
or U40949 (N_40949,N_32081,N_37566);
nor U40950 (N_40950,N_33418,N_34189);
xnor U40951 (N_40951,N_34062,N_38443);
nor U40952 (N_40952,N_34795,N_30566);
or U40953 (N_40953,N_31876,N_34608);
and U40954 (N_40954,N_38141,N_30961);
and U40955 (N_40955,N_39523,N_37708);
and U40956 (N_40956,N_30513,N_32495);
and U40957 (N_40957,N_34412,N_34414);
nor U40958 (N_40958,N_38569,N_30447);
or U40959 (N_40959,N_38973,N_31717);
or U40960 (N_40960,N_34644,N_36389);
nor U40961 (N_40961,N_31272,N_39893);
nor U40962 (N_40962,N_38614,N_32694);
nor U40963 (N_40963,N_39563,N_31487);
nand U40964 (N_40964,N_35341,N_35769);
nand U40965 (N_40965,N_31040,N_36939);
nor U40966 (N_40966,N_36386,N_37641);
nor U40967 (N_40967,N_39328,N_34878);
nand U40968 (N_40968,N_31918,N_30242);
xnor U40969 (N_40969,N_33261,N_33657);
nor U40970 (N_40970,N_36683,N_39317);
nor U40971 (N_40971,N_39004,N_32648);
nand U40972 (N_40972,N_36402,N_34306);
and U40973 (N_40973,N_31043,N_37562);
or U40974 (N_40974,N_35099,N_35419);
nor U40975 (N_40975,N_32046,N_38908);
nor U40976 (N_40976,N_39960,N_32831);
nand U40977 (N_40977,N_33390,N_37073);
and U40978 (N_40978,N_30736,N_37153);
nand U40979 (N_40979,N_31781,N_37544);
or U40980 (N_40980,N_36585,N_31641);
and U40981 (N_40981,N_32565,N_37726);
nand U40982 (N_40982,N_33102,N_36536);
nand U40983 (N_40983,N_39651,N_32135);
nand U40984 (N_40984,N_32207,N_32809);
nand U40985 (N_40985,N_34168,N_35894);
and U40986 (N_40986,N_36730,N_33322);
or U40987 (N_40987,N_31269,N_35701);
and U40988 (N_40988,N_33935,N_33701);
and U40989 (N_40989,N_32363,N_38826);
and U40990 (N_40990,N_30239,N_34142);
and U40991 (N_40991,N_30553,N_30644);
or U40992 (N_40992,N_34301,N_38499);
or U40993 (N_40993,N_39368,N_36232);
nor U40994 (N_40994,N_39799,N_34077);
or U40995 (N_40995,N_37189,N_38418);
and U40996 (N_40996,N_36113,N_34267);
nor U40997 (N_40997,N_39082,N_39994);
nand U40998 (N_40998,N_34901,N_34285);
and U40999 (N_40999,N_36744,N_33396);
or U41000 (N_41000,N_37823,N_36821);
and U41001 (N_41001,N_30234,N_30518);
and U41002 (N_41002,N_38403,N_31604);
and U41003 (N_41003,N_36023,N_33469);
nand U41004 (N_41004,N_37659,N_31587);
or U41005 (N_41005,N_30287,N_35371);
nand U41006 (N_41006,N_35861,N_36557);
nand U41007 (N_41007,N_39890,N_39310);
and U41008 (N_41008,N_36190,N_39215);
xnor U41009 (N_41009,N_35819,N_36524);
and U41010 (N_41010,N_33640,N_39288);
nand U41011 (N_41011,N_36071,N_37191);
nand U41012 (N_41012,N_38426,N_32551);
nand U41013 (N_41013,N_33879,N_32556);
xnor U41014 (N_41014,N_39341,N_30648);
and U41015 (N_41015,N_37569,N_31941);
nand U41016 (N_41016,N_30159,N_31565);
nand U41017 (N_41017,N_38509,N_32454);
nand U41018 (N_41018,N_36902,N_30271);
and U41019 (N_41019,N_37586,N_39454);
or U41020 (N_41020,N_30632,N_34938);
or U41021 (N_41021,N_37444,N_35123);
and U41022 (N_41022,N_39315,N_30319);
or U41023 (N_41023,N_37797,N_32056);
xnor U41024 (N_41024,N_33795,N_31827);
nand U41025 (N_41025,N_33547,N_30674);
nor U41026 (N_41026,N_36984,N_34064);
xnor U41027 (N_41027,N_35577,N_39739);
nor U41028 (N_41028,N_35852,N_35075);
nor U41029 (N_41029,N_32509,N_31630);
nor U41030 (N_41030,N_32855,N_32808);
or U41031 (N_41031,N_36336,N_33977);
and U41032 (N_41032,N_31655,N_38308);
nor U41033 (N_41033,N_31667,N_35784);
or U41034 (N_41034,N_30929,N_38195);
and U41035 (N_41035,N_30173,N_33763);
nand U41036 (N_41036,N_31090,N_30441);
and U41037 (N_41037,N_33915,N_34512);
or U41038 (N_41038,N_32010,N_32599);
and U41039 (N_41039,N_32212,N_33267);
and U41040 (N_41040,N_31299,N_31444);
nor U41041 (N_41041,N_30727,N_32947);
nor U41042 (N_41042,N_36317,N_36985);
or U41043 (N_41043,N_37223,N_32353);
nor U41044 (N_41044,N_35826,N_30711);
and U41045 (N_41045,N_39696,N_39268);
and U41046 (N_41046,N_32756,N_33504);
and U41047 (N_41047,N_37960,N_32674);
and U41048 (N_41048,N_38047,N_32228);
or U41049 (N_41049,N_35905,N_34371);
nand U41050 (N_41050,N_35621,N_39961);
nand U41051 (N_41051,N_33778,N_36951);
nor U41052 (N_41052,N_38660,N_37145);
and U41053 (N_41053,N_37721,N_31166);
or U41054 (N_41054,N_37422,N_37303);
nand U41055 (N_41055,N_32158,N_34247);
or U41056 (N_41056,N_30195,N_38389);
xor U41057 (N_41057,N_34607,N_34551);
nor U41058 (N_41058,N_38756,N_35258);
nand U41059 (N_41059,N_31946,N_32009);
or U41060 (N_41060,N_34906,N_31180);
nor U41061 (N_41061,N_33958,N_32663);
nor U41062 (N_41062,N_38261,N_33709);
or U41063 (N_41063,N_38977,N_38477);
nor U41064 (N_41064,N_34257,N_32788);
nand U41065 (N_41065,N_39101,N_36776);
nor U41066 (N_41066,N_32649,N_34573);
nor U41067 (N_41067,N_37334,N_30985);
and U41068 (N_41068,N_36109,N_33377);
and U41069 (N_41069,N_32737,N_35240);
nand U41070 (N_41070,N_31268,N_32204);
or U41071 (N_41071,N_31471,N_34130);
and U41072 (N_41072,N_33178,N_33107);
and U41073 (N_41073,N_33304,N_30956);
or U41074 (N_41074,N_37803,N_35184);
or U41075 (N_41075,N_38760,N_35505);
nand U41076 (N_41076,N_35086,N_35939);
or U41077 (N_41077,N_30582,N_39859);
nand U41078 (N_41078,N_30115,N_30010);
or U41079 (N_41079,N_30770,N_31688);
xor U41080 (N_41080,N_35698,N_34749);
or U41081 (N_41081,N_37131,N_35412);
nand U41082 (N_41082,N_38119,N_33452);
nand U41083 (N_41083,N_37982,N_31196);
and U41084 (N_41084,N_36331,N_38744);
nor U41085 (N_41085,N_34789,N_31648);
xor U41086 (N_41086,N_32976,N_33786);
or U41087 (N_41087,N_31897,N_39611);
xnor U41088 (N_41088,N_34129,N_39726);
nor U41089 (N_41089,N_36136,N_37694);
nor U41090 (N_41090,N_33962,N_38382);
nor U41091 (N_41091,N_33909,N_36920);
nor U41092 (N_41092,N_36672,N_35380);
or U41093 (N_41093,N_30623,N_34633);
nor U41094 (N_41094,N_31136,N_39441);
nand U41095 (N_41095,N_30558,N_34864);
or U41096 (N_41096,N_32142,N_32252);
or U41097 (N_41097,N_37392,N_33719);
nor U41098 (N_41098,N_31162,N_30660);
nand U41099 (N_41099,N_34328,N_39005);
nand U41100 (N_41100,N_33104,N_38874);
nor U41101 (N_41101,N_35463,N_36319);
nor U41102 (N_41102,N_35817,N_35946);
or U41103 (N_41103,N_30572,N_38597);
and U41104 (N_41104,N_32473,N_32578);
nor U41105 (N_41105,N_31302,N_32667);
nand U41106 (N_41106,N_30997,N_34725);
or U41107 (N_41107,N_35441,N_30184);
nand U41108 (N_41108,N_31226,N_36971);
nand U41109 (N_41109,N_38531,N_32314);
nor U41110 (N_41110,N_33495,N_39634);
or U41111 (N_41111,N_38624,N_32871);
or U41112 (N_41112,N_37418,N_30362);
and U41113 (N_41113,N_30822,N_38526);
nor U41114 (N_41114,N_39351,N_33829);
nor U41115 (N_41115,N_37165,N_36882);
or U41116 (N_41116,N_38966,N_38113);
nand U41117 (N_41117,N_32195,N_39114);
nor U41118 (N_41118,N_38306,N_39219);
or U41119 (N_41119,N_33673,N_32594);
nand U41120 (N_41120,N_39169,N_33624);
or U41121 (N_41121,N_31087,N_36916);
nor U41122 (N_41122,N_36398,N_30329);
or U41123 (N_41123,N_33251,N_36313);
nor U41124 (N_41124,N_34097,N_38228);
nand U41125 (N_41125,N_36530,N_34731);
or U41126 (N_41126,N_37782,N_36306);
and U41127 (N_41127,N_34701,N_30310);
or U41128 (N_41128,N_36928,N_32261);
nand U41129 (N_41129,N_30118,N_35550);
or U41130 (N_41130,N_38176,N_30489);
xor U41131 (N_41131,N_31342,N_39808);
or U41132 (N_41132,N_39531,N_31184);
or U41133 (N_41133,N_36768,N_38456);
nor U41134 (N_41134,N_38216,N_39939);
nor U41135 (N_41135,N_35756,N_36379);
nand U41136 (N_41136,N_37324,N_39117);
and U41137 (N_41137,N_38125,N_30520);
nand U41138 (N_41138,N_33479,N_31083);
nor U41139 (N_41139,N_33641,N_37023);
nor U41140 (N_41140,N_34986,N_35113);
and U41141 (N_41141,N_31887,N_35214);
nor U41142 (N_41142,N_33100,N_39512);
and U41143 (N_41143,N_33433,N_32262);
or U41144 (N_41144,N_33644,N_35636);
and U41145 (N_41145,N_39199,N_39170);
nor U41146 (N_41146,N_30989,N_34997);
and U41147 (N_41147,N_33878,N_32276);
nor U41148 (N_41148,N_39797,N_32607);
nor U41149 (N_41149,N_35549,N_39534);
nor U41150 (N_41150,N_33929,N_34905);
nand U41151 (N_41151,N_34817,N_37831);
or U41152 (N_41152,N_37095,N_34839);
nor U41153 (N_41153,N_36808,N_30345);
and U41154 (N_41154,N_32169,N_34686);
xnor U41155 (N_41155,N_36561,N_32413);
or U41156 (N_41156,N_30611,N_37612);
nor U41157 (N_41157,N_32595,N_39952);
nand U41158 (N_41158,N_31462,N_33544);
nor U41159 (N_41159,N_35633,N_30540);
xor U41160 (N_41160,N_30604,N_30743);
nand U41161 (N_41161,N_34465,N_36237);
or U41162 (N_41162,N_32011,N_30398);
nand U41163 (N_41163,N_34796,N_38722);
nand U41164 (N_41164,N_33046,N_35867);
or U41165 (N_41165,N_35286,N_34131);
nand U41166 (N_41166,N_36181,N_35742);
nand U41167 (N_41167,N_32146,N_34122);
and U41168 (N_41168,N_32541,N_32773);
and U41169 (N_41169,N_31371,N_32646);
and U41170 (N_41170,N_31783,N_33764);
nand U41171 (N_41171,N_38512,N_34353);
or U41172 (N_41172,N_35369,N_35684);
nor U41173 (N_41173,N_39109,N_37609);
nor U41174 (N_41174,N_37874,N_36073);
or U41175 (N_41175,N_34879,N_34463);
or U41176 (N_41176,N_37356,N_31450);
and U41177 (N_41177,N_34302,N_36670);
and U41178 (N_41178,N_35702,N_33903);
nor U41179 (N_41179,N_36851,N_32466);
or U41180 (N_41180,N_32071,N_31561);
and U41181 (N_41181,N_34854,N_36990);
or U41182 (N_41182,N_39416,N_32000);
nand U41183 (N_41183,N_37777,N_39419);
nand U41184 (N_41184,N_36773,N_31107);
xnor U41185 (N_41185,N_38297,N_34055);
nor U41186 (N_41186,N_35669,N_37435);
nor U41187 (N_41187,N_33493,N_32598);
and U41188 (N_41188,N_38893,N_33464);
nand U41189 (N_41189,N_30772,N_35145);
or U41190 (N_41190,N_35000,N_37044);
nand U41191 (N_41191,N_32068,N_37895);
and U41192 (N_41192,N_38198,N_32223);
nand U41193 (N_41193,N_34523,N_31743);
nor U41194 (N_41194,N_39234,N_32045);
nand U41195 (N_41195,N_31711,N_33678);
or U41196 (N_41196,N_35932,N_34081);
and U41197 (N_41197,N_30030,N_34912);
or U41198 (N_41198,N_38959,N_31956);
nand U41199 (N_41199,N_33317,N_30725);
nand U41200 (N_41200,N_38945,N_37190);
or U41201 (N_41201,N_39089,N_39607);
nor U41202 (N_41202,N_32270,N_32060);
or U41203 (N_41203,N_38365,N_30457);
and U41204 (N_41204,N_38227,N_36855);
and U41205 (N_41205,N_39597,N_36955);
or U41206 (N_41206,N_38375,N_34001);
or U41207 (N_41207,N_36404,N_38770);
nand U41208 (N_41208,N_37679,N_33955);
nor U41209 (N_41209,N_30601,N_37604);
nor U41210 (N_41210,N_37056,N_36866);
or U41211 (N_41211,N_39162,N_38452);
nand U41212 (N_41212,N_32590,N_30748);
nand U41213 (N_41213,N_37248,N_33845);
nor U41214 (N_41214,N_37793,N_31515);
and U41215 (N_41215,N_31646,N_34944);
or U41216 (N_41216,N_37653,N_34592);
nand U41217 (N_41217,N_30119,N_33529);
and U41218 (N_41218,N_34411,N_38736);
nand U41219 (N_41219,N_33925,N_37854);
nand U41220 (N_41220,N_38591,N_35136);
nor U41221 (N_41221,N_38341,N_34061);
or U41222 (N_41222,N_33959,N_36783);
xor U41223 (N_41223,N_36434,N_37143);
xor U41224 (N_41224,N_39864,N_37342);
xnor U41225 (N_41225,N_34005,N_39452);
nor U41226 (N_41226,N_37376,N_31734);
xor U41227 (N_41227,N_30186,N_33368);
and U41228 (N_41228,N_39072,N_39383);
nand U41229 (N_41229,N_34327,N_31390);
nand U41230 (N_41230,N_39226,N_33964);
and U41231 (N_41231,N_32805,N_35927);
nand U41232 (N_41232,N_39759,N_34932);
nor U41233 (N_41233,N_37361,N_30714);
or U41234 (N_41234,N_38540,N_34507);
nor U41235 (N_41235,N_35929,N_39852);
and U41236 (N_41236,N_33604,N_39793);
nand U41237 (N_41237,N_39045,N_36762);
nand U41238 (N_41238,N_34390,N_36853);
nor U41239 (N_41239,N_31150,N_39308);
and U41240 (N_41240,N_35236,N_32587);
or U41241 (N_41241,N_31210,N_33871);
nand U41242 (N_41242,N_34884,N_38801);
nor U41243 (N_41243,N_38575,N_30220);
xor U41244 (N_41244,N_33996,N_30664);
xor U41245 (N_41245,N_34036,N_35603);
xnor U41246 (N_41246,N_39325,N_39066);
nand U41247 (N_41247,N_30794,N_36965);
and U41248 (N_41248,N_31582,N_37371);
nor U41249 (N_41249,N_30396,N_38700);
and U41250 (N_41250,N_38488,N_37990);
or U41251 (N_41251,N_33120,N_31339);
nor U41252 (N_41252,N_34112,N_34850);
and U41253 (N_41253,N_33897,N_33182);
nand U41254 (N_41254,N_36004,N_32442);
and U41255 (N_41255,N_34505,N_39513);
or U41256 (N_41256,N_30806,N_36635);
nand U41257 (N_41257,N_34706,N_32718);
nand U41258 (N_41258,N_31776,N_39516);
xnor U41259 (N_41259,N_30192,N_37009);
and U41260 (N_41260,N_38278,N_33117);
nor U41261 (N_41261,N_36827,N_31737);
and U41262 (N_41262,N_32558,N_34545);
and U41263 (N_41263,N_36069,N_32999);
and U41264 (N_41264,N_36415,N_37017);
or U41265 (N_41265,N_32184,N_30222);
and U41266 (N_41266,N_35105,N_33877);
nor U41267 (N_41267,N_32916,N_33606);
or U41268 (N_41268,N_31904,N_36958);
xnor U41269 (N_41269,N_31970,N_30915);
and U41270 (N_41270,N_34471,N_32977);
nor U41271 (N_41271,N_38975,N_39480);
nor U41272 (N_41272,N_35098,N_32596);
or U41273 (N_41273,N_38128,N_32182);
and U41274 (N_41274,N_33998,N_35891);
nor U41275 (N_41275,N_32079,N_34697);
nand U41276 (N_41276,N_38942,N_30013);
and U41277 (N_41277,N_35738,N_32299);
and U41278 (N_41278,N_31883,N_39846);
nor U41279 (N_41279,N_33062,N_30137);
nand U41280 (N_41280,N_31988,N_30958);
nor U41281 (N_41281,N_34872,N_39141);
and U41282 (N_41282,N_36661,N_35843);
nand U41283 (N_41283,N_38686,N_31705);
and U41284 (N_41284,N_32507,N_37592);
nor U41285 (N_41285,N_37476,N_32927);
nor U41286 (N_41286,N_33674,N_35146);
nand U41287 (N_41287,N_37296,N_34531);
nand U41288 (N_41288,N_36940,N_32214);
or U41289 (N_41289,N_32108,N_36142);
nand U41290 (N_41290,N_35606,N_30006);
and U41291 (N_41291,N_38828,N_31616);
nand U41292 (N_41292,N_39174,N_31258);
or U41293 (N_41293,N_30459,N_33150);
nor U41294 (N_41294,N_31094,N_32099);
and U41295 (N_41295,N_34330,N_31351);
and U41296 (N_41296,N_38464,N_31502);
xor U41297 (N_41297,N_39842,N_36650);
and U41298 (N_41298,N_35460,N_32455);
and U41299 (N_41299,N_39501,N_30884);
and U41300 (N_41300,N_37663,N_35680);
or U41301 (N_41301,N_31221,N_31205);
nand U41302 (N_41302,N_33927,N_32311);
or U41303 (N_41303,N_33578,N_34292);
nor U41304 (N_41304,N_38046,N_33245);
nor U41305 (N_41305,N_35115,N_39806);
or U41306 (N_41306,N_38718,N_38743);
nand U41307 (N_41307,N_30783,N_35882);
or U41308 (N_41308,N_39496,N_30797);
and U41309 (N_41309,N_30891,N_38738);
and U41310 (N_41310,N_31706,N_37292);
nor U41311 (N_41311,N_38741,N_36957);
and U41312 (N_41312,N_32677,N_30657);
or U41313 (N_41313,N_30659,N_33344);
nand U41314 (N_41314,N_30373,N_35217);
xor U41315 (N_41315,N_30777,N_35162);
or U41316 (N_41316,N_38388,N_32941);
or U41317 (N_41317,N_34930,N_33042);
nand U41318 (N_41318,N_35665,N_38687);
nand U41319 (N_41319,N_37531,N_39724);
and U41320 (N_41320,N_34933,N_30379);
and U41321 (N_41321,N_30904,N_33870);
nor U41322 (N_41322,N_35651,N_31422);
nand U41323 (N_41323,N_35662,N_33975);
nor U41324 (N_41324,N_31893,N_37107);
and U41325 (N_41325,N_31112,N_32035);
nand U41326 (N_41326,N_39895,N_39477);
or U41327 (N_41327,N_30523,N_34897);
and U41328 (N_41328,N_38987,N_32790);
or U41329 (N_41329,N_36999,N_32543);
or U41330 (N_41330,N_32849,N_35825);
nor U41331 (N_41331,N_39140,N_39687);
or U41332 (N_41332,N_31085,N_39486);
xor U41333 (N_41333,N_32123,N_36361);
nor U41334 (N_41334,N_30666,N_37123);
and U41335 (N_41335,N_30264,N_34069);
nor U41336 (N_41336,N_30171,N_30551);
nand U41337 (N_41337,N_36950,N_38805);
xor U41338 (N_41338,N_31773,N_33225);
nor U41339 (N_41339,N_32529,N_35531);
and U41340 (N_41340,N_39723,N_36060);
nand U41341 (N_41341,N_36016,N_35377);
xor U41342 (N_41342,N_39847,N_35057);
nor U41343 (N_41343,N_33246,N_38864);
nand U41344 (N_41344,N_39576,N_30647);
or U41345 (N_41345,N_36342,N_30423);
nand U41346 (N_41346,N_37385,N_37207);
nand U41347 (N_41347,N_38146,N_34958);
nor U41348 (N_41348,N_34439,N_32942);
nor U41349 (N_41349,N_31724,N_36699);
nand U41350 (N_41350,N_31759,N_34100);
and U41351 (N_41351,N_33070,N_39812);
nor U41352 (N_41352,N_39124,N_36759);
and U41353 (N_41353,N_31836,N_33713);
nand U41354 (N_41354,N_31579,N_35087);
nor U41355 (N_41355,N_36103,N_34428);
or U41356 (N_41356,N_34895,N_34232);
and U41357 (N_41357,N_39648,N_33706);
or U41358 (N_41358,N_35988,N_35791);
or U41359 (N_41359,N_38402,N_35609);
or U41360 (N_41360,N_37081,N_37289);
xnor U41361 (N_41361,N_38064,N_34448);
or U41362 (N_41362,N_36824,N_34716);
nor U41363 (N_41363,N_37574,N_32577);
nand U41364 (N_41364,N_32361,N_32092);
nor U41365 (N_41365,N_37284,N_30172);
or U41366 (N_41366,N_38241,N_38255);
xnor U41367 (N_41367,N_37206,N_37934);
nand U41368 (N_41368,N_33553,N_35639);
and U41369 (N_41369,N_37581,N_36745);
and U41370 (N_41370,N_30846,N_31101);
or U41371 (N_41371,N_35498,N_36753);
or U41372 (N_41372,N_33253,N_31533);
nor U41373 (N_41373,N_30095,N_34915);
and U41374 (N_41374,N_34076,N_38562);
and U41375 (N_41375,N_33684,N_35587);
xnor U41376 (N_41376,N_36447,N_36996);
nor U41377 (N_41377,N_39303,N_35890);
or U41378 (N_41378,N_33463,N_33774);
nand U41379 (N_41379,N_34251,N_32014);
nor U41380 (N_41380,N_39122,N_32845);
and U41381 (N_41381,N_32029,N_33843);
nor U41382 (N_41382,N_33106,N_32161);
nand U41383 (N_41383,N_30316,N_30543);
or U41384 (N_41384,N_36261,N_38024);
xnor U41385 (N_41385,N_34848,N_39471);
and U41386 (N_41386,N_36265,N_38788);
or U41387 (N_41387,N_31488,N_35089);
and U41388 (N_41388,N_37826,N_36535);
xnor U41389 (N_41389,N_34156,N_32571);
nand U41390 (N_41390,N_33936,N_38631);
nor U41391 (N_41391,N_39972,N_39150);
or U41392 (N_41392,N_34125,N_35242);
nor U41393 (N_41393,N_34585,N_39336);
or U41394 (N_41394,N_32387,N_38169);
nand U41395 (N_41395,N_31417,N_38827);
nand U41396 (N_41396,N_33836,N_33012);
nand U41397 (N_41397,N_33051,N_34691);
and U41398 (N_41398,N_30381,N_32581);
nor U41399 (N_41399,N_30392,N_31612);
nor U41400 (N_41400,N_35977,N_37271);
and U41401 (N_41401,N_39612,N_39321);
or U41402 (N_41402,N_38029,N_33015);
nor U41403 (N_41403,N_39750,N_30614);
and U41404 (N_41404,N_39627,N_31164);
and U41405 (N_41405,N_32028,N_38637);
nor U41406 (N_41406,N_38963,N_36618);
nand U41407 (N_41407,N_36093,N_39293);
nand U41408 (N_41408,N_30957,N_37542);
xor U41409 (N_41409,N_34577,N_32434);
xnor U41410 (N_41410,N_38236,N_38201);
nand U41411 (N_41411,N_34233,N_31793);
nand U41412 (N_41412,N_32890,N_37638);
nand U41413 (N_41413,N_35812,N_39229);
nor U41414 (N_41414,N_34273,N_30339);
nor U41415 (N_41415,N_37584,N_35195);
or U41416 (N_41416,N_32851,N_33579);
nand U41417 (N_41417,N_38106,N_30774);
nand U41418 (N_41418,N_34658,N_32512);
xnor U41419 (N_41419,N_33146,N_38785);
nand U41420 (N_41420,N_38914,N_35612);
nand U41421 (N_41421,N_34894,N_34091);
and U41422 (N_41422,N_30454,N_30160);
xor U41423 (N_41423,N_36738,N_36669);
and U41424 (N_41424,N_31024,N_30525);
or U41425 (N_41425,N_36709,N_37579);
or U41426 (N_41426,N_34182,N_36642);
and U41427 (N_41427,N_36282,N_30839);
nand U41428 (N_41428,N_39228,N_32774);
nor U41429 (N_41429,N_31131,N_30141);
and U41430 (N_41430,N_31807,N_33944);
nor U41431 (N_41431,N_31473,N_32100);
nor U41432 (N_41432,N_30275,N_39077);
nand U41433 (N_41433,N_30547,N_38534);
or U41434 (N_41434,N_33413,N_39683);
xnor U41435 (N_41435,N_33358,N_32502);
or U41436 (N_41436,N_39704,N_36307);
nor U41437 (N_41437,N_33184,N_32894);
or U41438 (N_41438,N_31182,N_35955);
and U41439 (N_41439,N_38765,N_36375);
nor U41440 (N_41440,N_33810,N_36370);
and U41441 (N_41441,N_39502,N_39906);
and U41442 (N_41442,N_34536,N_39171);
xnor U41443 (N_41443,N_39107,N_38774);
nand U41444 (N_41444,N_30941,N_35154);
nand U41445 (N_41445,N_34175,N_30607);
and U41446 (N_41446,N_30043,N_33781);
and U41447 (N_41447,N_30414,N_35127);
nor U41448 (N_41448,N_38666,N_30156);
nor U41449 (N_41449,N_31831,N_38752);
nor U41450 (N_41450,N_37273,N_36648);
or U41451 (N_41451,N_31599,N_32138);
nand U41452 (N_41452,N_30485,N_33951);
xor U41453 (N_41453,N_34229,N_36042);
nand U41454 (N_41454,N_31726,N_30413);
and U41455 (N_41455,N_31319,N_35629);
or U41456 (N_41456,N_32828,N_32199);
nand U41457 (N_41457,N_32811,N_37227);
nor U41458 (N_41458,N_30621,N_34436);
and U41459 (N_41459,N_32823,N_38559);
nor U41460 (N_41460,N_33071,N_33020);
nor U41461 (N_41461,N_34350,N_33642);
nand U41462 (N_41462,N_35021,N_34497);
xor U41463 (N_41463,N_32007,N_32224);
or U41464 (N_41464,N_35049,N_39381);
xnor U41465 (N_41465,N_33662,N_37745);
nor U41466 (N_41466,N_35827,N_30762);
and U41467 (N_41467,N_36668,N_38476);
and U41468 (N_41468,N_36324,N_38897);
or U41469 (N_41469,N_37336,N_37459);
nor U41470 (N_41470,N_39624,N_39901);
and U41471 (N_41471,N_34646,N_35595);
and U41472 (N_41472,N_34220,N_35161);
nor U41473 (N_41473,N_38066,N_35119);
nand U41474 (N_41474,N_37375,N_33084);
xor U41475 (N_41475,N_39781,N_30289);
nand U41476 (N_41476,N_34972,N_31821);
nor U41477 (N_41477,N_33236,N_32043);
and U41478 (N_41478,N_39202,N_32692);
or U41479 (N_41479,N_34871,N_36664);
nand U41480 (N_41480,N_30268,N_34099);
and U41481 (N_41481,N_31297,N_38664);
nor U41482 (N_41482,N_34782,N_34372);
nand U41483 (N_41483,N_37900,N_34479);
xor U41484 (N_41484,N_34567,N_38051);
nor U41485 (N_41485,N_39254,N_36461);
nand U41486 (N_41486,N_38412,N_38712);
and U41487 (N_41487,N_39448,N_39422);
xor U41488 (N_41488,N_32452,N_31603);
or U41489 (N_41489,N_36993,N_34649);
and U41490 (N_41490,N_30944,N_32904);
nand U41491 (N_41491,N_32170,N_36211);
nand U41492 (N_41492,N_30341,N_31858);
nand U41493 (N_41493,N_38008,N_33921);
nand U41494 (N_41494,N_38505,N_37242);
and U41495 (N_41495,N_33710,N_33999);
nand U41496 (N_41496,N_33832,N_36137);
nand U41497 (N_41497,N_37358,N_30750);
and U41498 (N_41498,N_38819,N_30049);
nand U41499 (N_41499,N_37958,N_35112);
nor U41500 (N_41500,N_36911,N_34276);
nand U41501 (N_41501,N_31036,N_38110);
or U41502 (N_41502,N_32527,N_36716);
nor U41503 (N_41503,N_36854,N_33979);
or U41504 (N_41504,N_34810,N_36408);
nand U41505 (N_41505,N_39468,N_35634);
nor U41506 (N_41506,N_30859,N_36935);
or U41507 (N_41507,N_39880,N_34826);
and U41508 (N_41508,N_37776,N_32486);
and U41509 (N_41509,N_31930,N_34741);
nand U41510 (N_41510,N_37473,N_37692);
nand U41511 (N_41511,N_33492,N_34637);
or U41512 (N_41512,N_39526,N_30599);
nand U41513 (N_41513,N_37811,N_35530);
and U41514 (N_41514,N_32125,N_37665);
xor U41515 (N_41515,N_37018,N_34426);
nand U41516 (N_41516,N_34710,N_34831);
nand U41517 (N_41517,N_37687,N_34177);
nor U41518 (N_41518,N_38147,N_34597);
nor U41519 (N_41519,N_31310,N_32560);
nor U41520 (N_41520,N_34777,N_34352);
nand U41521 (N_41521,N_38417,N_37505);
nand U41522 (N_41522,N_37736,N_35866);
nor U41523 (N_41523,N_30651,N_32470);
or U41524 (N_41524,N_38572,N_33783);
nand U41525 (N_41525,N_37888,N_36320);
nor U41526 (N_41526,N_31401,N_38153);
or U41527 (N_41527,N_38018,N_34868);
nor U41528 (N_41528,N_36814,N_36173);
nand U41529 (N_41529,N_31311,N_37022);
nand U41530 (N_41530,N_30819,N_32200);
and U41531 (N_41531,N_34787,N_39113);
nor U41532 (N_41532,N_39052,N_33683);
nand U41533 (N_41533,N_35069,N_39092);
nand U41534 (N_41534,N_39804,N_36464);
and U41535 (N_41535,N_30179,N_32033);
nand U41536 (N_41536,N_30076,N_36100);
nor U41537 (N_41537,N_36055,N_37154);
nor U41538 (N_41538,N_33135,N_35667);
and U41539 (N_41539,N_31345,N_39787);
nand U41540 (N_41540,N_37806,N_36987);
nand U41541 (N_41541,N_35068,N_39121);
nor U41542 (N_41542,N_37374,N_38479);
or U41543 (N_41543,N_37136,N_33742);
or U41544 (N_41544,N_34812,N_32624);
or U41545 (N_41545,N_31324,N_39725);
nor U41546 (N_41546,N_38124,N_36159);
nor U41547 (N_41547,N_32175,N_37199);
nand U41548 (N_41548,N_30368,N_34863);
xor U41549 (N_41549,N_30522,N_37217);
nand U41550 (N_41550,N_33519,N_39476);
nor U41551 (N_41551,N_31492,N_32506);
and U41552 (N_41552,N_36522,N_35536);
and U41553 (N_41553,N_30960,N_36251);
or U41554 (N_41554,N_31906,N_31144);
or U41555 (N_41555,N_37168,N_34671);
or U41556 (N_41556,N_32891,N_30914);
nand U41557 (N_41557,N_32869,N_32439);
or U41558 (N_41558,N_37208,N_34842);
and U41559 (N_41559,N_30477,N_36329);
or U41560 (N_41560,N_38500,N_33739);
nand U41561 (N_41561,N_39751,N_32848);
nand U41562 (N_41562,N_35192,N_33765);
xor U41563 (N_41563,N_39949,N_38551);
or U41564 (N_41564,N_39055,N_32715);
or U41565 (N_41565,N_31911,N_31857);
nor U41566 (N_41566,N_36312,N_33467);
nor U41567 (N_41567,N_30636,N_30571);
or U41568 (N_41568,N_38387,N_31589);
or U41569 (N_41569,N_31141,N_37919);
nand U41570 (N_41570,N_35798,N_36000);
xor U41571 (N_41571,N_30468,N_31791);
nor U41572 (N_41572,N_30484,N_31921);
xor U41573 (N_41573,N_32500,N_33061);
xor U41574 (N_41574,N_30246,N_39173);
and U41575 (N_41575,N_39519,N_32384);
and U41576 (N_41576,N_31429,N_35426);
and U41577 (N_41577,N_31019,N_32682);
nand U41578 (N_41578,N_36289,N_38924);
xnor U41579 (N_41579,N_36280,N_34881);
nor U41580 (N_41580,N_34343,N_30886);
nand U41581 (N_41581,N_36886,N_32642);
nand U41582 (N_41582,N_37405,N_32516);
and U41583 (N_41583,N_32600,N_32111);
and U41584 (N_41584,N_30293,N_32937);
nor U41585 (N_41585,N_39307,N_32775);
nand U41586 (N_41586,N_35800,N_31133);
or U41587 (N_41587,N_32751,N_31999);
and U41588 (N_41588,N_35758,N_39291);
nand U41589 (N_41589,N_31733,N_30419);
xnor U41590 (N_41590,N_32568,N_37560);
or U41591 (N_41591,N_30017,N_39260);
or U41592 (N_41592,N_36439,N_38248);
or U41593 (N_41593,N_32282,N_39549);
or U41594 (N_41594,N_39258,N_32546);
nand U41595 (N_41595,N_30548,N_32930);
nor U41596 (N_41596,N_37047,N_32793);
nand U41597 (N_41597,N_33548,N_36788);
or U41598 (N_41598,N_31795,N_35973);
and U41599 (N_41599,N_39539,N_34222);
nand U41600 (N_41600,N_35823,N_33264);
or U41601 (N_41601,N_34587,N_35465);
nor U41602 (N_41602,N_38727,N_33405);
and U41603 (N_41603,N_38681,N_37622);
nand U41604 (N_41604,N_30923,N_33380);
nor U41605 (N_41605,N_35317,N_38270);
and U41606 (N_41606,N_36245,N_39505);
and U41607 (N_41607,N_32644,N_34054);
nand U41608 (N_41608,N_35688,N_36135);
nand U41609 (N_41609,N_38359,N_36576);
nor U41610 (N_41610,N_30312,N_32404);
nor U41611 (N_41611,N_35974,N_39822);
nor U41612 (N_41612,N_34751,N_37819);
nor U41613 (N_41613,N_35038,N_38676);
nand U41614 (N_41614,N_38427,N_32485);
nand U41615 (N_41615,N_30771,N_37230);
nor U41616 (N_41616,N_32669,N_31239);
xor U41617 (N_41617,N_36805,N_30668);
nand U41618 (N_41618,N_33449,N_38734);
xnor U41619 (N_41619,N_38305,N_39458);
nor U41620 (N_41620,N_32973,N_32240);
and U41621 (N_41621,N_39559,N_39555);
nand U41622 (N_41622,N_34447,N_39032);
and U41623 (N_41623,N_31578,N_34525);
nand U41624 (N_41624,N_32504,N_35006);
and U41625 (N_41625,N_37698,N_36825);
nand U41626 (N_41626,N_36554,N_32243);
and U41627 (N_41627,N_31004,N_34693);
and U41628 (N_41628,N_30467,N_36079);
nor U41629 (N_41629,N_32683,N_32759);
nand U41630 (N_41630,N_34635,N_31610);
or U41631 (N_41631,N_39186,N_32422);
nand U41632 (N_41632,N_37716,N_37084);
nand U41633 (N_41633,N_37929,N_38162);
and U41634 (N_41634,N_32778,N_33443);
or U41635 (N_41635,N_31522,N_39644);
nand U41636 (N_41636,N_37388,N_32844);
and U41637 (N_41637,N_38592,N_35884);
nand U41638 (N_41638,N_38620,N_31296);
nor U41639 (N_41639,N_35225,N_30042);
nor U41640 (N_41640,N_39366,N_31484);
nor U41641 (N_41641,N_34723,N_34928);
and U41642 (N_41642,N_35965,N_39921);
nor U41643 (N_41643,N_32548,N_31464);
nor U41644 (N_41644,N_34155,N_35764);
nand U41645 (N_41645,N_33976,N_33731);
and U41646 (N_41646,N_31703,N_39168);
nand U41647 (N_41647,N_30816,N_38810);
and U41648 (N_41648,N_34164,N_34326);
nor U41649 (N_41649,N_39673,N_39104);
or U41650 (N_41650,N_35185,N_34319);
and U41651 (N_41651,N_33250,N_31974);
nand U41652 (N_41652,N_31027,N_39517);
nand U41653 (N_41653,N_34070,N_35315);
nand U41654 (N_41654,N_35998,N_39868);
or U41655 (N_41655,N_39900,N_31252);
and U41656 (N_41656,N_36632,N_38773);
nor U41657 (N_41657,N_35967,N_30315);
and U41658 (N_41658,N_38397,N_30707);
nor U41659 (N_41659,N_36104,N_36708);
xor U41660 (N_41660,N_37234,N_37457);
nor U41661 (N_41661,N_36871,N_35428);
or U41662 (N_41662,N_35715,N_37252);
and U41663 (N_41663,N_31597,N_34781);
or U41664 (N_41664,N_39943,N_33485);
nor U41665 (N_41665,N_39028,N_35546);
xnor U41666 (N_41666,N_36367,N_33172);
nand U41667 (N_41667,N_33227,N_30812);
and U41668 (N_41668,N_32967,N_30820);
and U41669 (N_41669,N_32107,N_39591);
or U41670 (N_41670,N_36870,N_32190);
and U41671 (N_41671,N_38936,N_34459);
or U41672 (N_41672,N_39135,N_35706);
nor U41673 (N_41673,N_39672,N_30031);
nand U41674 (N_41674,N_39924,N_33784);
nand U41675 (N_41675,N_36311,N_37915);
nand U41676 (N_41676,N_34829,N_39460);
or U41677 (N_41677,N_39213,N_31022);
nand U41678 (N_41678,N_37926,N_38015);
nand U41679 (N_41679,N_31761,N_36019);
or U41680 (N_41680,N_36595,N_33067);
xor U41681 (N_41681,N_31605,N_39421);
or U41682 (N_41682,N_31227,N_32877);
and U41683 (N_41683,N_32547,N_34948);
nor U41684 (N_41684,N_35259,N_33123);
xor U41685 (N_41685,N_34489,N_34280);
and U41686 (N_41686,N_34814,N_37899);
or U41687 (N_41687,N_30842,N_31082);
nor U41688 (N_41688,N_38878,N_34078);
or U41689 (N_41689,N_30012,N_37872);
nor U41690 (N_41690,N_30785,N_34274);
or U41691 (N_41691,N_37967,N_36344);
nand U41692 (N_41692,N_33597,N_34294);
or U41693 (N_41693,N_38052,N_31208);
and U41694 (N_41694,N_35607,N_37011);
or U41695 (N_41695,N_37486,N_34314);
or U41696 (N_41696,N_32591,N_37064);
or U41697 (N_41697,N_32119,N_32860);
or U41698 (N_41698,N_31668,N_32063);
xnor U41699 (N_41699,N_33410,N_33259);
nand U41700 (N_41700,N_36989,N_35309);
xor U41701 (N_41701,N_34875,N_34400);
nor U41702 (N_41702,N_36545,N_30738);
xnor U41703 (N_41703,N_32887,N_32985);
nand U41704 (N_41704,N_33573,N_30875);
and U41705 (N_41705,N_30615,N_32949);
or U41706 (N_41706,N_37272,N_32286);
nor U41707 (N_41707,N_34532,N_39978);
and U41708 (N_41708,N_35032,N_33526);
nor U41709 (N_41709,N_37835,N_37768);
and U41710 (N_41710,N_36994,N_39620);
and U41711 (N_41711,N_31432,N_35912);
or U41712 (N_41712,N_34593,N_35391);
nor U41713 (N_41713,N_34000,N_33385);
xnor U41714 (N_41714,N_35834,N_33095);
nor U41715 (N_41715,N_38609,N_33203);
or U41716 (N_41716,N_39507,N_37349);
and U41717 (N_41717,N_37209,N_37995);
and U41718 (N_41718,N_34549,N_35470);
or U41719 (N_41719,N_38472,N_30322);
nand U41720 (N_41720,N_34385,N_31100);
nor U41721 (N_41721,N_32924,N_34763);
and U41722 (N_41722,N_34217,N_34625);
and U41723 (N_41723,N_35398,N_35376);
nor U41724 (N_41724,N_34338,N_36898);
nand U41725 (N_41725,N_30394,N_35484);
and U41726 (N_41726,N_30458,N_38795);
and U41727 (N_41727,N_37219,N_30191);
or U41728 (N_41728,N_36005,N_30146);
nor U41729 (N_41729,N_30058,N_34431);
or U41730 (N_41730,N_37778,N_39482);
or U41731 (N_41731,N_37137,N_31980);
nand U41732 (N_41732,N_34225,N_37734);
or U41733 (N_41733,N_38086,N_36622);
nand U41734 (N_41734,N_37387,N_32394);
and U41735 (N_41735,N_31244,N_33356);
and U41736 (N_41736,N_39190,N_36234);
nand U41737 (N_41737,N_30881,N_30384);
nand U41738 (N_41738,N_38480,N_33725);
nor U41739 (N_41739,N_32797,N_35624);
nand U41740 (N_41740,N_34424,N_37492);
nand U41741 (N_41741,N_36366,N_37800);
or U41742 (N_41742,N_39916,N_38410);
nor U41743 (N_41743,N_34031,N_36761);
xnor U41744 (N_41744,N_35005,N_38870);
xor U41745 (N_41745,N_33131,N_32738);
nor U41746 (N_41746,N_30429,N_36905);
nor U41747 (N_41747,N_36775,N_30440);
and U41748 (N_41748,N_38919,N_33145);
and U41749 (N_41749,N_37634,N_30733);
nand U41750 (N_41750,N_33153,N_37559);
or U41751 (N_41751,N_37534,N_31660);
nand U41752 (N_41752,N_30527,N_37918);
or U41753 (N_41753,N_30499,N_32235);
or U41754 (N_41754,N_38136,N_32149);
xor U41755 (N_41755,N_33716,N_33730);
nand U41756 (N_41756,N_39000,N_37120);
or U41757 (N_41757,N_33881,N_34476);
or U41758 (N_41758,N_33950,N_35874);
and U41759 (N_41759,N_33787,N_32206);
nand U41760 (N_41760,N_35401,N_38887);
nand U41761 (N_41761,N_38358,N_38421);
nor U41762 (N_41762,N_32836,N_30024);
nor U41763 (N_41763,N_32128,N_36250);
xnor U41764 (N_41764,N_31230,N_36817);
and U41765 (N_41765,N_32820,N_34490);
nand U41766 (N_41766,N_36888,N_32024);
nor U41767 (N_41767,N_36921,N_34851);
xnor U41768 (N_41768,N_33417,N_38415);
xnor U41769 (N_41769,N_34223,N_34333);
or U41770 (N_41770,N_37620,N_32726);
or U41771 (N_41771,N_35053,N_39263);
nor U41772 (N_41772,N_31411,N_37725);
nand U41773 (N_41773,N_34602,N_38628);
nor U41774 (N_41774,N_33371,N_37506);
or U41775 (N_41775,N_37482,N_39791);
and U41776 (N_41776,N_32398,N_37354);
nor U41777 (N_41777,N_34117,N_31176);
nor U41778 (N_41778,N_39552,N_30760);
or U41779 (N_41779,N_35432,N_32552);
nand U41780 (N_41780,N_37304,N_35747);
or U41781 (N_41781,N_34702,N_34345);
and U41782 (N_41782,N_39886,N_37328);
or U41783 (N_41783,N_33942,N_34244);
and U41784 (N_41784,N_31550,N_35306);
or U41785 (N_41785,N_33326,N_34946);
nand U41786 (N_41786,N_37514,N_31091);
xnor U41787 (N_41787,N_31055,N_37928);
or U41788 (N_41788,N_35492,N_39256);
or U41789 (N_41789,N_34035,N_35360);
nor U41790 (N_41790,N_38222,N_36832);
nor U41791 (N_41791,N_33030,N_37399);
or U41792 (N_41792,N_32001,N_33237);
or U41793 (N_41793,N_34043,N_31062);
or U41794 (N_41794,N_38935,N_35403);
nand U41795 (N_41795,N_39216,N_33876);
or U41796 (N_41796,N_33022,N_33114);
xnor U41797 (N_41797,N_36820,N_35990);
xnor U41798 (N_41798,N_36772,N_36740);
xnor U41799 (N_41799,N_32196,N_38693);
nor U41800 (N_41800,N_32266,N_32042);
or U41801 (N_41801,N_32133,N_37678);
nor U41802 (N_41802,N_32960,N_39142);
nand U41803 (N_41803,N_38833,N_35481);
or U41804 (N_41804,N_30025,N_37911);
and U41805 (N_41805,N_30335,N_30824);
nand U41806 (N_41806,N_36836,N_30545);
and U41807 (N_41807,N_36728,N_31195);
or U41808 (N_41808,N_36525,N_31653);
xor U41809 (N_41809,N_32896,N_31352);
and U41810 (N_41810,N_36362,N_35210);
nor U41811 (N_41811,N_33907,N_37496);
nor U41812 (N_41812,N_35452,N_38587);
and U41813 (N_41813,N_38495,N_30483);
nor U41814 (N_41814,N_33639,N_31682);
nand U41815 (N_41815,N_33660,N_34529);
nand U41816 (N_41816,N_32583,N_35729);
nand U41817 (N_41817,N_33398,N_30562);
or U41818 (N_41818,N_38781,N_37522);
or U41819 (N_41819,N_32407,N_35610);
nand U41820 (N_41820,N_35373,N_32172);
or U41821 (N_41821,N_35310,N_33470);
nor U41822 (N_41822,N_35194,N_35575);
nand U41823 (N_41823,N_33219,N_32080);
nor U41824 (N_41824,N_33771,N_30890);
and U41825 (N_41825,N_39712,N_38882);
or U41826 (N_41826,N_35714,N_33983);
or U41827 (N_41827,N_34900,N_34050);
nor U41828 (N_41828,N_37129,N_35390);
nor U41829 (N_41829,N_39022,N_31114);
nor U41830 (N_41830,N_30248,N_34337);
and U41831 (N_41831,N_35125,N_33758);
and U41832 (N_41832,N_30364,N_35216);
nor U41833 (N_41833,N_37718,N_31775);
nand U41834 (N_41834,N_37237,N_31913);
or U41835 (N_41835,N_35968,N_35506);
nor U41836 (N_41836,N_31879,N_38558);
nand U41837 (N_41837,N_39177,N_30092);
and U41838 (N_41838,N_33724,N_30032);
and U41839 (N_41839,N_31744,N_33183);
and U41840 (N_41840,N_30856,N_37251);
xor U41841 (N_41841,N_34714,N_31295);
nand U41842 (N_41842,N_38309,N_37630);
nand U41843 (N_41843,N_37499,N_37623);
nor U41844 (N_41844,N_34500,N_34270);
nor U41845 (N_41845,N_34588,N_33455);
nand U41846 (N_41846,N_34820,N_33090);
or U41847 (N_41847,N_39982,N_33806);
xnor U41848 (N_41848,N_31752,N_36572);
nor U41849 (N_41849,N_30697,N_35835);
or U41850 (N_41850,N_36907,N_33682);
nor U41851 (N_41851,N_33872,N_33099);
nor U41852 (N_41852,N_33080,N_31388);
nand U41853 (N_41853,N_30053,N_31798);
nand U41854 (N_41854,N_30925,N_30905);
or U41855 (N_41855,N_38643,N_36663);
and U41856 (N_41856,N_37987,N_30574);
and U41857 (N_41857,N_36202,N_39405);
and U41858 (N_41858,N_35173,N_38101);
xnor U41859 (N_41859,N_38372,N_30054);
nand U41860 (N_41860,N_36723,N_30311);
or U41861 (N_41861,N_30532,N_38871);
and U41862 (N_41862,N_39372,N_33018);
nor U41863 (N_41863,N_38150,N_31096);
or U41864 (N_41864,N_38707,N_32940);
nand U41865 (N_41865,N_39915,N_34834);
nor U41866 (N_41866,N_33271,N_35941);
nor U41867 (N_41867,N_30509,N_34397);
nand U41868 (N_41868,N_38782,N_39575);
xnor U41869 (N_41869,N_31786,N_34840);
nand U41870 (N_41870,N_38204,N_34289);
nand U41871 (N_41871,N_31383,N_30919);
nand U41872 (N_41872,N_35299,N_31505);
and U41873 (N_41873,N_31362,N_39125);
and U41874 (N_41874,N_36452,N_35643);
or U41875 (N_41875,N_35399,N_30700);
xor U41876 (N_41876,N_33162,N_32397);
and U41877 (N_41877,N_31113,N_39856);
nand U41878 (N_41878,N_30998,N_34511);
nand U41879 (N_41879,N_33052,N_36091);
nor U41880 (N_41880,N_30181,N_37658);
xnor U41881 (N_41881,N_30235,N_33825);
nand U41882 (N_41882,N_39490,N_30205);
nor U41883 (N_41883,N_35448,N_38187);
and U41884 (N_41884,N_33838,N_30307);
or U41885 (N_41885,N_36710,N_32517);
or U41886 (N_41886,N_34719,N_35215);
and U41887 (N_41887,N_35135,N_39394);
xor U41888 (N_41888,N_35730,N_37316);
and U41889 (N_41889,N_39596,N_33584);
or U41890 (N_41890,N_38554,N_34694);
nor U41891 (N_41891,N_36119,N_31802);
or U41892 (N_41892,N_37218,N_33801);
nand U41893 (N_41893,N_37111,N_37617);
xor U41894 (N_41894,N_31910,N_36588);
nand U41895 (N_41895,N_30101,N_39249);
and U41896 (N_41896,N_31326,N_33378);
xnor U41897 (N_41897,N_37573,N_38994);
nor U41898 (N_41898,N_34502,N_36354);
or U41899 (N_41899,N_37063,N_37526);
xnor U41900 (N_41900,N_32802,N_36040);
nand U41901 (N_41901,N_32757,N_35677);
nand U41902 (N_41902,N_30340,N_31978);
xor U41903 (N_41903,N_38154,N_32338);
or U41904 (N_41904,N_30763,N_33346);
or U41905 (N_41905,N_39489,N_30491);
xnor U41906 (N_41906,N_34998,N_31925);
nand U41907 (N_41907,N_34013,N_30444);
nor U41908 (N_41908,N_35438,N_30654);
or U41909 (N_41909,N_32467,N_36243);
nor U41910 (N_41910,N_31900,N_30687);
and U41911 (N_41911,N_30992,N_36341);
xnor U41912 (N_41912,N_30061,N_39646);
xnor U41913 (N_41913,N_33116,N_30662);
nand U41914 (N_41914,N_38118,N_30098);
and U41915 (N_41915,N_38471,N_34121);
or U41916 (N_41916,N_34191,N_31168);
and U41917 (N_41917,N_32364,N_38055);
xor U41918 (N_41918,N_39756,N_32330);
or U41919 (N_41919,N_34437,N_35668);
nand U41920 (N_41920,N_36238,N_32796);
nor U41921 (N_41921,N_32484,N_39326);
or U41922 (N_41922,N_30655,N_37240);
nand U41923 (N_41923,N_36641,N_38132);
or U41924 (N_41924,N_32524,N_30557);
nand U41925 (N_41925,N_34259,N_35831);
nand U41926 (N_41926,N_36355,N_39866);
xor U41927 (N_41927,N_39358,N_36423);
nor U41928 (N_41928,N_37954,N_34470);
nor U41929 (N_41929,N_36393,N_37662);
nand U41930 (N_41930,N_35027,N_36401);
nor U41931 (N_41931,N_33568,N_37939);
or U41932 (N_41932,N_34140,N_37034);
or U41933 (N_41933,N_37686,N_36932);
and U41934 (N_41934,N_36657,N_31763);
xor U41935 (N_41935,N_37945,N_37576);
nor U41936 (N_41936,N_36227,N_37973);
and U41937 (N_41937,N_38682,N_34449);
xor U41938 (N_41938,N_39318,N_36659);
xnor U41939 (N_41939,N_34561,N_33049);
or U41940 (N_41940,N_38271,N_37450);
nor U41941 (N_41941,N_35384,N_30380);
nand U41942 (N_41942,N_38690,N_34340);
nor U41943 (N_41943,N_36956,N_32908);
or U41944 (N_41944,N_31551,N_39297);
nand U41945 (N_41945,N_31349,N_35165);
nand U41946 (N_41946,N_30011,N_31438);
and U41947 (N_41947,N_33638,N_34403);
nor U41948 (N_41948,N_30550,N_37563);
nand U41949 (N_41949,N_37783,N_38202);
or U41950 (N_41950,N_31343,N_39201);
nand U41951 (N_41951,N_35981,N_31556);
xnor U41952 (N_41952,N_36381,N_35440);
and U41953 (N_41953,N_38084,N_33244);
and U41954 (N_41954,N_35670,N_39628);
nand U41955 (N_41955,N_38941,N_39965);
nor U41956 (N_41956,N_37816,N_33472);
or U41957 (N_41957,N_37186,N_31698);
and U41958 (N_41958,N_31028,N_31950);
nand U41959 (N_41959,N_35964,N_33496);
nor U41960 (N_41960,N_30021,N_38595);
nand U41961 (N_41961,N_31177,N_32640);
and U41962 (N_41962,N_31463,N_34772);
xor U41963 (N_41963,N_37909,N_37269);
and U41964 (N_41964,N_37428,N_36242);
or U41965 (N_41965,N_39588,N_36193);
and U41966 (N_41966,N_37455,N_34171);
and U41967 (N_41967,N_36791,N_39993);
nand U41968 (N_41968,N_32739,N_34227);
or U41969 (N_41969,N_38050,N_35312);
or U41970 (N_41970,N_32576,N_35858);
nand U41971 (N_41971,N_39158,N_39955);
nor U41972 (N_41972,N_39080,N_37773);
and U41973 (N_41973,N_39973,N_33008);
or U41974 (N_41974,N_32336,N_37883);
and U41975 (N_41975,N_33016,N_34336);
and U41976 (N_41976,N_32765,N_30661);
and U41977 (N_41977,N_34484,N_37152);
xor U41978 (N_41978,N_37907,N_38596);
or U41979 (N_41979,N_31846,N_30624);
nand U41980 (N_41980,N_32378,N_32606);
nand U41981 (N_41981,N_35991,N_33540);
and U41982 (N_41982,N_36639,N_30125);
and U41983 (N_41983,N_39025,N_36376);
nand U41984 (N_41984,N_33221,N_34761);
nand U41985 (N_41985,N_32493,N_30178);
or U41986 (N_41986,N_32083,N_38717);
xnor U41987 (N_41987,N_35787,N_32723);
and U41988 (N_41988,N_32505,N_34386);
nand U41989 (N_41989,N_35857,N_31198);
or U41990 (N_41990,N_36431,N_34740);
nor U41991 (N_41991,N_34911,N_36970);
and U41992 (N_41992,N_38754,N_34095);
nor U41993 (N_41993,N_38256,N_33650);
nor U41994 (N_41994,N_36954,N_32332);
and U41995 (N_41995,N_32850,N_39232);
nand U41996 (N_41996,N_30194,N_36207);
nand U41997 (N_41997,N_36743,N_30645);
and U41998 (N_41998,N_33209,N_39128);
and U41999 (N_41999,N_31320,N_36621);
and U42000 (N_42000,N_30625,N_35500);
nand U42001 (N_42001,N_35445,N_32482);
xnor U42002 (N_42002,N_34506,N_39379);
and U42003 (N_42003,N_34815,N_37182);
or U42004 (N_42004,N_37389,N_35249);
xor U42005 (N_42005,N_36226,N_32988);
or U42006 (N_42006,N_39869,N_30947);
or U42007 (N_42007,N_38416,N_32574);
nor U42008 (N_42008,N_36107,N_38398);
xnor U42009 (N_42009,N_35878,N_34708);
and U42010 (N_42010,N_39968,N_39884);
nand U42011 (N_42011,N_32259,N_36123);
xor U42012 (N_42012,N_31217,N_30466);
nor U42013 (N_42013,N_35580,N_31658);
and U42014 (N_42014,N_35118,N_38662);
nor U42015 (N_42015,N_37498,N_35518);
nor U42016 (N_42016,N_30775,N_39782);
nor U42017 (N_42017,N_33687,N_38138);
nand U42018 (N_42018,N_39820,N_35188);
and U42019 (N_42019,N_34951,N_31683);
and U42020 (N_42020,N_39667,N_33372);
and U42021 (N_42021,N_30292,N_34893);
or U42022 (N_42022,N_37013,N_37791);
nor U42023 (N_42023,N_33541,N_37955);
or U42024 (N_42024,N_35871,N_30600);
xor U42025 (N_42025,N_36631,N_39889);
nand U42026 (N_42026,N_39763,N_37565);
xor U42027 (N_42027,N_34325,N_36804);
or U42028 (N_42028,N_35327,N_39925);
nor U42029 (N_42029,N_30245,N_30845);
and U42030 (N_42030,N_35287,N_36880);
xnor U42031 (N_42031,N_36443,N_33898);
and U42032 (N_42032,N_33308,N_32545);
nor U42033 (N_42033,N_39222,N_30629);
xnor U42034 (N_42034,N_37923,N_32987);
or U42035 (N_42035,N_35675,N_39314);
or U42036 (N_42036,N_35359,N_39292);
nor U42037 (N_42037,N_34886,N_36922);
xor U42038 (N_42038,N_35477,N_39157);
nor U42039 (N_42039,N_33081,N_37212);
and U42040 (N_42040,N_32220,N_30056);
or U42041 (N_42041,N_30273,N_31421);
nand U42042 (N_42042,N_34406,N_31111);
nor U42043 (N_42043,N_37372,N_31852);
nor U42044 (N_42044,N_37362,N_32798);
nand U42045 (N_42045,N_30430,N_38192);
nor U42046 (N_42046,N_33707,N_35719);
xor U42047 (N_42047,N_32792,N_37067);
nand U42048 (N_42048,N_32575,N_35836);
nor U42049 (N_42049,N_38860,N_36020);
nand U42050 (N_42050,N_35552,N_32409);
nand U42051 (N_42051,N_36028,N_33766);
nand U42052 (N_42052,N_35017,N_34425);
nor U42053 (N_42053,N_31428,N_37126);
nand U42054 (N_42054,N_32813,N_32951);
nor U42055 (N_42055,N_30678,N_30442);
nand U42056 (N_42056,N_33805,N_30078);
nor U42057 (N_42057,N_33695,N_36587);
or U42058 (N_42058,N_36335,N_38669);
nor U42059 (N_42059,N_33552,N_33007);
nand U42060 (N_42060,N_38674,N_34844);
nand U42061 (N_42061,N_32094,N_31032);
nor U42062 (N_42062,N_31712,N_30167);
nor U42063 (N_42063,N_39834,N_39894);
and U42064 (N_42064,N_34162,N_35378);
or U42065 (N_42065,N_33668,N_37495);
or U42066 (N_42066,N_30560,N_30653);
or U42067 (N_42067,N_39593,N_39148);
nor U42068 (N_42068,N_35459,N_39139);
and U42069 (N_42069,N_37184,N_35841);
nor U42070 (N_42070,N_38440,N_31161);
nand U42071 (N_42071,N_36544,N_39642);
nand U42072 (N_42072,N_30747,N_32406);
nor U42073 (N_42073,N_37857,N_36465);
and U42074 (N_42074,N_39592,N_36458);
or U42075 (N_42075,N_31293,N_38964);
nor U42076 (N_42076,N_39536,N_32345);
xor U42077 (N_42077,N_31495,N_35342);
nor U42078 (N_42078,N_39920,N_31389);
or U42079 (N_42079,N_33079,N_31455);
nand U42080 (N_42080,N_38199,N_36409);
and U42081 (N_42081,N_37951,N_32897);
nand U42082 (N_42082,N_37994,N_38335);
nor U42083 (N_42083,N_39976,N_33055);
nor U42084 (N_42084,N_38523,N_36025);
and U42085 (N_42085,N_37002,N_35801);
and U42086 (N_42086,N_37441,N_37468);
and U42087 (N_42087,N_38636,N_34271);
or U42088 (N_42088,N_33826,N_38320);
xnor U42089 (N_42089,N_36983,N_38317);
nor U42090 (N_42090,N_35844,N_39876);
or U42091 (N_42091,N_39520,N_30602);
xnor U42092 (N_42092,N_36429,N_36027);
nand U42093 (N_42093,N_37843,N_34513);
nand U42094 (N_42094,N_30211,N_38904);
nand U42095 (N_42095,N_33490,N_37487);
xnor U42096 (N_42096,N_34445,N_31394);
nand U42097 (N_42097,N_34387,N_36862);
or U42098 (N_42098,N_39816,N_36926);
and U42099 (N_42099,N_30782,N_37382);
nor U42100 (N_42100,N_31278,N_38470);
or U42101 (N_42101,N_32862,N_32290);
and U42102 (N_42102,N_35449,N_31656);
and U42103 (N_42103,N_37832,N_35655);
and U42104 (N_42104,N_30344,N_34673);
or U42105 (N_42105,N_35354,N_36937);
or U42106 (N_42106,N_30983,N_39603);
nor U42107 (N_42107,N_39706,N_33585);
nor U42108 (N_42108,N_32755,N_38282);
and U42109 (N_42109,N_36467,N_33112);
and U42110 (N_42110,N_37326,N_37548);
nand U42111 (N_42111,N_33241,N_34002);
nor U42112 (N_42112,N_34376,N_32074);
nor U42113 (N_42113,N_32238,N_33249);
nand U42114 (N_42114,N_36995,N_38759);
nor U42115 (N_42115,N_31267,N_37575);
and U42116 (N_42116,N_30638,N_35704);
or U42117 (N_42117,N_36550,N_39775);
and U42118 (N_42118,N_34768,N_36944);
or U42119 (N_42119,N_33849,N_35292);
nand U42120 (N_42120,N_38604,N_32210);
nor U42121 (N_42121,N_35983,N_37233);
nand U42122 (N_42122,N_36045,N_37447);
or U42123 (N_42123,N_38091,N_37291);
nor U42124 (N_42124,N_35431,N_37402);
or U42125 (N_42125,N_30597,N_36275);
nor U42126 (N_42126,N_31915,N_31190);
nand U42127 (N_42127,N_37037,N_32098);
nor U42128 (N_42128,N_36363,N_30151);
nor U42129 (N_42129,N_30965,N_34762);
or U42130 (N_42130,N_39146,N_33593);
and U42131 (N_42131,N_37458,N_31071);
nor U42132 (N_42132,N_36704,N_38665);
nor U42133 (N_42133,N_30144,N_33434);
nor U42134 (N_42134,N_34699,N_37187);
or U42135 (N_42135,N_36244,N_34733);
or U42136 (N_42136,N_38943,N_31305);
nand U42137 (N_42137,N_37164,N_32408);
or U42138 (N_42138,N_39503,N_39274);
xor U42139 (N_42139,N_31218,N_32277);
nor U42140 (N_42140,N_33109,N_36690);
and U42141 (N_42141,N_38337,N_37821);
and U42142 (N_42142,N_31713,N_37847);
nor U42143 (N_42143,N_34208,N_31932);
and U42144 (N_42144,N_31246,N_35572);
and U42145 (N_42145,N_37481,N_32776);
or U42146 (N_42146,N_30040,N_38340);
nor U42147 (N_42147,N_36843,N_31884);
or U42148 (N_42148,N_39479,N_37841);
nand U42149 (N_42149,N_39070,N_36719);
nand U42150 (N_42150,N_30999,N_38645);
nand U42151 (N_42151,N_31370,N_39977);
or U42152 (N_42152,N_37423,N_39670);
nand U42153 (N_42153,N_37598,N_31926);
and U42154 (N_42154,N_30503,N_32350);
or U42155 (N_42155,N_32450,N_30692);
or U42156 (N_42156,N_39188,N_34953);
or U42157 (N_42157,N_38808,N_37697);
and U42158 (N_42158,N_31993,N_36435);
and U42159 (N_42159,N_38783,N_30498);
or U42160 (N_42160,N_32480,N_34830);
nand U42161 (N_42161,N_37749,N_31232);
nand U42162 (N_42162,N_35762,N_32040);
nor U42163 (N_42163,N_39369,N_33137);
and U42164 (N_42164,N_35700,N_35396);
nor U42165 (N_42165,N_33632,N_31066);
nand U42166 (N_42166,N_33963,N_37156);
nand U42167 (N_42167,N_32309,N_33361);
and U42168 (N_42168,N_33923,N_36977);
nand U42169 (N_42169,N_31490,N_38895);
or U42170 (N_42170,N_32316,N_32864);
or U42171 (N_42171,N_30698,N_39580);
or U42172 (N_42172,N_34934,N_39815);
nor U42173 (N_42173,N_36623,N_30204);
nand U42174 (N_42174,N_32936,N_37246);
and U42175 (N_42175,N_33612,N_37345);
or U42176 (N_42176,N_39679,N_39630);
xor U42177 (N_42177,N_33995,N_39601);
nand U42178 (N_42178,N_32167,N_35796);
nor U42179 (N_42179,N_35131,N_35768);
nand U42180 (N_42180,N_33207,N_39747);
xor U42181 (N_42181,N_30270,N_33543);
and U42182 (N_42182,N_30046,N_39839);
xnor U42183 (N_42183,N_39205,N_35862);
or U42184 (N_42184,N_39465,N_30885);
nor U42185 (N_42185,N_38753,N_32085);
and U42186 (N_42186,N_39508,N_33036);
and U42187 (N_42187,N_39462,N_39707);
or U42188 (N_42188,N_36201,N_32026);
xnor U42189 (N_42189,N_37323,N_32858);
and U42190 (N_42190,N_34052,N_31398);
xnor U42191 (N_42191,N_33223,N_38948);
and U42192 (N_42192,N_31825,N_33222);
xnor U42193 (N_42193,N_33446,N_31498);
nor U42194 (N_42194,N_38319,N_35562);
or U42195 (N_42195,N_30620,N_36010);
nor U42196 (N_42196,N_35711,N_39764);
nand U42197 (N_42197,N_32365,N_30243);
nor U42198 (N_42198,N_37597,N_33558);
and U42199 (N_42199,N_39346,N_37194);
and U42200 (N_42200,N_33594,N_32722);
or U42201 (N_42201,N_39030,N_37413);
nor U42202 (N_42202,N_34664,N_39882);
xor U42203 (N_42203,N_35583,N_37753);
and U42204 (N_42204,N_39273,N_33862);
and U42205 (N_42205,N_35482,N_32475);
nand U42206 (N_42206,N_37094,N_34568);
nand U42207 (N_42207,N_37670,N_37366);
or U42208 (N_42208,N_30139,N_33761);
or U42209 (N_42209,N_32051,N_36264);
nand U42210 (N_42210,N_39981,N_30934);
nand U42211 (N_42211,N_30299,N_38865);
and U42212 (N_42212,N_36407,N_30183);
or U42213 (N_42213,N_36819,N_35453);
nand U42214 (N_42214,N_31209,N_36054);
nand U42215 (N_42215,N_35018,N_32724);
or U42216 (N_42216,N_30606,N_34213);
and U42217 (N_42217,N_34488,N_32818);
and U42218 (N_42218,N_39086,N_34408);
and U42219 (N_42219,N_34967,N_37717);
and U42220 (N_42220,N_37901,N_33060);
or U42221 (N_42221,N_34628,N_32717);
nand U42222 (N_42222,N_31826,N_31137);
nand U42223 (N_42223,N_36333,N_37779);
or U42224 (N_42224,N_31327,N_35374);
and U42225 (N_42225,N_39183,N_31148);
and U42226 (N_42226,N_33595,N_35731);
or U42227 (N_42227,N_37400,N_36593);
xor U42228 (N_42228,N_31174,N_38287);
or U42229 (N_42229,N_36476,N_34982);
or U42230 (N_42230,N_34253,N_37668);
nand U42231 (N_42231,N_35579,N_39602);
nor U42232 (N_42232,N_34559,N_38991);
and U42233 (N_42233,N_32807,N_30037);
and U42234 (N_42234,N_30237,N_35480);
nor U42235 (N_42235,N_31965,N_37646);
or U42236 (N_42236,N_39495,N_31325);
nor U42237 (N_42237,N_36844,N_31203);
nor U42238 (N_42238,N_31982,N_36826);
xor U42239 (N_42239,N_32339,N_38532);
xnor U42240 (N_42240,N_33224,N_39658);
or U42241 (N_42241,N_36564,N_30175);
nor U42242 (N_42242,N_30693,N_35767);
nand U42243 (N_42243,N_38322,N_32258);
or U42244 (N_42244,N_36421,N_34407);
xnor U42245 (N_42245,N_33532,N_37898);
and U42246 (N_42246,N_36392,N_39585);
or U42247 (N_42247,N_36724,N_31536);
or U42248 (N_42248,N_34747,N_33029);
and U42249 (N_42249,N_30059,N_37140);
xor U42250 (N_42250,N_35155,N_31818);
and U42251 (N_42251,N_38343,N_34755);
nand U42252 (N_42252,N_31957,N_32746);
or U42253 (N_42253,N_35171,N_39875);
nand U42254 (N_42254,N_37132,N_34899);
nand U42255 (N_42255,N_34684,N_35560);
nor U42256 (N_42256,N_33430,N_36146);
nor U42257 (N_42257,N_31314,N_31517);
nor U42258 (N_42258,N_33360,N_39694);
and U42259 (N_42259,N_35352,N_33307);
nor U42260 (N_42260,N_33569,N_32698);
nand U42261 (N_42261,N_30207,N_32567);
nor U42262 (N_42262,N_30096,N_36179);
and U42263 (N_42263,N_38844,N_30710);
or U42264 (N_42264,N_39927,N_33714);
xor U42265 (N_42265,N_37780,N_34205);
nor U42266 (N_42266,N_32120,N_30589);
xor U42267 (N_42267,N_36438,N_30821);
xnor U42268 (N_42268,N_30044,N_33885);
nor U42269 (N_42269,N_39966,N_31476);
nand U42270 (N_42270,N_34538,N_39103);
or U42271 (N_42271,N_31584,N_33752);
and U42272 (N_42272,N_32883,N_34771);
nor U42273 (N_42273,N_34365,N_31901);
nor U42274 (N_42274,N_37201,N_30378);
and U42275 (N_42275,N_30834,N_35078);
or U42276 (N_42276,N_36348,N_35364);
nor U42277 (N_42277,N_38563,N_34922);
and U42278 (N_42278,N_38832,N_35182);
or U42279 (N_42279,N_38737,N_31165);
xor U42280 (N_42280,N_34041,N_36315);
nor U42281 (N_42281,N_35094,N_31212);
nor U42282 (N_42282,N_37431,N_34634);
xnor U42283 (N_42283,N_35751,N_37279);
and U42284 (N_42284,N_37941,N_37596);
or U42285 (N_42285,N_35958,N_34996);
or U42286 (N_42286,N_33523,N_34985);
nand U42287 (N_42287,N_31569,N_31672);
and U42288 (N_42288,N_38286,N_30052);
nand U42289 (N_42289,N_38082,N_38139);
and U42290 (N_42290,N_38059,N_35814);
nand U42291 (N_42291,N_37188,N_39068);
or U42292 (N_42292,N_39709,N_38275);
and U42293 (N_42293,N_35532,N_30962);
nor U42294 (N_42294,N_39009,N_32433);
or U42295 (N_42295,N_38780,N_30113);
nand U42296 (N_42296,N_32208,N_38921);
nand U42297 (N_42297,N_39375,N_33128);
or U42298 (N_42298,N_30713,N_32617);
and U42299 (N_42299,N_38005,N_30145);
nand U42300 (N_42300,N_38599,N_38291);
and U42301 (N_42301,N_39877,N_36626);
and U42302 (N_42302,N_38657,N_39304);
or U42303 (N_42303,N_37817,N_38980);
nand U42304 (N_42304,N_39099,N_35130);
and U42305 (N_42305,N_32308,N_38405);
or U42306 (N_42306,N_33032,N_37116);
nor U42307 (N_42307,N_35220,N_35860);
and U42308 (N_42308,N_33149,N_37446);
and U42309 (N_42309,N_31619,N_36948);
nor U42310 (N_42310,N_33859,N_31318);
xor U42311 (N_42311,N_36556,N_35418);
nor U42312 (N_42312,N_36188,N_31924);
and U42313 (N_42313,N_39309,N_36601);
nor U42314 (N_42314,N_39378,N_31403);
or U42315 (N_42315,N_33824,N_37731);
and U42316 (N_42316,N_35638,N_33348);
and U42317 (N_42317,N_30765,N_30412);
nand U42318 (N_42318,N_36444,N_39504);
or U42319 (N_42319,N_31330,N_33288);
nand U42320 (N_42320,N_31261,N_31119);
nor U42321 (N_42321,N_39618,N_39560);
or U42322 (N_42322,N_38239,N_36997);
or U42323 (N_42323,N_34823,N_31972);
and U42324 (N_42324,N_33837,N_37359);
nand U42325 (N_42325,N_32082,N_37231);
xnor U42326 (N_42326,N_38380,N_38993);
nor U42327 (N_42327,N_36829,N_38063);
or U42328 (N_42328,N_31991,N_38527);
and U42329 (N_42329,N_37879,N_39330);
nor U42330 (N_42330,N_38792,N_31316);
nand U42331 (N_42331,N_35648,N_38719);
nor U42332 (N_42332,N_38629,N_37606);
nand U42333 (N_42333,N_39833,N_32481);
and U42334 (N_42334,N_35765,N_38771);
or U42335 (N_42335,N_35585,N_30746);
or U42336 (N_42336,N_32358,N_38713);
nand U42337 (N_42337,N_31822,N_37637);
or U42338 (N_42338,N_38338,N_31127);
nor U42339 (N_42339,N_31358,N_32444);
nand U42340 (N_42340,N_34937,N_35186);
nand U42341 (N_42341,N_31891,N_32034);
and U42342 (N_42342,N_36968,N_30739);
and U42343 (N_42343,N_38911,N_34105);
and U42344 (N_42344,N_30950,N_36390);
and U42345 (N_42345,N_37602,N_30825);
and U42346 (N_42346,N_34046,N_30497);
and U42347 (N_42347,N_33000,N_38965);
nor U42348 (N_42348,N_38431,N_38448);
nand U42349 (N_42349,N_33797,N_30873);
nor U42350 (N_42350,N_39324,N_34989);
and U42351 (N_42351,N_37329,N_37166);
and U42352 (N_42352,N_32842,N_39899);
or U42353 (N_42353,N_31797,N_30034);
nand U42354 (N_42354,N_38567,N_36674);
nand U42355 (N_42355,N_34214,N_39259);
nor U42356 (N_42356,N_38092,N_33156);
and U42357 (N_42357,N_39243,N_36933);
and U42358 (N_42358,N_35172,N_33610);
or U42359 (N_42359,N_38588,N_35040);
and U42360 (N_42360,N_34141,N_39825);
or U42361 (N_42361,N_30939,N_31805);
and U42362 (N_42362,N_31361,N_33861);
nor U42363 (N_42363,N_36860,N_37226);
and U42364 (N_42364,N_35062,N_31270);
nor U42365 (N_42365,N_30828,N_39294);
xnor U42366 (N_42366,N_32625,N_39857);
xnor U42367 (N_42367,N_31564,N_39903);
nand U42368 (N_42368,N_37310,N_35568);
nor U42369 (N_42369,N_33867,N_36039);
xor U42370 (N_42370,N_39571,N_34260);
and U42371 (N_42371,N_37999,N_35140);
and U42372 (N_42372,N_33176,N_36035);
nand U42373 (N_42373,N_35294,N_34956);
nor U42374 (N_42374,N_36857,N_30495);
nand U42375 (N_42375,N_32803,N_39076);
nor U42376 (N_42376,N_34357,N_36258);
nand U42377 (N_42377,N_33489,N_39870);
or U42378 (N_42378,N_35944,N_38394);
nor U42379 (N_42379,N_38391,N_34522);
xor U42380 (N_42380,N_36120,N_33970);
and U42381 (N_42381,N_37728,N_31969);
nor U42382 (N_42382,N_32003,N_31039);
nor U42383 (N_42383,N_33400,N_34102);
nand U42384 (N_42384,N_32347,N_31702);
nor U42385 (N_42385,N_32510,N_35016);
nand U42386 (N_42386,N_32122,N_36534);
nor U42387 (N_42387,N_34430,N_36961);
nor U42388 (N_42388,N_36080,N_39352);
or U42389 (N_42389,N_36953,N_34486);
and U42390 (N_42390,N_39203,N_36813);
or U42391 (N_42391,N_37179,N_34416);
nand U42392 (N_42392,N_33954,N_30758);
and U42393 (N_42393,N_38581,N_39208);
nor U42394 (N_42394,N_37570,N_38978);
or U42395 (N_42395,N_35110,N_37845);
nand U42396 (N_42396,N_32688,N_34080);
or U42397 (N_42397,N_32643,N_37146);
nand U42398 (N_42398,N_38463,N_36432);
nand U42399 (N_42399,N_32464,N_35733);
nor U42400 (N_42400,N_38755,N_35386);
or U42401 (N_42401,N_33790,N_31659);
nand U42402 (N_42402,N_39653,N_31093);
or U42403 (N_42403,N_37429,N_38330);
and U42404 (N_42404,N_32084,N_31378);
or U42405 (N_42405,N_31348,N_33680);
nand U42406 (N_42406,N_34015,N_36737);
nand U42407 (N_42407,N_34309,N_32909);
xnor U42408 (N_42408,N_39329,N_32601);
nor U42409 (N_42409,N_31526,N_35637);
nand U42410 (N_42410,N_31350,N_31841);
nand U42411 (N_42411,N_37908,N_36915);
and U42412 (N_42412,N_38068,N_38804);
nor U42413 (N_42413,N_37322,N_36162);
and U42414 (N_42414,N_35246,N_31472);
and U42415 (N_42415,N_38556,N_30029);
nand U42416 (N_42416,N_39579,N_35181);
nor U42417 (N_42417,N_39741,N_37277);
and U42418 (N_42418,N_30318,N_31360);
nor U42419 (N_42419,N_32917,N_37151);
or U42420 (N_42420,N_38173,N_34916);
xnor U42421 (N_42421,N_37139,N_39181);
nand U42422 (N_42422,N_35797,N_36269);
nand U42423 (N_42423,N_37167,N_38060);
and U42424 (N_42424,N_37350,N_32411);
and U42425 (N_42425,N_35402,N_33564);
nand U42426 (N_42426,N_36636,N_34419);
or U42427 (N_42427,N_34066,N_33097);
and U42428 (N_42428,N_31801,N_30535);
and U42429 (N_42429,N_36794,N_35288);
or U42430 (N_42430,N_36884,N_38776);
or U42431 (N_42431,N_34342,N_33056);
and U42432 (N_42432,N_33439,N_38758);
or U42433 (N_42433,N_35395,N_31696);
or U42434 (N_42434,N_36616,N_39558);
nand U42435 (N_42435,N_39016,N_36163);
nand U42436 (N_42436,N_33853,N_33807);
nor U42437 (N_42437,N_31871,N_32088);
or U42438 (N_42438,N_37301,N_37158);
nand U42439 (N_42439,N_33753,N_32279);
nand U42440 (N_42440,N_31089,N_32931);
nand U42441 (N_42441,N_34103,N_35601);
or U42442 (N_42442,N_32285,N_33737);
nor U42443 (N_42443,N_33700,N_34379);
and U42444 (N_42444,N_34266,N_35727);
xor U42445 (N_42445,N_31685,N_38603);
or U42446 (N_42446,N_38449,N_37079);
xor U42447 (N_42447,N_38384,N_30511);
nand U42448 (N_42448,N_31820,N_32402);
or U42449 (N_42449,N_30786,N_33803);
nor U42450 (N_42450,N_30488,N_39562);
nor U42451 (N_42451,N_30291,N_36816);
or U42452 (N_42452,N_35446,N_35803);
and U42453 (N_42453,N_36424,N_37192);
xnor U42454 (N_42454,N_34468,N_34101);
nand U42455 (N_42455,N_39240,N_37180);
and U42456 (N_42456,N_37798,N_30973);
or U42457 (N_42457,N_34543,N_39550);
or U42458 (N_42458,N_36297,N_38634);
xor U42459 (N_42459,N_36637,N_33833);
and U42460 (N_42460,N_37507,N_31687);
nand U42461 (N_42461,N_36346,N_37722);
nor U42462 (N_42462,N_33555,N_38214);
nand U42463 (N_42463,N_30366,N_32918);
nor U42464 (N_42464,N_33474,N_37564);
nor U42465 (N_42465,N_36962,N_38983);
and U42466 (N_42466,N_36963,N_37058);
and U42467 (N_42467,N_36495,N_31898);
and U42468 (N_42468,N_32911,N_38279);
or U42469 (N_42469,N_34542,N_34242);
or U42470 (N_42470,N_39269,N_34993);
xnor U42471 (N_42471,N_39302,N_30400);
and U42472 (N_42472,N_35778,N_32106);
nor U42473 (N_42473,N_38656,N_36919);
nor U42474 (N_42474,N_32761,N_33265);
or U42475 (N_42475,N_30695,N_31814);
nor U42476 (N_42476,N_31481,N_37229);
and U42477 (N_42477,N_35340,N_37097);
and U42478 (N_42478,N_38568,N_30456);
and U42479 (N_42479,N_38961,N_35679);
or U42480 (N_42480,N_33685,N_33835);
nand U42481 (N_42481,N_35090,N_34660);
or U42482 (N_42482,N_35840,N_35223);
nand U42483 (N_42483,N_34245,N_32131);
nor U42484 (N_42484,N_37290,N_33494);
and U42485 (N_42485,N_39393,N_38251);
nand U42486 (N_42486,N_32801,N_36893);
and U42487 (N_42487,N_34791,N_31546);
nand U42488 (N_42488,N_34224,N_33336);
nand U42489 (N_42489,N_35493,N_32734);
nor U42490 (N_42490,N_39786,N_39320);
and U42491 (N_42491,N_31224,N_33511);
nor U42492 (N_42492,N_33864,N_38602);
or U42493 (N_42493,N_32443,N_38390);
nand U42494 (N_42494,N_30809,N_31832);
nor U42495 (N_42495,N_30751,N_39606);
and U42496 (N_42496,N_39376,N_35910);
nor U42497 (N_42497,N_30244,N_31882);
nand U42498 (N_42498,N_36726,N_34926);
xor U42499 (N_42499,N_30099,N_36385);
and U42500 (N_42500,N_33192,N_30752);
nor U42501 (N_42501,N_33525,N_37502);
or U42502 (N_42502,N_37561,N_37873);
and U42503 (N_42503,N_35415,N_36849);
nor U42504 (N_42504,N_37959,N_33865);
or U42505 (N_42505,N_38951,N_36473);
nor U42506 (N_42506,N_30951,N_38182);
or U42507 (N_42507,N_31092,N_39527);
and U42508 (N_42508,N_36172,N_32826);
or U42509 (N_42509,N_30598,N_31738);
nor U42510 (N_42510,N_33986,N_36219);
and U42511 (N_42511,N_36811,N_32076);
and U42512 (N_42512,N_38419,N_30460);
or U42513 (N_42513,N_31732,N_30267);
or U42514 (N_42514,N_34758,N_35200);
and U42515 (N_42515,N_36752,N_31315);
and U42516 (N_42516,N_39831,N_35918);
and U42517 (N_42517,N_34615,N_39988);
or U42518 (N_42518,N_30136,N_35276);
nor U42519 (N_42519,N_32303,N_37203);
and U42520 (N_42520,N_35728,N_39948);
or U42521 (N_42521,N_30549,N_33609);
and U42522 (N_42522,N_33082,N_34197);
and U42523 (N_42523,N_30831,N_34305);
or U42524 (N_42524,N_32499,N_37861);
nor U42525 (N_42525,N_34480,N_37282);
nand U42526 (N_42526,N_32367,N_37325);
xnor U42527 (N_42527,N_30208,N_30130);
nor U42528 (N_42528,N_36085,N_34802);
xor U42529 (N_42529,N_32549,N_34323);
nand U42530 (N_42530,N_35212,N_37957);
and U42531 (N_42531,N_34935,N_36501);
nor U42532 (N_42532,N_39837,N_30690);
and U42533 (N_42533,N_30007,N_35096);
and U42534 (N_42534,N_36203,N_30199);
or U42535 (N_42535,N_36755,N_33089);
nand U42536 (N_42536,N_39564,N_35003);
nand U42537 (N_42537,N_35642,N_38081);
nor U42538 (N_42538,N_37946,N_39251);
nor U42539 (N_42539,N_30496,N_34452);
nand U42540 (N_42540,N_33509,N_31405);
nor U42541 (N_42541,N_35268,N_34116);
nor U42542 (N_42542,N_32459,N_34738);
or U42543 (N_42543,N_33769,N_33914);
and U42544 (N_42544,N_39743,N_37270);
or U42545 (N_42545,N_32748,N_31544);
and U42546 (N_42546,N_39946,N_37518);
xor U42547 (N_42547,N_36897,N_38344);
nor U42548 (N_42548,N_33571,N_31959);
nand U42549 (N_42549,N_35816,N_30646);
and U42550 (N_42550,N_35082,N_31146);
nor U42551 (N_42551,N_30388,N_38539);
nand U42552 (N_42552,N_37420,N_35264);
and U42553 (N_42553,N_30143,N_32735);
or U42554 (N_42554,N_38537,N_39212);
or U42555 (N_42555,N_32109,N_33988);
nor U42556 (N_42556,N_31899,N_34258);
xor U42557 (N_42557,N_38378,N_34564);
nor U42558 (N_42558,N_39085,N_38253);
nor U42559 (N_42559,N_37298,N_35736);
nand U42560 (N_42560,N_30435,N_33503);
or U42561 (N_42561,N_32832,N_38099);
or U42562 (N_42562,N_33270,N_37972);
or U42563 (N_42563,N_30618,N_30103);
xor U42564 (N_42564,N_30251,N_35755);
and U42565 (N_42565,N_39283,N_33164);
nor U42566 (N_42566,N_32645,N_35253);
nor U42567 (N_42567,N_37050,N_32639);
nand U42568 (N_42568,N_35774,N_36865);
and U42569 (N_42569,N_32518,N_33373);
or U42570 (N_42570,N_36715,N_32714);
and U42571 (N_42571,N_32016,N_35382);
and U42572 (N_42572,N_38175,N_33357);
nor U42573 (N_42573,N_31015,N_32087);
xor U42574 (N_42574,N_38536,N_31163);
nor U42575 (N_42575,N_39385,N_37477);
nand U42576 (N_42576,N_33101,N_38907);
nor U42577 (N_42577,N_35241,N_31507);
or U42578 (N_42578,N_34398,N_32017);
or U42579 (N_42579,N_36013,N_38775);
nor U42580 (N_42580,N_32181,N_32689);
nand U42581 (N_42581,N_39398,N_30586);
and U42582 (N_42582,N_36011,N_32248);
xnor U42583 (N_42583,N_33645,N_31173);
or U42584 (N_42584,N_31005,N_38446);
or U42585 (N_42585,N_34939,N_33110);
nor U42586 (N_42586,N_39664,N_38492);
nor U42587 (N_42587,N_38013,N_36254);
or U42588 (N_42588,N_39849,N_32189);
and U42589 (N_42589,N_39155,N_38130);
and U42590 (N_42590,N_33776,N_37965);
and U42591 (N_42591,N_33468,N_31010);
nor U42592 (N_42592,N_35070,N_38067);
xnor U42593 (N_42593,N_30810,N_30903);
nor U42594 (N_42594,N_32925,N_39147);
nand U42595 (N_42595,N_30112,N_33522);
nand U42596 (N_42596,N_33419,N_30421);
or U42597 (N_42597,N_37115,N_38304);
or U42598 (N_42598,N_30790,N_32462);
nand U42599 (N_42599,N_35205,N_39851);
xnor U42600 (N_42600,N_32573,N_35013);
nor U42601 (N_42601,N_38854,N_39221);
nor U42602 (N_42602,N_36592,N_37263);
nand U42603 (N_42603,N_37709,N_39451);
and U42604 (N_42604,N_30294,N_31277);
nand U42605 (N_42605,N_37543,N_37671);
xor U42606 (N_42606,N_34927,N_37730);
and U42607 (N_42607,N_34241,N_36652);
or U42608 (N_42608,N_30940,N_35265);
or U42609 (N_42609,N_32267,N_39266);
nand U42610 (N_42610,N_34238,N_36166);
nor U42611 (N_42611,N_34970,N_33860);
nand U42612 (N_42612,N_33527,N_36441);
or U42613 (N_42613,N_31007,N_32664);
and U42614 (N_42614,N_35233,N_34373);
and U42615 (N_42615,N_34377,N_30836);
nand U42616 (N_42616,N_32392,N_31238);
and U42617 (N_42617,N_35349,N_30546);
or U42618 (N_42618,N_32957,N_37060);
or U42619 (N_42619,N_33633,N_38972);
nor U42620 (N_42620,N_39042,N_32660);
nand U42621 (N_42621,N_38633,N_30978);
nor U42622 (N_42622,N_30346,N_37947);
nand U42623 (N_42623,N_33017,N_36766);
and U42624 (N_42624,N_36828,N_35538);
nand U42625 (N_42625,N_36263,N_39821);
and U42626 (N_42626,N_39912,N_33421);
or U42627 (N_42627,N_34724,N_35124);
nor U42628 (N_42628,N_32800,N_32536);
or U42629 (N_42629,N_32915,N_33817);
and U42630 (N_42630,N_30924,N_33144);
nand U42631 (N_42631,N_39440,N_36607);
nor U42632 (N_42632,N_39594,N_33535);
or U42633 (N_42633,N_34288,N_36978);
xor U42634 (N_42634,N_35947,N_36026);
or U42635 (N_42635,N_37723,N_34736);
nand U42636 (N_42636,N_34784,N_32166);
nor U42637 (N_42637,N_36267,N_31080);
xor U42638 (N_42638,N_36643,N_36712);
xnor U42639 (N_42639,N_31202,N_30902);
nand U42640 (N_42640,N_33514,N_33670);
nand U42641 (N_42641,N_37794,N_38749);
or U42642 (N_42642,N_39515,N_31823);
nand U42643 (N_42643,N_35134,N_33045);
nor U42644 (N_42644,N_30082,N_30863);
nor U42645 (N_42645,N_33672,N_30482);
nor U42646 (N_42646,N_34843,N_34469);
nand U42647 (N_42647,N_35510,N_31191);
nand U42648 (N_42648,N_33234,N_33518);
and U42649 (N_42649,N_38672,N_34028);
nor U42650 (N_42650,N_39979,N_33453);
and U42651 (N_42651,N_33818,N_35106);
and U42652 (N_42652,N_32489,N_33931);
and U42653 (N_42653,N_30754,N_33119);
nor U42654 (N_42654,N_33789,N_36578);
nand U42655 (N_42655,N_39923,N_34022);
nor U42656 (N_42656,N_30588,N_36239);
nand U42657 (N_42657,N_34955,N_36440);
or U42658 (N_42658,N_30224,N_34349);
and U42659 (N_42659,N_37882,N_36372);
and U42660 (N_42660,N_35081,N_34580);
or U42661 (N_42661,N_38922,N_33388);
or U42662 (N_42662,N_39632,N_34896);
xnor U42663 (N_42663,N_34876,N_33198);
and U42664 (N_42664,N_38950,N_36303);
or U42665 (N_42665,N_38247,N_35045);
and U42666 (N_42666,N_38167,N_36873);
nand U42667 (N_42667,N_37991,N_39137);
xor U42668 (N_42668,N_39083,N_36182);
nand U42669 (N_42669,N_36600,N_32589);
and U42670 (N_42670,N_31572,N_37836);
or U42671 (N_42671,N_31070,N_38112);
xor U42672 (N_42672,N_33588,N_30124);
nor U42673 (N_42673,N_35248,N_31199);
and U42674 (N_42674,N_37216,N_30452);
nand U42675 (N_42675,N_36357,N_33282);
nand U42676 (N_42676,N_33165,N_33210);
nand U42677 (N_42677,N_36287,N_34450);
or U42678 (N_42678,N_37705,N_39891);
and U42679 (N_42679,N_37601,N_39123);
xnor U42680 (N_42680,N_31936,N_35839);
nand U42681 (N_42681,N_34307,N_31391);
or U42682 (N_42682,N_37299,N_37256);
nor U42683 (N_42683,N_35406,N_34636);
and U42684 (N_42684,N_39449,N_34145);
or U42685 (N_42685,N_36231,N_34838);
nand U42686 (N_42686,N_37894,N_33406);
nor U42687 (N_42687,N_32647,N_36164);
or U42688 (N_42688,N_36233,N_30212);
or U42689 (N_42689,N_34788,N_32784);
nand U42690 (N_42690,N_37693,N_33896);
nor U42691 (N_42691,N_38929,N_39339);
nand U42692 (N_42692,N_31485,N_36132);
and U42693 (N_42693,N_31410,N_38837);
and U42694 (N_42694,N_30297,N_37093);
xor U42695 (N_42695,N_34678,N_31072);
and U42696 (N_42696,N_37997,N_35320);
nor U42697 (N_42697,N_33740,N_33075);
nand U42698 (N_42698,N_34067,N_33602);
xor U42699 (N_42699,N_38493,N_31661);
nor U42700 (N_42700,N_30218,N_34186);
nor U42701 (N_42701,N_34071,N_39044);
and U42702 (N_42702,N_35479,N_38134);
and U42703 (N_42703,N_30590,N_36351);
nor U42704 (N_42704,N_39353,N_32655);
nor U42705 (N_42705,N_33744,N_36640);
and U42706 (N_42706,N_35631,N_30826);
nand U42707 (N_42707,N_39074,N_35347);
and U42708 (N_42708,N_33611,N_37711);
nor U42709 (N_42709,N_37262,N_30121);
or U42710 (N_42710,N_36697,N_31997);
and U42711 (N_42711,N_34313,N_38769);
or U42712 (N_42712,N_30257,N_35924);
and U42713 (N_42713,N_36972,N_35266);
nor U42714 (N_42714,N_30663,N_34807);
and U42715 (N_42715,N_31699,N_30443);
nand U42716 (N_42716,N_31620,N_33770);
and U42717 (N_42717,N_38033,N_35280);
nor U42718 (N_42718,N_34219,N_35422);
nand U42719 (N_42719,N_35748,N_34566);
nand U42720 (N_42720,N_30569,N_36731);
nor U42721 (N_42721,N_38230,N_35141);
nand U42722 (N_42722,N_31143,N_30968);
or U42723 (N_42723,N_37494,N_37452);
nor U42724 (N_42724,N_32331,N_38594);
nor U42725 (N_42725,N_35496,N_35653);
and U42726 (N_42726,N_34058,N_36586);
or U42727 (N_42727,N_36795,N_37135);
nor U42728 (N_42728,N_39227,N_37036);
nor U42729 (N_42729,N_31643,N_39180);
or U42730 (N_42730,N_36834,N_32760);
or U42731 (N_42731,N_37198,N_33918);
and U42732 (N_42732,N_36815,N_39382);
nand U42733 (N_42733,N_37614,N_33096);
nand U42734 (N_42734,N_35211,N_39054);
nand U42735 (N_42735,N_35196,N_33278);
nor U42736 (N_42736,N_35908,N_36598);
nand U42737 (N_42737,N_33928,N_36488);
nand U42738 (N_42738,N_36009,N_30982);
or U42739 (N_42739,N_37090,N_39098);
nand U42740 (N_42740,N_37651,N_39483);
xnor U42741 (N_42741,N_33617,N_38401);
or U42742 (N_42742,N_36305,N_32522);
and U42743 (N_42743,N_37091,N_35543);
nand U42744 (N_42744,N_31372,N_30209);
nor U42745 (N_42745,N_39126,N_35916);
and U42746 (N_42746,N_34799,N_37555);
nand U42747 (N_42747,N_30201,N_33880);
and U42748 (N_42748,N_36236,N_34303);
nor U42749 (N_42749,N_37790,N_33379);
and U42750 (N_42750,N_39985,N_34609);
nand U42751 (N_42751,N_32152,N_32271);
xor U42752 (N_42752,N_33592,N_36876);
xnor U42753 (N_42753,N_37870,N_32963);
and U42754 (N_42754,N_36082,N_38970);
nor U42755 (N_42755,N_38985,N_38469);
nand U42756 (N_42756,N_33607,N_37150);
and U42757 (N_42757,N_35558,N_33154);
nor U42758 (N_42758,N_39296,N_37281);
nor U42759 (N_42759,N_38455,N_34215);
or U42760 (N_42760,N_35683,N_35565);
nor U42761 (N_42761,N_32998,N_30872);
nand U42762 (N_42762,N_38668,N_38952);
nor U42763 (N_42763,N_38583,N_39633);
or U42764 (N_42764,N_37829,N_37513);
or U42765 (N_42765,N_32104,N_38933);
nor U42766 (N_42766,N_30851,N_39438);
or U42767 (N_42767,N_38346,N_39938);
and U42768 (N_42768,N_30490,N_33619);
and U42769 (N_42769,N_32520,N_38528);
nor U42770 (N_42770,N_30474,N_39193);
and U42771 (N_42771,N_30004,N_36033);
nor U42772 (N_42772,N_39532,N_34263);
nand U42773 (N_42773,N_35540,N_31700);
nand U42774 (N_42774,N_34661,N_33961);
nand U42775 (N_42775,N_39623,N_34109);
and U42776 (N_42776,N_36204,N_39641);
and U42777 (N_42777,N_31220,N_33235);
or U42778 (N_42778,N_33777,N_30908);
or U42779 (N_42779,N_38172,N_35338);
and U42780 (N_42780,N_37080,N_37655);
nand U42781 (N_42781,N_35389,N_33427);
xor U42782 (N_42782,N_30969,N_38285);
or U42783 (N_42783,N_37041,N_30734);
nor U42784 (N_42784,N_34558,N_31274);
nand U42785 (N_42785,N_31103,N_36841);
nand U42786 (N_42786,N_32438,N_39093);
nor U42787 (N_42787,N_36542,N_33622);
and U42788 (N_42788,N_31731,N_39951);
or U42789 (N_42789,N_33133,N_30524);
nor U42790 (N_42790,N_31571,N_37042);
nor U42791 (N_42791,N_39950,N_34950);
and U42792 (N_42792,N_37075,N_39164);
and U42793 (N_42793,N_32171,N_38252);
nand U42794 (N_42794,N_35108,N_37859);
or U42795 (N_42795,N_37539,N_31606);
or U42796 (N_42796,N_39908,N_30407);
xor U42797 (N_42797,N_31067,N_31747);
or U42798 (N_42798,N_38165,N_33839);
nand U42799 (N_42799,N_33635,N_31204);
nand U42800 (N_42800,N_38272,N_37986);
and U42801 (N_42801,N_31804,N_38916);
nor U42802 (N_42802,N_33002,N_32008);
and U42803 (N_42803,N_36092,N_32870);
or U42804 (N_42804,N_34632,N_39418);
nor U42805 (N_42805,N_30132,N_35856);
xor U42806 (N_42806,N_35737,N_32728);
or U42807 (N_42807,N_30161,N_38140);
and U42808 (N_42808,N_36417,N_32670);
nor U42809 (N_42809,N_36490,N_32448);
or U42810 (N_42810,N_39001,N_36198);
xor U42811 (N_42811,N_37763,N_38168);
xor U42812 (N_42812,N_31341,N_39581);
nor U42813 (N_42813,N_31684,N_30867);
and U42814 (N_42814,N_32241,N_34980);
or U42815 (N_42815,N_31916,N_37408);
and U42816 (N_42816,N_33690,N_35490);
xnor U42817 (N_42817,N_36015,N_32015);
nand U42818 (N_42818,N_32254,N_32979);
and U42819 (N_42819,N_34367,N_33478);
nor U42820 (N_42820,N_33159,N_37501);
xor U42821 (N_42821,N_31837,N_39650);
nand U42822 (N_42822,N_32921,N_34757);
nand U42823 (N_42823,N_32249,N_38732);
or U42824 (N_42824,N_35771,N_32929);
nor U42825 (N_42825,N_38679,N_37142);
and U42826 (N_42826,N_32226,N_37014);
nor U42827 (N_42827,N_32910,N_38045);
nand U42828 (N_42828,N_33933,N_33314);
and U42829 (N_42829,N_35193,N_34248);
nor U42830 (N_42830,N_30942,N_38226);
or U42831 (N_42831,N_30128,N_37657);
nor U42832 (N_42832,N_30391,N_38396);
or U42833 (N_42833,N_34127,N_38163);
and U42834 (N_42834,N_30675,N_35777);
or U42835 (N_42835,N_37159,N_30536);
or U42836 (N_42836,N_36713,N_36770);
nand U42837 (N_42837,N_31998,N_31106);
nand U42838 (N_42838,N_33088,N_32865);
nand U42839 (N_42839,N_39435,N_30202);
nor U42840 (N_42840,N_31336,N_38617);
and U42841 (N_42841,N_38514,N_35556);
nand U42842 (N_42842,N_39858,N_38875);
nor U42843 (N_42843,N_33366,N_35083);
and U42844 (N_42844,N_37893,N_38550);
or U42845 (N_42845,N_31902,N_33945);
or U42846 (N_42846,N_34009,N_34196);
xor U42847 (N_42847,N_30330,N_34118);
and U42848 (N_42848,N_30091,N_33960);
nor U42849 (N_42849,N_33151,N_31214);
nor U42850 (N_42850,N_31729,N_33364);
and U42851 (N_42851,N_38224,N_39048);
nand U42852 (N_42852,N_36577,N_36833);
nand U42853 (N_42853,N_30420,N_31583);
or U42854 (N_42854,N_38062,N_37181);
or U42855 (N_42855,N_31779,N_36259);
nand U42856 (N_42856,N_35143,N_36608);
nor U42857 (N_42857,N_31723,N_39400);
or U42858 (N_42858,N_32580,N_31806);
nand U42859 (N_42859,N_35010,N_32964);
xor U42860 (N_42860,N_32876,N_36904);
nor U42861 (N_42861,N_39827,N_35114);
xnor U42862 (N_42862,N_33376,N_39771);
and U42863 (N_42863,N_39262,N_30893);
nand U42864 (N_42864,N_36792,N_33858);
or U42865 (N_42865,N_39217,N_37628);
and U42866 (N_42866,N_31134,N_39131);
and U42867 (N_42867,N_31927,N_39198);
nand U42868 (N_42868,N_30946,N_36518);
and U42869 (N_42869,N_36751,N_31029);
or U42870 (N_42870,N_36807,N_36171);
and U42871 (N_42871,N_39587,N_36131);
and U42872 (N_42872,N_38888,N_34268);
nand U42873 (N_42873,N_34668,N_36470);
nor U42874 (N_42874,N_31966,N_37862);
and U42875 (N_42875,N_33200,N_38859);
and U42876 (N_42876,N_36031,N_39613);
nor U42877 (N_42877,N_31117,N_34378);
or U42878 (N_42878,N_37031,N_39334);
or U42879 (N_42879,N_37061,N_39657);
nand U42880 (N_42880,N_30164,N_38635);
and U42881 (N_42881,N_32946,N_36273);
xor U42882 (N_42882,N_39060,N_38200);
and U42883 (N_42883,N_37072,N_30705);
xnor U42884 (N_42884,N_37028,N_31625);
and U42885 (N_42885,N_32154,N_35614);
xor U42886 (N_42886,N_36044,N_32326);
or U42887 (N_42887,N_34924,N_35277);
nor U42888 (N_42888,N_30512,N_37409);
and U42889 (N_42889,N_36883,N_30685);
or U42890 (N_42890,N_32768,N_35741);
and U42891 (N_42891,N_38058,N_38855);
nor U42892 (N_42892,N_30959,N_33757);
xor U42893 (N_42893,N_30376,N_38684);
nand U42894 (N_42894,N_39037,N_39682);
xor U42895 (N_42895,N_32702,N_32616);
nor U42896 (N_42896,N_36929,N_37942);
nand U42897 (N_42897,N_36980,N_35417);
xor U42898 (N_42898,N_34017,N_33389);
nor U42899 (N_42899,N_33247,N_34857);
nand U42900 (N_42900,N_35535,N_32091);
and U42901 (N_42901,N_39059,N_39755);
nand U42902 (N_42902,N_32147,N_38007);
and U42903 (N_42903,N_34808,N_36436);
nor U42904 (N_42904,N_36513,N_38853);
xor U42905 (N_42905,N_30343,N_32329);
or U42906 (N_42906,N_36098,N_34481);
and U42907 (N_42907,N_34745,N_38564);
and U42908 (N_42908,N_31586,N_39261);
xor U42909 (N_42909,N_39802,N_34329);
xnor U42910 (N_42910,N_34717,N_34575);
nor U42911 (N_42911,N_31078,N_37403);
nand U42912 (N_42912,N_36532,N_39969);
nor U42913 (N_42913,N_38103,N_34822);
nand U42914 (N_42914,N_32906,N_33174);
nor U42915 (N_42915,N_36475,N_39331);
and U42916 (N_42916,N_38815,N_32115);
or U42917 (N_42917,N_30755,N_39524);
nor U42918 (N_42918,N_34874,N_32023);
and U42919 (N_42919,N_31357,N_30306);
xor U42920 (N_42920,N_35250,N_39690);
nor U42921 (N_42921,N_33440,N_31418);
xnor U42922 (N_42922,N_38073,N_31213);
or U42923 (N_42923,N_34992,N_31128);
nand U42924 (N_42924,N_36584,N_33340);
or U42925 (N_42925,N_31045,N_38310);
or U42926 (N_42926,N_34873,N_34072);
xnor U42927 (N_42927,N_39248,N_38017);
nor U42928 (N_42928,N_38254,N_38404);
nor U42929 (N_42929,N_33855,N_34188);
nor U42930 (N_42930,N_30561,N_37772);
nand U42931 (N_42931,N_35542,N_31016);
or U42932 (N_42932,N_38506,N_39322);
nand U42933 (N_42933,N_35793,N_39407);
nor U42934 (N_42934,N_34521,N_39300);
or U42935 (N_42935,N_35337,N_36270);
and U42936 (N_42936,N_34640,N_36975);
and U42937 (N_42937,N_38979,N_33703);
nand U42938 (N_42938,N_33613,N_30387);
xor U42939 (N_42939,N_35591,N_30475);
nor U42940 (N_42940,N_31008,N_31809);
or U42941 (N_42941,N_31845,N_38355);
or U42942 (N_42942,N_33482,N_39629);
nor U42943 (N_42943,N_37860,N_33521);
nor U42944 (N_42944,N_37802,N_38778);
and U42945 (N_42945,N_37176,N_31989);
or U42946 (N_42946,N_39665,N_34194);
or U42947 (N_42947,N_30871,N_32945);
and U42948 (N_42948,N_33274,N_37453);
or U42949 (N_42949,N_37676,N_34971);
and U42950 (N_42950,N_32095,N_35379);
or U42951 (N_42951,N_31511,N_33796);
or U42952 (N_42952,N_30567,N_30066);
or U42953 (N_42953,N_31521,N_34296);
and U42954 (N_42954,N_30910,N_33537);
nor U42955 (N_42955,N_32376,N_37701);
nand U42956 (N_42956,N_32368,N_33086);
nor U42957 (N_42957,N_34713,N_33572);
nor U42958 (N_42958,N_35466,N_36114);
nor U42959 (N_42959,N_30241,N_33746);
nor U42960 (N_42960,N_33688,N_36105);
xor U42961 (N_42961,N_35051,N_37117);
xnor U42962 (N_42962,N_37804,N_31298);
or U42963 (N_42963,N_38508,N_33476);
or U42964 (N_42964,N_37412,N_34859);
nor U42965 (N_42965,N_36095,N_37351);
xor U42966 (N_42966,N_36509,N_33363);
nand U42967 (N_42967,N_36894,N_37524);
nor U42968 (N_42968,N_35427,N_38982);
nor U42969 (N_42969,N_30085,N_30446);
and U42970 (N_42970,N_34462,N_32605);
and U42971 (N_42971,N_30728,N_30952);
nor U42972 (N_42972,N_39577,N_32292);
or U42973 (N_42973,N_39335,N_30913);
nor U42974 (N_42974,N_35776,N_32335);
or U42975 (N_42975,N_38695,N_36666);
nor U42976 (N_42976,N_36646,N_31943);
and U42977 (N_42977,N_34578,N_34508);
nand U42978 (N_42978,N_34410,N_36567);
nor U42979 (N_42979,N_37197,N_31860);
xnor U42980 (N_42980,N_31139,N_39999);
or U42981 (N_42981,N_30067,N_37892);
or U42982 (N_42982,N_39391,N_33750);
nand U42983 (N_42983,N_33091,N_32280);
nand U42984 (N_42984,N_33217,N_39830);
nand U42985 (N_42985,N_35985,N_38898);
nor U42986 (N_42986,N_33767,N_31404);
nand U42987 (N_42987,N_33031,N_32218);
xor U42988 (N_42988,N_33024,N_37992);
nand U42989 (N_42989,N_30639,N_38817);
nand U42990 (N_42990,N_31292,N_39064);
and U42991 (N_42991,N_37519,N_35169);
nor U42992 (N_42992,N_38677,N_33799);
and U42993 (N_42993,N_37558,N_32018);
and U42994 (N_42994,N_37172,N_36147);
nand U42995 (N_42995,N_33013,N_32284);
xnor U42996 (N_42996,N_35433,N_38042);
and U42997 (N_42997,N_37410,N_35640);
or U42998 (N_42998,N_36680,N_39470);
and U42999 (N_42999,N_31396,N_30494);
nor U43000 (N_43000,N_39355,N_35047);
or U43001 (N_43001,N_35553,N_34075);
or U43002 (N_43002,N_37766,N_32049);
and U43003 (N_43003,N_38347,N_32992);
nor U43004 (N_43004,N_36008,N_37010);
xor U43005 (N_43005,N_34742,N_36504);
nor U43006 (N_43006,N_36062,N_39399);
nor U43007 (N_43007,N_36106,N_38552);
nand U43008 (N_43008,N_34534,N_34595);
or U43009 (N_43009,N_33906,N_34432);
xnor U43010 (N_43010,N_37257,N_36627);
nor U43011 (N_43011,N_39411,N_39838);
nor U43012 (N_43012,N_31535,N_31153);
nor U43013 (N_43013,N_33546,N_37700);
nand U43014 (N_43014,N_36864,N_34200);
and U43015 (N_43015,N_35997,N_39542);
and U43016 (N_43016,N_30844,N_38056);
or U43017 (N_43017,N_39663,N_37938);
xor U43018 (N_43018,N_32762,N_35919);
nand U43019 (N_43019,N_32162,N_32709);
or U43020 (N_43020,N_36789,N_30829);
and U43021 (N_43021,N_36718,N_38849);
and U43022 (N_43022,N_31816,N_30964);
or U43023 (N_43023,N_30789,N_31229);
nand U43024 (N_43024,N_37981,N_32764);
nor U43025 (N_43025,N_39057,N_36838);
xnor U43026 (N_43026,N_36779,N_31283);
nand U43027 (N_43027,N_35388,N_39233);
nand U43028 (N_43028,N_32632,N_35806);
nand U43029 (N_43029,N_34908,N_31424);
or U43030 (N_43030,N_34293,N_38873);
xnor U43031 (N_43031,N_38938,N_30866);
or U43032 (N_43032,N_33516,N_32430);
and U43033 (N_43033,N_34581,N_35926);
and U43034 (N_43034,N_30676,N_30280);
xor U43035 (N_43035,N_33201,N_32972);
or U43036 (N_43036,N_38625,N_37313);
or U43037 (N_43037,N_38962,N_38296);
and U43038 (N_43038,N_39206,N_31129);
and U43039 (N_43039,N_33382,N_32704);
nor U43040 (N_43040,N_31651,N_38750);
or U43041 (N_43041,N_35898,N_37515);
nor U43042 (N_43042,N_33411,N_39116);
or U43043 (N_43043,N_38116,N_33335);
nand U43044 (N_43044,N_33816,N_35028);
or U43045 (N_43045,N_38011,N_30249);
and U43046 (N_43046,N_34239,N_30250);
nand U43047 (N_43047,N_37523,N_30068);
nand U43048 (N_43048,N_34456,N_31624);
or U43049 (N_43049,N_34750,N_33268);
nand U43050 (N_43050,N_39094,N_30369);
nor U43051 (N_43051,N_37253,N_35625);
and U43052 (N_43052,N_38956,N_33605);
or U43053 (N_43053,N_34136,N_36111);
xor U43054 (N_43054,N_38072,N_35632);
or U43055 (N_43055,N_30088,N_33043);
or U43056 (N_43056,N_36604,N_32817);
nor U43057 (N_43057,N_30342,N_36982);
or U43058 (N_43058,N_37533,N_33768);
or U43059 (N_43059,N_35917,N_34264);
and U43060 (N_43060,N_32668,N_39671);
or U43061 (N_43061,N_36150,N_35467);
xor U43062 (N_43062,N_31061,N_33941);
nand U43063 (N_43063,N_39829,N_37222);
nor U43064 (N_43064,N_32712,N_32396);
nor U43065 (N_43065,N_34180,N_32213);
or U43066 (N_43066,N_34460,N_30744);
xnor U43067 (N_43067,N_31636,N_37297);
nor U43068 (N_43068,N_36186,N_31084);
and U43069 (N_43069,N_39754,N_38710);
nor U43070 (N_43070,N_36846,N_39843);
nor U43071 (N_43071,N_33050,N_34825);
nor U43072 (N_43072,N_39947,N_36018);
nand U43073 (N_43073,N_35450,N_35903);
nand U43074 (N_43074,N_39535,N_38217);
nor U43075 (N_43075,N_30065,N_36081);
or U43076 (N_43076,N_33432,N_33948);
or U43077 (N_43077,N_31186,N_35158);
nand U43078 (N_43078,N_35883,N_38623);
nand U43079 (N_43079,N_39953,N_33423);
nor U43080 (N_43080,N_36848,N_35600);
or U43081 (N_43081,N_39668,N_35703);
nor U43082 (N_43082,N_32569,N_31621);
and U43083 (N_43083,N_31570,N_31588);
and U43084 (N_43084,N_39937,N_31954);
nand U43085 (N_43085,N_35167,N_30759);
or U43086 (N_43086,N_35303,N_32393);
or U43087 (N_43087,N_33033,N_31849);
nor U43088 (N_43088,N_32902,N_30735);
or U43089 (N_43089,N_30781,N_37367);
or U43090 (N_43090,N_36235,N_34068);
or U43091 (N_43091,N_34929,N_37648);
nor U43092 (N_43092,N_32829,N_37214);
xnor U43093 (N_43093,N_35888,N_32216);
nor U43094 (N_43094,N_35156,N_35818);
xnor U43095 (N_43095,N_31301,N_39810);
nand U43096 (N_43096,N_39740,N_33076);
and U43097 (N_43097,N_31870,N_32217);
nand U43098 (N_43098,N_35628,N_34570);
or U43099 (N_43099,N_31523,N_38988);
nor U43100 (N_43100,N_37394,N_38001);
and U43101 (N_43101,N_31650,N_37618);
or U43102 (N_43102,N_35491,N_39492);
or U43103 (N_43103,N_34621,N_32405);
or U43104 (N_43104,N_37461,N_38333);
and U43105 (N_43105,N_31271,N_38661);
xor U43106 (N_43106,N_32685,N_35886);
or U43107 (N_43107,N_32782,N_35107);
and U43108 (N_43108,N_35066,N_36803);
or U43109 (N_43109,N_36223,N_34674);
nor U43110 (N_43110,N_30365,N_37092);
or U43111 (N_43111,N_35328,N_36583);
and U43112 (N_43112,N_38912,N_36924);
nand U43113 (N_43113,N_39282,N_38839);
nor U43114 (N_43114,N_39919,N_36531);
nand U43115 (N_43115,N_33087,N_32458);
xor U43116 (N_43116,N_35887,N_30779);
or U43117 (N_43117,N_35824,N_31552);
xor U43118 (N_43118,N_34553,N_35290);
and U43119 (N_43119,N_30135,N_39312);
nand U43120 (N_43120,N_34586,N_37864);
or U43121 (N_43121,N_32615,N_31366);
nand U43122 (N_43122,N_38133,N_39789);
and U43123 (N_43123,N_32075,N_30720);
nand U43124 (N_43124,N_30075,N_36533);
nand U43125 (N_43125,N_32766,N_31768);
and U43126 (N_43126,N_39659,N_31433);
or U43127 (N_43127,N_30247,N_35656);
nor U43128 (N_43128,N_38671,N_35725);
or U43129 (N_43129,N_32371,N_37680);
xnor U43130 (N_43130,N_33204,N_37739);
and U43131 (N_43131,N_31730,N_30351);
nand U43132 (N_43132,N_33659,N_35658);
or U43133 (N_43133,N_39285,N_31947);
nand U43134 (N_43134,N_35938,N_39917);
or U43135 (N_43135,N_35011,N_38730);
nand U43136 (N_43136,N_34477,N_32614);
and U43137 (N_43137,N_39720,N_34012);
nand U43138 (N_43138,N_38114,N_30123);
nor U43139 (N_43139,N_37850,N_30564);
nor U43140 (N_43140,N_37952,N_32232);
and U43141 (N_43141,N_30079,N_34295);
and U43142 (N_43142,N_34493,N_36778);
or U43143 (N_43143,N_36373,N_36321);
nand U43144 (N_43144,N_36155,N_32582);
or U43145 (N_43145,N_33772,N_38161);
nor U43146 (N_43146,N_34317,N_32070);
and U43147 (N_43147,N_37840,N_37672);
xor U43148 (N_43148,N_31147,N_32777);
xnor U43149 (N_43149,N_33058,N_30906);
and U43150 (N_43150,N_34665,N_32306);
nor U43151 (N_43151,N_33281,N_35456);
nand U43152 (N_43152,N_37761,N_33481);
and U43153 (N_43153,N_31159,N_32794);
nor U43154 (N_43154,N_36257,N_33702);
nand U43155 (N_43155,N_32257,N_34149);
nand U43156 (N_43156,N_33140,N_33946);
nand U43157 (N_43157,N_39127,N_30837);
nor U43158 (N_43158,N_30878,N_36090);
nor U43159 (N_43159,N_34803,N_34272);
nand U43160 (N_43160,N_39434,N_39795);
and U43161 (N_43161,N_36271,N_33393);
nand U43162 (N_43162,N_39660,N_34528);
nand U43163 (N_43163,N_31566,N_38917);
or U43164 (N_43164,N_35847,N_35293);
nand U43165 (N_43165,N_34383,N_37810);
or U43166 (N_43166,N_34138,N_33851);
nor U43167 (N_43167,N_32375,N_33277);
or U43168 (N_43168,N_30808,N_32436);
xor U43169 (N_43169,N_31048,N_37249);
or U43170 (N_43170,N_35455,N_38021);
nand U43171 (N_43171,N_35499,N_33697);
nand U43172 (N_43172,N_36555,N_36133);
and U43173 (N_43173,N_36359,N_36112);
nor U43174 (N_43174,N_32498,N_32381);
or U43175 (N_43175,N_32047,N_30138);
nor U43176 (N_43176,N_32969,N_36671);
or U43177 (N_43177,N_30931,N_35128);
or U43178 (N_43178,N_37215,N_39873);
nor U43179 (N_43179,N_30977,N_31034);
or U43180 (N_43180,N_38680,N_39674);
or U43181 (N_43181,N_31681,N_30849);
or U43182 (N_43182,N_39845,N_31207);
and U43183 (N_43183,N_36340,N_33310);
or U43184 (N_43184,N_31912,N_34667);
xor U43185 (N_43185,N_34351,N_33813);
or U43186 (N_43186,N_38986,N_31657);
nand U43187 (N_43187,N_39785,N_33727);
nor U43188 (N_43188,N_39881,N_31256);
and U43189 (N_43189,N_39348,N_32913);
or U43190 (N_43190,N_37100,N_37373);
or U43191 (N_43191,N_30563,N_33497);
nor U43192 (N_43192,N_38435,N_35120);
or U43193 (N_43193,N_35969,N_37852);
nor U43194 (N_43194,N_34816,N_32555);
and U43195 (N_43195,N_39090,N_30107);
or U43196 (N_43196,N_33129,N_36684);
nand U43197 (N_43197,N_37756,N_38246);
or U43198 (N_43198,N_33113,N_39693);
nor U43199 (N_43199,N_36145,N_39401);
nand U43200 (N_43200,N_33094,N_34331);
nor U43201 (N_43201,N_35521,N_33138);
nor U43202 (N_43202,N_34969,N_34557);
and U43203 (N_43203,N_35504,N_35177);
or U43204 (N_43204,N_39404,N_35117);
nor U43205 (N_43205,N_31939,N_37377);
xor U43206 (N_43206,N_35899,N_33387);
nand U43207 (N_43207,N_32176,N_30689);
nand U43208 (N_43208,N_34681,N_34910);
or U43209 (N_43209,N_35275,N_34841);
nor U43210 (N_43210,N_39305,N_33827);
and U43211 (N_43211,N_33275,N_37295);
nor U43212 (N_43212,N_31741,N_37855);
nand U43213 (N_43213,N_35476,N_30231);
or U43214 (N_43214,N_37493,N_32468);
xnor U43215 (N_43215,N_31009,N_33655);
or U43216 (N_43216,N_31873,N_31875);
or U43217 (N_43217,N_35676,N_35247);
nand U43218 (N_43218,N_35761,N_37479);
and U43219 (N_43219,N_31135,N_38944);
xor U43220 (N_43220,N_31785,N_38764);
nor U43221 (N_43221,N_38301,N_34024);
nand U43222 (N_43222,N_34287,N_35783);
xor U43223 (N_43223,N_33671,N_38220);
nor U43224 (N_43224,N_35079,N_38868);
or U43225 (N_43225,N_35593,N_33010);
or U43226 (N_43226,N_32093,N_35920);
or U43227 (N_43227,N_31709,N_37983);
nand U43228 (N_43228,N_35041,N_36691);
nor U43229 (N_43229,N_32471,N_37443);
nor U43230 (N_43230,N_36537,N_31861);
or U43231 (N_43231,N_30464,N_34806);
nand U43232 (N_43232,N_32769,N_31627);
nor U43233 (N_43233,N_36856,N_32975);
xor U43234 (N_43234,N_34994,N_39554);
or U43235 (N_43235,N_33169,N_30035);
or U43236 (N_43236,N_35889,N_39685);
nor U43237 (N_43237,N_36624,N_33126);
nand U43238 (N_43238,N_31397,N_30500);
nand U43239 (N_43239,N_30005,N_36891);
or U43240 (N_43240,N_38806,N_39051);
nand U43241 (N_43241,N_38553,N_39414);
or U43242 (N_43242,N_39767,N_39790);
nor U43243 (N_43243,N_39964,N_34947);
nor U43244 (N_43244,N_31430,N_33118);
nand U43245 (N_43245,N_31757,N_34029);
and U43246 (N_43246,N_38940,N_30408);
nor U43247 (N_43247,N_38696,N_34423);
nand U43248 (N_43248,N_33782,N_33533);
and U43249 (N_43249,N_38100,N_34170);
nand U43250 (N_43250,N_35468,N_36949);
and U43251 (N_43251,N_31673,N_34552);
nand U43252 (N_43252,N_35300,N_31676);
and U43253 (N_43253,N_34169,N_33374);
or U43254 (N_43254,N_37109,N_30868);
and U43255 (N_43255,N_34252,N_39412);
or U43256 (N_43256,N_37673,N_33233);
xor U43257 (N_43257,N_32563,N_33734);
and U43258 (N_43258,N_39636,N_30402);
xor U43259 (N_43259,N_35611,N_39299);
nand U43260 (N_43260,N_34132,N_37236);
nor U43261 (N_43261,N_32188,N_39445);
nor U43262 (N_43262,N_38880,N_30918);
nor U43263 (N_43263,N_38352,N_30579);
or U43264 (N_43264,N_30521,N_32341);
and U43265 (N_43265,N_30262,N_37339);
nor U43266 (N_43266,N_36653,N_33735);
nand U43267 (N_43267,N_31377,N_31952);
nand U43268 (N_43268,N_30303,N_31504);
nand U43269 (N_43269,N_33819,N_36047);
and U43270 (N_43270,N_31453,N_36296);
and U43271 (N_43271,N_32771,N_31102);
and U43272 (N_43272,N_30162,N_36083);
nor U43273 (N_43273,N_34048,N_37866);
and U43274 (N_43274,N_32150,N_36427);
nor U43275 (N_43275,N_30077,N_32933);
or U43276 (N_43276,N_39231,N_36260);
nor U43277 (N_43277,N_37436,N_33220);
nor U43278 (N_43278,N_39455,N_38971);
and U43279 (N_43279,N_32720,N_32490);
xnor U43280 (N_43280,N_39257,N_37989);
or U43281 (N_43281,N_39484,N_38219);
nor U43282 (N_43282,N_31323,N_37213);
nor U43283 (N_43283,N_36786,N_38057);
nor U43284 (N_43284,N_39752,N_34866);
xnor U43285 (N_43285,N_31506,N_35693);
nor U43286 (N_43286,N_38881,N_36685);
or U43287 (N_43287,N_34918,N_32168);
and U43288 (N_43288,N_30409,N_32370);
nor U43289 (N_43289,N_36224,N_36494);
and U43290 (N_43290,N_30975,N_32412);
nor U43291 (N_43291,N_37876,N_37757);
xor U43292 (N_43292,N_31992,N_32222);
nand U43293 (N_43293,N_31189,N_30539);
nor U43294 (N_43294,N_30595,N_33444);
nor U43295 (N_43295,N_33721,N_38053);
and U43296 (N_43296,N_32584,N_38179);
nand U43297 (N_43297,N_34032,N_35394);
nand U43298 (N_43298,N_32593,N_31356);
nand U43299 (N_43299,N_38646,N_30967);
and U43300 (N_43300,N_38816,N_39081);
nor U43301 (N_43301,N_34154,N_39153);
or U43302 (N_43302,N_35960,N_30699);
nor U43303 (N_43303,N_33369,N_31097);
nand U43304 (N_43304,N_36934,N_31574);
nand U43305 (N_43305,N_36868,N_37309);
and U43306 (N_43306,N_39598,N_32064);
or U43307 (N_43307,N_37491,N_35487);
or U43308 (N_43308,N_32508,N_30896);
and U43309 (N_43309,N_31241,N_36507);
nand U43310 (N_43310,N_36218,N_32386);
nand U43311 (N_43311,N_34318,N_37076);
nor U43312 (N_43312,N_32237,N_33919);
nor U43313 (N_43313,N_37956,N_36638);
nand U43314 (N_43314,N_31766,N_37704);
nor U43315 (N_43315,N_30537,N_34178);
nand U43316 (N_43316,N_31555,N_38038);
nor U43317 (N_43317,N_36658,N_30133);
nor U43318 (N_43318,N_39184,N_38877);
or U43319 (N_43319,N_39800,N_34974);
or U43320 (N_43320,N_36758,N_33027);
nor U43321 (N_43321,N_37530,N_37440);
nor U43322 (N_43322,N_34284,N_39662);
nor U43323 (N_43323,N_36220,N_33038);
nand U43324 (N_43324,N_32952,N_31440);
and U43325 (N_43325,N_38905,N_38237);
nand U43326 (N_43326,N_34976,N_38481);
nor U43327 (N_43327,N_31300,N_33166);
and U43328 (N_43328,N_32597,N_37675);
nor U43329 (N_43329,N_38570,N_31075);
and U43330 (N_43330,N_30930,N_34440);
and U43331 (N_43331,N_32713,N_34025);
nor U43332 (N_43332,N_33911,N_38659);
nand U43333 (N_43333,N_38886,N_34010);
and U43334 (N_43334,N_32143,N_30672);
and U43335 (N_43335,N_32349,N_32307);
nand U43336 (N_43336,N_34865,N_38314);
and U43337 (N_43337,N_36516,N_36874);
or U43338 (N_43338,N_39474,N_38032);
or U43339 (N_43339,N_38233,N_35945);
or U43340 (N_43340,N_30898,N_36822);
and U43341 (N_43341,N_33039,N_37472);
or U43342 (N_43342,N_37535,N_35050);
or U43343 (N_43343,N_35635,N_35563);
nor U43344 (N_43344,N_36057,N_30628);
nor U43345 (N_43345,N_32863,N_38830);
xor U43346 (N_43346,N_33414,N_38444);
and U43347 (N_43347,N_33828,N_32431);
and U43348 (N_43348,N_37417,N_37462);
or U43349 (N_43349,N_34389,N_30619);
nor U43350 (N_43350,N_32839,N_34957);
nor U43351 (N_43351,N_37950,N_32886);
nand U43352 (N_43352,N_31865,N_31099);
nor U43353 (N_43353,N_34981,N_30718);
nand U43354 (N_43354,N_32401,N_31355);
or U43355 (N_43355,N_38144,N_38889);
or U43356 (N_43356,N_30196,N_36909);
and U43357 (N_43357,N_31469,N_32414);
nor U43358 (N_43358,N_31105,N_37465);
or U43359 (N_43359,N_37639,N_32435);
and U43360 (N_43360,N_33556,N_34413);
nand U43361 (N_43361,N_36656,N_37770);
nand U43362 (N_43362,N_35329,N_38458);
nor U43363 (N_43363,N_33077,N_32934);
or U43364 (N_43364,N_38866,N_39420);
xor U43365 (N_43365,N_39931,N_39194);
or U43366 (N_43366,N_31609,N_34824);
nor U43367 (N_43367,N_31265,N_32539);
nand U43368 (N_43368,N_36976,N_37885);
nand U43369 (N_43369,N_31590,N_33093);
nor U43370 (N_43370,N_32654,N_34752);
and U43371 (N_43371,N_30658,N_32219);
nand U43372 (N_43372,N_39410,N_34020);
nor U43373 (N_43373,N_30858,N_36262);
or U43374 (N_43374,N_35795,N_35475);
nor U43375 (N_43375,N_31780,N_37684);
and U43376 (N_43376,N_33181,N_31638);
xnor U43377 (N_43377,N_32570,N_38105);
or U43378 (N_43378,N_32519,N_31680);
and U43379 (N_43379,N_38349,N_38845);
and U43380 (N_43380,N_34151,N_38843);
and U43381 (N_43381,N_35392,N_31895);
nand U43382 (N_43382,N_34297,N_35175);
and U43383 (N_43383,N_30117,N_37582);
nor U43384 (N_43384,N_34656,N_36061);
nor U43385 (N_43385,N_31940,N_34682);
nand U43386 (N_43386,N_38014,N_39854);
and U43387 (N_43387,N_39774,N_39002);
or U43388 (N_43388,N_32050,N_37353);
and U43389 (N_43389,N_34516,N_32513);
and U43390 (N_43390,N_35238,N_30559);
nand U43391 (N_43391,N_38768,N_30372);
nand U43392 (N_43392,N_30608,N_31847);
nor U43393 (N_43393,N_38142,N_36842);
or U43394 (N_43394,N_37268,N_31211);
or U43395 (N_43395,N_30519,N_32521);
xor U43396 (N_43396,N_35752,N_32426);
or U43397 (N_43397,N_31537,N_39311);
nand U43398 (N_43398,N_34728,N_35934);
and U43399 (N_43399,N_31510,N_32840);
nor U43400 (N_43400,N_37391,N_30862);
nand U43401 (N_43401,N_39853,N_35204);
or U43402 (N_43402,N_30935,N_39933);
and U43403 (N_43403,N_37250,N_30630);
nand U43404 (N_43404,N_31376,N_37975);
or U43405 (N_43405,N_39548,N_36096);
nand U43406 (N_43406,N_36609,N_33422);
and U43407 (N_43407,N_36022,N_37347);
nor U43408 (N_43408,N_32984,N_30334);
nor U43409 (N_43409,N_38517,N_30492);
or U43410 (N_43410,N_38883,N_39075);
and U43411 (N_43411,N_38533,N_36050);
or U43412 (N_43412,N_34104,N_30428);
and U43413 (N_43413,N_39015,N_32072);
nand U43414 (N_43414,N_36952,N_39011);
and U43415 (N_43415,N_31607,N_31151);
nor U43416 (N_43416,N_37948,N_37397);
nand U43417 (N_43417,N_39444,N_39997);
nand U43418 (N_43418,N_31054,N_38535);
nor U43419 (N_43419,N_35339,N_36338);
xor U43420 (N_43420,N_38504,N_37285);
and U43421 (N_43421,N_32373,N_32857);
and U43422 (N_43422,N_31628,N_34051);
nor U43423 (N_43423,N_36720,N_37774);
nand U43424 (N_43424,N_30283,N_34499);
nand U43425 (N_43425,N_39377,N_32744);
and U43426 (N_43426,N_31185,N_34198);
nor U43427 (N_43427,N_31896,N_38423);
nand U43428 (N_43428,N_35923,N_36148);
and U43429 (N_43429,N_34018,N_36526);
or U43430 (N_43430,N_39835,N_34228);
nand U43431 (N_43431,N_32419,N_31600);
and U43432 (N_43432,N_33550,N_31704);
xor U43433 (N_43433,N_36614,N_37943);
nor U43434 (N_43434,N_36326,N_37677);
nand U43435 (N_43435,N_39275,N_36141);
xor U43436 (N_43436,N_32995,N_36153);
or U43437 (N_43437,N_34262,N_37814);
nand U43438 (N_43438,N_33044,N_33652);
or U43439 (N_43439,N_33301,N_36225);
nor U43440 (N_43440,N_34382,N_31172);
and U43441 (N_43441,N_38885,N_37688);
nand U43442 (N_43442,N_39878,N_30994);
or U43443 (N_43443,N_33185,N_37737);
or U43444 (N_43444,N_34949,N_30988);
and U43445 (N_43445,N_36384,N_37038);
nand U43446 (N_43446,N_35838,N_34688);
nor U43447 (N_43447,N_32447,N_32019);
nor U43448 (N_43448,N_39959,N_37340);
or U43449 (N_43449,N_35524,N_31393);
nand U43450 (N_43450,N_38174,N_31594);
nand U43451 (N_43451,N_37963,N_37421);
xor U43452 (N_43452,N_37463,N_39826);
or U43453 (N_43453,N_33409,N_36412);
and U43454 (N_43454,N_31695,N_31435);
nand U43455 (N_43455,N_37125,N_39078);
nor U43456 (N_43456,N_34094,N_38379);
and U43457 (N_43457,N_33186,N_32814);
or U43458 (N_43458,N_33712,N_30643);
nand U43459 (N_43459,N_38283,N_35252);
or U43460 (N_43460,N_31608,N_39796);
or U43461 (N_43461,N_35065,N_38076);
nor U43462 (N_43462,N_38491,N_32491);
and U43463 (N_43463,N_33785,N_31026);
nand U43464 (N_43464,N_33167,N_32752);
nand U43465 (N_43465,N_30374,N_39129);
nor U43466 (N_43466,N_32346,N_33272);
nor U43467 (N_43467,N_38872,N_31126);
and U43468 (N_43468,N_30116,N_32501);
or U43469 (N_43469,N_37916,N_31284);
nand U43470 (N_43470,N_33932,N_32525);
nand U43471 (N_43471,N_37280,N_36774);
and U43472 (N_43472,N_38041,N_34461);
or U43473 (N_43473,N_37225,N_38259);
and U43474 (N_43474,N_32078,N_31922);
nand U43475 (N_43475,N_37331,N_39914);
nand U43476 (N_43476,N_35870,N_35984);
nand U43477 (N_43477,N_34346,N_33759);
nor U43478 (N_43478,N_36892,N_32037);
nor U43479 (N_43479,N_36687,N_33132);
nand U43480 (N_43480,N_34040,N_37483);
nor U43481 (N_43481,N_32201,N_31132);
nor U43482 (N_43482,N_39544,N_35564);
or U43483 (N_43483,N_35132,N_32938);
nor U43484 (N_43484,N_34526,N_34358);
nand U43485 (N_43485,N_39255,N_37775);
and U43486 (N_43486,N_32055,N_36830);
and U43487 (N_43487,N_34527,N_31602);
nand U43488 (N_43488,N_36615,N_32127);
nor U43489 (N_43489,N_37935,N_35030);
nor U43490 (N_43490,N_37255,N_33788);
nor U43491 (N_43491,N_37318,N_39984);
nor U43492 (N_43492,N_34631,N_31637);
xnor U43493 (N_43493,N_30057,N_30309);
nor U43494 (N_43494,N_30180,N_30986);
and U43495 (N_43495,N_38089,N_38336);
and U43496 (N_43496,N_37603,N_35723);
nand U43497 (N_43497,N_38890,N_30084);
and U43498 (N_43498,N_30382,N_30225);
nand U43499 (N_43499,N_31714,N_35750);
nand U43500 (N_43500,N_33034,N_36187);
or U43501 (N_43501,N_32980,N_31652);
nand U43502 (N_43502,N_32446,N_35289);
nand U43503 (N_43503,N_31467,N_35526);
nor U43504 (N_43504,N_37193,N_30033);
xnor U43505 (N_43505,N_39427,N_31513);
or U43506 (N_43506,N_32348,N_35760);
nor U43507 (N_43507,N_30328,N_38351);
nand U43508 (N_43508,N_36872,N_30290);
and U43509 (N_43509,N_32884,N_33331);
and U43510 (N_43510,N_36410,N_31465);
and U43511 (N_43511,N_30767,N_34393);
nor U43512 (N_43512,N_37666,N_32603);
and U43513 (N_43513,N_36030,N_36908);
nand U43514 (N_43514,N_32157,N_31765);
xnor U43515 (N_43515,N_37414,N_39684);
nor U43516 (N_43516,N_34098,N_31508);
or U43517 (N_43517,N_37754,N_31739);
nor U43518 (N_43518,N_38193,N_34721);
and U43519 (N_43519,N_31149,N_30802);
nand U43520 (N_43520,N_34226,N_31379);
or U43521 (N_43521,N_32553,N_39698);
xor U43522 (N_43522,N_38459,N_38277);
nor U43523 (N_43523,N_31038,N_39498);
nor U43524 (N_43524,N_39540,N_30350);
and U43525 (N_43525,N_37608,N_30932);
nor U43526 (N_43526,N_34518,N_31253);
nor U43527 (N_43527,N_34846,N_32209);
xor U43528 (N_43528,N_32604,N_37594);
and U43529 (N_43529,N_39029,N_34715);
or U43530 (N_43530,N_34648,N_39433);
or U43531 (N_43531,N_32173,N_38400);
or U43532 (N_43532,N_38867,N_30981);
and U43533 (N_43533,N_39040,N_39867);
or U43534 (N_43534,N_38414,N_38170);
nand U43535 (N_43535,N_38622,N_34085);
nand U43536 (N_43536,N_39898,N_32637);
or U43537 (N_43537,N_31425,N_36869);
nor U43538 (N_43538,N_33894,N_39087);
and U43539 (N_43539,N_31856,N_33450);
xor U43540 (N_43540,N_37616,N_31663);
xor U43541 (N_43541,N_31260,N_32658);
or U43542 (N_43542,N_39313,N_32030);
and U43543 (N_43543,N_35443,N_38022);
or U43544 (N_43544,N_32140,N_39863);
and U43545 (N_43545,N_36041,N_35462);
or U43546 (N_43546,N_34680,N_34049);
or U43547 (N_43547,N_30427,N_33232);
nand U43548 (N_43548,N_34348,N_38565);
xor U43549 (N_43549,N_30451,N_36278);
nand U43550 (N_43550,N_35766,N_33292);
nor U43551 (N_43551,N_39003,N_36191);
nand U43552 (N_43552,N_33567,N_35987);
nor U43553 (N_43553,N_35740,N_33580);
nor U43554 (N_43554,N_32695,N_38838);
nor U43555 (N_43555,N_38640,N_37346);
and U43556 (N_43556,N_39100,N_32052);
or U43557 (N_43557,N_36088,N_32612);
or U43558 (N_43558,N_36463,N_34209);
nor U43559 (N_43559,N_37712,N_33857);
nand U43560 (N_43560,N_33886,N_30324);
and U43561 (N_43561,N_32421,N_33004);
nand U43562 (N_43562,N_33327,N_37599);
nand U43563 (N_43563,N_33319,N_31735);
nand U43564 (N_43564,N_32706,N_39700);
nand U43565 (N_43565,N_30370,N_38590);
nor U43566 (N_43566,N_37319,N_39780);
nand U43567 (N_43567,N_30401,N_35474);
and U43568 (N_43568,N_36077,N_38411);
or U43569 (N_43569,N_36437,N_37333);
and U43570 (N_43570,N_35661,N_31228);
or U43571 (N_43571,N_37868,N_39067);
nor U43572 (N_43572,N_32295,N_35149);
nand U43573 (N_43573,N_37474,N_33260);
nand U43574 (N_43574,N_31242,N_38350);
and U43575 (N_43575,N_36185,N_32532);
or U43576 (N_43576,N_38436,N_37619);
nand U43577 (N_43577,N_34021,N_37504);
nand U43578 (N_43578,N_33108,N_31046);
nor U43579 (N_43579,N_31985,N_38292);
or U43580 (N_43580,N_33749,N_37685);
and U43581 (N_43581,N_38468,N_39270);
nor U43582 (N_43582,N_37702,N_33290);
and U43583 (N_43583,N_36484,N_38260);
nor U43584 (N_43584,N_35578,N_32389);
nor U43585 (N_43585,N_39705,N_33665);
nand U43586 (N_43586,N_33800,N_38746);
and U43587 (N_43587,N_39944,N_32174);
and U43588 (N_43588,N_33471,N_36700);
and U43589 (N_43589,N_35251,N_36689);
or U43590 (N_43590,N_38610,N_32866);
or U43591 (N_43591,N_32825,N_34847);
nand U43592 (N_43592,N_38178,N_31155);
nand U43593 (N_43593,N_33352,N_34945);
nor U43594 (N_43594,N_35351,N_35956);
or U43595 (N_43595,N_33403,N_32020);
nand U43596 (N_43596,N_37649,N_34973);
nor U43597 (N_43597,N_34794,N_36420);
or U43598 (N_43598,N_39638,N_37378);
nor U43599 (N_43599,N_38238,N_39729);
or U43600 (N_43600,N_39862,N_32298);
nand U43601 (N_43601,N_38706,N_33882);
nand U43602 (N_43602,N_35516,N_32264);
and U43603 (N_43603,N_35365,N_31439);
and U43604 (N_43604,N_38002,N_33969);
xnor U43605 (N_43605,N_36538,N_36469);
nor U43606 (N_43606,N_31903,N_35650);
nor U43607 (N_43607,N_38557,N_39485);
or U43608 (N_43608,N_31368,N_35514);
nand U43609 (N_43609,N_38098,N_39210);
or U43610 (N_43610,N_37445,N_33412);
nand U43611 (N_43611,N_37308,N_30326);
nand U43612 (N_43612,N_32608,N_38210);
nor U43613 (N_43613,N_30219,N_33809);
or U43614 (N_43614,N_36101,N_39932);
xor U43615 (N_43615,N_30215,N_39298);
nor U43616 (N_43616,N_34256,N_32846);
and U43617 (N_43617,N_35164,N_32868);
nor U43618 (N_43618,N_36552,N_38957);
nor U43619 (N_43619,N_30187,N_30277);
xor U43620 (N_43620,N_38767,N_34647);
and U43621 (N_43621,N_33984,N_38802);
or U43622 (N_43622,N_35942,N_37568);
and U43623 (N_43623,N_33480,N_33590);
xnor U43624 (N_43624,N_30386,N_38678);
nor U43625 (N_43625,N_39097,N_37500);
and U43626 (N_43626,N_39691,N_31829);
or U43627 (N_43627,N_31877,N_39637);
nor U43628 (N_43628,N_30793,N_33549);
xor U43629 (N_43629,N_33691,N_32086);
or U43630 (N_43630,N_37407,N_39024);
xnor U43631 (N_43631,N_33616,N_30823);
nor U43632 (N_43632,N_37511,N_31784);
xnor U43633 (N_43633,N_34676,N_32425);
nor U43634 (N_43634,N_39244,N_35269);
or U43635 (N_43635,N_39631,N_37865);
nand U43636 (N_43636,N_30995,N_30285);
xor U43637 (N_43637,N_39481,N_31736);
nor U43638 (N_43638,N_36293,N_35657);
nand U43639 (N_43639,N_35074,N_39178);
nand U43640 (N_43640,N_36566,N_35507);
and U43641 (N_43641,N_34623,N_35745);
or U43642 (N_43642,N_34042,N_31188);
and U43643 (N_43643,N_39488,N_39746);
and U43644 (N_43644,N_39556,N_34683);
or U43645 (N_43645,N_39472,N_35413);
xor U43646 (N_43646,N_33756,N_35026);
nand U43647 (N_43647,N_38513,N_32416);
and U43648 (N_43648,N_36078,N_36695);
and U43649 (N_43649,N_30897,N_33177);
xor U43650 (N_43650,N_31347,N_32672);
nand U43651 (N_43651,N_34925,N_32662);
nor U43652 (N_43652,N_34157,N_34174);
nand U43653 (N_43653,N_30302,N_34396);
nor U43654 (N_43654,N_37259,N_38039);
and U43655 (N_43655,N_36125,N_36406);
and U43656 (N_43656,N_36388,N_36867);
nor U43657 (N_43657,N_39413,N_33743);
and U43658 (N_43658,N_32294,N_30504);
or U43659 (N_43659,N_39406,N_33228);
nor U43660 (N_43660,N_39614,N_38786);
nand U43661 (N_43661,N_31548,N_30949);
nor U43662 (N_43662,N_32700,N_31160);
nand U43663 (N_43663,N_35461,N_30649);
and U43664 (N_43664,N_34744,N_39277);
and U43665 (N_43665,N_36268,N_35660);
or U43666 (N_43666,N_31799,N_39676);
xor U43667 (N_43667,N_36349,N_36058);
nand U43668 (N_43668,N_34011,N_34639);
nand U43669 (N_43669,N_34026,N_32586);
nor U43670 (N_43670,N_32993,N_30228);
nand U43671 (N_43671,N_32134,N_38715);
nor U43672 (N_43672,N_35594,N_34618);
and U43673 (N_43673,N_39798,N_32620);
nor U43674 (N_43674,N_30580,N_34144);
nor U43675 (N_43675,N_36617,N_37074);
nand U43676 (N_43676,N_34442,N_39695);
nor U43677 (N_43677,N_30920,N_36741);
nor U43678 (N_43678,N_37497,N_33512);
xor U43679 (N_43679,N_32542,N_35304);
xor U43680 (N_43680,N_32885,N_35785);
and U43681 (N_43681,N_33484,N_38688);
nor U43682 (N_43682,N_30356,N_38824);
nand U43683 (N_43683,N_31079,N_34056);
and U43684 (N_43684,N_38345,N_33465);
xor U43685 (N_43685,N_32265,N_36161);
and U43686 (N_43686,N_38651,N_34073);
nor U43687 (N_43687,N_32437,N_33284);
xor U43688 (N_43688,N_31098,N_30256);
nand U43689 (N_43689,N_35694,N_31381);
or U43690 (N_43690,N_31671,N_37715);
or U43691 (N_43691,N_34855,N_38698);
nand U43692 (N_43692,N_30894,N_36277);
and U43693 (N_43693,N_35111,N_30148);
nand U43694 (N_43694,N_38121,N_30514);
and U43695 (N_43695,N_36547,N_31593);
and U43696 (N_43696,N_33435,N_32289);
nand U43697 (N_43697,N_33255,N_36352);
nand U43698 (N_43698,N_39635,N_38354);
or U43699 (N_43699,N_34088,N_35901);
xor U43700 (N_43700,N_37160,N_34743);
nor U43701 (N_43701,N_38803,N_34569);
or U43702 (N_43702,N_36128,N_39728);
nand U43703 (N_43703,N_39749,N_33968);
or U43704 (N_43704,N_37890,N_30051);
nand U43705 (N_43705,N_36739,N_31525);
and U43706 (N_43706,N_34108,N_38127);
and U43707 (N_43707,N_35190,N_33517);
nor U43708 (N_43708,N_34086,N_35773);
nand U43709 (N_43709,N_36702,N_34279);
nand U43710 (N_43710,N_33370,N_32787);
and U43711 (N_43711,N_36167,N_38927);
or U43712 (N_43712,N_36767,N_34861);
and U43713 (N_43713,N_31304,N_34627);
or U43714 (N_43714,N_36517,N_38561);
and U43715 (N_43715,N_31059,N_39616);
nor U43716 (N_43716,N_33830,N_32899);
nor U43717 (N_43717,N_39736,N_37169);
nor U43718 (N_43718,N_31014,N_35503);
or U43719 (N_43719,N_30288,N_30911);
xor U43720 (N_43720,N_36143,N_31478);
xor U43721 (N_43721,N_36394,N_37364);
nor U43722 (N_43722,N_31437,N_31206);
or U43723 (N_43723,N_37760,N_30083);
nor U43724 (N_43724,N_38494,N_31862);
or U43725 (N_43725,N_35554,N_31044);
nand U43726 (N_43726,N_36127,N_38442);
and U43727 (N_43727,N_31145,N_38235);
nor U43728 (N_43728,N_30433,N_30681);
nor U43729 (N_43729,N_37904,N_32830);
xor U43730 (N_43730,N_39073,N_35842);
nand U43731 (N_43731,N_30833,N_34571);
nor U43732 (N_43732,N_34783,N_30278);
or U43733 (N_43733,N_39290,N_39586);
and U43734 (N_43734,N_36456,N_33693);
and U43735 (N_43735,N_37104,N_34663);
nand U43736 (N_43736,N_32483,N_30300);
nand U43737 (N_43737,N_34690,N_39494);
or U43738 (N_43738,N_36591,N_38171);
or U43739 (N_43739,N_31613,N_39457);
and U43740 (N_43740,N_30020,N_36863);
or U43741 (N_43741,N_30060,N_35744);
or U43742 (N_43742,N_39850,N_34113);
or U43743 (N_43743,N_31753,N_36969);
nand U43744 (N_43744,N_38158,N_34619);
nor U43745 (N_43745,N_31885,N_34159);
nand U43746 (N_43746,N_32533,N_36121);
nor U43747 (N_43747,N_37627,N_34033);
and U43748 (N_43748,N_36581,N_30406);
nand U43749 (N_43749,N_37276,N_33539);
and U43750 (N_43750,N_34065,N_37335);
nand U43751 (N_43751,N_35495,N_37024);
and U43752 (N_43752,N_31855,N_35262);
nor U43753 (N_43753,N_33289,N_32707);
and U43754 (N_43754,N_31503,N_34984);
nand U43755 (N_43755,N_37532,N_33451);
nand U43756 (N_43756,N_34960,N_35859);
nor U43757 (N_43757,N_31408,N_33189);
nor U43758 (N_43758,N_30455,N_32165);
and U43759 (N_43759,N_35949,N_34269);
nor U43760 (N_43760,N_33794,N_32641);
nor U43761 (N_43761,N_37059,N_34962);
or U43762 (N_43762,N_38549,N_33438);
nand U43763 (N_43763,N_35770,N_33431);
nor U43764 (N_43764,N_36241,N_34563);
and U43765 (N_43765,N_33934,N_32888);
nor U43766 (N_43766,N_33718,N_31415);
and U43767 (N_43767,N_39286,N_36721);
or U43768 (N_43768,N_30404,N_32651);
or U43769 (N_43769,N_32736,N_31794);
or U43770 (N_43770,N_33545,N_38197);
and U43771 (N_43771,N_38123,N_30712);
nor U43772 (N_43772,N_32889,N_33939);
xnor U43773 (N_43773,N_35555,N_38913);
nor U43774 (N_43774,N_30377,N_34604);
and U43775 (N_43775,N_36519,N_34153);
or U43776 (N_43776,N_30729,N_34827);
and U43777 (N_43777,N_33708,N_33582);
or U43778 (N_43778,N_36184,N_35059);
nand U43779 (N_43779,N_39813,N_33895);
nor U43780 (N_43780,N_38010,N_31064);
or U43781 (N_43781,N_36228,N_37878);
nand U43782 (N_43782,N_31722,N_31197);
nand U43783 (N_43783,N_37110,N_38619);
or U43784 (N_43784,N_30889,N_31400);
xor U43785 (N_43785,N_37654,N_39466);
nor U43786 (N_43786,N_30403,N_36780);
nand U43787 (N_43787,N_32758,N_35966);
nand U43788 (N_43788,N_37849,N_35970);
or U43789 (N_43789,N_33351,N_31375);
nand U43790 (N_43790,N_36734,N_35641);
or U43791 (N_43791,N_36529,N_31889);
or U43792 (N_43792,N_39120,N_38724);
nand U43793 (N_43793,N_31788,N_39807);
xnor U43794 (N_43794,N_38909,N_30776);
or U43795 (N_43795,N_34698,N_36012);
xnor U43796 (N_43796,N_35429,N_32686);
and U43797 (N_43797,N_36478,N_38180);
nor U43798 (N_43798,N_35331,N_34315);
nor U43799 (N_43799,N_35222,N_39619);
nor U43800 (N_43800,N_36304,N_32961);
nand U43801 (N_43801,N_32328,N_33196);
nand U43802 (N_43802,N_39145,N_31994);
xnor U43803 (N_43803,N_30955,N_36998);
nor U43804 (N_43804,N_37077,N_33001);
nor U43805 (N_43805,N_30155,N_32799);
xor U43806 (N_43806,N_36457,N_32873);
or U43807 (N_43807,N_31815,N_39525);
or U43808 (N_43808,N_39509,N_37846);
or U43809 (N_43809,N_37572,N_33461);
and U43810 (N_43810,N_30768,N_34185);
nor U43811 (N_43811,N_34466,N_36175);
or U43812 (N_43812,N_36602,N_35393);
and U43813 (N_43813,N_34275,N_38543);
nand U43814 (N_43814,N_34765,N_36413);
xor U43815 (N_43815,N_39703,N_35522);
nor U43816 (N_43816,N_34964,N_39008);
xor U43817 (N_43817,N_31000,N_32233);
nand U43818 (N_43818,N_30631,N_38207);
or U43819 (N_43819,N_38478,N_37307);
nand U43820 (N_43820,N_32250,N_37931);
nand U43821 (N_43821,N_36629,N_32062);
nand U43822 (N_43822,N_35002,N_31169);
and U43823 (N_43823,N_37557,N_38269);
xnor U43824 (N_43824,N_30694,N_39828);
nand U43825 (N_43825,N_38992,N_33179);
or U43826 (N_43826,N_34907,N_36562);
or U43827 (N_43827,N_32789,N_34629);
nor U43828 (N_43828,N_36812,N_34221);
nand U43829 (N_43829,N_36325,N_37379);
nor U43830 (N_43830,N_37751,N_34727);
nor U43831 (N_43831,N_30110,N_33459);
and U43832 (N_43832,N_34047,N_32160);
nor U43833 (N_43833,N_30534,N_33775);
and U43834 (N_43834,N_31937,N_37590);
nand U43835 (N_43835,N_33888,N_39902);
or U43836 (N_43836,N_32456,N_38692);
nor U43837 (N_43837,N_38367,N_30214);
or U43838 (N_43838,N_37650,N_39063);
nor U43839 (N_43839,N_39237,N_34384);
nor U43840 (N_43840,N_36230,N_36823);
and U43841 (N_43841,N_34882,N_33334);
nand U43842 (N_43842,N_33991,N_37078);
xor U43843 (N_43843,N_35869,N_39279);
nor U43844 (N_43844,N_36256,N_35405);
and U43845 (N_43845,N_30028,N_30063);
or U43846 (N_43846,N_32193,N_30938);
or U43847 (N_43847,N_32234,N_30800);
nor U43848 (N_43848,N_36485,N_38012);
or U43849 (N_43849,N_30193,N_36885);
nand U43850 (N_43850,N_31353,N_35948);
nor U43851 (N_43851,N_32673,N_39779);
nand U43852 (N_43852,N_30102,N_39428);
or U43853 (N_43853,N_38083,N_36014);
and U43854 (N_43854,N_35439,N_38496);
or U43855 (N_43855,N_37007,N_38639);
nor U43856 (N_43856,N_35576,N_37437);
nand U43857 (N_43857,N_31013,N_37577);
nand U43858 (N_43858,N_34977,N_38638);
nand U43859 (N_43859,N_30479,N_34212);
nor U43860 (N_43860,N_35980,N_34760);
nand U43861 (N_43861,N_36693,N_32898);
or U43862 (N_43862,N_38325,N_37540);
nor U43863 (N_43863,N_31240,N_33686);
xnor U43864 (N_43864,N_31708,N_36144);
nand U43865 (N_43865,N_38183,N_36850);
xnor U43866 (N_43866,N_30308,N_31497);
nor U43867 (N_43867,N_39179,N_35142);
and U43868 (N_43868,N_39553,N_31748);
and U43869 (N_43869,N_30305,N_33508);
nand U43870 (N_43870,N_35284,N_34544);
nand U43871 (N_43871,N_37520,N_36353);
nor U43872 (N_43872,N_33349,N_35166);
nor U43873 (N_43873,N_31601,N_30127);
or U43874 (N_43874,N_38028,N_36831);
and U43875 (N_43875,N_39319,N_33240);
nand U43876 (N_43876,N_32783,N_33063);
or U43877 (N_43877,N_35080,N_39306);
and U43878 (N_43878,N_30463,N_34093);
and U43879 (N_43879,N_35685,N_33831);
nand U43880 (N_43880,N_38185,N_39758);
nor U43881 (N_43881,N_39566,N_38701);
and U43882 (N_43882,N_31933,N_39761);
or U43883 (N_43883,N_31629,N_39423);
nand U43884 (N_43884,N_35447,N_32337);
and U43885 (N_43885,N_36698,N_38607);
and U43886 (N_43886,N_32151,N_38797);
nand U43887 (N_43887,N_39990,N_38447);
nand U43888 (N_43888,N_32747,N_32526);
xnor U43889 (N_43889,N_33155,N_37605);
and U43890 (N_43890,N_33850,N_33663);
and U43891 (N_43891,N_35559,N_32812);
nor U43892 (N_43892,N_30706,N_36736);
or U43893 (N_43893,N_33229,N_30686);
or U43894 (N_43894,N_33997,N_30169);
nor U43895 (N_43895,N_32302,N_31598);
and U43896 (N_43896,N_38544,N_39661);
or U43897 (N_43897,N_34236,N_36266);
or U43898 (N_43898,N_30093,N_38926);
and U43899 (N_43899,N_37266,N_31962);
nor U43900 (N_43900,N_32895,N_36890);
nand U43901 (N_43901,N_31442,N_38615);
and U43902 (N_43902,N_37043,N_32274);
nor U43903 (N_43903,N_32566,N_31512);
or U43904 (N_43904,N_30323,N_37177);
xnor U43905 (N_43905,N_34234,N_39006);
nor U43906 (N_43906,N_30850,N_39768);
and U43907 (N_43907,N_31961,N_30281);
xnor U43908 (N_43908,N_37809,N_38903);
nand U43909 (N_43909,N_39187,N_37769);
nand U43910 (N_43910,N_31255,N_30907);
nand U43911 (N_43911,N_38703,N_34250);
nor U43912 (N_43912,N_33208,N_30936);
and U43913 (N_43913,N_34281,N_32511);
or U43914 (N_43914,N_31264,N_38205);
and U43915 (N_43915,N_34983,N_35829);
and U43916 (N_43916,N_37512,N_35209);
nor U43917 (N_43917,N_32531,N_32245);
nand U43918 (N_43918,N_36992,N_37528);
nand U43919 (N_43919,N_30709,N_33554);
nand U43920 (N_43920,N_37607,N_33717);
nor U43921 (N_43921,N_35588,N_36645);
and U43922 (N_43922,N_36151,N_31872);
nor U43923 (N_43923,N_37863,N_31025);
and U43924 (N_43924,N_31003,N_39095);
nand U43925 (N_43925,N_38109,N_33815);
or U43926 (N_43926,N_39541,N_36733);
and U43927 (N_43927,N_36487,N_32440);
nand U43928 (N_43928,N_33647,N_30265);
and U43929 (N_43929,N_36403,N_38762);
nor U43930 (N_43930,N_32025,N_39271);
and U43931 (N_43931,N_34202,N_32379);
and U43932 (N_43932,N_31545,N_32318);
nand U43933 (N_43933,N_35646,N_33654);
and U43934 (N_43934,N_33023,N_35291);
nor U43935 (N_43935,N_38545,N_31529);
or U43936 (N_43936,N_38094,N_33466);
xor U43937 (N_43937,N_34165,N_39415);
and U43938 (N_43938,N_35689,N_37265);
or U43939 (N_43939,N_32136,N_38876);
or U43940 (N_43940,N_30461,N_35064);
nand U43941 (N_43941,N_35515,N_30544);
nand U43942 (N_43942,N_32319,N_33634);
and U43943 (N_43943,N_32634,N_31986);
or U43944 (N_43944,N_33808,N_34790);
and U43945 (N_43945,N_37460,N_36676);
nor U43946 (N_43946,N_39621,N_39026);
and U43947 (N_43947,N_38311,N_36511);
and U43948 (N_43948,N_36160,N_36290);
xor U43949 (N_43949,N_38484,N_30980);
or U43950 (N_43950,N_31803,N_35709);
nor U43951 (N_43951,N_31866,N_39573);
or U43952 (N_43952,N_31181,N_39342);
nor U43953 (N_43953,N_36746,N_31560);
nand U43954 (N_43954,N_37933,N_34503);
nand U43955 (N_43955,N_30301,N_35256);
or U43956 (N_43956,N_35381,N_35936);
and U43957 (N_43957,N_35039,N_37664);
nor U43958 (N_43958,N_37629,N_32197);
nor U43959 (N_43959,N_31392,N_39610);
and U43960 (N_43960,N_35345,N_37724);
nor U43961 (N_43961,N_34818,N_31156);
and U43962 (N_43962,N_34711,N_32880);
nor U43963 (N_43963,N_36400,N_30008);
xor U43964 (N_43964,N_38606,N_33981);
nand U43965 (N_43965,N_39855,N_33631);
nand U43966 (N_43966,N_38653,N_38020);
or U43967 (N_43967,N_33583,N_37488);
and U43968 (N_43968,N_36756,N_33365);
nand U43969 (N_43969,N_38413,N_32610);
and U43970 (N_43970,N_39818,N_31138);
or U43971 (N_43971,N_34860,N_39224);
or U43972 (N_43972,N_34574,N_30972);
nand U43973 (N_43973,N_32324,N_32333);
or U43974 (N_43974,N_34923,N_37978);
xor U43975 (N_43975,N_30622,N_33681);
or U43976 (N_43976,N_34237,N_30963);
and U43977 (N_43977,N_39778,N_38621);
and U43978 (N_43978,N_35024,N_37433);
nand U43979 (N_43979,N_34887,N_36763);
nand U43980 (N_43980,N_31945,N_34137);
nor U43981 (N_43981,N_36798,N_33125);
nor U43982 (N_43982,N_33748,N_33195);
nand U43983 (N_43983,N_38049,N_38923);
nand U43984 (N_43984,N_30592,N_33462);
nor U43985 (N_43985,N_37529,N_31745);
nand U43986 (N_43986,N_34443,N_36606);
and U43987 (N_43987,N_39589,N_32990);
nand U43988 (N_43988,N_34190,N_35811);
or U43989 (N_43989,N_37099,N_34821);
and U43990 (N_43990,N_36240,N_33486);
or U43991 (N_43991,N_37365,N_34548);
nor U43992 (N_43992,N_37993,N_39247);
or U43993 (N_43993,N_33065,N_36084);
or U43994 (N_43994,N_38196,N_36579);
and U43995 (N_43995,N_38406,N_37108);
nand U43996 (N_43996,N_38184,N_31920);
and U43997 (N_43997,N_39154,N_30385);
and U43998 (N_43998,N_32012,N_34453);
or U43999 (N_43999,N_31458,N_38486);
and U44000 (N_44000,N_33188,N_35855);
xnor U44001 (N_44001,N_36565,N_32730);
or U44002 (N_44002,N_38004,N_34146);
nor U44003 (N_44003,N_30976,N_36455);
nand U44004 (N_44004,N_33651,N_38697);
nand U44005 (N_44005,N_32065,N_31835);
nand U44006 (N_44006,N_38151,N_33994);
and U44007 (N_44007,N_34458,N_32031);
or U44008 (N_44008,N_31501,N_39242);
nand U44009 (N_44009,N_33269,N_32684);
or U44010 (N_44010,N_33943,N_37510);
or U44011 (N_44011,N_38188,N_32693);
or U44012 (N_44012,N_31850,N_34060);
or U44013 (N_44013,N_38135,N_39547);
nor U44014 (N_44014,N_38931,N_36212);
and U44015 (N_44015,N_39792,N_36662);
nand U44016 (N_44016,N_37669,N_33844);
or U44017 (N_44017,N_36208,N_35666);
or U44018 (N_44018,N_38361,N_36274);
nor U44019 (N_44019,N_38821,N_34420);
nor U44020 (N_44020,N_34246,N_36673);
nand U44021 (N_44021,N_34255,N_38348);
or U44022 (N_44022,N_38025,N_38906);
nor U44023 (N_44023,N_38107,N_35782);
or U44024 (N_44024,N_35103,N_34139);
nand U44025 (N_44025,N_31130,N_38474);
and U44026 (N_44026,N_37415,N_36063);
nor U44027 (N_44027,N_39185,N_39975);
nand U44028 (N_44028,N_37254,N_34774);
nand U44029 (N_44029,N_35219,N_33560);
nor U44030 (N_44030,N_34422,N_36790);
and U44031 (N_44031,N_35691,N_38264);
nor U44032 (N_44032,N_31677,N_30399);
and U44033 (N_44033,N_31216,N_30439);
nor U44034 (N_44034,N_32004,N_37903);
nor U44035 (N_44035,N_30815,N_39105);
and U44036 (N_44036,N_32779,N_37727);
nand U44037 (N_44037,N_34966,N_38851);
and U44038 (N_44038,N_36906,N_39537);
and U44039 (N_44039,N_33992,N_36068);
and U44040 (N_44040,N_32618,N_32144);
xor U44041 (N_44041,N_36510,N_33025);
or U44042 (N_44042,N_39836,N_33054);
nand U44043 (N_44043,N_31448,N_34161);
or U44044 (N_44044,N_35368,N_31317);
or U44045 (N_44045,N_39463,N_38811);
or U44046 (N_44046,N_39942,N_36677);
or U44047 (N_44047,N_31519,N_32124);
or U44048 (N_44048,N_34809,N_32260);
or U44049 (N_44049,N_37049,N_37828);
and U44050 (N_44050,N_30584,N_33437);
nor U44051 (N_44051,N_37106,N_30515);
xor U44052 (N_44052,N_33661,N_30001);
and U44053 (N_44053,N_35809,N_39874);
nand U44054 (N_44054,N_37977,N_33152);
nor U44055 (N_44055,N_32357,N_39370);
and U44056 (N_44056,N_35971,N_31419);
nor U44057 (N_44057,N_30367,N_37103);
nand U44058 (N_44058,N_37795,N_37469);
nand U44059 (N_44059,N_35387,N_35573);
or U44060 (N_44060,N_37914,N_36692);
nor U44061 (N_44061,N_31632,N_31851);
or U44062 (N_44062,N_39359,N_38149);
nand U44063 (N_44063,N_37877,N_31790);
or U44064 (N_44064,N_31626,N_39987);
nand U44065 (N_44065,N_39047,N_33401);
or U44066 (N_44066,N_36426,N_37121);
and U44067 (N_44067,N_32420,N_30418);
or U44068 (N_44068,N_38989,N_38566);
xor U44069 (N_44069,N_32666,N_30106);
nand U44070 (N_44070,N_33848,N_30168);
nor U44071 (N_44071,N_31461,N_39023);
xor U44072 (N_44072,N_31331,N_34304);
xnor U44073 (N_44073,N_32882,N_30047);
and U44074 (N_44074,N_32791,N_32155);
and U44075 (N_44075,N_39133,N_36806);
nand U44076 (N_44076,N_34890,N_32733);
nor U44077 (N_44077,N_38126,N_32247);
nor U44078 (N_44078,N_31243,N_37327);
nor U44079 (N_44079,N_31286,N_37032);
and U44080 (N_44080,N_35551,N_30798);
and U44081 (N_44081,N_37815,N_36914);
and U44082 (N_44082,N_30258,N_34004);
and U44083 (N_44083,N_35950,N_38763);
nand U44084 (N_44084,N_33355,N_39615);
or U44085 (N_44085,N_34919,N_32255);
and U44086 (N_44086,N_36126,N_34482);
or U44087 (N_44087,N_38689,N_36925);
and U44088 (N_44088,N_32523,N_38555);
xnor U44089 (N_44089,N_31518,N_38720);
and U44090 (N_44090,N_37343,N_39018);
nor U44091 (N_44091,N_33729,N_31581);
or U44092 (N_44092,N_39936,N_35605);
nand U44093 (N_44093,N_33563,N_33330);
and U44094 (N_44094,N_36052,N_31740);
nor U44095 (N_44095,N_38339,N_33689);
nand U44096 (N_44096,N_37839,N_34106);
nor U44097 (N_44097,N_37856,N_36899);
or U44098 (N_44098,N_36210,N_31041);
nor U44099 (N_44099,N_32305,N_36611);
and U44100 (N_44100,N_39102,N_30583);
nand U44101 (N_44101,N_30236,N_30478);
nor U44102 (N_44102,N_35234,N_32854);
or U44103 (N_44103,N_30114,N_34540);
or U44104 (N_44104,N_34438,N_31280);
and U44105 (N_44105,N_37258,N_34560);
nor U44106 (N_44106,N_30971,N_39584);
nand U44107 (N_44107,N_33841,N_38211);
nor U44108 (N_44108,N_36433,N_35281);
or U44109 (N_44109,N_38995,N_30578);
xnor U44110 (N_44110,N_36896,N_35283);
and U44111 (N_44111,N_36067,N_35695);
and U44112 (N_44112,N_31944,N_34514);
nand U44113 (N_44113,N_31742,N_38399);
nand U44114 (N_44114,N_31017,N_33242);
nor U44115 (N_44115,N_34801,N_32494);
nand U44116 (N_44116,N_39904,N_31810);
nor U44117 (N_44117,N_31095,N_32041);
or U44118 (N_44118,N_36991,N_35781);
nor U44119 (N_44119,N_39500,N_30530);
and U44120 (N_44120,N_39371,N_37682);
nor U44121 (N_44121,N_31854,N_35044);
or U44122 (N_44122,N_35567,N_34504);
nand U44123 (N_44123,N_38937,N_37235);
and U44124 (N_44124,N_39380,N_33922);
and U44125 (N_44125,N_33078,N_36471);
xor U44126 (N_44126,N_36477,N_35925);
nor U44127 (N_44127,N_33531,N_30493);
nor U44128 (N_44128,N_39459,N_31633);
nand U44129 (N_44129,N_33913,N_35330);
nor U44130 (N_44130,N_32301,N_38721);
xor U44131 (N_44131,N_33747,N_35434);
nand U44132 (N_44132,N_38461,N_38318);
and U44133 (N_44133,N_31426,N_35828);
nand U44134 (N_44134,N_33675,N_33248);
nor U44135 (N_44135,N_37585,N_32383);
nand U44136 (N_44136,N_36818,N_35473);
or U44137 (N_44137,N_36881,N_37549);
nor U44138 (N_44138,N_33280,N_36334);
or U44139 (N_44139,N_38117,N_35100);
xnor U44140 (N_44140,N_34498,N_33141);
nor U44141 (N_44141,N_39115,N_35085);
nand U44142 (N_44142,N_33362,N_33350);
xor U44143 (N_44143,N_35355,N_34685);
nor U44144 (N_44144,N_35072,N_39360);
and U44145 (N_44145,N_31719,N_38295);
nand U44146 (N_44146,N_30450,N_30926);
and U44147 (N_44147,N_37985,N_32926);
nor U44148 (N_44148,N_34216,N_35323);
nand U44149 (N_44149,N_31108,N_39590);
and U44150 (N_44150,N_30026,N_37984);
or U44151 (N_44151,N_39250,N_31109);
and U44152 (N_44152,N_38299,N_39211);
xnor U44153 (N_44153,N_34645,N_39617);
nor U44154 (N_44154,N_39801,N_33603);
xnor U44155 (N_44155,N_38326,N_36917);
xnor U44156 (N_44156,N_31567,N_36399);
nand U44157 (N_44157,N_34598,N_39926);
nor U44158 (N_44158,N_35201,N_31423);
or U44159 (N_44159,N_38807,N_31514);
nand U44160 (N_44160,N_32503,N_31750);
nand U44161 (N_44161,N_30279,N_37396);
and U44162 (N_44162,N_35356,N_30198);
nor U44163 (N_44163,N_34845,N_38298);
or U44164 (N_44164,N_31848,N_34184);
or U44165 (N_44165,N_33536,N_39645);
xor U44166 (N_44166,N_39239,N_38502);
or U44167 (N_44167,N_33883,N_37538);
or U44168 (N_44168,N_30437,N_32129);
nor U44169 (N_44169,N_33596,N_34434);
nand U44170 (N_44170,N_35458,N_34014);
or U44171 (N_44171,N_34359,N_33551);
nand U44172 (N_44172,N_36858,N_37998);
or U44173 (N_44173,N_36497,N_36528);
or U44174 (N_44174,N_34019,N_34562);
or U44175 (N_44175,N_30274,N_36918);
and U44176 (N_44176,N_32725,N_36116);
and U44177 (N_44177,N_39473,N_33291);
or U44178 (N_44178,N_31337,N_30097);
xor U44179 (N_44179,N_39225,N_31399);
or U44180 (N_44180,N_36489,N_35178);
or U44181 (N_44181,N_36793,N_31281);
xnor U44182 (N_44182,N_38035,N_38393);
or U44183 (N_44183,N_36765,N_35267);
and U44184 (N_44184,N_37713,N_37055);
or U44185 (N_44185,N_31234,N_39088);
or U44186 (N_44186,N_38267,N_38009);
nor U44187 (N_44187,N_35619,N_30593);
nand U44188 (N_44188,N_34240,N_38430);
or U44189 (N_44189,N_36964,N_35739);
nor U44190 (N_44190,N_39655,N_33924);
nand U44191 (N_44191,N_37173,N_30086);
xor U44192 (N_44192,N_36879,N_31058);
xor U44193 (N_44193,N_37891,N_36466);
nor U44194 (N_44194,N_38884,N_32867);
nor U44195 (N_44195,N_34614,N_33974);
nand U44196 (N_44196,N_34892,N_37485);
nand U44197 (N_44197,N_35092,N_32293);
nor U44198 (N_44198,N_35029,N_31193);
nor U44199 (N_44199,N_34492,N_35385);
and U44200 (N_44200,N_33618,N_36974);
and U44201 (N_44201,N_31460,N_38953);
nand U44202 (N_44202,N_36391,N_36322);
or U44203 (N_44203,N_35202,N_39207);
nand U44204 (N_44204,N_36610,N_35598);
and U44205 (N_44205,N_31288,N_37053);
or U44206 (N_44206,N_37521,N_31322);
and U44207 (N_44207,N_39447,N_35407);
nand U44208 (N_44208,N_30927,N_36835);
nor U44209 (N_44209,N_32067,N_30954);
and U44210 (N_44210,N_37083,N_32320);
nand U44211 (N_44211,N_36502,N_32822);
xor U44212 (N_44212,N_30333,N_38467);
or U44213 (N_44213,N_34638,N_30177);
and U44214 (N_44214,N_33938,N_30395);
nor U44215 (N_44215,N_30642,N_34793);
nand U44216 (N_44216,N_31958,N_33581);
and U44217 (N_44217,N_36445,N_30470);
and U44218 (N_44218,N_35788,N_38915);
nand U44219 (N_44219,N_32781,N_32374);
and U44220 (N_44220,N_32905,N_37464);
nor U44221 (N_44221,N_33773,N_33276);
and U44222 (N_44222,N_35749,N_39715);
nor U44223 (N_44223,N_32354,N_36138);
or U44224 (N_44224,N_38498,N_38735);
and U44225 (N_44225,N_37211,N_35877);
or U44226 (N_44226,N_31142,N_30331);
nor U44227 (N_44227,N_35226,N_31285);
and U44228 (N_44228,N_38422,N_35148);
nor U44229 (N_44229,N_35257,N_39967);
and U44230 (N_44230,N_37820,N_34059);
or U44231 (N_44231,N_33014,N_33557);
and U44232 (N_44232,N_39272,N_30528);
or U44233 (N_44233,N_38601,N_30048);
or U44234 (N_44234,N_34124,N_33901);
xor U44235 (N_44235,N_30501,N_30691);
and U44236 (N_44236,N_34520,N_38846);
or U44237 (N_44237,N_30506,N_36308);
and U44238 (N_44238,N_30970,N_37786);
nor U44239 (N_44239,N_34703,N_34889);
or U44240 (N_44240,N_30991,N_31559);
or U44241 (N_44241,N_39112,N_38974);
or U44242 (N_44242,N_31665,N_30269);
and U44243 (N_44243,N_33653,N_35627);
nand U44244 (N_44244,N_33587,N_33559);
or U44245 (N_44245,N_33305,N_35545);
nand U44246 (N_44246,N_32991,N_38027);
nand U44247 (N_44247,N_37311,N_39345);
and U44248 (N_44248,N_38829,N_31287);
and U44249 (N_44249,N_35848,N_37161);
nor U44250 (N_44250,N_35822,N_34572);
nor U44251 (N_44251,N_32919,N_32948);
and U44252 (N_44252,N_39395,N_30650);
and U44253 (N_44253,N_34265,N_30359);
nor U44254 (N_44254,N_38901,N_33905);
nor U44255 (N_44255,N_37706,N_38156);
or U44256 (N_44256,N_34853,N_36301);
nand U44257 (N_44257,N_39907,N_34457);
and U44258 (N_44258,N_39731,N_31869);
xor U44259 (N_44259,N_32156,N_37825);
nand U44260 (N_44260,N_31445,N_34455);
or U44261 (N_44261,N_33035,N_32021);
or U44262 (N_44262,N_30818,N_35716);
and U44263 (N_44263,N_36986,N_35537);
or U44264 (N_44264,N_35244,N_38445);
xor U44265 (N_44265,N_35690,N_30732);
nand U44266 (N_44266,N_32602,N_30715);
or U44267 (N_44267,N_37000,N_37195);
and U44268 (N_44268,N_37434,N_33212);
nor U44269 (N_44269,N_30656,N_33205);
or U44270 (N_44270,N_35208,N_35830);
or U44271 (N_44271,N_31170,N_35717);
or U44272 (N_44272,N_37370,N_30677);
or U44273 (N_44273,N_31618,N_37033);
xnor U44274 (N_44274,N_38155,N_35093);
nand U44275 (N_44275,N_35592,N_39475);
or U44276 (N_44276,N_30357,N_36281);
nor U44277 (N_44277,N_37238,N_34653);
nor U44278 (N_44278,N_31516,N_39910);
nand U44279 (N_44279,N_38731,N_34921);
and U44280 (N_44280,N_37691,N_37644);
xor U44281 (N_44281,N_31088,N_39557);
or U44282 (N_44282,N_39132,N_33623);
or U44283 (N_44283,N_37886,N_35159);
nand U44284 (N_44284,N_39922,N_34150);
nand U44285 (N_44285,N_34975,N_31340);
and U44286 (N_44286,N_35959,N_35697);
nor U44287 (N_44287,N_30852,N_38667);
nand U44288 (N_44288,N_31414,N_34207);
and U44289 (N_44289,N_36288,N_36134);
nand U44290 (N_44290,N_39811,N_30039);
and U44291 (N_44291,N_34057,N_37875);
nand U44292 (N_44292,N_33293,N_38641);
nor U44293 (N_44293,N_36797,N_32965);
nor U44294 (N_44294,N_33121,N_36156);
nand U44295 (N_44295,N_31645,N_37927);
nand U44296 (N_44296,N_39361,N_34903);
nand U44297 (N_44297,N_31344,N_35994);
nand U44298 (N_44298,N_36747,N_31953);
or U44299 (N_44299,N_35846,N_38723);
or U44300 (N_44300,N_37547,N_30814);
xnor U44301 (N_44301,N_32362,N_31077);
nor U44302 (N_44302,N_32966,N_32833);
and U44303 (N_44303,N_37283,N_34143);
and U44304 (N_44304,N_34652,N_33426);
and U44305 (N_44305,N_34617,N_30272);
nand U44306 (N_44306,N_33947,N_31049);
and U44307 (N_44307,N_32534,N_39529);
or U44308 (N_44308,N_37647,N_32749);
and U44309 (N_44309,N_35713,N_37767);
or U44310 (N_44310,N_32903,N_38203);
or U44311 (N_44311,N_37489,N_39569);
xnor U44312 (N_44312,N_30142,N_36574);
xor U44313 (N_44313,N_34192,N_37380);
nand U44314 (N_44314,N_39604,N_37134);
nor U44315 (N_44315,N_35046,N_30529);
nand U44316 (N_44316,N_34203,N_35911);
or U44317 (N_44317,N_39238,N_34395);
nor U44318 (N_44318,N_36612,N_39518);
nand U44319 (N_44319,N_32697,N_35020);
or U44320 (N_44320,N_39945,N_38840);
nor U44321 (N_44321,N_36575,N_32579);
and U44322 (N_44322,N_38453,N_39134);
and U44323 (N_44323,N_31152,N_30838);
xnor U44324 (N_44324,N_37293,N_38061);
or U44325 (N_44325,N_31183,N_38334);
or U44326 (N_44326,N_36679,N_34201);
and U44327 (N_44327,N_30158,N_37157);
or U44328 (N_44328,N_33273,N_34748);
and U44329 (N_44329,N_31819,N_30314);
and U44330 (N_44330,N_38997,N_38360);
or U44331 (N_44331,N_38605,N_36108);
nand U44332 (N_44332,N_35978,N_38148);
and U44333 (N_44333,N_35199,N_33982);
xnor U44334 (N_44334,N_31020,N_32340);
nand U44335 (N_44335,N_30445,N_39963);
and U44336 (N_44336,N_35122,N_34366);
and U44337 (N_44337,N_31222,N_36309);
nand U44338 (N_44338,N_34167,N_31905);
nand U44339 (N_44339,N_31679,N_37427);
or U44340 (N_44340,N_37812,N_35895);
nand U44341 (N_44341,N_32164,N_34172);
nand U44342 (N_44342,N_35170,N_33066);
nand U44343 (N_44343,N_33381,N_38626);
nand U44344 (N_44344,N_38497,N_38268);
and U44345 (N_44345,N_34427,N_39722);
nand U44346 (N_44346,N_34677,N_32492);
or U44347 (N_44347,N_33005,N_33621);
nand U44348 (N_44348,N_33341,N_33216);
xnor U44349 (N_44349,N_34849,N_30723);
or U44350 (N_44350,N_38208,N_31689);
or U44351 (N_44351,N_32269,N_39338);
or U44352 (N_44352,N_38048,N_36936);
nor U44353 (N_44353,N_32982,N_31542);
nand U44354 (N_44354,N_36895,N_34626);
or U44355 (N_44355,N_39934,N_34773);
nand U44356 (N_44356,N_35008,N_39362);
and U44357 (N_44357,N_34008,N_34759);
xor U44358 (N_44358,N_34739,N_35963);
and U44359 (N_44359,N_33230,N_37406);
or U44360 (N_44360,N_35451,N_39144);
nor U44361 (N_44361,N_38694,N_35613);
nor U44362 (N_44362,N_39928,N_34483);
and U44363 (N_44363,N_35547,N_33505);
nor U44364 (N_44364,N_30510,N_32861);
nor U44365 (N_44365,N_38589,N_31175);
nor U44366 (N_44366,N_37089,N_35313);
nor U44367 (N_44367,N_34555,N_30538);
or U44368 (N_44368,N_35319,N_36875);
nor U44369 (N_44369,N_30637,N_39013);
nor U44370 (N_44370,N_39364,N_30870);
xnor U44371 (N_44371,N_32321,N_38274);
or U44372 (N_44372,N_35144,N_39436);
nand U44373 (N_44373,N_38579,N_31975);
or U44374 (N_44374,N_35218,N_37788);
and U44375 (N_44375,N_38796,N_37906);
and U44376 (N_44376,N_39192,N_31541);
xor U44377 (N_44377,N_38425,N_35726);
xnor U44378 (N_44378,N_34166,N_39918);
or U44379 (N_44379,N_37170,N_32540);
nor U44380 (N_44380,N_38257,N_35023);
or U44381 (N_44381,N_33917,N_30317);
nand U44382 (N_44382,N_34034,N_32630);
nand U44383 (N_44383,N_33711,N_33542);
nor U44384 (N_44384,N_39456,N_35227);
and U44385 (N_44385,N_35721,N_35902);
nor U44386 (N_44386,N_34756,N_39149);
nor U44387 (N_44387,N_35617,N_38302);
xor U44388 (N_44388,N_34206,N_38739);
xnor U44389 (N_44389,N_33856,N_36177);
or U44390 (N_44390,N_38215,N_32609);
nand U44391 (N_44391,N_32676,N_36176);
nand U44392 (N_44392,N_37796,N_39680);
nand U44393 (N_44393,N_35851,N_36596);
nor U44394 (N_44394,N_31789,N_31642);
nor U44395 (N_44395,N_31977,N_39773);
nand U44396 (N_44396,N_35645,N_35832);
nand U44397 (N_44397,N_32986,N_39284);
nand U44398 (N_44398,N_39397,N_37071);
or U44399 (N_44399,N_31248,N_35295);
and U44400 (N_44400,N_37758,N_33488);
and U44401 (N_44401,N_31664,N_38191);
nand U44402 (N_44402,N_35992,N_32477);
nand U44403 (N_44403,N_31187,N_35232);
nand U44404 (N_44404,N_39431,N_37260);
nand U44405 (N_44405,N_32472,N_31531);
or U44406 (N_44406,N_35261,N_31563);
and U44407 (N_44407,N_31811,N_31192);
and U44408 (N_44408,N_38642,N_30371);
nor U44409 (N_44409,N_31499,N_39892);
or U44410 (N_44410,N_38842,N_35511);
or U44411 (N_44411,N_35009,N_34474);
nand U44412 (N_44412,N_31576,N_37021);
nand U44413 (N_44413,N_30684,N_38429);
and U44414 (N_44414,N_34837,N_35004);
and U44415 (N_44415,N_35999,N_34836);
nand U44416 (N_44416,N_35972,N_35962);
and U44417 (N_44417,N_34828,N_38280);
nor U44418 (N_44418,N_30594,N_37747);
and U44419 (N_44419,N_39765,N_30855);
and U44420 (N_44420,N_32550,N_36493);
or U44421 (N_44421,N_36508,N_32113);
xor U44422 (N_44422,N_33180,N_32058);
nand U44423 (N_44423,N_38244,N_38899);
or U44424 (N_44424,N_37070,N_33019);
and U44425 (N_44425,N_32487,N_34657);
xnor U44426 (N_44426,N_35596,N_38584);
nor U44427 (N_44427,N_35724,N_30165);
or U44428 (N_44428,N_34038,N_39788);
nand U44429 (N_44429,N_30347,N_32554);
or U44430 (N_44430,N_33483,N_35896);
or U44431 (N_44431,N_35520,N_30568);
nand U44432 (N_44432,N_39885,N_37746);
nand U44433 (N_44433,N_35031,N_30945);
and U44434 (N_44434,N_34968,N_34858);
nor U44435 (N_44435,N_38632,N_34082);
nor U44436 (N_44436,N_39911,N_39301);
or U44437 (N_44437,N_39007,N_37098);
and U44438 (N_44438,N_38999,N_36541);
and U44439 (N_44439,N_38364,N_35187);
nand U44440 (N_44440,N_32137,N_37300);
nand U44441 (N_44441,N_35815,N_37583);
and U44442 (N_44442,N_35746,N_33359);
and U44443 (N_44443,N_37787,N_31868);
and U44444 (N_44444,N_36877,N_36350);
nand U44445 (N_44445,N_36560,N_35735);
or U44446 (N_44446,N_35133,N_35813);
nand U44447 (N_44447,N_33762,N_35849);
and U44448 (N_44448,N_30062,N_39757);
nor U44449 (N_44449,N_32463,N_32313);
xnor U44450 (N_44450,N_30221,N_33575);
and U44451 (N_44451,N_37789,N_30073);
or U44452 (N_44452,N_34565,N_39337);
or U44453 (N_44453,N_37525,N_32710);
nor U44454 (N_44454,N_38245,N_38023);
nand U44455 (N_44455,N_35138,N_35928);
and U44456 (N_44456,N_35150,N_31622);
or U44457 (N_44457,N_31474,N_35348);
and U44458 (N_44458,N_35048,N_32036);
or U44459 (N_44459,N_30349,N_38003);
and U44460 (N_44460,N_36043,N_35206);
nand U44461 (N_44461,N_30295,N_37287);
xor U44462 (N_44462,N_33347,N_34308);
xor U44463 (N_44463,N_34089,N_32621);
nand U44464 (N_44464,N_37905,N_39929);
xnor U44465 (N_44465,N_37454,N_39896);
nor U44466 (N_44466,N_33728,N_36339);
or U44467 (N_44467,N_38613,N_39079);
nor U44468 (N_44468,N_33846,N_32619);
xnor U44469 (N_44469,N_32110,N_38108);
or U44470 (N_44470,N_31257,N_34045);
or U44471 (N_44471,N_34730,N_31384);
and U44472 (N_44472,N_39940,N_36943);
and U44473 (N_44473,N_37052,N_31995);
nor U44474 (N_44474,N_35366,N_30987);
nand U44475 (N_44475,N_31110,N_37312);
or U44476 (N_44476,N_34672,N_38177);
and U44477 (N_44477,N_34541,N_31289);
nand U44478 (N_44478,N_33965,N_33912);
or U44479 (N_44479,N_36332,N_36543);
nand U44480 (N_44480,N_38814,N_32390);
or U44481 (N_44481,N_34204,N_33491);
or U44482 (N_44482,N_35982,N_33972);
nor U44483 (N_44483,N_32588,N_30869);
nor U44484 (N_44484,N_34176,N_32096);
and U44485 (N_44485,N_36474,N_31402);
or U44486 (N_44486,N_36206,N_34833);
or U44487 (N_44487,N_32048,N_35260);
and U44488 (N_44488,N_31769,N_34107);
nand U44489 (N_44489,N_36910,N_37920);
nand U44490 (N_44490,N_34990,N_39223);
xnor U44491 (N_44491,N_36777,N_38618);
and U44492 (N_44492,N_31167,N_30943);
and U44493 (N_44493,N_36149,N_34952);
nor U44494 (N_44494,N_32231,N_34754);
or U44495 (N_44495,N_32859,N_39499);
nand U44496 (N_44496,N_36110,N_38374);
and U44497 (N_44497,N_33952,N_36981);
nor U44498 (N_44498,N_37113,N_38409);
nand U44499 (N_44499,N_35254,N_32077);
nand U44500 (N_44500,N_30701,N_38329);
nand U44501 (N_44501,N_30937,N_31250);
or U44502 (N_44502,N_37118,N_37801);
or U44503 (N_44503,N_39745,N_30416);
nand U44504 (N_44504,N_30916,N_38918);
xnor U44505 (N_44505,N_32750,N_32912);
nand U44506 (N_44506,N_31359,N_37393);
xor U44507 (N_44507,N_33940,N_38370);
or U44508 (N_44508,N_35775,N_38519);
or U44509 (N_44509,N_32687,N_35263);
or U44510 (N_44510,N_39714,N_39439);
xor U44511 (N_44511,N_35307,N_33980);
and U44512 (N_44512,N_39027,N_35718);
and U44513 (N_44513,N_38627,N_37750);
or U44514 (N_44514,N_37587,N_31549);
nand U44515 (N_44515,N_33614,N_35845);
nor U44516 (N_44516,N_35370,N_36749);
and U44517 (N_44517,N_39583,N_38122);
and U44518 (N_44518,N_35383,N_31547);
nand U44519 (N_44519,N_32638,N_30788);
nor U44520 (N_44520,N_38685,N_37683);
nand U44521 (N_44521,N_37732,N_38580);
xor U44522 (N_44522,N_33342,N_35513);
and U44523 (N_44523,N_37807,N_35892);
nor U44524 (N_44524,N_32117,N_33332);
and U44525 (N_44525,N_38307,N_37048);
nor U44526 (N_44526,N_35557,N_30182);
nand U44527 (N_44527,N_39609,N_31259);
and U44528 (N_44528,N_35416,N_30612);
nand U44529 (N_44529,N_30737,N_37348);
nor U44530 (N_44530,N_31707,N_33904);
and U44531 (N_44531,N_32334,N_38159);
nor U44532 (N_44532,N_32650,N_35864);
xor U44533 (N_44533,N_37470,N_32538);
and U44534 (N_44534,N_37690,N_34007);
or U44535 (N_44535,N_31909,N_37842);
or U44536 (N_44536,N_33792,N_35993);
nand U44537 (N_44537,N_32922,N_37314);
nor U44538 (N_44538,N_30585,N_35001);
or U44539 (N_44539,N_37243,N_39384);
or U44540 (N_44540,N_34576,N_39106);
or U44541 (N_44541,N_37781,N_37030);
nor U44542 (N_44542,N_32671,N_30680);
nand U44543 (N_44543,N_35071,N_39432);
and U44544 (N_44544,N_37937,N_31121);
nand U44545 (N_44545,N_33656,N_39675);
nor U44546 (N_44546,N_34904,N_33629);
nor U44547 (N_44547,N_36725,N_35687);
and U44548 (N_44548,N_39841,N_36124);
nand U44549 (N_44549,N_33303,N_30122);
nor U44550 (N_44550,N_36086,N_35597);
xor U44551 (N_44551,N_34654,N_39118);
or U44552 (N_44552,N_33726,N_36300);
nor U44553 (N_44553,N_38186,N_36603);
xor U44554 (N_44554,N_39182,N_31817);
nand U44555 (N_44555,N_34467,N_38071);
xor U44556 (N_44556,N_31068,N_31777);
nor U44557 (N_44557,N_35794,N_37288);
nand U44558 (N_44558,N_39887,N_30531);
and U44559 (N_44559,N_35581,N_30126);
or U44560 (N_44560,N_38432,N_37681);
nand U44561 (N_44561,N_37381,N_31457);
and U44562 (N_44562,N_36703,N_31520);
nand U44563 (N_44563,N_35935,N_30190);
nand U44564 (N_44564,N_32013,N_38363);
nand U44565 (N_44565,N_36630,N_31720);
or U44566 (N_44566,N_35608,N_37922);
nand U44567 (N_44567,N_38462,N_32893);
and U44568 (N_44568,N_37390,N_34995);
or U44569 (N_44569,N_34344,N_38862);
xnor U44570 (N_44570,N_39565,N_33755);
nor U44571 (N_44571,N_37147,N_30353);
nor U44572 (N_44572,N_38385,N_36847);
or U44573 (N_44573,N_39236,N_32629);
nor U44574 (N_44574,N_37344,N_34092);
nor U44575 (N_44575,N_34472,N_35574);
nand U44576 (N_44576,N_31050,N_38799);
nand U44577 (N_44577,N_33601,N_32956);
and U44578 (N_44578,N_36059,N_39453);
and U44579 (N_44579,N_38969,N_35056);
nand U44580 (N_44580,N_32192,N_36945);
or U44581 (N_44581,N_35539,N_32754);
nand U44582 (N_44582,N_32323,N_30120);
nand U44583 (N_44583,N_37026,N_31290);
and U44584 (N_44584,N_31063,N_35058);
xnor U44585 (N_44585,N_33218,N_35301);
nand U44586 (N_44586,N_33312,N_38879);
nand U44587 (N_44587,N_33168,N_30426);
nor U44588 (N_44588,N_36748,N_31021);
and U44589 (N_44589,N_32636,N_35121);
and U44590 (N_44590,N_32185,N_39386);
nor U44591 (N_44591,N_38451,N_34601);
nand U44592 (N_44592,N_31380,N_34324);
or U44593 (N_44593,N_30200,N_39930);
nand U44594 (N_44594,N_30487,N_37714);
nand U44595 (N_44595,N_30922,N_34283);
and U44596 (N_44596,N_33780,N_37133);
or U44597 (N_44597,N_35102,N_30438);
or U44598 (N_44598,N_35357,N_30431);
nor U44599 (N_44599,N_30286,N_36397);
nor U44600 (N_44600,N_31690,N_31122);
nand U44601 (N_44601,N_36405,N_34494);
nor U44602 (N_44602,N_37085,N_31585);
and U44603 (N_44603,N_30895,N_31276);
and U44604 (N_44604,N_31235,N_35868);
and U44605 (N_44605,N_39197,N_30864);
xnor U44606 (N_44606,N_33966,N_39784);
xnor U44607 (N_44607,N_36314,N_31931);
and U44608 (N_44608,N_36099,N_30486);
and U44609 (N_44609,N_31669,N_36764);
nor U44610 (N_44610,N_38327,N_32044);
nor U44611 (N_44611,N_31374,N_32403);
nor U44612 (N_44612,N_35589,N_30480);
nor U44613 (N_44613,N_32032,N_37383);
nor U44614 (N_44614,N_30667,N_35302);
or U44615 (N_44615,N_34811,N_35907);
or U44616 (N_44616,N_39493,N_34959);
and U44617 (N_44617,N_33069,N_31843);
or U44618 (N_44618,N_36364,N_30811);
and U44619 (N_44619,N_35618,N_37818);
nor U44620 (N_44620,N_34767,N_32907);
and U44621 (N_44621,N_31833,N_37204);
nand U44622 (N_44622,N_39730,N_39742);
nand U44623 (N_44623,N_30140,N_32708);
and U44624 (N_44624,N_39719,N_34277);
nand U44625 (N_44625,N_30671,N_38524);
or U44626 (N_44626,N_33397,N_39062);
nand U44627 (N_44627,N_39913,N_37141);
nand U44628 (N_44628,N_38709,N_34600);
or U44629 (N_44629,N_37516,N_34123);
xor U44630 (N_44630,N_33705,N_32457);
or U44631 (N_44631,N_33458,N_33147);
nand U44632 (N_44632,N_33620,N_38747);
nor U44633 (N_44633,N_39711,N_34119);
and U44634 (N_44634,N_34491,N_36197);
nand U44635 (N_44635,N_34290,N_39069);
nor U44636 (N_44636,N_34805,N_31073);
nor U44637 (N_44637,N_33299,N_35255);
xor U44638 (N_44638,N_32281,N_37838);
xnor U44639 (N_44639,N_36694,N_38790);
nand U44640 (N_44640,N_38077,N_36512);
nor U44641 (N_44641,N_32696,N_38728);
nor U44642 (N_44642,N_30761,N_35231);
xor U44643 (N_44643,N_35897,N_38800);
nor U44644 (N_44644,N_32806,N_34722);
or U44645 (N_44645,N_35361,N_39136);
or U44646 (N_44646,N_39769,N_35362);
nor U44647 (N_44647,N_30673,N_38342);
and U44648 (N_44648,N_38932,N_32955);
and U44649 (N_44649,N_36450,N_36249);
and U44650 (N_44650,N_37425,N_38996);
nand U44651 (N_44651,N_32703,N_31701);
nand U44652 (N_44652,N_31828,N_36255);
or U44653 (N_44653,N_33318,N_31179);
nor U44654 (N_44654,N_35464,N_37848);
and U44655 (N_44655,N_35424,N_33745);
or U44656 (N_44656,N_34792,N_33193);
xnor U44657 (N_44657,N_34278,N_38070);
nor U44658 (N_44658,N_31838,N_34599);
nor U44659 (N_44659,N_36298,N_32244);
nand U44660 (N_44660,N_36613,N_31960);
and U44661 (N_44661,N_36003,N_35953);
nor U44662 (N_44662,N_38960,N_32971);
nor U44663 (N_44663,N_37478,N_35904);
nor U44664 (N_44664,N_30230,N_38813);
xnor U44665 (N_44665,N_33500,N_37338);
and U44666 (N_44666,N_39974,N_35221);
and U44667 (N_44667,N_37996,N_35497);
nor U44668 (N_44668,N_35802,N_33441);
and U44669 (N_44669,N_34037,N_30104);
nand U44670 (N_44670,N_35501,N_34158);
nor U44671 (N_44671,N_37112,N_35696);
or U44672 (N_44672,N_30354,N_30383);
nor U44673 (N_44673,N_31385,N_31929);
nor U44674 (N_44674,N_35873,N_34160);
and U44675 (N_44675,N_32741,N_31917);
or U44676 (N_44676,N_33425,N_30741);
nor U44677 (N_44677,N_33323,N_39021);
nor U44678 (N_44678,N_39491,N_31483);
nor U44679 (N_44679,N_37571,N_33134);
nor U44680 (N_44680,N_39425,N_32623);
nor U44681 (N_44681,N_31233,N_39983);
or U44682 (N_44682,N_33266,N_30792);
nand U44683 (N_44683,N_35274,N_32275);
or U44684 (N_44684,N_35025,N_34778);
xnor U44685 (N_44685,N_31907,N_34530);
or U44686 (N_44686,N_37128,N_30111);
and U44687 (N_44687,N_33679,N_30363);
nor U44688 (N_44688,N_32460,N_35989);
nand U44689 (N_44689,N_32114,N_34641);
and U44690 (N_44690,N_37944,N_37029);
and U44691 (N_44691,N_34394,N_35436);
nand U44692 (N_44692,N_30722,N_38194);
or U44693 (N_44693,N_34547,N_37968);
nor U44694 (N_44694,N_35820,N_31670);
or U44695 (N_44695,N_35425,N_32359);
nand U44696 (N_44696,N_38520,N_34163);
or U44697 (N_44697,N_35805,N_30670);
nor U44698 (N_44698,N_35067,N_31577);
or U44699 (N_44699,N_35664,N_34347);
nor U44700 (N_44700,N_32312,N_38120);
nor U44701 (N_44701,N_30688,N_30610);
or U44702 (N_44702,N_31666,N_30000);
or U44703 (N_44703,N_35367,N_39514);
nand U44704 (N_44704,N_38654,N_32953);
nand U44705 (N_44705,N_36169,N_39289);
and U44706 (N_44706,N_32203,N_30252);
nor U44707 (N_44707,N_35061,N_32958);
and U44708 (N_44708,N_32139,N_39159);
nand U44709 (N_44709,N_33751,N_30425);
nor U44710 (N_44710,N_32729,N_32841);
or U44711 (N_44711,N_36927,N_31215);
nor U44712 (N_44712,N_34798,N_37046);
nand U44713 (N_44713,N_32423,N_33677);
xor U44714 (N_44714,N_36140,N_39387);
or U44715 (N_44715,N_36422,N_30570);
nor U44716 (N_44716,N_37689,N_34087);
or U44717 (N_44717,N_31782,N_30348);
and U44718 (N_44718,N_30683,N_33142);
or U44719 (N_44719,N_31120,N_30716);
nand U44720 (N_44720,N_31065,N_32944);
nand U44721 (N_44721,N_35197,N_34533);
nand U44722 (N_44722,N_35885,N_36634);
or U44723 (N_44723,N_32954,N_39278);
nor U44724 (N_44724,N_37114,N_39652);
or U44725 (N_44725,N_36065,N_33615);
and U44726 (N_44726,N_35326,N_33842);
or U44727 (N_44727,N_33320,N_31200);
and U44728 (N_44728,N_37624,N_36681);
and U44729 (N_44729,N_33510,N_34800);
or U44730 (N_44730,N_33507,N_34027);
xor U44731 (N_44731,N_33328,N_36696);
nand U44732 (N_44732,N_30261,N_37155);
or U44733 (N_44733,N_35630,N_39817);
and U44734 (N_44734,N_35541,N_39998);
nor U44735 (N_44735,N_37475,N_34401);
nor U44736 (N_44736,N_35400,N_30626);
nand U44737 (N_44737,N_32631,N_37912);
or U44738 (N_44738,N_36292,N_30702);
nand U44739 (N_44739,N_38946,N_36966);
nand U44740 (N_44740,N_30556,N_36590);
or U44741 (N_44741,N_32027,N_36337);
nand U44742 (N_44742,N_33566,N_39713);
and U44743 (N_44743,N_31718,N_34651);
and U44744 (N_44744,N_31382,N_35853);
and U44745 (N_44745,N_31363,N_38571);
or U44746 (N_44746,N_30472,N_34700);
nand U44747 (N_44747,N_38439,N_35191);
and U44748 (N_44748,N_37442,N_30730);
nor U44749 (N_44749,N_31491,N_31456);
or U44750 (N_44750,N_39390,N_34988);
or U44751 (N_44751,N_35153,N_38857);
xnor U44752 (N_44752,N_31591,N_30100);
or U44753 (N_44753,N_38229,N_34978);
nor U44754 (N_44754,N_39805,N_38356);
or U44755 (N_44755,N_35940,N_38733);
nor U44756 (N_44756,N_30542,N_32680);
or U44757 (N_44757,N_35976,N_32721);
or U44758 (N_44758,N_33630,N_39084);
xor U44759 (N_44759,N_34362,N_36369);
or U44760 (N_44760,N_38328,N_37320);
nand U44761 (N_44761,N_30948,N_38934);
nand U44762 (N_44762,N_34111,N_35336);
nor U44763 (N_44763,N_33814,N_39605);
and U44764 (N_44764,N_38852,N_39041);
nand U44765 (N_44765,N_32874,N_35649);
nor U44766 (N_44766,N_38784,N_36129);
nor U44767 (N_44767,N_36852,N_34539);
or U44768 (N_44768,N_31808,N_37917);
or U44769 (N_44769,N_31279,N_36430);
xnor U44770 (N_44770,N_34509,N_36711);
nor U44771 (N_44771,N_31951,N_31282);
and U44772 (N_44772,N_38249,N_34877);
or U44773 (N_44773,N_38030,N_34299);
or U44774 (N_44774,N_33987,N_37068);
nor U44775 (N_44775,N_34712,N_38483);
nor U44776 (N_44776,N_31446,N_33161);
or U44777 (N_44777,N_32399,N_34596);
nand U44778 (N_44778,N_36380,N_33021);
or U44779 (N_44779,N_30575,N_35931);
nor U44780 (N_44780,N_33257,N_35324);
or U44781 (N_44781,N_31266,N_33315);
or U44782 (N_44782,N_30210,N_34931);
and U44783 (N_44783,N_32920,N_36299);
nand U44784 (N_44784,N_39119,N_36923);
and U44785 (N_44785,N_33239,N_34110);
or U44786 (N_44786,N_31824,N_35183);
nand U44787 (N_44787,N_34339,N_35472);
nand U44788 (N_44788,N_36365,N_37517);
and U44789 (N_44789,N_33704,N_33254);
nand U44790 (N_44790,N_31834,N_37720);
and U44791 (N_44791,N_36667,N_38779);
or U44792 (N_44792,N_39111,N_37228);
and U44793 (N_44793,N_37851,N_38331);
and U44794 (N_44794,N_37127,N_32061);
nor U44795 (N_44795,N_37449,N_32743);
nand U44796 (N_44796,N_39163,N_36360);
nor U44797 (N_44797,N_31367,N_31976);
nor U44798 (N_44798,N_39200,N_33738);
and U44799 (N_44799,N_39568,N_35414);
nor U44800 (N_44800,N_34550,N_34515);
or U44801 (N_44801,N_33798,N_39031);
and U44802 (N_44802,N_39176,N_31328);
and U44803 (N_44803,N_38016,N_35914);
and U44804 (N_44804,N_38856,N_31052);
or U44805 (N_44805,N_33085,N_34063);
and U44806 (N_44806,N_35213,N_37196);
or U44807 (N_44807,N_35763,N_38560);
nor U44808 (N_44808,N_30827,N_37274);
or U44809 (N_44809,N_31840,N_32322);
nor U44810 (N_44810,N_39195,N_35674);
or U44811 (N_44811,N_30266,N_32441);
and U44812 (N_44812,N_35478,N_34133);
and U44813 (N_44813,N_34381,N_36900);
or U44814 (N_44814,N_35954,N_34415);
nor U44815 (N_44815,N_34316,N_39626);
or U44816 (N_44816,N_34775,N_33733);
nor U44817 (N_44817,N_35616,N_30813);
nor U44818 (N_44818,N_31647,N_32804);
nor U44819 (N_44819,N_31042,N_31386);
nor U44820 (N_44820,N_30134,N_30764);
or U44821 (N_44821,N_32391,N_32429);
or U44822 (N_44822,N_38976,N_30917);
nor U44823 (N_44823,N_33287,N_35686);
or U44824 (N_44824,N_30974,N_39403);
or U44825 (N_44825,N_39167,N_38586);
nor U44826 (N_44826,N_38787,N_33625);
xnor U44827 (N_44827,N_35076,N_33215);
and U44828 (N_44828,N_35485,N_30216);
nor U44829 (N_44829,N_33973,N_37966);
and U44830 (N_44830,N_34913,N_37546);
nor U44831 (N_44831,N_34495,N_31056);
xnor U44832 (N_44832,N_34006,N_30803);
nand U44833 (N_44833,N_35512,N_32273);
or U44834 (N_44834,N_31890,N_32180);
nor U44835 (N_44835,N_36199,N_37315);
nor U44836 (N_44836,N_30804,N_31231);
or U44837 (N_44837,N_35772,N_32415);
nor U44838 (N_44838,N_38031,N_36442);
or U44839 (N_44839,N_31057,N_33811);
nand U44840 (N_44840,N_34334,N_33840);
or U44841 (N_44841,N_30390,N_32879);
nor U44842 (N_44842,N_30801,N_30417);
and U44843 (N_44843,N_38243,N_37588);
nand U44844 (N_44844,N_37016,N_35471);
and U44845 (N_44845,N_33589,N_36064);
nand U44846 (N_44846,N_39865,N_31412);
or U44847 (N_44847,N_31494,N_39608);
nand U44848 (N_44848,N_36192,N_39733);
and U44849 (N_44849,N_35951,N_35363);
and U44850 (N_44850,N_32372,N_36628);
nand U44851 (N_44851,N_36479,N_30170);
or U44852 (N_44852,N_37792,N_35019);
and U44853 (N_44853,N_33754,N_38600);
nand U44854 (N_44854,N_31540,N_37695);
nand U44855 (N_44855,N_31575,N_39897);
nor U44856 (N_44856,N_38289,N_30071);
xor U44857 (N_44857,N_38212,N_38525);
or U44858 (N_44858,N_34435,N_35720);
and U44859 (N_44859,N_38818,N_35444);
or U44860 (N_44860,N_37799,N_30336);
or U44861 (N_44861,N_35821,N_37748);
nand U44862 (N_44862,N_38383,N_35321);
xnor U44863 (N_44863,N_39058,N_37275);
and U44864 (N_44864,N_37707,N_39962);
nand U44865 (N_44865,N_39727,N_36903);
or U44866 (N_44866,N_37069,N_38675);
nor U44867 (N_44867,N_32351,N_31035);
xnor U44868 (N_44868,N_38262,N_33157);
nor U44869 (N_44869,N_31644,N_38751);
nand U44870 (N_44870,N_36416,N_34218);
nand U44871 (N_44871,N_38408,N_37202);
and U44872 (N_44872,N_39970,N_33173);
xnor U44873 (N_44873,N_35586,N_35245);
nor U44874 (N_44874,N_32145,N_34429);
or U44875 (N_44875,N_37759,N_38894);
or U44876 (N_44876,N_35272,N_30213);
and U44877 (N_44877,N_36428,N_30874);
xor U44878 (N_44878,N_34417,N_34620);
nand U44879 (N_44879,N_38998,N_36802);
and U44880 (N_44880,N_30152,N_37703);
and U44881 (N_44881,N_32544,N_30332);
nand U44882 (N_44882,N_32102,N_37640);
or U44883 (N_44883,N_35671,N_33854);
or U44884 (N_44884,N_36500,N_34720);
nor U44885 (N_44885,N_36523,N_37183);
or U44886 (N_44886,N_31033,N_34517);
or U44887 (N_44887,N_37087,N_38284);
and U44888 (N_44888,N_32427,N_37949);
and U44889 (N_44889,N_39056,N_34421);
or U44890 (N_44890,N_39823,N_36387);
nand U44891 (N_44891,N_30703,N_39467);
nand U44892 (N_44892,N_36498,N_32763);
nor U44893 (N_44893,N_30773,N_36347);
or U44894 (N_44894,N_36034,N_34737);
or U44895 (N_44895,N_36839,N_34187);
and U44896 (N_44896,N_32453,N_33600);
nor U44897 (N_44897,N_36722,N_38218);
or U44898 (N_44898,N_34231,N_35116);
nand U44899 (N_44899,N_36706,N_31774);
or U44900 (N_44900,N_33890,N_39350);
xnor U44901 (N_44901,N_30471,N_37337);
or U44902 (N_44902,N_34311,N_38546);
nand U44903 (N_44903,N_35033,N_31573);
nor U44904 (N_44904,N_30298,N_36527);
or U44905 (N_44905,N_31459,N_38460);
and U44906 (N_44906,N_31580,N_36454);
nand U44907 (N_44907,N_36941,N_38434);
and U44908 (N_44908,N_36859,N_33127);
or U44909 (N_44909,N_33206,N_38160);
nor U44910 (N_44910,N_30719,N_30397);
and U44911 (N_44911,N_39253,N_31787);
xnor U44912 (N_44912,N_38521,N_32656);
or U44913 (N_44913,N_35699,N_31001);
nor U44914 (N_44914,N_39430,N_32496);
or U44915 (N_44915,N_37247,N_36947);
xnor U44916 (N_44916,N_38850,N_35077);
nor U44917 (N_44917,N_38392,N_37467);
nand U44918 (N_44918,N_36620,N_33386);
nor U44919 (N_44919,N_37550,N_32179);
xor U44920 (N_44920,N_39954,N_38085);
xor U44921 (N_44921,N_35906,N_35224);
nand U44922 (N_44922,N_36070,N_35678);
nand U44923 (N_44923,N_31715,N_32272);
and U44924 (N_44924,N_33891,N_32287);
nand U44925 (N_44925,N_39772,N_38258);
and U44926 (N_44926,N_37808,N_38848);
xor U44927 (N_44927,N_31118,N_38967);
nor U44928 (N_44928,N_37306,N_31178);
and U44929 (N_44929,N_32356,N_37674);
nor U44930 (N_44930,N_38075,N_32053);
xnor U44931 (N_44931,N_33416,N_38465);
nor U44932 (N_44932,N_31312,N_30360);
or U44933 (N_44933,N_32242,N_35239);
and U44934 (N_44934,N_36285,N_32183);
or U44935 (N_44935,N_37398,N_37384);
nand U44936 (N_44936,N_38920,N_34662);
or U44937 (N_44937,N_33454,N_39511);
nor U44938 (N_44938,N_32943,N_31031);
nand U44939 (N_44939,N_38529,N_31489);
nor U44940 (N_44940,N_32681,N_37456);
and U44941 (N_44941,N_38593,N_31942);
nand U44942 (N_44942,N_35333,N_30163);
nand U44943 (N_44943,N_37988,N_31928);
nor U44944 (N_44944,N_30990,N_30321);
or U44945 (N_44945,N_38095,N_38164);
or U44946 (N_44946,N_37278,N_37645);
xor U44947 (N_44947,N_34147,N_31615);
and U44948 (N_44948,N_34300,N_34729);
or U44949 (N_44949,N_30206,N_34655);
nand U44950 (N_44950,N_30284,N_31294);
and U44951 (N_44951,N_34999,N_31990);
nor U44952 (N_44952,N_36183,N_30502);
nand U44953 (N_44953,N_37509,N_36492);
nor U44954 (N_44954,N_35137,N_31338);
nor U44955 (N_44955,N_30921,N_33404);
nor U44956 (N_44956,N_38714,N_33666);
or U44957 (N_44957,N_30554,N_36291);
nand U44958 (N_44958,N_32066,N_31030);
nand U44959 (N_44959,N_31948,N_34368);
nor U44960 (N_44960,N_38482,N_36328);
or U44961 (N_44961,N_32514,N_31623);
xor U44962 (N_44962,N_35151,N_31125);
and U44963 (N_44963,N_38265,N_31558);
or U44964 (N_44964,N_35097,N_31158);
or U44965 (N_44965,N_35486,N_32198);
and U44966 (N_44966,N_30415,N_38925);
or U44967 (N_44967,N_31758,N_31012);
nor U44968 (N_44968,N_36087,N_37244);
nor U44969 (N_44969,N_32821,N_36276);
or U44970 (N_44970,N_31728,N_34485);
xor U44971 (N_44971,N_33333,N_35430);
and U44972 (N_44972,N_34835,N_39220);
nor U44973 (N_44973,N_33820,N_35786);
nor U44974 (N_44974,N_35590,N_37580);
xnor U44975 (N_44975,N_37416,N_34074);
or U44976 (N_44976,N_35804,N_32785);
and U44977 (N_44977,N_34361,N_36395);
or U44978 (N_44978,N_33692,N_30481);
nor U44979 (N_44979,N_30254,N_37424);
and U44980 (N_44980,N_31963,N_37015);
or U44981 (N_44981,N_34183,N_31332);
nor U44982 (N_44982,N_35180,N_31888);
or U44983 (N_44983,N_34211,N_35534);
or U44984 (N_44984,N_39241,N_38658);
or U44985 (N_44985,N_36491,N_32824);
nor U44986 (N_44986,N_32935,N_38630);
nand U44987 (N_44987,N_36619,N_30526);
nand U44988 (N_44988,N_33057,N_33698);
and U44989 (N_44989,N_33279,N_39522);
or U44990 (N_44990,N_36861,N_34891);
nor U44991 (N_44991,N_38896,N_32834);
nor U44992 (N_44992,N_35237,N_38143);
or U44993 (N_44993,N_32369,N_39189);
nand U44994 (N_44994,N_36570,N_39417);
or U44995 (N_44995,N_36665,N_32101);
or U44996 (N_44996,N_38433,N_32856);
xor U44997 (N_44997,N_34630,N_38300);
or U44998 (N_44998,N_38573,N_31406);
nor U44999 (N_44999,N_31251,N_38485);
nor U45000 (N_45000,N_38131,N_32549);
and U45001 (N_45001,N_31713,N_34626);
or U45002 (N_45002,N_39021,N_33468);
nor U45003 (N_45003,N_39088,N_35853);
and U45004 (N_45004,N_31928,N_30678);
xor U45005 (N_45005,N_35109,N_30095);
nand U45006 (N_45006,N_33933,N_39932);
or U45007 (N_45007,N_30557,N_37359);
and U45008 (N_45008,N_38667,N_35212);
nand U45009 (N_45009,N_33542,N_32828);
xor U45010 (N_45010,N_39971,N_32689);
nand U45011 (N_45011,N_36547,N_30258);
and U45012 (N_45012,N_39116,N_39322);
xnor U45013 (N_45013,N_35490,N_38546);
and U45014 (N_45014,N_35899,N_35567);
or U45015 (N_45015,N_31087,N_37235);
or U45016 (N_45016,N_32537,N_37743);
or U45017 (N_45017,N_35412,N_39466);
nand U45018 (N_45018,N_37670,N_36965);
nor U45019 (N_45019,N_37643,N_39945);
or U45020 (N_45020,N_30936,N_36459);
or U45021 (N_45021,N_35939,N_33736);
xor U45022 (N_45022,N_30693,N_33132);
xor U45023 (N_45023,N_32805,N_32885);
and U45024 (N_45024,N_33504,N_32959);
or U45025 (N_45025,N_30522,N_33034);
xnor U45026 (N_45026,N_31272,N_36228);
nor U45027 (N_45027,N_38947,N_32248);
or U45028 (N_45028,N_31226,N_38278);
or U45029 (N_45029,N_35684,N_38227);
nand U45030 (N_45030,N_33652,N_39790);
nand U45031 (N_45031,N_31672,N_32102);
or U45032 (N_45032,N_38615,N_35220);
and U45033 (N_45033,N_34901,N_36930);
and U45034 (N_45034,N_36420,N_31823);
or U45035 (N_45035,N_39455,N_34514);
or U45036 (N_45036,N_36076,N_34808);
nor U45037 (N_45037,N_31640,N_37541);
and U45038 (N_45038,N_31658,N_33719);
xor U45039 (N_45039,N_33645,N_38012);
or U45040 (N_45040,N_35889,N_34496);
or U45041 (N_45041,N_31501,N_31767);
or U45042 (N_45042,N_35890,N_35078);
or U45043 (N_45043,N_35166,N_35071);
or U45044 (N_45044,N_32843,N_33277);
or U45045 (N_45045,N_38401,N_39788);
nor U45046 (N_45046,N_33147,N_30768);
and U45047 (N_45047,N_31272,N_38745);
and U45048 (N_45048,N_39068,N_38723);
or U45049 (N_45049,N_38138,N_34242);
or U45050 (N_45050,N_33090,N_31164);
and U45051 (N_45051,N_39688,N_34771);
nand U45052 (N_45052,N_34631,N_38218);
nand U45053 (N_45053,N_34031,N_35686);
xor U45054 (N_45054,N_31243,N_39616);
nand U45055 (N_45055,N_35218,N_35633);
nand U45056 (N_45056,N_38223,N_30120);
nor U45057 (N_45057,N_36192,N_38050);
or U45058 (N_45058,N_37228,N_33910);
xor U45059 (N_45059,N_35808,N_34106);
nor U45060 (N_45060,N_38570,N_30716);
or U45061 (N_45061,N_32917,N_38179);
and U45062 (N_45062,N_32650,N_34684);
or U45063 (N_45063,N_32101,N_30743);
and U45064 (N_45064,N_32609,N_36875);
nor U45065 (N_45065,N_34304,N_32501);
or U45066 (N_45066,N_39760,N_37069);
nand U45067 (N_45067,N_35616,N_32204);
and U45068 (N_45068,N_35695,N_39822);
xnor U45069 (N_45069,N_32373,N_35259);
and U45070 (N_45070,N_35241,N_37014);
nand U45071 (N_45071,N_32069,N_33129);
and U45072 (N_45072,N_37495,N_38539);
and U45073 (N_45073,N_39474,N_36233);
nor U45074 (N_45074,N_36647,N_35506);
nand U45075 (N_45075,N_30986,N_36081);
and U45076 (N_45076,N_39086,N_35782);
nor U45077 (N_45077,N_32967,N_31733);
or U45078 (N_45078,N_38429,N_38618);
nor U45079 (N_45079,N_30550,N_34266);
nor U45080 (N_45080,N_38845,N_31724);
and U45081 (N_45081,N_32865,N_33751);
nor U45082 (N_45082,N_39206,N_36903);
and U45083 (N_45083,N_30572,N_34237);
nand U45084 (N_45084,N_38181,N_34842);
and U45085 (N_45085,N_35373,N_37166);
and U45086 (N_45086,N_31273,N_34389);
nand U45087 (N_45087,N_32465,N_30383);
nand U45088 (N_45088,N_35830,N_37600);
or U45089 (N_45089,N_32282,N_39161);
or U45090 (N_45090,N_37245,N_39469);
nand U45091 (N_45091,N_31873,N_38305);
nor U45092 (N_45092,N_31165,N_33531);
nand U45093 (N_45093,N_39826,N_32045);
or U45094 (N_45094,N_30772,N_36386);
nand U45095 (N_45095,N_33694,N_37907);
and U45096 (N_45096,N_35378,N_39621);
or U45097 (N_45097,N_35701,N_33957);
nand U45098 (N_45098,N_30742,N_39063);
xnor U45099 (N_45099,N_37803,N_37240);
xnor U45100 (N_45100,N_35515,N_34071);
nand U45101 (N_45101,N_33936,N_30957);
and U45102 (N_45102,N_39950,N_31637);
nand U45103 (N_45103,N_38699,N_34169);
or U45104 (N_45104,N_39685,N_30942);
xor U45105 (N_45105,N_39853,N_39204);
and U45106 (N_45106,N_36793,N_35284);
or U45107 (N_45107,N_32622,N_33118);
xnor U45108 (N_45108,N_34994,N_31269);
nor U45109 (N_45109,N_32283,N_31901);
xnor U45110 (N_45110,N_35571,N_30474);
nand U45111 (N_45111,N_37118,N_38257);
xor U45112 (N_45112,N_32782,N_36852);
xor U45113 (N_45113,N_35668,N_30348);
nor U45114 (N_45114,N_36545,N_39069);
nand U45115 (N_45115,N_31581,N_36288);
nor U45116 (N_45116,N_38917,N_30335);
or U45117 (N_45117,N_34931,N_39878);
or U45118 (N_45118,N_37484,N_39884);
and U45119 (N_45119,N_34221,N_38972);
nor U45120 (N_45120,N_37696,N_34246);
nand U45121 (N_45121,N_35824,N_35312);
nor U45122 (N_45122,N_34596,N_31037);
or U45123 (N_45123,N_38066,N_31219);
and U45124 (N_45124,N_31746,N_33821);
nor U45125 (N_45125,N_35861,N_32705);
or U45126 (N_45126,N_32751,N_36766);
nand U45127 (N_45127,N_36154,N_39443);
nor U45128 (N_45128,N_32006,N_36458);
and U45129 (N_45129,N_36778,N_35904);
nor U45130 (N_45130,N_39741,N_35079);
or U45131 (N_45131,N_30001,N_37065);
nor U45132 (N_45132,N_33411,N_30259);
xnor U45133 (N_45133,N_32775,N_38411);
or U45134 (N_45134,N_33080,N_33055);
and U45135 (N_45135,N_31706,N_38122);
nor U45136 (N_45136,N_32575,N_31545);
nand U45137 (N_45137,N_31310,N_36357);
and U45138 (N_45138,N_33453,N_37321);
nand U45139 (N_45139,N_30758,N_31304);
and U45140 (N_45140,N_38366,N_38730);
nor U45141 (N_45141,N_31241,N_38198);
xor U45142 (N_45142,N_38476,N_33692);
and U45143 (N_45143,N_37144,N_36917);
nor U45144 (N_45144,N_30514,N_37804);
or U45145 (N_45145,N_33808,N_32353);
nor U45146 (N_45146,N_37176,N_39533);
and U45147 (N_45147,N_33721,N_35441);
and U45148 (N_45148,N_33318,N_34580);
nand U45149 (N_45149,N_33439,N_35768);
nand U45150 (N_45150,N_35446,N_33084);
or U45151 (N_45151,N_39885,N_36844);
nand U45152 (N_45152,N_38354,N_35713);
nand U45153 (N_45153,N_32174,N_37162);
and U45154 (N_45154,N_32630,N_36335);
and U45155 (N_45155,N_31013,N_36513);
xnor U45156 (N_45156,N_36300,N_38873);
or U45157 (N_45157,N_36085,N_35130);
or U45158 (N_45158,N_38406,N_31467);
xnor U45159 (N_45159,N_31739,N_34673);
nor U45160 (N_45160,N_36565,N_34731);
nor U45161 (N_45161,N_30929,N_32011);
or U45162 (N_45162,N_37189,N_38586);
nand U45163 (N_45163,N_39546,N_33602);
nor U45164 (N_45164,N_30362,N_32229);
nor U45165 (N_45165,N_39690,N_38010);
or U45166 (N_45166,N_32211,N_38635);
or U45167 (N_45167,N_39273,N_33869);
and U45168 (N_45168,N_36086,N_39134);
and U45169 (N_45169,N_34066,N_31996);
or U45170 (N_45170,N_35856,N_32224);
nand U45171 (N_45171,N_35730,N_39786);
or U45172 (N_45172,N_35695,N_32067);
xor U45173 (N_45173,N_32715,N_36056);
and U45174 (N_45174,N_31896,N_32818);
nor U45175 (N_45175,N_32639,N_32441);
or U45176 (N_45176,N_38178,N_34446);
nor U45177 (N_45177,N_30184,N_38952);
or U45178 (N_45178,N_38859,N_37240);
xnor U45179 (N_45179,N_30603,N_39760);
or U45180 (N_45180,N_39956,N_34000);
nand U45181 (N_45181,N_35891,N_37072);
or U45182 (N_45182,N_30225,N_35800);
nand U45183 (N_45183,N_39101,N_39202);
nand U45184 (N_45184,N_30414,N_34392);
nor U45185 (N_45185,N_31646,N_35845);
and U45186 (N_45186,N_32321,N_39172);
xnor U45187 (N_45187,N_30128,N_38453);
and U45188 (N_45188,N_36475,N_36332);
nand U45189 (N_45189,N_36614,N_36526);
and U45190 (N_45190,N_31094,N_35005);
or U45191 (N_45191,N_32826,N_30030);
and U45192 (N_45192,N_37530,N_33939);
and U45193 (N_45193,N_36869,N_38595);
and U45194 (N_45194,N_30252,N_33988);
xnor U45195 (N_45195,N_35205,N_39352);
nand U45196 (N_45196,N_33099,N_35555);
or U45197 (N_45197,N_30113,N_31722);
nor U45198 (N_45198,N_33824,N_35326);
nor U45199 (N_45199,N_31536,N_31203);
and U45200 (N_45200,N_38474,N_39905);
or U45201 (N_45201,N_39437,N_36326);
nand U45202 (N_45202,N_30322,N_39763);
or U45203 (N_45203,N_37661,N_30495);
xnor U45204 (N_45204,N_35626,N_31191);
nor U45205 (N_45205,N_35577,N_38633);
nand U45206 (N_45206,N_39623,N_39975);
nor U45207 (N_45207,N_30182,N_38783);
nand U45208 (N_45208,N_37923,N_31102);
or U45209 (N_45209,N_34555,N_30559);
and U45210 (N_45210,N_36088,N_37801);
and U45211 (N_45211,N_34721,N_38883);
or U45212 (N_45212,N_35955,N_35127);
nand U45213 (N_45213,N_36844,N_38395);
nor U45214 (N_45214,N_39739,N_30406);
xor U45215 (N_45215,N_38138,N_33038);
or U45216 (N_45216,N_33304,N_39205);
and U45217 (N_45217,N_30245,N_37241);
and U45218 (N_45218,N_35616,N_34541);
nor U45219 (N_45219,N_36573,N_37757);
and U45220 (N_45220,N_32135,N_31377);
and U45221 (N_45221,N_35233,N_31364);
or U45222 (N_45222,N_36762,N_37866);
or U45223 (N_45223,N_36365,N_31370);
or U45224 (N_45224,N_39988,N_35364);
and U45225 (N_45225,N_38874,N_39838);
nor U45226 (N_45226,N_33128,N_33555);
and U45227 (N_45227,N_35672,N_33619);
or U45228 (N_45228,N_35164,N_39329);
nand U45229 (N_45229,N_31123,N_31746);
or U45230 (N_45230,N_31744,N_35026);
and U45231 (N_45231,N_39083,N_30465);
and U45232 (N_45232,N_30143,N_34581);
or U45233 (N_45233,N_35319,N_32481);
and U45234 (N_45234,N_36939,N_35375);
and U45235 (N_45235,N_30542,N_38417);
nand U45236 (N_45236,N_39845,N_34940);
and U45237 (N_45237,N_36624,N_31058);
or U45238 (N_45238,N_38531,N_31253);
nor U45239 (N_45239,N_38768,N_31653);
xor U45240 (N_45240,N_31530,N_37828);
nor U45241 (N_45241,N_33978,N_35636);
nand U45242 (N_45242,N_35280,N_36333);
nand U45243 (N_45243,N_34448,N_38603);
or U45244 (N_45244,N_34295,N_31953);
and U45245 (N_45245,N_32082,N_35268);
or U45246 (N_45246,N_33758,N_36605);
and U45247 (N_45247,N_38183,N_33558);
and U45248 (N_45248,N_32019,N_31632);
xor U45249 (N_45249,N_39154,N_34618);
or U45250 (N_45250,N_36369,N_38136);
xnor U45251 (N_45251,N_35553,N_34984);
or U45252 (N_45252,N_39458,N_31412);
or U45253 (N_45253,N_37049,N_30472);
or U45254 (N_45254,N_35352,N_31484);
and U45255 (N_45255,N_36340,N_36398);
nand U45256 (N_45256,N_35826,N_31247);
nand U45257 (N_45257,N_31774,N_35568);
xor U45258 (N_45258,N_34246,N_35280);
or U45259 (N_45259,N_30822,N_36200);
nand U45260 (N_45260,N_30844,N_33902);
nand U45261 (N_45261,N_32059,N_38586);
nand U45262 (N_45262,N_38039,N_30766);
nand U45263 (N_45263,N_34795,N_32284);
nor U45264 (N_45264,N_33065,N_38158);
and U45265 (N_45265,N_36272,N_30224);
and U45266 (N_45266,N_35037,N_39687);
and U45267 (N_45267,N_34026,N_35530);
xor U45268 (N_45268,N_39273,N_37839);
nor U45269 (N_45269,N_35848,N_31805);
nor U45270 (N_45270,N_34918,N_36443);
and U45271 (N_45271,N_39528,N_34819);
nand U45272 (N_45272,N_37154,N_31797);
nor U45273 (N_45273,N_35272,N_38621);
or U45274 (N_45274,N_39364,N_32207);
nor U45275 (N_45275,N_39813,N_36874);
or U45276 (N_45276,N_38266,N_34037);
or U45277 (N_45277,N_30692,N_35495);
nand U45278 (N_45278,N_36873,N_36640);
or U45279 (N_45279,N_30467,N_32062);
and U45280 (N_45280,N_39694,N_34988);
or U45281 (N_45281,N_31872,N_35222);
or U45282 (N_45282,N_36614,N_36146);
and U45283 (N_45283,N_37443,N_39555);
and U45284 (N_45284,N_38466,N_32234);
or U45285 (N_45285,N_39695,N_39521);
and U45286 (N_45286,N_30403,N_30846);
and U45287 (N_45287,N_39771,N_34606);
xnor U45288 (N_45288,N_35698,N_30085);
or U45289 (N_45289,N_33240,N_37840);
nor U45290 (N_45290,N_34097,N_30912);
nand U45291 (N_45291,N_35281,N_30362);
xor U45292 (N_45292,N_32390,N_32777);
nand U45293 (N_45293,N_34227,N_39300);
nor U45294 (N_45294,N_31824,N_33075);
and U45295 (N_45295,N_38129,N_31276);
nor U45296 (N_45296,N_31803,N_31243);
nor U45297 (N_45297,N_31362,N_32916);
and U45298 (N_45298,N_31231,N_39243);
nor U45299 (N_45299,N_37525,N_38096);
and U45300 (N_45300,N_37269,N_30431);
nand U45301 (N_45301,N_37772,N_39070);
and U45302 (N_45302,N_37511,N_37630);
and U45303 (N_45303,N_34333,N_36317);
and U45304 (N_45304,N_37942,N_34234);
nor U45305 (N_45305,N_39812,N_36094);
or U45306 (N_45306,N_38782,N_32013);
xnor U45307 (N_45307,N_38464,N_31441);
or U45308 (N_45308,N_35731,N_33628);
and U45309 (N_45309,N_33447,N_39352);
nand U45310 (N_45310,N_32019,N_34397);
and U45311 (N_45311,N_39225,N_35792);
nand U45312 (N_45312,N_36929,N_35045);
and U45313 (N_45313,N_37055,N_30834);
nor U45314 (N_45314,N_35331,N_30359);
or U45315 (N_45315,N_33624,N_39451);
or U45316 (N_45316,N_38618,N_38797);
nand U45317 (N_45317,N_30215,N_39776);
nand U45318 (N_45318,N_33513,N_34412);
nand U45319 (N_45319,N_30626,N_35475);
and U45320 (N_45320,N_34138,N_36249);
nor U45321 (N_45321,N_30296,N_36642);
nand U45322 (N_45322,N_34610,N_32527);
nand U45323 (N_45323,N_33969,N_38153);
or U45324 (N_45324,N_37488,N_39350);
nand U45325 (N_45325,N_38022,N_34294);
nand U45326 (N_45326,N_37769,N_37241);
nor U45327 (N_45327,N_30508,N_33429);
and U45328 (N_45328,N_31938,N_33716);
nand U45329 (N_45329,N_31190,N_37223);
nor U45330 (N_45330,N_33405,N_34084);
xor U45331 (N_45331,N_31515,N_30363);
or U45332 (N_45332,N_37767,N_30273);
nor U45333 (N_45333,N_35090,N_39192);
and U45334 (N_45334,N_36938,N_32331);
nand U45335 (N_45335,N_38738,N_31433);
nand U45336 (N_45336,N_33293,N_38004);
nor U45337 (N_45337,N_30183,N_33183);
or U45338 (N_45338,N_36398,N_36266);
xor U45339 (N_45339,N_32332,N_38042);
nor U45340 (N_45340,N_39255,N_32887);
nand U45341 (N_45341,N_32340,N_38726);
nand U45342 (N_45342,N_37548,N_34086);
or U45343 (N_45343,N_30616,N_30799);
or U45344 (N_45344,N_39581,N_32159);
or U45345 (N_45345,N_38937,N_30518);
xor U45346 (N_45346,N_30183,N_30216);
nand U45347 (N_45347,N_31659,N_35170);
or U45348 (N_45348,N_38083,N_33345);
xnor U45349 (N_45349,N_34791,N_34208);
and U45350 (N_45350,N_36867,N_37196);
or U45351 (N_45351,N_32963,N_30392);
nand U45352 (N_45352,N_36465,N_31963);
nand U45353 (N_45353,N_34240,N_35482);
nor U45354 (N_45354,N_30281,N_33396);
nor U45355 (N_45355,N_39711,N_36713);
nand U45356 (N_45356,N_39769,N_31402);
nor U45357 (N_45357,N_39713,N_39537);
nand U45358 (N_45358,N_34296,N_33311);
nand U45359 (N_45359,N_39328,N_37475);
nand U45360 (N_45360,N_30845,N_30874);
and U45361 (N_45361,N_39133,N_33367);
and U45362 (N_45362,N_34525,N_31370);
and U45363 (N_45363,N_36467,N_39661);
nor U45364 (N_45364,N_34039,N_34070);
or U45365 (N_45365,N_38809,N_39706);
or U45366 (N_45366,N_36380,N_35343);
nor U45367 (N_45367,N_30713,N_36291);
and U45368 (N_45368,N_37211,N_31645);
or U45369 (N_45369,N_39581,N_30392);
nand U45370 (N_45370,N_34929,N_37203);
xor U45371 (N_45371,N_34544,N_32091);
or U45372 (N_45372,N_30472,N_38322);
or U45373 (N_45373,N_37150,N_31159);
nor U45374 (N_45374,N_39311,N_33690);
and U45375 (N_45375,N_39118,N_30300);
nor U45376 (N_45376,N_33971,N_37831);
nor U45377 (N_45377,N_36702,N_33339);
xnor U45378 (N_45378,N_33381,N_31947);
nand U45379 (N_45379,N_30996,N_39165);
nor U45380 (N_45380,N_35398,N_37647);
nand U45381 (N_45381,N_39454,N_38240);
nand U45382 (N_45382,N_38461,N_33844);
and U45383 (N_45383,N_39070,N_34163);
or U45384 (N_45384,N_34880,N_34619);
and U45385 (N_45385,N_32034,N_37422);
nor U45386 (N_45386,N_30464,N_34826);
and U45387 (N_45387,N_35690,N_31231);
nor U45388 (N_45388,N_33874,N_31122);
xor U45389 (N_45389,N_31903,N_34037);
and U45390 (N_45390,N_37731,N_39633);
xnor U45391 (N_45391,N_30008,N_34160);
xor U45392 (N_45392,N_30323,N_33010);
and U45393 (N_45393,N_30969,N_37081);
nand U45394 (N_45394,N_32596,N_31836);
or U45395 (N_45395,N_37216,N_38194);
nand U45396 (N_45396,N_38569,N_30657);
nand U45397 (N_45397,N_30013,N_33388);
and U45398 (N_45398,N_31182,N_31546);
nand U45399 (N_45399,N_38494,N_30544);
nor U45400 (N_45400,N_34684,N_38455);
nand U45401 (N_45401,N_31399,N_39951);
nand U45402 (N_45402,N_38221,N_34576);
nor U45403 (N_45403,N_33635,N_33613);
and U45404 (N_45404,N_31462,N_39729);
and U45405 (N_45405,N_37012,N_38735);
and U45406 (N_45406,N_32875,N_32211);
xnor U45407 (N_45407,N_39709,N_30005);
or U45408 (N_45408,N_34845,N_33664);
nor U45409 (N_45409,N_38680,N_37684);
nor U45410 (N_45410,N_30495,N_32371);
nor U45411 (N_45411,N_36722,N_30701);
or U45412 (N_45412,N_33737,N_34573);
nor U45413 (N_45413,N_35053,N_33448);
or U45414 (N_45414,N_37799,N_39362);
and U45415 (N_45415,N_35480,N_39810);
xor U45416 (N_45416,N_30347,N_34180);
nor U45417 (N_45417,N_37671,N_33467);
nand U45418 (N_45418,N_35430,N_38384);
or U45419 (N_45419,N_32743,N_36820);
and U45420 (N_45420,N_36552,N_30361);
and U45421 (N_45421,N_32339,N_37983);
and U45422 (N_45422,N_33551,N_33757);
nand U45423 (N_45423,N_35459,N_37180);
and U45424 (N_45424,N_36525,N_33412);
or U45425 (N_45425,N_39236,N_38133);
and U45426 (N_45426,N_30755,N_32765);
and U45427 (N_45427,N_31261,N_38034);
and U45428 (N_45428,N_39581,N_35446);
and U45429 (N_45429,N_35554,N_37075);
or U45430 (N_45430,N_32869,N_38397);
and U45431 (N_45431,N_33366,N_37239);
xor U45432 (N_45432,N_39635,N_36934);
nand U45433 (N_45433,N_39760,N_38866);
nand U45434 (N_45434,N_30544,N_38890);
or U45435 (N_45435,N_31637,N_36498);
nor U45436 (N_45436,N_37938,N_34902);
or U45437 (N_45437,N_37925,N_38380);
or U45438 (N_45438,N_39889,N_37790);
and U45439 (N_45439,N_39442,N_31054);
nand U45440 (N_45440,N_31075,N_31204);
nand U45441 (N_45441,N_36431,N_33935);
nor U45442 (N_45442,N_37428,N_33785);
and U45443 (N_45443,N_35369,N_39120);
xor U45444 (N_45444,N_35630,N_31156);
nand U45445 (N_45445,N_35271,N_30519);
and U45446 (N_45446,N_31894,N_36896);
and U45447 (N_45447,N_37637,N_32826);
nand U45448 (N_45448,N_30807,N_31538);
or U45449 (N_45449,N_30334,N_30090);
nor U45450 (N_45450,N_33481,N_36399);
nor U45451 (N_45451,N_30201,N_39808);
and U45452 (N_45452,N_32739,N_36456);
nand U45453 (N_45453,N_32605,N_35726);
nand U45454 (N_45454,N_37398,N_38242);
or U45455 (N_45455,N_31741,N_38057);
xor U45456 (N_45456,N_34434,N_33404);
or U45457 (N_45457,N_34639,N_39869);
nand U45458 (N_45458,N_38188,N_38690);
nand U45459 (N_45459,N_33382,N_36110);
nand U45460 (N_45460,N_36928,N_33327);
xor U45461 (N_45461,N_37283,N_30610);
nand U45462 (N_45462,N_38126,N_39532);
or U45463 (N_45463,N_36911,N_38737);
or U45464 (N_45464,N_38775,N_39108);
nand U45465 (N_45465,N_39111,N_30865);
xnor U45466 (N_45466,N_39534,N_37514);
nand U45467 (N_45467,N_39602,N_36844);
nor U45468 (N_45468,N_38739,N_34963);
nor U45469 (N_45469,N_35114,N_31112);
nor U45470 (N_45470,N_35963,N_38118);
nand U45471 (N_45471,N_30942,N_39597);
and U45472 (N_45472,N_35610,N_35322);
nand U45473 (N_45473,N_33944,N_39657);
or U45474 (N_45474,N_31732,N_33602);
xor U45475 (N_45475,N_37717,N_30484);
and U45476 (N_45476,N_36072,N_30334);
nand U45477 (N_45477,N_36198,N_35783);
nand U45478 (N_45478,N_34867,N_37199);
or U45479 (N_45479,N_33348,N_30920);
nand U45480 (N_45480,N_33428,N_38063);
nand U45481 (N_45481,N_33017,N_31517);
xor U45482 (N_45482,N_34779,N_36379);
or U45483 (N_45483,N_32558,N_38051);
or U45484 (N_45484,N_34386,N_39539);
nor U45485 (N_45485,N_31299,N_30887);
and U45486 (N_45486,N_33359,N_37259);
and U45487 (N_45487,N_38500,N_33057);
or U45488 (N_45488,N_35592,N_31368);
nor U45489 (N_45489,N_35695,N_33128);
nor U45490 (N_45490,N_31754,N_35619);
nand U45491 (N_45491,N_33902,N_36779);
and U45492 (N_45492,N_33873,N_34373);
xnor U45493 (N_45493,N_34670,N_31171);
nand U45494 (N_45494,N_31580,N_38338);
nor U45495 (N_45495,N_39823,N_33500);
and U45496 (N_45496,N_37741,N_36247);
nor U45497 (N_45497,N_32609,N_33189);
or U45498 (N_45498,N_38407,N_34564);
and U45499 (N_45499,N_30367,N_36073);
and U45500 (N_45500,N_35965,N_36637);
nor U45501 (N_45501,N_33491,N_32868);
and U45502 (N_45502,N_34758,N_31660);
or U45503 (N_45503,N_35953,N_32399);
nor U45504 (N_45504,N_32734,N_30875);
nand U45505 (N_45505,N_35454,N_38181);
or U45506 (N_45506,N_34487,N_39692);
and U45507 (N_45507,N_30149,N_31841);
and U45508 (N_45508,N_33042,N_37653);
and U45509 (N_45509,N_38181,N_31466);
or U45510 (N_45510,N_32541,N_33878);
or U45511 (N_45511,N_32912,N_30469);
or U45512 (N_45512,N_35309,N_36970);
or U45513 (N_45513,N_30746,N_31775);
xnor U45514 (N_45514,N_35558,N_34288);
nand U45515 (N_45515,N_35754,N_30781);
nor U45516 (N_45516,N_39409,N_37904);
nor U45517 (N_45517,N_39001,N_39160);
nor U45518 (N_45518,N_36773,N_33135);
xnor U45519 (N_45519,N_35538,N_31825);
nand U45520 (N_45520,N_31930,N_38595);
xnor U45521 (N_45521,N_32043,N_30253);
nor U45522 (N_45522,N_35788,N_31497);
or U45523 (N_45523,N_30394,N_34253);
nand U45524 (N_45524,N_32710,N_32873);
nand U45525 (N_45525,N_32360,N_31470);
and U45526 (N_45526,N_32747,N_30810);
nand U45527 (N_45527,N_36216,N_38359);
and U45528 (N_45528,N_32568,N_35153);
and U45529 (N_45529,N_37411,N_39898);
and U45530 (N_45530,N_37904,N_30023);
nand U45531 (N_45531,N_37790,N_30231);
xnor U45532 (N_45532,N_33746,N_30145);
nor U45533 (N_45533,N_37930,N_33210);
nor U45534 (N_45534,N_30743,N_37396);
or U45535 (N_45535,N_33088,N_30856);
xnor U45536 (N_45536,N_34769,N_37164);
and U45537 (N_45537,N_30073,N_36180);
and U45538 (N_45538,N_34865,N_32977);
and U45539 (N_45539,N_34152,N_31632);
nand U45540 (N_45540,N_37611,N_34916);
nor U45541 (N_45541,N_30481,N_34443);
nand U45542 (N_45542,N_36106,N_39840);
nor U45543 (N_45543,N_33961,N_36465);
and U45544 (N_45544,N_31771,N_38651);
nand U45545 (N_45545,N_32143,N_39549);
or U45546 (N_45546,N_38641,N_34589);
nand U45547 (N_45547,N_39718,N_36130);
or U45548 (N_45548,N_38160,N_31122);
nand U45549 (N_45549,N_31395,N_32326);
nor U45550 (N_45550,N_38623,N_30137);
nand U45551 (N_45551,N_38328,N_38414);
and U45552 (N_45552,N_30351,N_39901);
or U45553 (N_45553,N_35017,N_37078);
nand U45554 (N_45554,N_36918,N_34486);
and U45555 (N_45555,N_30870,N_36906);
or U45556 (N_45556,N_34200,N_32477);
xor U45557 (N_45557,N_37880,N_31908);
nand U45558 (N_45558,N_30499,N_30051);
nor U45559 (N_45559,N_33909,N_31869);
nand U45560 (N_45560,N_37703,N_39426);
or U45561 (N_45561,N_39929,N_38230);
nor U45562 (N_45562,N_30610,N_39755);
xor U45563 (N_45563,N_35355,N_34175);
and U45564 (N_45564,N_30030,N_32147);
nor U45565 (N_45565,N_32750,N_31313);
nor U45566 (N_45566,N_31541,N_39678);
or U45567 (N_45567,N_39045,N_37203);
and U45568 (N_45568,N_37535,N_31335);
nor U45569 (N_45569,N_31312,N_39002);
nor U45570 (N_45570,N_39350,N_33361);
or U45571 (N_45571,N_34194,N_35101);
nor U45572 (N_45572,N_34990,N_35290);
nand U45573 (N_45573,N_35529,N_38078);
nand U45574 (N_45574,N_33322,N_33977);
or U45575 (N_45575,N_30466,N_37299);
and U45576 (N_45576,N_38823,N_36195);
xor U45577 (N_45577,N_37066,N_35640);
nor U45578 (N_45578,N_34364,N_34535);
xor U45579 (N_45579,N_38075,N_33770);
nor U45580 (N_45580,N_35523,N_31293);
and U45581 (N_45581,N_30606,N_30008);
nand U45582 (N_45582,N_35412,N_34991);
nand U45583 (N_45583,N_34002,N_37536);
or U45584 (N_45584,N_30853,N_39917);
nand U45585 (N_45585,N_32311,N_31811);
and U45586 (N_45586,N_32590,N_34039);
or U45587 (N_45587,N_37885,N_33808);
nor U45588 (N_45588,N_38861,N_34737);
xor U45589 (N_45589,N_30377,N_36452);
xor U45590 (N_45590,N_31920,N_34360);
and U45591 (N_45591,N_31829,N_39770);
or U45592 (N_45592,N_32869,N_35495);
nand U45593 (N_45593,N_30082,N_33401);
nand U45594 (N_45594,N_34166,N_30188);
and U45595 (N_45595,N_30273,N_39636);
xor U45596 (N_45596,N_34021,N_36012);
nand U45597 (N_45597,N_30949,N_35210);
nor U45598 (N_45598,N_38731,N_32054);
nor U45599 (N_45599,N_36259,N_38706);
nor U45600 (N_45600,N_34109,N_39634);
nor U45601 (N_45601,N_31601,N_32589);
and U45602 (N_45602,N_33785,N_32414);
or U45603 (N_45603,N_34210,N_31552);
nor U45604 (N_45604,N_39300,N_38202);
nand U45605 (N_45605,N_30914,N_34259);
nand U45606 (N_45606,N_34955,N_39804);
nor U45607 (N_45607,N_34145,N_33147);
nand U45608 (N_45608,N_34903,N_32117);
nor U45609 (N_45609,N_32048,N_34268);
or U45610 (N_45610,N_35463,N_33519);
and U45611 (N_45611,N_36096,N_37183);
xor U45612 (N_45612,N_34641,N_36564);
nand U45613 (N_45613,N_32949,N_33714);
nor U45614 (N_45614,N_33324,N_39599);
or U45615 (N_45615,N_31765,N_31387);
nand U45616 (N_45616,N_31988,N_33302);
nor U45617 (N_45617,N_35028,N_31879);
and U45618 (N_45618,N_33708,N_32980);
and U45619 (N_45619,N_32077,N_33153);
nand U45620 (N_45620,N_34986,N_31640);
nor U45621 (N_45621,N_31289,N_37966);
or U45622 (N_45622,N_30422,N_39159);
nor U45623 (N_45623,N_39916,N_38399);
nand U45624 (N_45624,N_32972,N_36335);
nand U45625 (N_45625,N_34248,N_39861);
nand U45626 (N_45626,N_34426,N_33909);
xnor U45627 (N_45627,N_35053,N_38442);
or U45628 (N_45628,N_37317,N_36104);
and U45629 (N_45629,N_39906,N_32026);
and U45630 (N_45630,N_30209,N_33953);
or U45631 (N_45631,N_30713,N_34125);
and U45632 (N_45632,N_37396,N_39177);
nor U45633 (N_45633,N_32472,N_38866);
and U45634 (N_45634,N_30208,N_32781);
or U45635 (N_45635,N_35382,N_36159);
nor U45636 (N_45636,N_35811,N_30622);
nand U45637 (N_45637,N_33446,N_36043);
nor U45638 (N_45638,N_33750,N_33747);
or U45639 (N_45639,N_31199,N_36984);
and U45640 (N_45640,N_37946,N_32226);
nand U45641 (N_45641,N_30107,N_36711);
nor U45642 (N_45642,N_34255,N_33363);
and U45643 (N_45643,N_38526,N_38635);
and U45644 (N_45644,N_31645,N_31428);
nand U45645 (N_45645,N_39470,N_35880);
or U45646 (N_45646,N_32756,N_31626);
or U45647 (N_45647,N_39608,N_38858);
xnor U45648 (N_45648,N_34645,N_32816);
nand U45649 (N_45649,N_35477,N_38629);
nor U45650 (N_45650,N_30662,N_38530);
nand U45651 (N_45651,N_31107,N_39730);
and U45652 (N_45652,N_31500,N_37483);
nand U45653 (N_45653,N_33688,N_30483);
and U45654 (N_45654,N_37286,N_35604);
nor U45655 (N_45655,N_31307,N_33459);
nand U45656 (N_45656,N_35068,N_32857);
xor U45657 (N_45657,N_37609,N_35097);
and U45658 (N_45658,N_39764,N_30244);
or U45659 (N_45659,N_35310,N_35172);
and U45660 (N_45660,N_34389,N_33591);
nand U45661 (N_45661,N_32705,N_34360);
or U45662 (N_45662,N_36754,N_38550);
nand U45663 (N_45663,N_33390,N_32656);
and U45664 (N_45664,N_34899,N_37624);
nor U45665 (N_45665,N_37478,N_39870);
or U45666 (N_45666,N_33843,N_34395);
nand U45667 (N_45667,N_37700,N_36013);
or U45668 (N_45668,N_37663,N_38948);
and U45669 (N_45669,N_32797,N_35516);
and U45670 (N_45670,N_30426,N_31827);
and U45671 (N_45671,N_37859,N_31560);
and U45672 (N_45672,N_39057,N_37200);
and U45673 (N_45673,N_35279,N_30985);
or U45674 (N_45674,N_38006,N_39005);
nor U45675 (N_45675,N_35487,N_39798);
and U45676 (N_45676,N_34437,N_38325);
and U45677 (N_45677,N_39710,N_39186);
nand U45678 (N_45678,N_37707,N_35655);
nand U45679 (N_45679,N_30834,N_39222);
nand U45680 (N_45680,N_32984,N_30431);
and U45681 (N_45681,N_37335,N_31110);
and U45682 (N_45682,N_33825,N_34421);
xor U45683 (N_45683,N_31929,N_39390);
nand U45684 (N_45684,N_32494,N_37169);
nor U45685 (N_45685,N_31628,N_37258);
or U45686 (N_45686,N_30772,N_37495);
nand U45687 (N_45687,N_36313,N_30019);
and U45688 (N_45688,N_34032,N_34068);
or U45689 (N_45689,N_36910,N_39924);
or U45690 (N_45690,N_32246,N_39033);
or U45691 (N_45691,N_32519,N_34875);
nor U45692 (N_45692,N_33493,N_31454);
nand U45693 (N_45693,N_30975,N_39722);
and U45694 (N_45694,N_37549,N_32745);
nand U45695 (N_45695,N_34095,N_35070);
nor U45696 (N_45696,N_31166,N_35656);
and U45697 (N_45697,N_37432,N_33605);
and U45698 (N_45698,N_39130,N_37029);
nor U45699 (N_45699,N_31392,N_30017);
and U45700 (N_45700,N_39644,N_30051);
or U45701 (N_45701,N_37856,N_30648);
xor U45702 (N_45702,N_37588,N_37649);
and U45703 (N_45703,N_36054,N_36910);
nor U45704 (N_45704,N_35563,N_37211);
and U45705 (N_45705,N_38627,N_37106);
and U45706 (N_45706,N_33727,N_36781);
and U45707 (N_45707,N_37036,N_35712);
nor U45708 (N_45708,N_37109,N_33036);
nand U45709 (N_45709,N_34678,N_31089);
nor U45710 (N_45710,N_39004,N_30286);
or U45711 (N_45711,N_32579,N_35846);
nand U45712 (N_45712,N_31602,N_30947);
or U45713 (N_45713,N_31086,N_36591);
nor U45714 (N_45714,N_35977,N_33895);
nor U45715 (N_45715,N_31515,N_33517);
and U45716 (N_45716,N_31632,N_30689);
nor U45717 (N_45717,N_31896,N_39886);
and U45718 (N_45718,N_36049,N_39162);
nand U45719 (N_45719,N_30131,N_33687);
xnor U45720 (N_45720,N_36868,N_30193);
or U45721 (N_45721,N_38353,N_37939);
and U45722 (N_45722,N_39720,N_39460);
nor U45723 (N_45723,N_36827,N_39719);
nor U45724 (N_45724,N_34323,N_30959);
nor U45725 (N_45725,N_31151,N_33266);
xnor U45726 (N_45726,N_30471,N_34672);
or U45727 (N_45727,N_37718,N_34347);
or U45728 (N_45728,N_39381,N_35061);
nand U45729 (N_45729,N_30299,N_38015);
and U45730 (N_45730,N_35879,N_36784);
or U45731 (N_45731,N_35807,N_38136);
or U45732 (N_45732,N_37068,N_38168);
nand U45733 (N_45733,N_34130,N_38953);
nor U45734 (N_45734,N_32794,N_35458);
and U45735 (N_45735,N_32335,N_34827);
xnor U45736 (N_45736,N_31828,N_35513);
and U45737 (N_45737,N_30472,N_33404);
nand U45738 (N_45738,N_35675,N_33040);
nor U45739 (N_45739,N_32110,N_39183);
xnor U45740 (N_45740,N_39967,N_33246);
and U45741 (N_45741,N_32701,N_35024);
nand U45742 (N_45742,N_31759,N_31213);
nand U45743 (N_45743,N_34855,N_35078);
and U45744 (N_45744,N_31335,N_39811);
or U45745 (N_45745,N_35500,N_31906);
or U45746 (N_45746,N_38190,N_35283);
nand U45747 (N_45747,N_30608,N_31618);
nor U45748 (N_45748,N_35851,N_36748);
nand U45749 (N_45749,N_33752,N_35735);
nor U45750 (N_45750,N_37849,N_34844);
xnor U45751 (N_45751,N_35492,N_37468);
nor U45752 (N_45752,N_31686,N_35513);
nor U45753 (N_45753,N_39027,N_36673);
nor U45754 (N_45754,N_33627,N_30397);
or U45755 (N_45755,N_32419,N_37632);
nor U45756 (N_45756,N_30962,N_37851);
or U45757 (N_45757,N_37401,N_38607);
nand U45758 (N_45758,N_36780,N_30833);
nor U45759 (N_45759,N_35384,N_36529);
nor U45760 (N_45760,N_31829,N_30037);
and U45761 (N_45761,N_36465,N_36648);
nand U45762 (N_45762,N_39671,N_39044);
and U45763 (N_45763,N_36988,N_34047);
nor U45764 (N_45764,N_35104,N_34207);
or U45765 (N_45765,N_36175,N_35944);
nor U45766 (N_45766,N_38480,N_34665);
nand U45767 (N_45767,N_37311,N_35875);
or U45768 (N_45768,N_39100,N_38562);
nand U45769 (N_45769,N_31967,N_33200);
or U45770 (N_45770,N_33280,N_32604);
or U45771 (N_45771,N_37627,N_38885);
and U45772 (N_45772,N_30211,N_39620);
or U45773 (N_45773,N_35635,N_33068);
nand U45774 (N_45774,N_35983,N_33405);
and U45775 (N_45775,N_36782,N_37784);
nand U45776 (N_45776,N_33593,N_30013);
xnor U45777 (N_45777,N_32910,N_35040);
and U45778 (N_45778,N_36349,N_37543);
and U45779 (N_45779,N_33746,N_33471);
and U45780 (N_45780,N_36403,N_34404);
and U45781 (N_45781,N_32841,N_30960);
and U45782 (N_45782,N_34889,N_38865);
nor U45783 (N_45783,N_36403,N_36173);
xnor U45784 (N_45784,N_35412,N_30411);
and U45785 (N_45785,N_31683,N_34385);
or U45786 (N_45786,N_37130,N_30600);
nor U45787 (N_45787,N_39890,N_31752);
xnor U45788 (N_45788,N_33050,N_38916);
and U45789 (N_45789,N_35230,N_32711);
and U45790 (N_45790,N_39478,N_32463);
xor U45791 (N_45791,N_35256,N_31572);
and U45792 (N_45792,N_39193,N_37237);
nor U45793 (N_45793,N_36748,N_37726);
nand U45794 (N_45794,N_34140,N_32941);
nor U45795 (N_45795,N_33491,N_32171);
or U45796 (N_45796,N_35766,N_36689);
xor U45797 (N_45797,N_33391,N_34867);
nand U45798 (N_45798,N_35687,N_35189);
or U45799 (N_45799,N_37421,N_33838);
and U45800 (N_45800,N_33722,N_39491);
nor U45801 (N_45801,N_36531,N_35850);
nand U45802 (N_45802,N_33142,N_37921);
and U45803 (N_45803,N_38230,N_37629);
nor U45804 (N_45804,N_30818,N_39357);
nor U45805 (N_45805,N_36796,N_32095);
and U45806 (N_45806,N_35557,N_34863);
and U45807 (N_45807,N_31540,N_30446);
or U45808 (N_45808,N_31580,N_39416);
nor U45809 (N_45809,N_30040,N_31265);
xnor U45810 (N_45810,N_30024,N_30503);
nor U45811 (N_45811,N_34652,N_30148);
and U45812 (N_45812,N_30397,N_37716);
or U45813 (N_45813,N_33023,N_35218);
nor U45814 (N_45814,N_39099,N_38101);
and U45815 (N_45815,N_33131,N_35728);
and U45816 (N_45816,N_36567,N_36868);
or U45817 (N_45817,N_36097,N_39517);
nor U45818 (N_45818,N_38347,N_30197);
nand U45819 (N_45819,N_34967,N_38363);
xnor U45820 (N_45820,N_35639,N_38624);
or U45821 (N_45821,N_30870,N_35376);
xor U45822 (N_45822,N_31002,N_39724);
and U45823 (N_45823,N_36942,N_38124);
and U45824 (N_45824,N_30471,N_30659);
and U45825 (N_45825,N_36192,N_38416);
or U45826 (N_45826,N_38007,N_36565);
or U45827 (N_45827,N_32294,N_33370);
and U45828 (N_45828,N_38435,N_30843);
nand U45829 (N_45829,N_32717,N_36432);
nor U45830 (N_45830,N_39902,N_36874);
nor U45831 (N_45831,N_36813,N_33502);
xor U45832 (N_45832,N_37575,N_30350);
or U45833 (N_45833,N_39626,N_32790);
and U45834 (N_45834,N_38341,N_32354);
and U45835 (N_45835,N_34547,N_37086);
nor U45836 (N_45836,N_32548,N_36150);
nand U45837 (N_45837,N_34893,N_39912);
nand U45838 (N_45838,N_32332,N_30102);
nor U45839 (N_45839,N_32241,N_33041);
xor U45840 (N_45840,N_35746,N_31126);
nor U45841 (N_45841,N_33627,N_32013);
nor U45842 (N_45842,N_30689,N_39483);
xor U45843 (N_45843,N_35437,N_35855);
nor U45844 (N_45844,N_32429,N_37104);
or U45845 (N_45845,N_36087,N_31536);
nor U45846 (N_45846,N_32612,N_31753);
or U45847 (N_45847,N_34887,N_39631);
nor U45848 (N_45848,N_32232,N_37871);
xor U45849 (N_45849,N_36775,N_36463);
or U45850 (N_45850,N_33171,N_38471);
xnor U45851 (N_45851,N_36646,N_34706);
or U45852 (N_45852,N_30750,N_30330);
or U45853 (N_45853,N_32907,N_37812);
and U45854 (N_45854,N_35118,N_39243);
and U45855 (N_45855,N_35963,N_38718);
xor U45856 (N_45856,N_32299,N_39206);
nor U45857 (N_45857,N_31937,N_38505);
or U45858 (N_45858,N_33379,N_31496);
nand U45859 (N_45859,N_35940,N_32627);
or U45860 (N_45860,N_35069,N_39985);
nor U45861 (N_45861,N_37100,N_33808);
nand U45862 (N_45862,N_31957,N_39734);
nor U45863 (N_45863,N_33722,N_35536);
xor U45864 (N_45864,N_33767,N_37173);
xnor U45865 (N_45865,N_37064,N_36840);
nand U45866 (N_45866,N_30309,N_34417);
or U45867 (N_45867,N_34697,N_36430);
nand U45868 (N_45868,N_33917,N_36560);
nand U45869 (N_45869,N_30184,N_30866);
nor U45870 (N_45870,N_31066,N_31332);
and U45871 (N_45871,N_35652,N_38747);
xor U45872 (N_45872,N_33066,N_36797);
nor U45873 (N_45873,N_35559,N_30259);
and U45874 (N_45874,N_35224,N_35604);
nand U45875 (N_45875,N_30169,N_30662);
and U45876 (N_45876,N_33008,N_33423);
nand U45877 (N_45877,N_33533,N_33776);
nand U45878 (N_45878,N_37601,N_31521);
xnor U45879 (N_45879,N_32976,N_35122);
and U45880 (N_45880,N_38619,N_31171);
and U45881 (N_45881,N_33167,N_37399);
nor U45882 (N_45882,N_37336,N_32832);
or U45883 (N_45883,N_32809,N_36726);
and U45884 (N_45884,N_38985,N_38739);
nand U45885 (N_45885,N_38556,N_38956);
nand U45886 (N_45886,N_34627,N_38700);
or U45887 (N_45887,N_35148,N_32947);
nor U45888 (N_45888,N_30499,N_38244);
or U45889 (N_45889,N_37937,N_38447);
or U45890 (N_45890,N_39006,N_38503);
nor U45891 (N_45891,N_35022,N_37430);
or U45892 (N_45892,N_38050,N_30427);
nand U45893 (N_45893,N_37962,N_34800);
nor U45894 (N_45894,N_33521,N_39297);
or U45895 (N_45895,N_35521,N_39535);
and U45896 (N_45896,N_30138,N_39237);
and U45897 (N_45897,N_30971,N_32847);
and U45898 (N_45898,N_37284,N_32917);
nand U45899 (N_45899,N_33638,N_37561);
or U45900 (N_45900,N_33426,N_38359);
or U45901 (N_45901,N_30144,N_38284);
nor U45902 (N_45902,N_36545,N_36025);
and U45903 (N_45903,N_37988,N_39158);
and U45904 (N_45904,N_30894,N_36303);
and U45905 (N_45905,N_38576,N_35765);
or U45906 (N_45906,N_36912,N_34122);
or U45907 (N_45907,N_35362,N_33449);
and U45908 (N_45908,N_31696,N_36381);
nor U45909 (N_45909,N_34962,N_31681);
and U45910 (N_45910,N_38050,N_39022);
nor U45911 (N_45911,N_32981,N_39542);
nor U45912 (N_45912,N_39833,N_32203);
nor U45913 (N_45913,N_36858,N_38911);
xor U45914 (N_45914,N_35002,N_35201);
nand U45915 (N_45915,N_38110,N_35211);
nor U45916 (N_45916,N_39614,N_31036);
nor U45917 (N_45917,N_38043,N_36964);
nor U45918 (N_45918,N_31577,N_37399);
nor U45919 (N_45919,N_31571,N_32963);
nand U45920 (N_45920,N_31591,N_36839);
and U45921 (N_45921,N_35735,N_38573);
or U45922 (N_45922,N_38898,N_34202);
and U45923 (N_45923,N_36827,N_38864);
or U45924 (N_45924,N_39798,N_38496);
nand U45925 (N_45925,N_30084,N_39260);
and U45926 (N_45926,N_35693,N_31538);
and U45927 (N_45927,N_37707,N_33610);
xor U45928 (N_45928,N_37538,N_36325);
nand U45929 (N_45929,N_36861,N_33362);
or U45930 (N_45930,N_30969,N_32811);
nand U45931 (N_45931,N_35300,N_35996);
or U45932 (N_45932,N_36522,N_31196);
and U45933 (N_45933,N_34879,N_32169);
or U45934 (N_45934,N_33195,N_35973);
or U45935 (N_45935,N_30144,N_33783);
nor U45936 (N_45936,N_39156,N_37682);
and U45937 (N_45937,N_38565,N_37157);
and U45938 (N_45938,N_31070,N_37757);
and U45939 (N_45939,N_39288,N_35938);
nor U45940 (N_45940,N_36304,N_37950);
or U45941 (N_45941,N_36036,N_31235);
xor U45942 (N_45942,N_35315,N_33119);
xnor U45943 (N_45943,N_35848,N_36996);
nand U45944 (N_45944,N_30533,N_36125);
and U45945 (N_45945,N_37643,N_37387);
or U45946 (N_45946,N_34198,N_30769);
and U45947 (N_45947,N_33694,N_34034);
and U45948 (N_45948,N_38226,N_30219);
or U45949 (N_45949,N_30250,N_33409);
and U45950 (N_45950,N_34911,N_30204);
or U45951 (N_45951,N_31151,N_33800);
nand U45952 (N_45952,N_38266,N_36297);
nor U45953 (N_45953,N_36269,N_31224);
or U45954 (N_45954,N_36107,N_34964);
nand U45955 (N_45955,N_39997,N_39642);
xor U45956 (N_45956,N_32177,N_39113);
and U45957 (N_45957,N_35355,N_34702);
nor U45958 (N_45958,N_37660,N_35958);
or U45959 (N_45959,N_35118,N_37823);
nand U45960 (N_45960,N_37492,N_33110);
xor U45961 (N_45961,N_38431,N_32326);
nand U45962 (N_45962,N_34471,N_33956);
or U45963 (N_45963,N_30374,N_30880);
xnor U45964 (N_45964,N_34973,N_37712);
nor U45965 (N_45965,N_32159,N_31595);
and U45966 (N_45966,N_35054,N_30627);
xnor U45967 (N_45967,N_32983,N_36855);
and U45968 (N_45968,N_37491,N_31027);
and U45969 (N_45969,N_39222,N_36347);
nor U45970 (N_45970,N_31859,N_38730);
nand U45971 (N_45971,N_37196,N_35470);
xnor U45972 (N_45972,N_35246,N_35685);
nand U45973 (N_45973,N_32251,N_33251);
or U45974 (N_45974,N_38929,N_32647);
xor U45975 (N_45975,N_38123,N_31062);
nand U45976 (N_45976,N_38071,N_32473);
and U45977 (N_45977,N_30363,N_31479);
or U45978 (N_45978,N_37738,N_38102);
or U45979 (N_45979,N_33238,N_32545);
nor U45980 (N_45980,N_36407,N_31133);
and U45981 (N_45981,N_31424,N_37668);
nor U45982 (N_45982,N_33548,N_30827);
or U45983 (N_45983,N_37618,N_34339);
or U45984 (N_45984,N_35458,N_37227);
or U45985 (N_45985,N_31575,N_33213);
xnor U45986 (N_45986,N_35878,N_30560);
nor U45987 (N_45987,N_37162,N_36487);
or U45988 (N_45988,N_33547,N_31928);
nand U45989 (N_45989,N_35743,N_30586);
nor U45990 (N_45990,N_30623,N_30698);
and U45991 (N_45991,N_32934,N_33072);
or U45992 (N_45992,N_39366,N_38501);
and U45993 (N_45993,N_38755,N_31993);
nor U45994 (N_45994,N_31104,N_38833);
nor U45995 (N_45995,N_36509,N_38107);
and U45996 (N_45996,N_38577,N_32074);
nor U45997 (N_45997,N_37595,N_39251);
or U45998 (N_45998,N_34204,N_33380);
and U45999 (N_45999,N_32120,N_36609);
nor U46000 (N_46000,N_35547,N_30305);
or U46001 (N_46001,N_33870,N_37875);
and U46002 (N_46002,N_34224,N_35442);
nand U46003 (N_46003,N_34178,N_39640);
and U46004 (N_46004,N_38767,N_31523);
nand U46005 (N_46005,N_33207,N_35802);
or U46006 (N_46006,N_33183,N_39875);
nor U46007 (N_46007,N_39122,N_39501);
nand U46008 (N_46008,N_34874,N_32669);
nand U46009 (N_46009,N_32446,N_31729);
nand U46010 (N_46010,N_35305,N_33667);
nand U46011 (N_46011,N_33977,N_35973);
and U46012 (N_46012,N_37683,N_31056);
nor U46013 (N_46013,N_31871,N_38271);
nor U46014 (N_46014,N_33273,N_38482);
and U46015 (N_46015,N_39653,N_36274);
nand U46016 (N_46016,N_35995,N_34087);
xor U46017 (N_46017,N_35648,N_34760);
and U46018 (N_46018,N_33602,N_35998);
and U46019 (N_46019,N_39279,N_33534);
or U46020 (N_46020,N_31213,N_34885);
or U46021 (N_46021,N_35854,N_32808);
or U46022 (N_46022,N_34538,N_38988);
and U46023 (N_46023,N_33683,N_31262);
nand U46024 (N_46024,N_35917,N_31909);
nand U46025 (N_46025,N_32462,N_36869);
and U46026 (N_46026,N_33655,N_34731);
and U46027 (N_46027,N_30385,N_33406);
and U46028 (N_46028,N_38316,N_32785);
nor U46029 (N_46029,N_30008,N_34995);
nand U46030 (N_46030,N_30293,N_39961);
nor U46031 (N_46031,N_38636,N_34755);
or U46032 (N_46032,N_36315,N_39639);
or U46033 (N_46033,N_37155,N_36572);
nand U46034 (N_46034,N_30319,N_36819);
or U46035 (N_46035,N_36878,N_37669);
nor U46036 (N_46036,N_35016,N_36764);
or U46037 (N_46037,N_34154,N_35373);
nand U46038 (N_46038,N_34566,N_39523);
and U46039 (N_46039,N_39126,N_32313);
or U46040 (N_46040,N_39678,N_38059);
nor U46041 (N_46041,N_38197,N_33637);
and U46042 (N_46042,N_32502,N_34417);
or U46043 (N_46043,N_35691,N_30769);
and U46044 (N_46044,N_31813,N_32407);
nor U46045 (N_46045,N_31031,N_31641);
nand U46046 (N_46046,N_36814,N_35321);
nor U46047 (N_46047,N_33167,N_34800);
nand U46048 (N_46048,N_36458,N_39688);
xnor U46049 (N_46049,N_39819,N_30134);
or U46050 (N_46050,N_32686,N_35380);
xnor U46051 (N_46051,N_34084,N_30773);
or U46052 (N_46052,N_36729,N_35168);
nand U46053 (N_46053,N_38908,N_39482);
nand U46054 (N_46054,N_39450,N_38622);
or U46055 (N_46055,N_37728,N_35906);
nand U46056 (N_46056,N_30692,N_33807);
nand U46057 (N_46057,N_31732,N_37151);
and U46058 (N_46058,N_35288,N_35641);
or U46059 (N_46059,N_36213,N_37656);
nand U46060 (N_46060,N_39664,N_34210);
and U46061 (N_46061,N_38995,N_31444);
and U46062 (N_46062,N_35637,N_31574);
and U46063 (N_46063,N_33505,N_35068);
nor U46064 (N_46064,N_30568,N_33066);
or U46065 (N_46065,N_35446,N_35925);
or U46066 (N_46066,N_39686,N_33180);
nand U46067 (N_46067,N_37268,N_34680);
and U46068 (N_46068,N_39043,N_39621);
and U46069 (N_46069,N_33122,N_32923);
nand U46070 (N_46070,N_32270,N_31413);
xor U46071 (N_46071,N_37163,N_32869);
nor U46072 (N_46072,N_34692,N_34875);
nor U46073 (N_46073,N_36901,N_31500);
nand U46074 (N_46074,N_38956,N_37761);
or U46075 (N_46075,N_33303,N_37319);
nor U46076 (N_46076,N_35318,N_30005);
nor U46077 (N_46077,N_39679,N_38518);
xnor U46078 (N_46078,N_35040,N_33773);
nand U46079 (N_46079,N_35985,N_37413);
xor U46080 (N_46080,N_32744,N_31358);
nor U46081 (N_46081,N_33781,N_33802);
and U46082 (N_46082,N_32471,N_31054);
nand U46083 (N_46083,N_33364,N_31250);
and U46084 (N_46084,N_35123,N_35162);
nor U46085 (N_46085,N_35002,N_30571);
nand U46086 (N_46086,N_31357,N_38136);
and U46087 (N_46087,N_39091,N_33870);
and U46088 (N_46088,N_34155,N_37042);
nand U46089 (N_46089,N_33645,N_35097);
or U46090 (N_46090,N_33679,N_37316);
xor U46091 (N_46091,N_32872,N_34929);
nor U46092 (N_46092,N_35427,N_33484);
and U46093 (N_46093,N_34754,N_31253);
or U46094 (N_46094,N_36689,N_36765);
or U46095 (N_46095,N_38940,N_36634);
nand U46096 (N_46096,N_39147,N_32345);
nor U46097 (N_46097,N_38422,N_35190);
or U46098 (N_46098,N_31537,N_30180);
and U46099 (N_46099,N_37351,N_36455);
nor U46100 (N_46100,N_32247,N_31912);
and U46101 (N_46101,N_36162,N_36001);
nor U46102 (N_46102,N_36755,N_33414);
nand U46103 (N_46103,N_37864,N_33235);
nand U46104 (N_46104,N_31438,N_37103);
or U46105 (N_46105,N_39869,N_32498);
xor U46106 (N_46106,N_31931,N_37070);
xor U46107 (N_46107,N_34253,N_39766);
nand U46108 (N_46108,N_36371,N_36702);
nand U46109 (N_46109,N_39010,N_39700);
xor U46110 (N_46110,N_30808,N_38252);
or U46111 (N_46111,N_38929,N_31798);
nor U46112 (N_46112,N_39699,N_35065);
or U46113 (N_46113,N_35708,N_32252);
nand U46114 (N_46114,N_31036,N_39312);
or U46115 (N_46115,N_36949,N_36789);
nor U46116 (N_46116,N_36463,N_35803);
nor U46117 (N_46117,N_36719,N_35948);
or U46118 (N_46118,N_30355,N_36777);
or U46119 (N_46119,N_34301,N_38054);
and U46120 (N_46120,N_32021,N_31128);
xnor U46121 (N_46121,N_36490,N_30377);
and U46122 (N_46122,N_30376,N_37395);
or U46123 (N_46123,N_36159,N_31312);
nor U46124 (N_46124,N_36227,N_39142);
or U46125 (N_46125,N_38540,N_38481);
and U46126 (N_46126,N_33944,N_34181);
or U46127 (N_46127,N_39544,N_31681);
and U46128 (N_46128,N_36515,N_35940);
xor U46129 (N_46129,N_39871,N_38326);
nor U46130 (N_46130,N_39068,N_36960);
nor U46131 (N_46131,N_37530,N_38499);
nor U46132 (N_46132,N_35739,N_34091);
and U46133 (N_46133,N_39487,N_31768);
xnor U46134 (N_46134,N_36017,N_33252);
nand U46135 (N_46135,N_35738,N_39693);
nand U46136 (N_46136,N_37407,N_36550);
and U46137 (N_46137,N_34356,N_39921);
nor U46138 (N_46138,N_36797,N_38719);
xnor U46139 (N_46139,N_33264,N_34580);
or U46140 (N_46140,N_33633,N_31944);
nand U46141 (N_46141,N_39444,N_34834);
nor U46142 (N_46142,N_35667,N_38646);
nor U46143 (N_46143,N_33762,N_39832);
nand U46144 (N_46144,N_37296,N_31583);
and U46145 (N_46145,N_33146,N_32877);
or U46146 (N_46146,N_30175,N_38338);
or U46147 (N_46147,N_37440,N_33328);
and U46148 (N_46148,N_36229,N_37883);
or U46149 (N_46149,N_30044,N_39623);
and U46150 (N_46150,N_32272,N_32538);
nor U46151 (N_46151,N_33188,N_33180);
nor U46152 (N_46152,N_38390,N_30725);
or U46153 (N_46153,N_36797,N_34309);
and U46154 (N_46154,N_30661,N_34787);
nor U46155 (N_46155,N_31995,N_34556);
nand U46156 (N_46156,N_36446,N_31347);
xnor U46157 (N_46157,N_34881,N_37476);
and U46158 (N_46158,N_30211,N_31919);
or U46159 (N_46159,N_36019,N_38692);
or U46160 (N_46160,N_30666,N_38564);
and U46161 (N_46161,N_34193,N_38730);
nor U46162 (N_46162,N_31966,N_38552);
nand U46163 (N_46163,N_30835,N_37120);
nor U46164 (N_46164,N_37259,N_33942);
nor U46165 (N_46165,N_36791,N_37508);
xor U46166 (N_46166,N_39096,N_38473);
nand U46167 (N_46167,N_31410,N_31595);
and U46168 (N_46168,N_34548,N_30157);
or U46169 (N_46169,N_33235,N_37151);
nand U46170 (N_46170,N_34931,N_34111);
and U46171 (N_46171,N_30953,N_30298);
and U46172 (N_46172,N_34186,N_39195);
and U46173 (N_46173,N_39356,N_33259);
or U46174 (N_46174,N_30058,N_34265);
xor U46175 (N_46175,N_36612,N_36721);
xor U46176 (N_46176,N_32939,N_34753);
nor U46177 (N_46177,N_34129,N_33447);
nand U46178 (N_46178,N_38189,N_33714);
or U46179 (N_46179,N_35630,N_39169);
nand U46180 (N_46180,N_37651,N_30505);
or U46181 (N_46181,N_36820,N_39944);
or U46182 (N_46182,N_37797,N_30891);
and U46183 (N_46183,N_34272,N_38647);
nand U46184 (N_46184,N_35405,N_35900);
nor U46185 (N_46185,N_35191,N_31124);
nand U46186 (N_46186,N_31236,N_32026);
xnor U46187 (N_46187,N_34197,N_37469);
nand U46188 (N_46188,N_35428,N_30029);
xnor U46189 (N_46189,N_38927,N_30246);
and U46190 (N_46190,N_36138,N_39139);
and U46191 (N_46191,N_35752,N_35080);
or U46192 (N_46192,N_39069,N_39630);
nand U46193 (N_46193,N_32505,N_35606);
nor U46194 (N_46194,N_31772,N_37076);
nor U46195 (N_46195,N_35302,N_39787);
and U46196 (N_46196,N_36049,N_34875);
and U46197 (N_46197,N_31454,N_37557);
or U46198 (N_46198,N_33016,N_30829);
or U46199 (N_46199,N_32590,N_34090);
nor U46200 (N_46200,N_36910,N_30400);
nor U46201 (N_46201,N_39083,N_32772);
nand U46202 (N_46202,N_36285,N_33539);
nor U46203 (N_46203,N_39335,N_39138);
nand U46204 (N_46204,N_35314,N_35700);
or U46205 (N_46205,N_32994,N_38489);
or U46206 (N_46206,N_31798,N_31489);
and U46207 (N_46207,N_33257,N_35462);
nor U46208 (N_46208,N_39883,N_30984);
xnor U46209 (N_46209,N_37540,N_33996);
xor U46210 (N_46210,N_31428,N_36453);
or U46211 (N_46211,N_37491,N_32104);
nor U46212 (N_46212,N_36967,N_34259);
nand U46213 (N_46213,N_34532,N_39261);
and U46214 (N_46214,N_38767,N_31574);
nor U46215 (N_46215,N_32900,N_31119);
and U46216 (N_46216,N_33506,N_32018);
nor U46217 (N_46217,N_39569,N_33200);
and U46218 (N_46218,N_30793,N_35038);
or U46219 (N_46219,N_39965,N_36979);
or U46220 (N_46220,N_30532,N_33656);
and U46221 (N_46221,N_36732,N_37847);
nand U46222 (N_46222,N_31176,N_36723);
and U46223 (N_46223,N_39012,N_32182);
and U46224 (N_46224,N_33860,N_37327);
or U46225 (N_46225,N_31751,N_32233);
nor U46226 (N_46226,N_38659,N_36067);
or U46227 (N_46227,N_31449,N_34300);
and U46228 (N_46228,N_32104,N_39304);
and U46229 (N_46229,N_38853,N_37800);
nand U46230 (N_46230,N_36280,N_32531);
nand U46231 (N_46231,N_32795,N_37901);
and U46232 (N_46232,N_36623,N_34034);
xnor U46233 (N_46233,N_30491,N_33788);
or U46234 (N_46234,N_35107,N_33928);
nand U46235 (N_46235,N_37932,N_32637);
nand U46236 (N_46236,N_34058,N_39089);
nand U46237 (N_46237,N_36801,N_38447);
nor U46238 (N_46238,N_32395,N_34189);
nor U46239 (N_46239,N_35558,N_37615);
nor U46240 (N_46240,N_33475,N_30345);
nor U46241 (N_46241,N_36967,N_34989);
or U46242 (N_46242,N_30114,N_34348);
nor U46243 (N_46243,N_34455,N_30069);
and U46244 (N_46244,N_31895,N_35332);
and U46245 (N_46245,N_31188,N_35200);
and U46246 (N_46246,N_30445,N_30360);
or U46247 (N_46247,N_36131,N_34134);
and U46248 (N_46248,N_35971,N_35001);
or U46249 (N_46249,N_39960,N_39062);
nor U46250 (N_46250,N_39946,N_32190);
and U46251 (N_46251,N_38658,N_39010);
or U46252 (N_46252,N_37332,N_33730);
and U46253 (N_46253,N_35345,N_34968);
nand U46254 (N_46254,N_31338,N_39954);
nand U46255 (N_46255,N_31805,N_31729);
and U46256 (N_46256,N_33301,N_37518);
or U46257 (N_46257,N_31640,N_37129);
or U46258 (N_46258,N_34031,N_30622);
or U46259 (N_46259,N_34610,N_37452);
or U46260 (N_46260,N_33827,N_33553);
nor U46261 (N_46261,N_38681,N_39708);
nor U46262 (N_46262,N_38896,N_36820);
nor U46263 (N_46263,N_30993,N_39355);
nand U46264 (N_46264,N_39004,N_37132);
or U46265 (N_46265,N_36844,N_38878);
and U46266 (N_46266,N_32351,N_32539);
nand U46267 (N_46267,N_33222,N_34400);
and U46268 (N_46268,N_37499,N_38256);
nand U46269 (N_46269,N_34466,N_39798);
nand U46270 (N_46270,N_37921,N_38450);
nor U46271 (N_46271,N_38300,N_38098);
nand U46272 (N_46272,N_30349,N_30308);
nor U46273 (N_46273,N_38445,N_35272);
nand U46274 (N_46274,N_35174,N_35097);
and U46275 (N_46275,N_34790,N_37346);
xor U46276 (N_46276,N_33154,N_33595);
nand U46277 (N_46277,N_35318,N_31368);
or U46278 (N_46278,N_36323,N_30583);
nand U46279 (N_46279,N_33844,N_39377);
nor U46280 (N_46280,N_39253,N_30182);
or U46281 (N_46281,N_31098,N_34548);
and U46282 (N_46282,N_35708,N_32066);
nor U46283 (N_46283,N_32915,N_38356);
nor U46284 (N_46284,N_35531,N_33050);
nor U46285 (N_46285,N_34640,N_32595);
nor U46286 (N_46286,N_31462,N_36552);
nor U46287 (N_46287,N_36325,N_30264);
xnor U46288 (N_46288,N_32833,N_35267);
and U46289 (N_46289,N_38998,N_34884);
or U46290 (N_46290,N_33839,N_37676);
and U46291 (N_46291,N_37113,N_33398);
and U46292 (N_46292,N_34625,N_30973);
nor U46293 (N_46293,N_39197,N_31193);
or U46294 (N_46294,N_36195,N_35486);
nor U46295 (N_46295,N_32010,N_33784);
xor U46296 (N_46296,N_32410,N_30032);
nand U46297 (N_46297,N_30247,N_30512);
nor U46298 (N_46298,N_36417,N_30852);
or U46299 (N_46299,N_35113,N_39549);
and U46300 (N_46300,N_30053,N_32119);
nand U46301 (N_46301,N_37012,N_33374);
xor U46302 (N_46302,N_31383,N_36034);
nand U46303 (N_46303,N_31186,N_30206);
xor U46304 (N_46304,N_32430,N_30741);
nand U46305 (N_46305,N_37679,N_30004);
or U46306 (N_46306,N_35392,N_37300);
nor U46307 (N_46307,N_32827,N_33961);
xor U46308 (N_46308,N_33178,N_39344);
nor U46309 (N_46309,N_34111,N_36345);
or U46310 (N_46310,N_37454,N_35122);
xnor U46311 (N_46311,N_34198,N_38854);
nand U46312 (N_46312,N_33235,N_38242);
or U46313 (N_46313,N_30024,N_37360);
xnor U46314 (N_46314,N_33575,N_32101);
and U46315 (N_46315,N_35187,N_38231);
and U46316 (N_46316,N_38391,N_38559);
nand U46317 (N_46317,N_35695,N_31933);
xor U46318 (N_46318,N_30970,N_33104);
and U46319 (N_46319,N_39834,N_37599);
or U46320 (N_46320,N_36732,N_39593);
nor U46321 (N_46321,N_36632,N_33212);
nand U46322 (N_46322,N_36830,N_32966);
or U46323 (N_46323,N_36629,N_30130);
and U46324 (N_46324,N_37723,N_34391);
or U46325 (N_46325,N_34879,N_39530);
or U46326 (N_46326,N_35799,N_33294);
nand U46327 (N_46327,N_35311,N_31689);
or U46328 (N_46328,N_35870,N_36756);
nand U46329 (N_46329,N_33927,N_33319);
nand U46330 (N_46330,N_33647,N_30368);
or U46331 (N_46331,N_33974,N_30641);
and U46332 (N_46332,N_37269,N_32372);
or U46333 (N_46333,N_30541,N_38258);
nand U46334 (N_46334,N_36242,N_32656);
nor U46335 (N_46335,N_32593,N_38683);
nand U46336 (N_46336,N_31419,N_33764);
xnor U46337 (N_46337,N_31932,N_32126);
nor U46338 (N_46338,N_37291,N_32346);
or U46339 (N_46339,N_35484,N_30347);
nand U46340 (N_46340,N_39053,N_39751);
or U46341 (N_46341,N_33629,N_39234);
and U46342 (N_46342,N_37276,N_39939);
and U46343 (N_46343,N_32703,N_31568);
nand U46344 (N_46344,N_38920,N_36553);
nor U46345 (N_46345,N_33350,N_37452);
or U46346 (N_46346,N_39889,N_32370);
nor U46347 (N_46347,N_36129,N_31009);
nand U46348 (N_46348,N_36721,N_30877);
and U46349 (N_46349,N_34394,N_33382);
nor U46350 (N_46350,N_33553,N_38556);
xor U46351 (N_46351,N_39212,N_35439);
or U46352 (N_46352,N_35450,N_38979);
or U46353 (N_46353,N_30808,N_30050);
or U46354 (N_46354,N_32358,N_35140);
or U46355 (N_46355,N_34125,N_38803);
or U46356 (N_46356,N_31579,N_39375);
nor U46357 (N_46357,N_30634,N_35785);
or U46358 (N_46358,N_33516,N_33427);
nand U46359 (N_46359,N_30480,N_31993);
nand U46360 (N_46360,N_38448,N_33197);
or U46361 (N_46361,N_34527,N_35112);
nand U46362 (N_46362,N_32593,N_34332);
and U46363 (N_46363,N_36133,N_36471);
nand U46364 (N_46364,N_34837,N_31692);
or U46365 (N_46365,N_34545,N_33623);
and U46366 (N_46366,N_35934,N_31098);
nor U46367 (N_46367,N_31114,N_34473);
and U46368 (N_46368,N_36129,N_34142);
nor U46369 (N_46369,N_37455,N_34386);
and U46370 (N_46370,N_36462,N_32537);
nand U46371 (N_46371,N_36786,N_32434);
and U46372 (N_46372,N_34317,N_34077);
and U46373 (N_46373,N_39364,N_33527);
nor U46374 (N_46374,N_34904,N_35586);
and U46375 (N_46375,N_33066,N_39768);
and U46376 (N_46376,N_31885,N_33828);
nor U46377 (N_46377,N_30602,N_37074);
nor U46378 (N_46378,N_31695,N_35209);
nand U46379 (N_46379,N_30373,N_39751);
or U46380 (N_46380,N_33639,N_32920);
nand U46381 (N_46381,N_32289,N_31745);
xnor U46382 (N_46382,N_32775,N_30671);
nand U46383 (N_46383,N_30776,N_31848);
xnor U46384 (N_46384,N_31627,N_35340);
nor U46385 (N_46385,N_32687,N_38850);
or U46386 (N_46386,N_36384,N_38700);
nand U46387 (N_46387,N_36195,N_34961);
and U46388 (N_46388,N_36140,N_35388);
or U46389 (N_46389,N_30589,N_32154);
and U46390 (N_46390,N_31344,N_38478);
nor U46391 (N_46391,N_31512,N_38184);
nor U46392 (N_46392,N_36981,N_34698);
or U46393 (N_46393,N_30137,N_32963);
or U46394 (N_46394,N_31624,N_37955);
and U46395 (N_46395,N_34422,N_34089);
nor U46396 (N_46396,N_33999,N_35224);
and U46397 (N_46397,N_36364,N_35314);
and U46398 (N_46398,N_39760,N_36394);
nor U46399 (N_46399,N_38703,N_32483);
or U46400 (N_46400,N_39512,N_36573);
and U46401 (N_46401,N_39900,N_37151);
or U46402 (N_46402,N_36486,N_30251);
nor U46403 (N_46403,N_31088,N_34296);
nor U46404 (N_46404,N_31378,N_31003);
nand U46405 (N_46405,N_34169,N_34506);
or U46406 (N_46406,N_36859,N_35784);
nor U46407 (N_46407,N_39998,N_38663);
and U46408 (N_46408,N_35439,N_39013);
nor U46409 (N_46409,N_34644,N_32877);
or U46410 (N_46410,N_30968,N_32860);
nor U46411 (N_46411,N_34753,N_32065);
nor U46412 (N_46412,N_32783,N_35225);
or U46413 (N_46413,N_38862,N_34900);
and U46414 (N_46414,N_36549,N_32746);
nor U46415 (N_46415,N_36760,N_32374);
nand U46416 (N_46416,N_33274,N_38790);
nand U46417 (N_46417,N_34671,N_32351);
nor U46418 (N_46418,N_38508,N_36989);
or U46419 (N_46419,N_35447,N_31160);
or U46420 (N_46420,N_33331,N_31755);
and U46421 (N_46421,N_37236,N_35810);
nor U46422 (N_46422,N_37899,N_32938);
or U46423 (N_46423,N_37273,N_36400);
nand U46424 (N_46424,N_30869,N_34000);
xor U46425 (N_46425,N_32078,N_36118);
nor U46426 (N_46426,N_30439,N_39141);
nand U46427 (N_46427,N_33694,N_34439);
xor U46428 (N_46428,N_32803,N_32019);
and U46429 (N_46429,N_36342,N_39393);
or U46430 (N_46430,N_39772,N_38210);
and U46431 (N_46431,N_36652,N_36120);
and U46432 (N_46432,N_35786,N_31623);
xnor U46433 (N_46433,N_37144,N_38264);
and U46434 (N_46434,N_35418,N_35276);
nor U46435 (N_46435,N_31624,N_33049);
and U46436 (N_46436,N_32511,N_39691);
xnor U46437 (N_46437,N_32990,N_37191);
nand U46438 (N_46438,N_36898,N_33006);
and U46439 (N_46439,N_31900,N_31296);
nand U46440 (N_46440,N_30311,N_33991);
or U46441 (N_46441,N_32267,N_33691);
or U46442 (N_46442,N_32969,N_30614);
or U46443 (N_46443,N_34543,N_30971);
nand U46444 (N_46444,N_33570,N_34758);
and U46445 (N_46445,N_33217,N_39040);
nor U46446 (N_46446,N_39111,N_34277);
nand U46447 (N_46447,N_33333,N_32095);
and U46448 (N_46448,N_31044,N_39637);
xor U46449 (N_46449,N_32603,N_37130);
or U46450 (N_46450,N_38878,N_30958);
or U46451 (N_46451,N_35811,N_39510);
nor U46452 (N_46452,N_33411,N_39144);
or U46453 (N_46453,N_38578,N_36102);
and U46454 (N_46454,N_33628,N_33538);
xnor U46455 (N_46455,N_37440,N_31408);
nor U46456 (N_46456,N_36956,N_37457);
and U46457 (N_46457,N_31841,N_38598);
nor U46458 (N_46458,N_34841,N_32767);
xnor U46459 (N_46459,N_38552,N_30686);
or U46460 (N_46460,N_35337,N_36332);
nand U46461 (N_46461,N_39136,N_37619);
nor U46462 (N_46462,N_32563,N_33459);
nand U46463 (N_46463,N_30508,N_30325);
and U46464 (N_46464,N_39069,N_36341);
nand U46465 (N_46465,N_39528,N_33197);
nand U46466 (N_46466,N_30433,N_30584);
or U46467 (N_46467,N_36100,N_38791);
nor U46468 (N_46468,N_35700,N_36346);
nand U46469 (N_46469,N_31397,N_38439);
nor U46470 (N_46470,N_35717,N_30862);
and U46471 (N_46471,N_30607,N_30992);
nand U46472 (N_46472,N_30380,N_39419);
or U46473 (N_46473,N_32682,N_31147);
nand U46474 (N_46474,N_38245,N_32244);
nor U46475 (N_46475,N_36735,N_32138);
and U46476 (N_46476,N_33385,N_35802);
and U46477 (N_46477,N_37943,N_38235);
and U46478 (N_46478,N_36171,N_33725);
nor U46479 (N_46479,N_35191,N_30386);
nor U46480 (N_46480,N_35424,N_36813);
or U46481 (N_46481,N_37828,N_34740);
nor U46482 (N_46482,N_31509,N_32531);
and U46483 (N_46483,N_34631,N_34739);
nor U46484 (N_46484,N_32820,N_31032);
nor U46485 (N_46485,N_34567,N_37340);
or U46486 (N_46486,N_30812,N_38334);
nand U46487 (N_46487,N_38913,N_33536);
nand U46488 (N_46488,N_38257,N_33194);
xor U46489 (N_46489,N_30123,N_31862);
or U46490 (N_46490,N_35613,N_31568);
nor U46491 (N_46491,N_35434,N_35997);
nor U46492 (N_46492,N_35799,N_31775);
and U46493 (N_46493,N_38684,N_33880);
nand U46494 (N_46494,N_31302,N_38963);
nor U46495 (N_46495,N_33086,N_35580);
xnor U46496 (N_46496,N_35350,N_30777);
nand U46497 (N_46497,N_36256,N_37383);
and U46498 (N_46498,N_34356,N_38096);
or U46499 (N_46499,N_31766,N_39596);
nand U46500 (N_46500,N_35147,N_38082);
and U46501 (N_46501,N_39913,N_32081);
or U46502 (N_46502,N_39481,N_35317);
and U46503 (N_46503,N_31279,N_38462);
or U46504 (N_46504,N_33744,N_37044);
nor U46505 (N_46505,N_39635,N_31013);
or U46506 (N_46506,N_36954,N_38341);
and U46507 (N_46507,N_35194,N_30143);
nand U46508 (N_46508,N_36496,N_30167);
and U46509 (N_46509,N_32283,N_30645);
and U46510 (N_46510,N_32181,N_32239);
nor U46511 (N_46511,N_37143,N_36213);
and U46512 (N_46512,N_39583,N_31210);
nor U46513 (N_46513,N_39291,N_30586);
nor U46514 (N_46514,N_32198,N_33682);
or U46515 (N_46515,N_35666,N_33873);
or U46516 (N_46516,N_39346,N_32700);
nor U46517 (N_46517,N_37789,N_31493);
nor U46518 (N_46518,N_39681,N_38709);
nor U46519 (N_46519,N_38082,N_30588);
or U46520 (N_46520,N_31701,N_31354);
nor U46521 (N_46521,N_34193,N_38843);
and U46522 (N_46522,N_33370,N_30628);
and U46523 (N_46523,N_36382,N_37114);
nand U46524 (N_46524,N_31957,N_39087);
or U46525 (N_46525,N_35816,N_30750);
nor U46526 (N_46526,N_36913,N_38581);
nand U46527 (N_46527,N_33460,N_30578);
or U46528 (N_46528,N_32984,N_39938);
and U46529 (N_46529,N_32487,N_38791);
nor U46530 (N_46530,N_33371,N_34682);
nor U46531 (N_46531,N_32484,N_37749);
nor U46532 (N_46532,N_34384,N_30278);
nand U46533 (N_46533,N_36465,N_38572);
or U46534 (N_46534,N_38072,N_38786);
nor U46535 (N_46535,N_36271,N_39313);
or U46536 (N_46536,N_39108,N_39569);
nand U46537 (N_46537,N_32628,N_39203);
nor U46538 (N_46538,N_38465,N_38828);
nand U46539 (N_46539,N_34557,N_32355);
nor U46540 (N_46540,N_37991,N_36753);
nand U46541 (N_46541,N_35786,N_38319);
and U46542 (N_46542,N_38043,N_37270);
nand U46543 (N_46543,N_31591,N_37775);
xor U46544 (N_46544,N_33858,N_31222);
and U46545 (N_46545,N_38528,N_33985);
nand U46546 (N_46546,N_39051,N_36484);
nand U46547 (N_46547,N_35970,N_39642);
and U46548 (N_46548,N_37148,N_38745);
or U46549 (N_46549,N_33064,N_34884);
and U46550 (N_46550,N_39579,N_30100);
or U46551 (N_46551,N_33844,N_35707);
or U46552 (N_46552,N_38025,N_33106);
nand U46553 (N_46553,N_36568,N_38422);
nor U46554 (N_46554,N_30731,N_32070);
and U46555 (N_46555,N_37242,N_37041);
nand U46556 (N_46556,N_32220,N_31777);
and U46557 (N_46557,N_30772,N_38913);
and U46558 (N_46558,N_38557,N_30533);
nand U46559 (N_46559,N_38343,N_31335);
xor U46560 (N_46560,N_31514,N_31030);
or U46561 (N_46561,N_38005,N_36239);
xor U46562 (N_46562,N_30739,N_31860);
and U46563 (N_46563,N_38102,N_39666);
and U46564 (N_46564,N_36163,N_34714);
nor U46565 (N_46565,N_32720,N_38021);
nor U46566 (N_46566,N_38580,N_38930);
nand U46567 (N_46567,N_37999,N_39292);
and U46568 (N_46568,N_35044,N_39064);
xnor U46569 (N_46569,N_31584,N_37494);
xor U46570 (N_46570,N_37689,N_35006);
nand U46571 (N_46571,N_34048,N_32084);
and U46572 (N_46572,N_36061,N_37404);
xnor U46573 (N_46573,N_35094,N_32745);
or U46574 (N_46574,N_32739,N_31464);
and U46575 (N_46575,N_32798,N_35438);
and U46576 (N_46576,N_39966,N_38005);
nand U46577 (N_46577,N_39599,N_34931);
nor U46578 (N_46578,N_36124,N_34581);
nor U46579 (N_46579,N_30350,N_39171);
nor U46580 (N_46580,N_34629,N_36860);
xnor U46581 (N_46581,N_38571,N_31386);
nor U46582 (N_46582,N_35043,N_32590);
xnor U46583 (N_46583,N_33412,N_34938);
nor U46584 (N_46584,N_32912,N_37587);
nor U46585 (N_46585,N_35474,N_33625);
nand U46586 (N_46586,N_39368,N_34046);
nor U46587 (N_46587,N_31240,N_38153);
and U46588 (N_46588,N_37917,N_37487);
nor U46589 (N_46589,N_30981,N_34661);
and U46590 (N_46590,N_32770,N_39713);
nand U46591 (N_46591,N_36988,N_38393);
and U46592 (N_46592,N_35186,N_33480);
xor U46593 (N_46593,N_31059,N_30104);
nor U46594 (N_46594,N_38966,N_34618);
nor U46595 (N_46595,N_34232,N_35737);
xor U46596 (N_46596,N_32550,N_37856);
nor U46597 (N_46597,N_38351,N_38540);
xnor U46598 (N_46598,N_30079,N_34151);
and U46599 (N_46599,N_34592,N_31614);
xnor U46600 (N_46600,N_39717,N_36027);
or U46601 (N_46601,N_38606,N_35558);
nor U46602 (N_46602,N_31083,N_36883);
or U46603 (N_46603,N_31256,N_31587);
and U46604 (N_46604,N_36113,N_39064);
and U46605 (N_46605,N_34302,N_30479);
xnor U46606 (N_46606,N_33219,N_34933);
or U46607 (N_46607,N_37196,N_31800);
nand U46608 (N_46608,N_31297,N_35878);
and U46609 (N_46609,N_36102,N_31232);
xnor U46610 (N_46610,N_34120,N_39039);
xor U46611 (N_46611,N_33872,N_35638);
nand U46612 (N_46612,N_37080,N_35096);
nand U46613 (N_46613,N_31446,N_37112);
and U46614 (N_46614,N_39432,N_32892);
xor U46615 (N_46615,N_36881,N_38534);
nand U46616 (N_46616,N_30855,N_31135);
and U46617 (N_46617,N_31094,N_31540);
nor U46618 (N_46618,N_36386,N_31958);
or U46619 (N_46619,N_37959,N_38287);
and U46620 (N_46620,N_33344,N_37385);
or U46621 (N_46621,N_31070,N_33657);
or U46622 (N_46622,N_33538,N_38591);
nor U46623 (N_46623,N_30391,N_31724);
nand U46624 (N_46624,N_35158,N_36540);
and U46625 (N_46625,N_31431,N_39431);
and U46626 (N_46626,N_35343,N_35773);
and U46627 (N_46627,N_39032,N_39849);
nand U46628 (N_46628,N_33439,N_32465);
nor U46629 (N_46629,N_38264,N_32984);
nor U46630 (N_46630,N_39556,N_37281);
or U46631 (N_46631,N_37699,N_30148);
or U46632 (N_46632,N_37462,N_31654);
xnor U46633 (N_46633,N_36773,N_39385);
or U46634 (N_46634,N_38370,N_37231);
and U46635 (N_46635,N_39140,N_37908);
or U46636 (N_46636,N_39270,N_31724);
nor U46637 (N_46637,N_39835,N_39535);
or U46638 (N_46638,N_35938,N_39679);
and U46639 (N_46639,N_33399,N_30343);
or U46640 (N_46640,N_34416,N_32841);
or U46641 (N_46641,N_38785,N_38797);
and U46642 (N_46642,N_39587,N_34760);
nand U46643 (N_46643,N_33536,N_35267);
and U46644 (N_46644,N_33217,N_32593);
and U46645 (N_46645,N_34178,N_30491);
and U46646 (N_46646,N_30278,N_30841);
nor U46647 (N_46647,N_35556,N_36859);
xnor U46648 (N_46648,N_35163,N_35993);
nor U46649 (N_46649,N_31171,N_36461);
or U46650 (N_46650,N_34014,N_30422);
or U46651 (N_46651,N_38696,N_36430);
xnor U46652 (N_46652,N_35756,N_36475);
nor U46653 (N_46653,N_33744,N_32570);
or U46654 (N_46654,N_36411,N_39748);
nand U46655 (N_46655,N_33464,N_35035);
nand U46656 (N_46656,N_37431,N_39535);
nor U46657 (N_46657,N_31420,N_37020);
or U46658 (N_46658,N_38369,N_34348);
nor U46659 (N_46659,N_31654,N_35640);
nand U46660 (N_46660,N_33990,N_39157);
or U46661 (N_46661,N_39346,N_36806);
or U46662 (N_46662,N_34402,N_33688);
and U46663 (N_46663,N_38009,N_35223);
nand U46664 (N_46664,N_32854,N_30908);
nor U46665 (N_46665,N_31887,N_38767);
nand U46666 (N_46666,N_38320,N_39924);
nor U46667 (N_46667,N_31654,N_31876);
xnor U46668 (N_46668,N_36981,N_31665);
nand U46669 (N_46669,N_37774,N_34576);
xnor U46670 (N_46670,N_39087,N_34169);
nor U46671 (N_46671,N_33395,N_37429);
nor U46672 (N_46672,N_35261,N_39624);
or U46673 (N_46673,N_38863,N_36645);
nor U46674 (N_46674,N_37813,N_39117);
xnor U46675 (N_46675,N_34111,N_34417);
and U46676 (N_46676,N_33624,N_36378);
and U46677 (N_46677,N_34082,N_39938);
and U46678 (N_46678,N_39866,N_38679);
nor U46679 (N_46679,N_31603,N_32503);
and U46680 (N_46680,N_33676,N_30283);
or U46681 (N_46681,N_33674,N_37378);
and U46682 (N_46682,N_39733,N_31799);
nor U46683 (N_46683,N_31603,N_31087);
and U46684 (N_46684,N_37315,N_38846);
and U46685 (N_46685,N_32132,N_39552);
nor U46686 (N_46686,N_33092,N_36692);
nand U46687 (N_46687,N_37561,N_30082);
nand U46688 (N_46688,N_31470,N_39615);
and U46689 (N_46689,N_38801,N_33666);
or U46690 (N_46690,N_32821,N_30789);
nor U46691 (N_46691,N_34713,N_31035);
and U46692 (N_46692,N_33238,N_32508);
and U46693 (N_46693,N_35793,N_37803);
nand U46694 (N_46694,N_36132,N_31283);
nor U46695 (N_46695,N_32133,N_39091);
nand U46696 (N_46696,N_32121,N_39355);
nor U46697 (N_46697,N_35561,N_32859);
nor U46698 (N_46698,N_30876,N_32655);
or U46699 (N_46699,N_36794,N_32643);
or U46700 (N_46700,N_34972,N_37596);
or U46701 (N_46701,N_39381,N_30105);
nor U46702 (N_46702,N_36273,N_36453);
and U46703 (N_46703,N_32528,N_39412);
or U46704 (N_46704,N_30899,N_34237);
or U46705 (N_46705,N_38783,N_36878);
or U46706 (N_46706,N_39246,N_38049);
nor U46707 (N_46707,N_36871,N_32940);
nand U46708 (N_46708,N_32383,N_32093);
nor U46709 (N_46709,N_33965,N_38447);
and U46710 (N_46710,N_33931,N_39581);
or U46711 (N_46711,N_34575,N_32087);
nand U46712 (N_46712,N_30340,N_35531);
or U46713 (N_46713,N_38669,N_31930);
or U46714 (N_46714,N_38928,N_31949);
or U46715 (N_46715,N_37192,N_33279);
and U46716 (N_46716,N_35061,N_32432);
nor U46717 (N_46717,N_34114,N_31296);
nor U46718 (N_46718,N_39277,N_33474);
nor U46719 (N_46719,N_30410,N_36510);
and U46720 (N_46720,N_35103,N_32495);
nor U46721 (N_46721,N_39169,N_36946);
nor U46722 (N_46722,N_33900,N_32818);
or U46723 (N_46723,N_34690,N_36886);
and U46724 (N_46724,N_31520,N_35377);
or U46725 (N_46725,N_30458,N_37329);
nor U46726 (N_46726,N_34597,N_39196);
nor U46727 (N_46727,N_39275,N_30441);
and U46728 (N_46728,N_30176,N_30041);
xor U46729 (N_46729,N_35425,N_32932);
nor U46730 (N_46730,N_39113,N_37531);
nand U46731 (N_46731,N_32407,N_37578);
or U46732 (N_46732,N_33987,N_31251);
or U46733 (N_46733,N_38588,N_34928);
nor U46734 (N_46734,N_35792,N_38957);
nor U46735 (N_46735,N_33882,N_30629);
xnor U46736 (N_46736,N_37815,N_33695);
and U46737 (N_46737,N_32335,N_30929);
and U46738 (N_46738,N_37886,N_39043);
nor U46739 (N_46739,N_33315,N_38732);
or U46740 (N_46740,N_34045,N_31765);
nand U46741 (N_46741,N_31781,N_39213);
and U46742 (N_46742,N_39009,N_34237);
nor U46743 (N_46743,N_30947,N_36368);
nand U46744 (N_46744,N_34502,N_38209);
nor U46745 (N_46745,N_36791,N_31783);
nor U46746 (N_46746,N_35250,N_31819);
or U46747 (N_46747,N_39768,N_34877);
nand U46748 (N_46748,N_39842,N_30900);
xnor U46749 (N_46749,N_30380,N_37829);
xnor U46750 (N_46750,N_38517,N_35966);
and U46751 (N_46751,N_37774,N_35987);
or U46752 (N_46752,N_38856,N_38459);
nand U46753 (N_46753,N_34800,N_38942);
nand U46754 (N_46754,N_36452,N_32664);
or U46755 (N_46755,N_34332,N_38457);
or U46756 (N_46756,N_34666,N_31374);
or U46757 (N_46757,N_30748,N_30694);
xnor U46758 (N_46758,N_31006,N_31023);
nand U46759 (N_46759,N_31284,N_39534);
and U46760 (N_46760,N_35878,N_32681);
nor U46761 (N_46761,N_30958,N_35221);
nand U46762 (N_46762,N_39238,N_30928);
nor U46763 (N_46763,N_36128,N_35158);
or U46764 (N_46764,N_34845,N_39541);
nand U46765 (N_46765,N_30440,N_38226);
nor U46766 (N_46766,N_34110,N_37738);
and U46767 (N_46767,N_35564,N_35470);
xor U46768 (N_46768,N_32044,N_32625);
xnor U46769 (N_46769,N_30055,N_35019);
and U46770 (N_46770,N_35111,N_32910);
nand U46771 (N_46771,N_38176,N_33962);
and U46772 (N_46772,N_37935,N_32073);
or U46773 (N_46773,N_35864,N_35398);
nand U46774 (N_46774,N_36114,N_39465);
and U46775 (N_46775,N_35128,N_30492);
nor U46776 (N_46776,N_36539,N_31840);
nor U46777 (N_46777,N_34171,N_36195);
or U46778 (N_46778,N_39798,N_34737);
nand U46779 (N_46779,N_34360,N_30722);
nor U46780 (N_46780,N_34737,N_33386);
nor U46781 (N_46781,N_31416,N_37813);
and U46782 (N_46782,N_39636,N_33465);
nand U46783 (N_46783,N_37736,N_30552);
and U46784 (N_46784,N_38454,N_31668);
or U46785 (N_46785,N_36899,N_36942);
nor U46786 (N_46786,N_35577,N_32709);
nand U46787 (N_46787,N_36361,N_31093);
nand U46788 (N_46788,N_34688,N_39210);
xnor U46789 (N_46789,N_37316,N_30514);
or U46790 (N_46790,N_32526,N_31826);
nor U46791 (N_46791,N_32433,N_31810);
nand U46792 (N_46792,N_38677,N_32176);
xnor U46793 (N_46793,N_33073,N_33222);
or U46794 (N_46794,N_36160,N_33716);
and U46795 (N_46795,N_38744,N_34213);
nor U46796 (N_46796,N_35190,N_35408);
nand U46797 (N_46797,N_33197,N_30838);
and U46798 (N_46798,N_32822,N_33705);
xor U46799 (N_46799,N_30196,N_37591);
nor U46800 (N_46800,N_37516,N_34731);
nand U46801 (N_46801,N_34779,N_36880);
nand U46802 (N_46802,N_30583,N_36696);
nor U46803 (N_46803,N_38089,N_30207);
nand U46804 (N_46804,N_39043,N_34816);
and U46805 (N_46805,N_34863,N_32233);
nor U46806 (N_46806,N_38739,N_37893);
nor U46807 (N_46807,N_38965,N_30025);
or U46808 (N_46808,N_34327,N_38533);
nand U46809 (N_46809,N_30027,N_36227);
or U46810 (N_46810,N_39123,N_38191);
and U46811 (N_46811,N_31162,N_32131);
nand U46812 (N_46812,N_30662,N_35204);
nand U46813 (N_46813,N_36851,N_39159);
nor U46814 (N_46814,N_30809,N_38009);
and U46815 (N_46815,N_33482,N_33138);
and U46816 (N_46816,N_38791,N_30191);
nand U46817 (N_46817,N_32592,N_34746);
nand U46818 (N_46818,N_39267,N_38769);
or U46819 (N_46819,N_37034,N_31208);
nand U46820 (N_46820,N_30681,N_38780);
or U46821 (N_46821,N_33402,N_35928);
and U46822 (N_46822,N_34482,N_31007);
and U46823 (N_46823,N_32930,N_33619);
and U46824 (N_46824,N_35975,N_33324);
nor U46825 (N_46825,N_31961,N_35455);
nor U46826 (N_46826,N_37821,N_37188);
or U46827 (N_46827,N_32741,N_32395);
or U46828 (N_46828,N_32826,N_33145);
nor U46829 (N_46829,N_39532,N_36505);
nor U46830 (N_46830,N_30799,N_35623);
nand U46831 (N_46831,N_33834,N_31224);
nand U46832 (N_46832,N_35920,N_34294);
or U46833 (N_46833,N_32112,N_30320);
nand U46834 (N_46834,N_32722,N_35775);
nand U46835 (N_46835,N_32006,N_37525);
nor U46836 (N_46836,N_39373,N_32333);
nor U46837 (N_46837,N_35739,N_35760);
nor U46838 (N_46838,N_37631,N_35268);
and U46839 (N_46839,N_35057,N_35563);
xnor U46840 (N_46840,N_37274,N_37171);
nor U46841 (N_46841,N_32846,N_32377);
and U46842 (N_46842,N_34626,N_31594);
and U46843 (N_46843,N_38256,N_39610);
and U46844 (N_46844,N_38982,N_34204);
nor U46845 (N_46845,N_38756,N_34874);
nor U46846 (N_46846,N_35141,N_30921);
nand U46847 (N_46847,N_37480,N_30070);
and U46848 (N_46848,N_33116,N_30956);
nand U46849 (N_46849,N_32758,N_38814);
and U46850 (N_46850,N_32388,N_34546);
and U46851 (N_46851,N_30915,N_38028);
nor U46852 (N_46852,N_38122,N_35103);
nor U46853 (N_46853,N_34083,N_33259);
and U46854 (N_46854,N_30469,N_38352);
or U46855 (N_46855,N_30330,N_37009);
xor U46856 (N_46856,N_36548,N_35051);
and U46857 (N_46857,N_36743,N_38097);
nand U46858 (N_46858,N_32117,N_35908);
or U46859 (N_46859,N_30467,N_35697);
nand U46860 (N_46860,N_38729,N_33195);
or U46861 (N_46861,N_38653,N_33629);
nand U46862 (N_46862,N_35298,N_37425);
nand U46863 (N_46863,N_34801,N_37480);
or U46864 (N_46864,N_39139,N_30416);
nand U46865 (N_46865,N_36095,N_30161);
or U46866 (N_46866,N_39044,N_38810);
nor U46867 (N_46867,N_33038,N_37220);
xor U46868 (N_46868,N_30273,N_37084);
nor U46869 (N_46869,N_30743,N_39564);
and U46870 (N_46870,N_37772,N_36155);
nand U46871 (N_46871,N_31438,N_34808);
nand U46872 (N_46872,N_33160,N_33260);
nand U46873 (N_46873,N_30824,N_34598);
xor U46874 (N_46874,N_39686,N_39378);
and U46875 (N_46875,N_34966,N_36381);
or U46876 (N_46876,N_38166,N_36188);
xnor U46877 (N_46877,N_35718,N_36123);
or U46878 (N_46878,N_37955,N_35131);
nand U46879 (N_46879,N_36741,N_35226);
nor U46880 (N_46880,N_37636,N_32151);
or U46881 (N_46881,N_33360,N_39460);
and U46882 (N_46882,N_38501,N_34870);
nor U46883 (N_46883,N_36814,N_32921);
and U46884 (N_46884,N_31581,N_34001);
nor U46885 (N_46885,N_30704,N_37805);
nand U46886 (N_46886,N_36199,N_37469);
nand U46887 (N_46887,N_37933,N_37352);
nor U46888 (N_46888,N_39850,N_33087);
or U46889 (N_46889,N_38421,N_38679);
nand U46890 (N_46890,N_32054,N_38726);
nand U46891 (N_46891,N_34357,N_35857);
nor U46892 (N_46892,N_30521,N_31382);
nand U46893 (N_46893,N_34812,N_36739);
xor U46894 (N_46894,N_32680,N_33445);
nor U46895 (N_46895,N_33670,N_38686);
nand U46896 (N_46896,N_39974,N_38850);
nor U46897 (N_46897,N_30444,N_31140);
and U46898 (N_46898,N_34073,N_30818);
xor U46899 (N_46899,N_31808,N_35110);
and U46900 (N_46900,N_38996,N_30503);
nor U46901 (N_46901,N_34105,N_30046);
nand U46902 (N_46902,N_39802,N_36407);
nand U46903 (N_46903,N_38551,N_39469);
nand U46904 (N_46904,N_36236,N_34264);
and U46905 (N_46905,N_36859,N_39149);
or U46906 (N_46906,N_33389,N_39893);
or U46907 (N_46907,N_39928,N_36310);
and U46908 (N_46908,N_37181,N_31874);
nor U46909 (N_46909,N_36230,N_33445);
nor U46910 (N_46910,N_33678,N_32555);
nor U46911 (N_46911,N_36801,N_31447);
nor U46912 (N_46912,N_38902,N_37134);
nor U46913 (N_46913,N_38861,N_32312);
nor U46914 (N_46914,N_33257,N_39549);
nand U46915 (N_46915,N_37592,N_32470);
and U46916 (N_46916,N_36204,N_32812);
and U46917 (N_46917,N_34513,N_32494);
nor U46918 (N_46918,N_31876,N_31970);
nand U46919 (N_46919,N_33789,N_34340);
nor U46920 (N_46920,N_39769,N_36200);
or U46921 (N_46921,N_35883,N_32111);
nand U46922 (N_46922,N_34126,N_38829);
nor U46923 (N_46923,N_39418,N_37115);
nor U46924 (N_46924,N_36351,N_31967);
or U46925 (N_46925,N_37362,N_36038);
or U46926 (N_46926,N_31613,N_35796);
nand U46927 (N_46927,N_37033,N_34572);
nor U46928 (N_46928,N_37924,N_30479);
or U46929 (N_46929,N_33640,N_37587);
or U46930 (N_46930,N_34549,N_35557);
and U46931 (N_46931,N_32252,N_34295);
and U46932 (N_46932,N_33840,N_37228);
nor U46933 (N_46933,N_30548,N_32729);
nor U46934 (N_46934,N_38659,N_37680);
nor U46935 (N_46935,N_34411,N_32608);
nor U46936 (N_46936,N_39614,N_32066);
or U46937 (N_46937,N_30285,N_37302);
and U46938 (N_46938,N_33448,N_31514);
nand U46939 (N_46939,N_35699,N_38789);
or U46940 (N_46940,N_38029,N_30007);
nand U46941 (N_46941,N_32357,N_31488);
and U46942 (N_46942,N_32147,N_35350);
nor U46943 (N_46943,N_32468,N_35158);
and U46944 (N_46944,N_30450,N_36893);
or U46945 (N_46945,N_36677,N_38255);
or U46946 (N_46946,N_35396,N_36559);
or U46947 (N_46947,N_35860,N_39993);
or U46948 (N_46948,N_35007,N_30141);
nand U46949 (N_46949,N_30311,N_35830);
and U46950 (N_46950,N_38933,N_39478);
nor U46951 (N_46951,N_39352,N_32440);
xor U46952 (N_46952,N_37361,N_30320);
and U46953 (N_46953,N_34683,N_30047);
nor U46954 (N_46954,N_38234,N_33494);
or U46955 (N_46955,N_30486,N_37638);
nand U46956 (N_46956,N_33971,N_38086);
and U46957 (N_46957,N_32153,N_37311);
nor U46958 (N_46958,N_32208,N_31548);
and U46959 (N_46959,N_37559,N_35337);
and U46960 (N_46960,N_36768,N_35865);
nor U46961 (N_46961,N_38340,N_31540);
nor U46962 (N_46962,N_36338,N_33288);
nor U46963 (N_46963,N_30150,N_38909);
or U46964 (N_46964,N_34971,N_35552);
and U46965 (N_46965,N_36332,N_39548);
nor U46966 (N_46966,N_38628,N_35953);
nor U46967 (N_46967,N_38230,N_33981);
and U46968 (N_46968,N_37827,N_38987);
and U46969 (N_46969,N_33651,N_39644);
xor U46970 (N_46970,N_30231,N_33266);
nand U46971 (N_46971,N_32373,N_32195);
or U46972 (N_46972,N_37620,N_30327);
and U46973 (N_46973,N_38800,N_39092);
nor U46974 (N_46974,N_31480,N_39437);
or U46975 (N_46975,N_36540,N_32396);
nand U46976 (N_46976,N_33794,N_33016);
nor U46977 (N_46977,N_30157,N_30217);
and U46978 (N_46978,N_37111,N_39334);
nand U46979 (N_46979,N_35147,N_37832);
and U46980 (N_46980,N_37644,N_33367);
nand U46981 (N_46981,N_33847,N_31764);
nor U46982 (N_46982,N_34237,N_38012);
or U46983 (N_46983,N_37023,N_36637);
or U46984 (N_46984,N_35411,N_30112);
nand U46985 (N_46985,N_39578,N_35315);
nand U46986 (N_46986,N_32715,N_31736);
nor U46987 (N_46987,N_33518,N_31772);
or U46988 (N_46988,N_37278,N_35826);
and U46989 (N_46989,N_34157,N_31978);
and U46990 (N_46990,N_36582,N_38503);
nand U46991 (N_46991,N_32089,N_30116);
or U46992 (N_46992,N_34555,N_35240);
and U46993 (N_46993,N_36573,N_30193);
or U46994 (N_46994,N_34705,N_37847);
or U46995 (N_46995,N_33908,N_36701);
and U46996 (N_46996,N_32410,N_31611);
nor U46997 (N_46997,N_30168,N_35162);
and U46998 (N_46998,N_34684,N_32899);
or U46999 (N_46999,N_32907,N_32936);
or U47000 (N_47000,N_38590,N_35893);
or U47001 (N_47001,N_37913,N_30856);
nor U47002 (N_47002,N_34428,N_34138);
nor U47003 (N_47003,N_38183,N_39371);
nand U47004 (N_47004,N_32625,N_39378);
and U47005 (N_47005,N_33585,N_31229);
nor U47006 (N_47006,N_38556,N_31783);
nor U47007 (N_47007,N_32603,N_32362);
or U47008 (N_47008,N_31660,N_39050);
nor U47009 (N_47009,N_30281,N_37154);
nand U47010 (N_47010,N_37116,N_33364);
nor U47011 (N_47011,N_39867,N_35875);
and U47012 (N_47012,N_37472,N_32091);
nor U47013 (N_47013,N_34057,N_31821);
nand U47014 (N_47014,N_35442,N_36490);
nor U47015 (N_47015,N_31126,N_30797);
nand U47016 (N_47016,N_39351,N_30054);
or U47017 (N_47017,N_31971,N_34640);
nand U47018 (N_47018,N_35460,N_33197);
nand U47019 (N_47019,N_30463,N_37848);
and U47020 (N_47020,N_33466,N_35389);
or U47021 (N_47021,N_32739,N_39517);
xnor U47022 (N_47022,N_36782,N_33030);
nand U47023 (N_47023,N_33923,N_35052);
nand U47024 (N_47024,N_37381,N_34425);
or U47025 (N_47025,N_35597,N_37742);
nand U47026 (N_47026,N_32805,N_30207);
and U47027 (N_47027,N_31189,N_34197);
xnor U47028 (N_47028,N_33228,N_33325);
or U47029 (N_47029,N_33302,N_32814);
xor U47030 (N_47030,N_33540,N_37439);
nor U47031 (N_47031,N_36831,N_35331);
or U47032 (N_47032,N_31471,N_32592);
and U47033 (N_47033,N_38390,N_32669);
or U47034 (N_47034,N_39187,N_31665);
or U47035 (N_47035,N_33934,N_35331);
nor U47036 (N_47036,N_38843,N_37886);
nand U47037 (N_47037,N_38722,N_33199);
nor U47038 (N_47038,N_38449,N_33831);
or U47039 (N_47039,N_37250,N_36380);
or U47040 (N_47040,N_34606,N_32145);
nand U47041 (N_47041,N_30596,N_37544);
and U47042 (N_47042,N_38772,N_34933);
nand U47043 (N_47043,N_39356,N_32052);
and U47044 (N_47044,N_39159,N_34976);
nor U47045 (N_47045,N_33711,N_30283);
or U47046 (N_47046,N_35370,N_36805);
or U47047 (N_47047,N_35087,N_31174);
and U47048 (N_47048,N_35328,N_30797);
xnor U47049 (N_47049,N_36265,N_32505);
and U47050 (N_47050,N_31164,N_32844);
and U47051 (N_47051,N_36107,N_33917);
and U47052 (N_47052,N_36502,N_35567);
or U47053 (N_47053,N_38571,N_32295);
nor U47054 (N_47054,N_36384,N_36329);
nand U47055 (N_47055,N_34368,N_38259);
nand U47056 (N_47056,N_37893,N_33778);
and U47057 (N_47057,N_32097,N_30938);
and U47058 (N_47058,N_32928,N_35855);
and U47059 (N_47059,N_35265,N_30054);
nor U47060 (N_47060,N_31078,N_33601);
or U47061 (N_47061,N_32637,N_30195);
or U47062 (N_47062,N_37107,N_34130);
nand U47063 (N_47063,N_37224,N_35109);
xor U47064 (N_47064,N_32012,N_30173);
nand U47065 (N_47065,N_32858,N_32281);
nand U47066 (N_47066,N_34464,N_31532);
nand U47067 (N_47067,N_35671,N_31438);
nand U47068 (N_47068,N_32635,N_38277);
or U47069 (N_47069,N_33562,N_38592);
nor U47070 (N_47070,N_36749,N_31351);
nor U47071 (N_47071,N_31304,N_35402);
nor U47072 (N_47072,N_36620,N_31899);
nand U47073 (N_47073,N_35736,N_37390);
nor U47074 (N_47074,N_31397,N_31333);
xor U47075 (N_47075,N_30748,N_36231);
nor U47076 (N_47076,N_33882,N_33019);
xnor U47077 (N_47077,N_34157,N_38029);
nor U47078 (N_47078,N_31897,N_35224);
or U47079 (N_47079,N_38588,N_30122);
or U47080 (N_47080,N_30426,N_39475);
and U47081 (N_47081,N_33552,N_38441);
nor U47082 (N_47082,N_34466,N_38393);
or U47083 (N_47083,N_33000,N_38209);
and U47084 (N_47084,N_33688,N_30363);
or U47085 (N_47085,N_39581,N_37107);
and U47086 (N_47086,N_31490,N_31425);
or U47087 (N_47087,N_31483,N_31154);
nor U47088 (N_47088,N_34960,N_31830);
nor U47089 (N_47089,N_30913,N_37102);
nor U47090 (N_47090,N_37519,N_32542);
or U47091 (N_47091,N_33843,N_30440);
and U47092 (N_47092,N_36008,N_37433);
nand U47093 (N_47093,N_33038,N_38384);
and U47094 (N_47094,N_30086,N_35170);
nand U47095 (N_47095,N_31498,N_38268);
and U47096 (N_47096,N_32828,N_37600);
and U47097 (N_47097,N_37338,N_36345);
or U47098 (N_47098,N_33194,N_38597);
or U47099 (N_47099,N_30975,N_32382);
or U47100 (N_47100,N_34713,N_37399);
nand U47101 (N_47101,N_38497,N_31761);
nand U47102 (N_47102,N_39157,N_35615);
nand U47103 (N_47103,N_30212,N_33773);
nand U47104 (N_47104,N_30831,N_31389);
nor U47105 (N_47105,N_32985,N_33532);
and U47106 (N_47106,N_35444,N_30696);
nand U47107 (N_47107,N_33606,N_32484);
nand U47108 (N_47108,N_30668,N_34417);
nor U47109 (N_47109,N_30845,N_37788);
nor U47110 (N_47110,N_30185,N_33098);
and U47111 (N_47111,N_35919,N_35846);
nor U47112 (N_47112,N_34549,N_39193);
xnor U47113 (N_47113,N_31243,N_34977);
and U47114 (N_47114,N_35522,N_39707);
and U47115 (N_47115,N_37132,N_33543);
or U47116 (N_47116,N_38349,N_38900);
nand U47117 (N_47117,N_30975,N_36992);
or U47118 (N_47118,N_32728,N_33070);
or U47119 (N_47119,N_34812,N_36879);
nor U47120 (N_47120,N_35267,N_31093);
and U47121 (N_47121,N_39115,N_39216);
xor U47122 (N_47122,N_30365,N_32271);
and U47123 (N_47123,N_33609,N_34668);
xnor U47124 (N_47124,N_31909,N_39155);
nor U47125 (N_47125,N_32020,N_38081);
nand U47126 (N_47126,N_35680,N_35810);
nand U47127 (N_47127,N_31730,N_37771);
and U47128 (N_47128,N_35816,N_32740);
or U47129 (N_47129,N_32796,N_35593);
or U47130 (N_47130,N_30024,N_39285);
and U47131 (N_47131,N_38277,N_36484);
or U47132 (N_47132,N_38893,N_34340);
and U47133 (N_47133,N_35567,N_34491);
nand U47134 (N_47134,N_35618,N_37337);
nand U47135 (N_47135,N_37754,N_37577);
nor U47136 (N_47136,N_36782,N_39415);
or U47137 (N_47137,N_39382,N_37820);
or U47138 (N_47138,N_34603,N_30736);
xor U47139 (N_47139,N_30309,N_38227);
or U47140 (N_47140,N_39376,N_39475);
and U47141 (N_47141,N_36807,N_35695);
nor U47142 (N_47142,N_36958,N_32641);
and U47143 (N_47143,N_32994,N_32291);
xor U47144 (N_47144,N_39185,N_30787);
and U47145 (N_47145,N_36402,N_35471);
nor U47146 (N_47146,N_31612,N_38747);
xnor U47147 (N_47147,N_34646,N_35931);
nor U47148 (N_47148,N_35685,N_39073);
and U47149 (N_47149,N_37799,N_36257);
nand U47150 (N_47150,N_38067,N_31740);
and U47151 (N_47151,N_35030,N_36329);
or U47152 (N_47152,N_32568,N_33312);
or U47153 (N_47153,N_39376,N_31908);
and U47154 (N_47154,N_37766,N_36812);
or U47155 (N_47155,N_31457,N_35241);
nor U47156 (N_47156,N_35895,N_38664);
and U47157 (N_47157,N_36042,N_37507);
or U47158 (N_47158,N_32615,N_36140);
nand U47159 (N_47159,N_38390,N_32618);
nand U47160 (N_47160,N_32692,N_36394);
or U47161 (N_47161,N_31951,N_39631);
and U47162 (N_47162,N_33876,N_39033);
nor U47163 (N_47163,N_33999,N_32378);
nor U47164 (N_47164,N_35094,N_35547);
nand U47165 (N_47165,N_35776,N_32743);
nand U47166 (N_47166,N_36808,N_35179);
or U47167 (N_47167,N_37003,N_34592);
and U47168 (N_47168,N_35099,N_30872);
or U47169 (N_47169,N_39054,N_32631);
nor U47170 (N_47170,N_32203,N_38818);
nand U47171 (N_47171,N_30402,N_36286);
and U47172 (N_47172,N_31373,N_39364);
or U47173 (N_47173,N_30158,N_30280);
nand U47174 (N_47174,N_35906,N_30238);
nor U47175 (N_47175,N_36371,N_32375);
and U47176 (N_47176,N_36758,N_37337);
xnor U47177 (N_47177,N_30044,N_34451);
xnor U47178 (N_47178,N_36079,N_35217);
or U47179 (N_47179,N_31286,N_34339);
or U47180 (N_47180,N_35865,N_31297);
nand U47181 (N_47181,N_38691,N_30421);
and U47182 (N_47182,N_34750,N_32316);
and U47183 (N_47183,N_35537,N_34703);
or U47184 (N_47184,N_32237,N_31054);
nand U47185 (N_47185,N_36761,N_32282);
or U47186 (N_47186,N_39501,N_35210);
nor U47187 (N_47187,N_36153,N_31925);
nand U47188 (N_47188,N_35467,N_37603);
or U47189 (N_47189,N_36794,N_38203);
and U47190 (N_47190,N_33674,N_33848);
or U47191 (N_47191,N_39193,N_36744);
or U47192 (N_47192,N_35830,N_32844);
or U47193 (N_47193,N_39047,N_38211);
nor U47194 (N_47194,N_33145,N_31419);
and U47195 (N_47195,N_34701,N_37087);
nor U47196 (N_47196,N_34781,N_36980);
and U47197 (N_47197,N_36794,N_39235);
xor U47198 (N_47198,N_37602,N_31243);
nand U47199 (N_47199,N_36834,N_38153);
nor U47200 (N_47200,N_39936,N_32853);
or U47201 (N_47201,N_36947,N_39209);
or U47202 (N_47202,N_32459,N_39952);
and U47203 (N_47203,N_35425,N_34756);
nand U47204 (N_47204,N_30019,N_30421);
or U47205 (N_47205,N_37091,N_33513);
xnor U47206 (N_47206,N_35317,N_31837);
xnor U47207 (N_47207,N_30339,N_37514);
and U47208 (N_47208,N_31072,N_35022);
or U47209 (N_47209,N_37799,N_31692);
nand U47210 (N_47210,N_30731,N_37902);
nor U47211 (N_47211,N_33565,N_36220);
or U47212 (N_47212,N_33150,N_33886);
nor U47213 (N_47213,N_32151,N_35143);
nor U47214 (N_47214,N_36025,N_36370);
nand U47215 (N_47215,N_35936,N_30445);
nor U47216 (N_47216,N_31279,N_34075);
and U47217 (N_47217,N_33700,N_32835);
or U47218 (N_47218,N_39257,N_33962);
nand U47219 (N_47219,N_35569,N_31577);
nand U47220 (N_47220,N_38514,N_33887);
nand U47221 (N_47221,N_31630,N_32751);
nand U47222 (N_47222,N_30677,N_35573);
nor U47223 (N_47223,N_39904,N_34090);
and U47224 (N_47224,N_36288,N_34839);
and U47225 (N_47225,N_37181,N_32639);
nand U47226 (N_47226,N_37596,N_31057);
nor U47227 (N_47227,N_30793,N_37260);
nand U47228 (N_47228,N_32793,N_31699);
and U47229 (N_47229,N_38752,N_38054);
nor U47230 (N_47230,N_37836,N_33009);
and U47231 (N_47231,N_36954,N_35599);
or U47232 (N_47232,N_30874,N_35640);
or U47233 (N_47233,N_31022,N_36811);
or U47234 (N_47234,N_38851,N_36095);
and U47235 (N_47235,N_35628,N_31415);
nor U47236 (N_47236,N_33780,N_35718);
nand U47237 (N_47237,N_36930,N_36715);
and U47238 (N_47238,N_32839,N_37608);
and U47239 (N_47239,N_36174,N_33434);
or U47240 (N_47240,N_33527,N_31213);
nand U47241 (N_47241,N_30577,N_37558);
or U47242 (N_47242,N_34919,N_34789);
and U47243 (N_47243,N_30256,N_31520);
nor U47244 (N_47244,N_36016,N_33455);
or U47245 (N_47245,N_38818,N_38320);
or U47246 (N_47246,N_32215,N_39668);
nand U47247 (N_47247,N_35519,N_30219);
or U47248 (N_47248,N_34646,N_32657);
nor U47249 (N_47249,N_34338,N_36708);
and U47250 (N_47250,N_37398,N_39013);
and U47251 (N_47251,N_38571,N_39326);
or U47252 (N_47252,N_36665,N_37572);
and U47253 (N_47253,N_31609,N_36409);
or U47254 (N_47254,N_30047,N_36398);
xor U47255 (N_47255,N_35370,N_34049);
xnor U47256 (N_47256,N_30871,N_35690);
and U47257 (N_47257,N_31390,N_37529);
nor U47258 (N_47258,N_32345,N_32855);
nand U47259 (N_47259,N_33158,N_33096);
nand U47260 (N_47260,N_30455,N_32295);
nor U47261 (N_47261,N_34545,N_36430);
xor U47262 (N_47262,N_37729,N_36638);
and U47263 (N_47263,N_38634,N_32663);
nand U47264 (N_47264,N_39383,N_38647);
nand U47265 (N_47265,N_35949,N_35231);
or U47266 (N_47266,N_33704,N_33388);
and U47267 (N_47267,N_38637,N_30654);
nor U47268 (N_47268,N_38560,N_37352);
and U47269 (N_47269,N_31828,N_37723);
nand U47270 (N_47270,N_30400,N_32044);
or U47271 (N_47271,N_34886,N_34090);
nand U47272 (N_47272,N_30064,N_32254);
nor U47273 (N_47273,N_35883,N_39417);
nand U47274 (N_47274,N_36424,N_36976);
and U47275 (N_47275,N_34088,N_34188);
nor U47276 (N_47276,N_32395,N_33918);
and U47277 (N_47277,N_36785,N_35216);
nor U47278 (N_47278,N_38299,N_33810);
or U47279 (N_47279,N_35299,N_36301);
nor U47280 (N_47280,N_35000,N_34314);
xor U47281 (N_47281,N_31577,N_36357);
and U47282 (N_47282,N_38482,N_35602);
xor U47283 (N_47283,N_33893,N_36753);
nor U47284 (N_47284,N_32563,N_35124);
or U47285 (N_47285,N_35004,N_36061);
xnor U47286 (N_47286,N_31631,N_39602);
nor U47287 (N_47287,N_33909,N_39014);
nor U47288 (N_47288,N_30324,N_36947);
and U47289 (N_47289,N_34448,N_32730);
or U47290 (N_47290,N_38701,N_31915);
or U47291 (N_47291,N_31764,N_34031);
or U47292 (N_47292,N_39941,N_32199);
nand U47293 (N_47293,N_32448,N_36386);
and U47294 (N_47294,N_39309,N_36943);
and U47295 (N_47295,N_38738,N_34391);
xor U47296 (N_47296,N_30145,N_37880);
nor U47297 (N_47297,N_37436,N_33041);
nor U47298 (N_47298,N_36258,N_31658);
nor U47299 (N_47299,N_33296,N_38169);
xnor U47300 (N_47300,N_32304,N_32661);
and U47301 (N_47301,N_30944,N_31332);
or U47302 (N_47302,N_32570,N_38026);
or U47303 (N_47303,N_30373,N_30423);
nor U47304 (N_47304,N_30079,N_31100);
or U47305 (N_47305,N_31047,N_39594);
nor U47306 (N_47306,N_33409,N_33403);
and U47307 (N_47307,N_37661,N_34511);
nor U47308 (N_47308,N_37226,N_33282);
nor U47309 (N_47309,N_35842,N_30182);
or U47310 (N_47310,N_39200,N_35098);
nor U47311 (N_47311,N_39583,N_34562);
or U47312 (N_47312,N_35580,N_36171);
nor U47313 (N_47313,N_33964,N_38299);
nor U47314 (N_47314,N_34580,N_39481);
xor U47315 (N_47315,N_39133,N_37273);
or U47316 (N_47316,N_38755,N_35887);
xor U47317 (N_47317,N_30868,N_34231);
nand U47318 (N_47318,N_30556,N_34105);
and U47319 (N_47319,N_32664,N_38862);
nand U47320 (N_47320,N_32090,N_36260);
xor U47321 (N_47321,N_36922,N_34263);
and U47322 (N_47322,N_36080,N_31253);
and U47323 (N_47323,N_31421,N_33493);
xor U47324 (N_47324,N_39639,N_38272);
and U47325 (N_47325,N_33749,N_35274);
and U47326 (N_47326,N_32343,N_32044);
nor U47327 (N_47327,N_35129,N_39303);
or U47328 (N_47328,N_35163,N_32730);
nand U47329 (N_47329,N_31727,N_31213);
and U47330 (N_47330,N_33461,N_39679);
and U47331 (N_47331,N_37173,N_35994);
and U47332 (N_47332,N_38094,N_36481);
and U47333 (N_47333,N_31285,N_32975);
nand U47334 (N_47334,N_33305,N_33988);
nand U47335 (N_47335,N_34918,N_30908);
or U47336 (N_47336,N_31643,N_33628);
nor U47337 (N_47337,N_33370,N_36340);
and U47338 (N_47338,N_37193,N_38102);
or U47339 (N_47339,N_35442,N_38288);
nand U47340 (N_47340,N_34542,N_31620);
nor U47341 (N_47341,N_30462,N_35168);
nor U47342 (N_47342,N_39574,N_37799);
nor U47343 (N_47343,N_35230,N_33086);
nor U47344 (N_47344,N_32634,N_39541);
nand U47345 (N_47345,N_30757,N_34327);
nor U47346 (N_47346,N_33859,N_31423);
xor U47347 (N_47347,N_37506,N_31140);
or U47348 (N_47348,N_39830,N_32699);
nand U47349 (N_47349,N_38732,N_30974);
nand U47350 (N_47350,N_35755,N_37353);
nand U47351 (N_47351,N_32967,N_31043);
nor U47352 (N_47352,N_35583,N_35497);
or U47353 (N_47353,N_31853,N_32017);
nor U47354 (N_47354,N_39513,N_35639);
nand U47355 (N_47355,N_32494,N_30610);
nand U47356 (N_47356,N_31129,N_32277);
or U47357 (N_47357,N_37978,N_30351);
or U47358 (N_47358,N_31686,N_39544);
nand U47359 (N_47359,N_33882,N_38705);
or U47360 (N_47360,N_31679,N_32220);
xnor U47361 (N_47361,N_39985,N_32577);
or U47362 (N_47362,N_37934,N_32779);
and U47363 (N_47363,N_31568,N_39054);
and U47364 (N_47364,N_38915,N_36568);
xor U47365 (N_47365,N_32201,N_30807);
and U47366 (N_47366,N_36782,N_39389);
and U47367 (N_47367,N_36110,N_39831);
or U47368 (N_47368,N_36856,N_32607);
and U47369 (N_47369,N_30623,N_31437);
xnor U47370 (N_47370,N_30178,N_38954);
and U47371 (N_47371,N_35333,N_37436);
nand U47372 (N_47372,N_33562,N_36757);
or U47373 (N_47373,N_37306,N_36106);
and U47374 (N_47374,N_34404,N_39163);
or U47375 (N_47375,N_31390,N_38827);
nor U47376 (N_47376,N_37988,N_36603);
nor U47377 (N_47377,N_37198,N_39066);
nor U47378 (N_47378,N_33578,N_33980);
nor U47379 (N_47379,N_38347,N_36814);
or U47380 (N_47380,N_35703,N_36046);
and U47381 (N_47381,N_38800,N_31062);
nand U47382 (N_47382,N_38977,N_34521);
xnor U47383 (N_47383,N_35828,N_33302);
nand U47384 (N_47384,N_33423,N_35875);
nor U47385 (N_47385,N_34839,N_36263);
nand U47386 (N_47386,N_31806,N_32736);
nor U47387 (N_47387,N_36458,N_39551);
or U47388 (N_47388,N_37882,N_34114);
nand U47389 (N_47389,N_39541,N_36296);
nand U47390 (N_47390,N_34652,N_33460);
nor U47391 (N_47391,N_33559,N_38521);
nand U47392 (N_47392,N_38919,N_31766);
nor U47393 (N_47393,N_38198,N_31267);
or U47394 (N_47394,N_37590,N_36804);
xnor U47395 (N_47395,N_31863,N_36512);
and U47396 (N_47396,N_36286,N_39403);
xnor U47397 (N_47397,N_33719,N_35321);
nand U47398 (N_47398,N_37795,N_35215);
nand U47399 (N_47399,N_35405,N_38379);
and U47400 (N_47400,N_35522,N_35542);
nor U47401 (N_47401,N_33186,N_34765);
nor U47402 (N_47402,N_36391,N_36779);
nor U47403 (N_47403,N_37333,N_35858);
nand U47404 (N_47404,N_33138,N_34351);
and U47405 (N_47405,N_35887,N_35107);
nand U47406 (N_47406,N_32316,N_34019);
and U47407 (N_47407,N_37082,N_31941);
and U47408 (N_47408,N_30766,N_37359);
nor U47409 (N_47409,N_37763,N_32743);
and U47410 (N_47410,N_33489,N_31661);
and U47411 (N_47411,N_39696,N_33039);
xnor U47412 (N_47412,N_36259,N_35614);
or U47413 (N_47413,N_38319,N_36394);
and U47414 (N_47414,N_39759,N_30678);
and U47415 (N_47415,N_33445,N_36513);
nor U47416 (N_47416,N_34079,N_37730);
nor U47417 (N_47417,N_30458,N_30226);
xnor U47418 (N_47418,N_31975,N_31227);
nand U47419 (N_47419,N_33450,N_35664);
nand U47420 (N_47420,N_30312,N_38460);
or U47421 (N_47421,N_36489,N_38159);
nor U47422 (N_47422,N_32130,N_33132);
nor U47423 (N_47423,N_30748,N_30326);
xnor U47424 (N_47424,N_31385,N_33211);
and U47425 (N_47425,N_35052,N_36382);
nor U47426 (N_47426,N_31583,N_37642);
or U47427 (N_47427,N_31951,N_35305);
xor U47428 (N_47428,N_30899,N_30758);
or U47429 (N_47429,N_36079,N_33986);
nand U47430 (N_47430,N_37436,N_33061);
nand U47431 (N_47431,N_35559,N_37319);
xor U47432 (N_47432,N_32617,N_35187);
and U47433 (N_47433,N_33725,N_33520);
nand U47434 (N_47434,N_34476,N_37984);
and U47435 (N_47435,N_31426,N_38371);
or U47436 (N_47436,N_31323,N_38401);
nor U47437 (N_47437,N_30689,N_38160);
or U47438 (N_47438,N_30934,N_38983);
xnor U47439 (N_47439,N_36433,N_39511);
or U47440 (N_47440,N_39602,N_32815);
xor U47441 (N_47441,N_32709,N_37213);
or U47442 (N_47442,N_39437,N_30026);
or U47443 (N_47443,N_33546,N_33677);
or U47444 (N_47444,N_31167,N_30680);
nor U47445 (N_47445,N_39092,N_39876);
nand U47446 (N_47446,N_39132,N_38708);
nor U47447 (N_47447,N_38024,N_36921);
or U47448 (N_47448,N_34504,N_35040);
or U47449 (N_47449,N_32846,N_37959);
and U47450 (N_47450,N_33856,N_36244);
and U47451 (N_47451,N_37703,N_39876);
and U47452 (N_47452,N_31368,N_37393);
nand U47453 (N_47453,N_35834,N_37088);
nand U47454 (N_47454,N_39390,N_33808);
nor U47455 (N_47455,N_33521,N_37327);
or U47456 (N_47456,N_34920,N_36911);
and U47457 (N_47457,N_34548,N_32424);
nor U47458 (N_47458,N_34153,N_31089);
nand U47459 (N_47459,N_34500,N_31749);
and U47460 (N_47460,N_38308,N_34242);
nor U47461 (N_47461,N_31672,N_38997);
and U47462 (N_47462,N_35114,N_38997);
or U47463 (N_47463,N_35616,N_31069);
nand U47464 (N_47464,N_36768,N_35342);
nor U47465 (N_47465,N_34924,N_38982);
xor U47466 (N_47466,N_31423,N_36655);
nor U47467 (N_47467,N_36785,N_33267);
or U47468 (N_47468,N_32653,N_30903);
or U47469 (N_47469,N_37644,N_35372);
or U47470 (N_47470,N_36627,N_30820);
or U47471 (N_47471,N_31763,N_36278);
nand U47472 (N_47472,N_38897,N_36488);
nor U47473 (N_47473,N_35843,N_33741);
nor U47474 (N_47474,N_30592,N_32057);
and U47475 (N_47475,N_31190,N_33713);
xnor U47476 (N_47476,N_36924,N_30420);
nor U47477 (N_47477,N_36949,N_35802);
or U47478 (N_47478,N_37571,N_32790);
nor U47479 (N_47479,N_31961,N_37736);
and U47480 (N_47480,N_33187,N_34246);
nand U47481 (N_47481,N_31177,N_39173);
and U47482 (N_47482,N_38414,N_35074);
or U47483 (N_47483,N_37675,N_33545);
or U47484 (N_47484,N_31189,N_38560);
and U47485 (N_47485,N_39199,N_37165);
or U47486 (N_47486,N_30897,N_37139);
or U47487 (N_47487,N_33368,N_34568);
nor U47488 (N_47488,N_34747,N_30430);
nor U47489 (N_47489,N_38016,N_31002);
nor U47490 (N_47490,N_38899,N_37987);
and U47491 (N_47491,N_36321,N_33341);
and U47492 (N_47492,N_31021,N_36178);
and U47493 (N_47493,N_32987,N_39933);
nor U47494 (N_47494,N_33204,N_39425);
and U47495 (N_47495,N_33270,N_31223);
or U47496 (N_47496,N_33974,N_33045);
nand U47497 (N_47497,N_37732,N_37222);
xor U47498 (N_47498,N_30698,N_37417);
or U47499 (N_47499,N_39774,N_36124);
nor U47500 (N_47500,N_37358,N_38903);
nor U47501 (N_47501,N_30048,N_38507);
or U47502 (N_47502,N_30175,N_34529);
nor U47503 (N_47503,N_31373,N_38304);
or U47504 (N_47504,N_33169,N_38507);
xor U47505 (N_47505,N_35692,N_36971);
nor U47506 (N_47506,N_36660,N_34076);
nor U47507 (N_47507,N_35457,N_38309);
or U47508 (N_47508,N_33288,N_38391);
or U47509 (N_47509,N_30468,N_32886);
or U47510 (N_47510,N_38673,N_31336);
nor U47511 (N_47511,N_33747,N_34048);
nand U47512 (N_47512,N_38418,N_39178);
and U47513 (N_47513,N_34776,N_38653);
or U47514 (N_47514,N_34473,N_36986);
or U47515 (N_47515,N_35385,N_39264);
nand U47516 (N_47516,N_33362,N_37973);
or U47517 (N_47517,N_33727,N_35943);
nand U47518 (N_47518,N_38440,N_39741);
and U47519 (N_47519,N_36907,N_34887);
nand U47520 (N_47520,N_33166,N_36381);
and U47521 (N_47521,N_39658,N_33919);
nand U47522 (N_47522,N_33436,N_34899);
nand U47523 (N_47523,N_34277,N_32555);
or U47524 (N_47524,N_30840,N_37272);
and U47525 (N_47525,N_32844,N_36941);
and U47526 (N_47526,N_37457,N_37043);
and U47527 (N_47527,N_32781,N_38274);
or U47528 (N_47528,N_36538,N_38140);
nor U47529 (N_47529,N_39435,N_30428);
nor U47530 (N_47530,N_36396,N_37804);
and U47531 (N_47531,N_36957,N_35878);
nor U47532 (N_47532,N_33354,N_32117);
xnor U47533 (N_47533,N_36717,N_39885);
and U47534 (N_47534,N_35961,N_34872);
or U47535 (N_47535,N_33061,N_37902);
and U47536 (N_47536,N_38648,N_33260);
nor U47537 (N_47537,N_33253,N_35896);
xnor U47538 (N_47538,N_39107,N_33516);
nor U47539 (N_47539,N_35012,N_31448);
nor U47540 (N_47540,N_36674,N_30419);
or U47541 (N_47541,N_30664,N_33552);
or U47542 (N_47542,N_33579,N_38456);
nand U47543 (N_47543,N_31176,N_35667);
nor U47544 (N_47544,N_33696,N_35597);
and U47545 (N_47545,N_35696,N_39126);
nand U47546 (N_47546,N_36575,N_32902);
nand U47547 (N_47547,N_33368,N_33433);
or U47548 (N_47548,N_39806,N_34185);
nand U47549 (N_47549,N_30490,N_34494);
nor U47550 (N_47550,N_31201,N_33379);
or U47551 (N_47551,N_30186,N_32498);
and U47552 (N_47552,N_33908,N_36565);
nand U47553 (N_47553,N_32643,N_31135);
or U47554 (N_47554,N_32189,N_39878);
nor U47555 (N_47555,N_35836,N_33633);
nand U47556 (N_47556,N_30900,N_36854);
and U47557 (N_47557,N_33712,N_39581);
and U47558 (N_47558,N_31695,N_38237);
or U47559 (N_47559,N_30614,N_35910);
and U47560 (N_47560,N_35950,N_33066);
and U47561 (N_47561,N_32076,N_39306);
nor U47562 (N_47562,N_38008,N_33355);
or U47563 (N_47563,N_38602,N_33056);
and U47564 (N_47564,N_33286,N_36835);
nor U47565 (N_47565,N_35037,N_38239);
or U47566 (N_47566,N_34561,N_39642);
and U47567 (N_47567,N_36159,N_34999);
and U47568 (N_47568,N_38098,N_38932);
or U47569 (N_47569,N_33495,N_31840);
or U47570 (N_47570,N_31133,N_38772);
or U47571 (N_47571,N_36943,N_31683);
or U47572 (N_47572,N_39837,N_35796);
nor U47573 (N_47573,N_34734,N_39971);
nor U47574 (N_47574,N_30717,N_30120);
and U47575 (N_47575,N_32122,N_32812);
nand U47576 (N_47576,N_31496,N_30602);
nor U47577 (N_47577,N_30285,N_38557);
or U47578 (N_47578,N_31546,N_33022);
nand U47579 (N_47579,N_35957,N_36240);
nor U47580 (N_47580,N_35960,N_37771);
nor U47581 (N_47581,N_31923,N_38149);
nand U47582 (N_47582,N_31985,N_31049);
nand U47583 (N_47583,N_32425,N_39106);
nand U47584 (N_47584,N_32961,N_36218);
nand U47585 (N_47585,N_33428,N_31991);
and U47586 (N_47586,N_31348,N_39262);
and U47587 (N_47587,N_35186,N_31150);
or U47588 (N_47588,N_38332,N_31011);
nor U47589 (N_47589,N_31905,N_34590);
nand U47590 (N_47590,N_37840,N_39654);
and U47591 (N_47591,N_35341,N_36269);
xor U47592 (N_47592,N_33853,N_30467);
or U47593 (N_47593,N_33322,N_34307);
or U47594 (N_47594,N_30030,N_37535);
nand U47595 (N_47595,N_38948,N_34812);
and U47596 (N_47596,N_37134,N_39912);
and U47597 (N_47597,N_38782,N_32858);
nand U47598 (N_47598,N_30320,N_30989);
nand U47599 (N_47599,N_38430,N_31327);
nor U47600 (N_47600,N_32906,N_38965);
and U47601 (N_47601,N_38842,N_36970);
nand U47602 (N_47602,N_34473,N_39214);
nor U47603 (N_47603,N_37661,N_32021);
nand U47604 (N_47604,N_35627,N_31548);
and U47605 (N_47605,N_34525,N_39256);
or U47606 (N_47606,N_30279,N_33297);
and U47607 (N_47607,N_39359,N_36418);
nor U47608 (N_47608,N_30993,N_34277);
or U47609 (N_47609,N_34710,N_33977);
nand U47610 (N_47610,N_34584,N_35081);
and U47611 (N_47611,N_34307,N_32092);
nand U47612 (N_47612,N_39656,N_34625);
nor U47613 (N_47613,N_30078,N_34431);
or U47614 (N_47614,N_37298,N_36208);
xnor U47615 (N_47615,N_33654,N_38672);
nand U47616 (N_47616,N_33096,N_39870);
nand U47617 (N_47617,N_33898,N_30157);
nor U47618 (N_47618,N_36652,N_33269);
xnor U47619 (N_47619,N_35614,N_39287);
nor U47620 (N_47620,N_34745,N_32705);
and U47621 (N_47621,N_39416,N_32200);
nor U47622 (N_47622,N_34383,N_32694);
and U47623 (N_47623,N_39842,N_32876);
and U47624 (N_47624,N_34943,N_34341);
xor U47625 (N_47625,N_32648,N_31616);
nor U47626 (N_47626,N_34981,N_30344);
nor U47627 (N_47627,N_36732,N_30873);
nand U47628 (N_47628,N_31628,N_39149);
or U47629 (N_47629,N_38341,N_32709);
and U47630 (N_47630,N_33423,N_35715);
or U47631 (N_47631,N_36662,N_36582);
and U47632 (N_47632,N_39572,N_37841);
and U47633 (N_47633,N_36678,N_32134);
and U47634 (N_47634,N_30510,N_31232);
nand U47635 (N_47635,N_35698,N_37357);
or U47636 (N_47636,N_39240,N_35268);
and U47637 (N_47637,N_39048,N_33236);
or U47638 (N_47638,N_32788,N_32263);
or U47639 (N_47639,N_36096,N_36022);
or U47640 (N_47640,N_38391,N_37755);
nand U47641 (N_47641,N_38009,N_30680);
or U47642 (N_47642,N_39986,N_37292);
and U47643 (N_47643,N_34409,N_35643);
and U47644 (N_47644,N_31865,N_35762);
nand U47645 (N_47645,N_38138,N_30961);
and U47646 (N_47646,N_31772,N_34963);
or U47647 (N_47647,N_36740,N_32689);
nor U47648 (N_47648,N_32608,N_32733);
nor U47649 (N_47649,N_37420,N_39085);
nand U47650 (N_47650,N_35735,N_34886);
and U47651 (N_47651,N_37635,N_38959);
or U47652 (N_47652,N_33625,N_38910);
and U47653 (N_47653,N_35198,N_32734);
nand U47654 (N_47654,N_35320,N_39143);
nor U47655 (N_47655,N_35341,N_38602);
and U47656 (N_47656,N_30776,N_38119);
nand U47657 (N_47657,N_35211,N_39491);
or U47658 (N_47658,N_36015,N_37103);
and U47659 (N_47659,N_31242,N_37556);
or U47660 (N_47660,N_33486,N_33043);
and U47661 (N_47661,N_33839,N_36866);
nand U47662 (N_47662,N_30605,N_32447);
or U47663 (N_47663,N_30447,N_34443);
and U47664 (N_47664,N_34749,N_37142);
nor U47665 (N_47665,N_33894,N_34067);
and U47666 (N_47666,N_30842,N_33716);
and U47667 (N_47667,N_34183,N_38706);
nor U47668 (N_47668,N_38374,N_39789);
or U47669 (N_47669,N_38028,N_30395);
and U47670 (N_47670,N_39233,N_30941);
or U47671 (N_47671,N_39936,N_38892);
or U47672 (N_47672,N_39034,N_37290);
nand U47673 (N_47673,N_35816,N_31716);
nor U47674 (N_47674,N_30781,N_37800);
or U47675 (N_47675,N_38996,N_39683);
and U47676 (N_47676,N_31124,N_35887);
nand U47677 (N_47677,N_36495,N_33111);
or U47678 (N_47678,N_35907,N_30534);
nor U47679 (N_47679,N_39388,N_39977);
and U47680 (N_47680,N_31778,N_34290);
nor U47681 (N_47681,N_34594,N_37661);
and U47682 (N_47682,N_37170,N_38908);
nand U47683 (N_47683,N_39245,N_38691);
nor U47684 (N_47684,N_32153,N_32630);
nand U47685 (N_47685,N_38239,N_33807);
nand U47686 (N_47686,N_34801,N_30281);
or U47687 (N_47687,N_33204,N_35612);
or U47688 (N_47688,N_30492,N_30708);
nor U47689 (N_47689,N_32168,N_34235);
or U47690 (N_47690,N_39862,N_31961);
or U47691 (N_47691,N_36765,N_38570);
nand U47692 (N_47692,N_33454,N_32884);
nand U47693 (N_47693,N_36050,N_35687);
nand U47694 (N_47694,N_37390,N_32342);
and U47695 (N_47695,N_39659,N_32227);
xnor U47696 (N_47696,N_32602,N_35159);
or U47697 (N_47697,N_31063,N_34506);
or U47698 (N_47698,N_30003,N_37358);
nor U47699 (N_47699,N_31624,N_37200);
or U47700 (N_47700,N_38812,N_37281);
nand U47701 (N_47701,N_32374,N_32981);
or U47702 (N_47702,N_30218,N_38350);
nor U47703 (N_47703,N_33046,N_32038);
or U47704 (N_47704,N_30258,N_33712);
nor U47705 (N_47705,N_39295,N_36873);
or U47706 (N_47706,N_37941,N_37593);
xnor U47707 (N_47707,N_35540,N_38865);
xor U47708 (N_47708,N_38758,N_31971);
and U47709 (N_47709,N_31156,N_37789);
xnor U47710 (N_47710,N_30886,N_35858);
or U47711 (N_47711,N_38900,N_33544);
nand U47712 (N_47712,N_35442,N_32522);
nand U47713 (N_47713,N_33034,N_37898);
xnor U47714 (N_47714,N_34457,N_32150);
nor U47715 (N_47715,N_33556,N_30015);
xor U47716 (N_47716,N_30011,N_30501);
nor U47717 (N_47717,N_33931,N_33887);
nor U47718 (N_47718,N_35302,N_35054);
nor U47719 (N_47719,N_33453,N_34420);
nand U47720 (N_47720,N_37868,N_39513);
and U47721 (N_47721,N_33542,N_33810);
nand U47722 (N_47722,N_34953,N_35357);
nor U47723 (N_47723,N_37728,N_39865);
or U47724 (N_47724,N_34883,N_33019);
nor U47725 (N_47725,N_36742,N_37372);
nand U47726 (N_47726,N_39019,N_38562);
nand U47727 (N_47727,N_36320,N_33781);
nor U47728 (N_47728,N_36672,N_36409);
nand U47729 (N_47729,N_34243,N_35423);
and U47730 (N_47730,N_30192,N_38543);
nand U47731 (N_47731,N_39192,N_35243);
and U47732 (N_47732,N_34371,N_36525);
and U47733 (N_47733,N_33544,N_32162);
nand U47734 (N_47734,N_34399,N_30396);
or U47735 (N_47735,N_37707,N_31176);
or U47736 (N_47736,N_30681,N_38921);
nor U47737 (N_47737,N_32065,N_35260);
nand U47738 (N_47738,N_34407,N_32305);
nand U47739 (N_47739,N_37113,N_38265);
nor U47740 (N_47740,N_30994,N_38942);
and U47741 (N_47741,N_31694,N_33316);
and U47742 (N_47742,N_32825,N_39320);
nor U47743 (N_47743,N_32534,N_32623);
and U47744 (N_47744,N_31241,N_34900);
nor U47745 (N_47745,N_32108,N_39224);
and U47746 (N_47746,N_31160,N_36428);
nor U47747 (N_47747,N_34885,N_33486);
and U47748 (N_47748,N_30652,N_30061);
nand U47749 (N_47749,N_31103,N_39957);
nand U47750 (N_47750,N_30541,N_38202);
nor U47751 (N_47751,N_35171,N_35262);
and U47752 (N_47752,N_33631,N_36324);
and U47753 (N_47753,N_39645,N_30608);
nor U47754 (N_47754,N_34099,N_32162);
nand U47755 (N_47755,N_32636,N_31153);
or U47756 (N_47756,N_35436,N_30882);
or U47757 (N_47757,N_33706,N_37451);
nand U47758 (N_47758,N_39119,N_30317);
nor U47759 (N_47759,N_35732,N_35538);
nand U47760 (N_47760,N_33817,N_37492);
nor U47761 (N_47761,N_31183,N_32180);
and U47762 (N_47762,N_31201,N_34710);
or U47763 (N_47763,N_39063,N_36819);
or U47764 (N_47764,N_35818,N_34717);
or U47765 (N_47765,N_34417,N_33860);
or U47766 (N_47766,N_33877,N_34240);
xnor U47767 (N_47767,N_33852,N_39525);
nand U47768 (N_47768,N_31552,N_36852);
nand U47769 (N_47769,N_37334,N_31698);
and U47770 (N_47770,N_32474,N_32547);
and U47771 (N_47771,N_35708,N_36184);
and U47772 (N_47772,N_34592,N_31209);
and U47773 (N_47773,N_35604,N_31852);
nor U47774 (N_47774,N_31678,N_31053);
xnor U47775 (N_47775,N_35842,N_33513);
and U47776 (N_47776,N_31206,N_38993);
or U47777 (N_47777,N_35966,N_39859);
and U47778 (N_47778,N_39664,N_32634);
nand U47779 (N_47779,N_38134,N_39730);
nor U47780 (N_47780,N_35258,N_34930);
nand U47781 (N_47781,N_33789,N_37311);
nand U47782 (N_47782,N_30093,N_34812);
and U47783 (N_47783,N_30355,N_34049);
nor U47784 (N_47784,N_32853,N_32565);
xor U47785 (N_47785,N_36840,N_32250);
and U47786 (N_47786,N_36708,N_36682);
nor U47787 (N_47787,N_31315,N_31381);
and U47788 (N_47788,N_30606,N_30332);
and U47789 (N_47789,N_30114,N_36789);
nor U47790 (N_47790,N_34258,N_34146);
nand U47791 (N_47791,N_38793,N_34765);
nor U47792 (N_47792,N_34565,N_38448);
or U47793 (N_47793,N_33045,N_38486);
or U47794 (N_47794,N_31190,N_35499);
nand U47795 (N_47795,N_32992,N_34122);
nor U47796 (N_47796,N_36165,N_37156);
nand U47797 (N_47797,N_31854,N_33365);
nor U47798 (N_47798,N_39934,N_32391);
or U47799 (N_47799,N_30974,N_32312);
and U47800 (N_47800,N_39452,N_34086);
or U47801 (N_47801,N_38283,N_31636);
or U47802 (N_47802,N_30546,N_32581);
and U47803 (N_47803,N_37331,N_32293);
nand U47804 (N_47804,N_33777,N_38380);
nand U47805 (N_47805,N_34311,N_33048);
nand U47806 (N_47806,N_35858,N_32709);
and U47807 (N_47807,N_32576,N_35328);
nor U47808 (N_47808,N_39792,N_33641);
nand U47809 (N_47809,N_38031,N_33450);
and U47810 (N_47810,N_33016,N_31330);
nor U47811 (N_47811,N_33050,N_36992);
nor U47812 (N_47812,N_36068,N_35900);
or U47813 (N_47813,N_37445,N_34161);
nand U47814 (N_47814,N_30046,N_38936);
xnor U47815 (N_47815,N_37544,N_34923);
nand U47816 (N_47816,N_33588,N_38844);
and U47817 (N_47817,N_30371,N_34260);
and U47818 (N_47818,N_30517,N_39591);
nor U47819 (N_47819,N_37328,N_36982);
nor U47820 (N_47820,N_33430,N_36682);
and U47821 (N_47821,N_36109,N_30357);
or U47822 (N_47822,N_36992,N_37780);
or U47823 (N_47823,N_39186,N_36749);
or U47824 (N_47824,N_32855,N_33301);
nor U47825 (N_47825,N_37715,N_33400);
and U47826 (N_47826,N_35889,N_37711);
or U47827 (N_47827,N_39995,N_39642);
and U47828 (N_47828,N_33656,N_33250);
xor U47829 (N_47829,N_31214,N_34673);
nor U47830 (N_47830,N_33122,N_32738);
or U47831 (N_47831,N_33449,N_31079);
nand U47832 (N_47832,N_34982,N_33410);
or U47833 (N_47833,N_33639,N_35611);
and U47834 (N_47834,N_35485,N_35243);
nand U47835 (N_47835,N_37390,N_39528);
xor U47836 (N_47836,N_35339,N_39012);
or U47837 (N_47837,N_33934,N_34753);
or U47838 (N_47838,N_39867,N_34182);
and U47839 (N_47839,N_39153,N_30105);
nor U47840 (N_47840,N_38830,N_34481);
xnor U47841 (N_47841,N_33493,N_32156);
nor U47842 (N_47842,N_35537,N_31791);
and U47843 (N_47843,N_31640,N_37155);
and U47844 (N_47844,N_35018,N_35252);
or U47845 (N_47845,N_38598,N_39239);
nand U47846 (N_47846,N_32032,N_37483);
and U47847 (N_47847,N_33566,N_37968);
and U47848 (N_47848,N_39072,N_39527);
and U47849 (N_47849,N_35756,N_35599);
and U47850 (N_47850,N_32870,N_36397);
or U47851 (N_47851,N_36236,N_39823);
or U47852 (N_47852,N_33206,N_36531);
xnor U47853 (N_47853,N_31587,N_33872);
nor U47854 (N_47854,N_36289,N_36019);
and U47855 (N_47855,N_39507,N_32569);
nand U47856 (N_47856,N_35205,N_35280);
or U47857 (N_47857,N_30310,N_31215);
and U47858 (N_47858,N_33981,N_35209);
xor U47859 (N_47859,N_37433,N_31257);
and U47860 (N_47860,N_31367,N_36741);
nand U47861 (N_47861,N_39449,N_32518);
nand U47862 (N_47862,N_33090,N_37114);
or U47863 (N_47863,N_33744,N_33753);
and U47864 (N_47864,N_39305,N_32372);
or U47865 (N_47865,N_33585,N_39472);
or U47866 (N_47866,N_31846,N_32221);
or U47867 (N_47867,N_31057,N_30762);
and U47868 (N_47868,N_30929,N_35656);
nand U47869 (N_47869,N_35884,N_31964);
nor U47870 (N_47870,N_38886,N_34596);
nand U47871 (N_47871,N_31800,N_36864);
and U47872 (N_47872,N_37457,N_39043);
nand U47873 (N_47873,N_39824,N_37768);
nor U47874 (N_47874,N_31646,N_32231);
xor U47875 (N_47875,N_32852,N_36856);
or U47876 (N_47876,N_38096,N_38251);
or U47877 (N_47877,N_32201,N_37859);
nor U47878 (N_47878,N_34802,N_35391);
or U47879 (N_47879,N_39208,N_37830);
and U47880 (N_47880,N_36756,N_36828);
nand U47881 (N_47881,N_37835,N_33338);
and U47882 (N_47882,N_35786,N_33252);
or U47883 (N_47883,N_30754,N_30930);
xor U47884 (N_47884,N_38047,N_34875);
or U47885 (N_47885,N_39003,N_39969);
nor U47886 (N_47886,N_34410,N_30057);
and U47887 (N_47887,N_34893,N_30829);
nor U47888 (N_47888,N_33361,N_32343);
and U47889 (N_47889,N_37123,N_31999);
and U47890 (N_47890,N_35357,N_38474);
nand U47891 (N_47891,N_38501,N_33389);
or U47892 (N_47892,N_30669,N_38013);
nand U47893 (N_47893,N_30792,N_33785);
or U47894 (N_47894,N_38395,N_34547);
and U47895 (N_47895,N_36077,N_36628);
nor U47896 (N_47896,N_33205,N_36987);
and U47897 (N_47897,N_38342,N_33592);
xor U47898 (N_47898,N_33436,N_36028);
or U47899 (N_47899,N_32230,N_38980);
xnor U47900 (N_47900,N_31585,N_38211);
nand U47901 (N_47901,N_32578,N_39873);
or U47902 (N_47902,N_36004,N_35295);
and U47903 (N_47903,N_33660,N_38065);
nand U47904 (N_47904,N_32823,N_35432);
xnor U47905 (N_47905,N_39241,N_37642);
nand U47906 (N_47906,N_32034,N_39693);
nand U47907 (N_47907,N_30866,N_32378);
nor U47908 (N_47908,N_33414,N_34597);
and U47909 (N_47909,N_36055,N_35236);
or U47910 (N_47910,N_34379,N_31780);
nor U47911 (N_47911,N_36985,N_34726);
xnor U47912 (N_47912,N_34343,N_30090);
and U47913 (N_47913,N_31912,N_35468);
nor U47914 (N_47914,N_36070,N_33047);
nor U47915 (N_47915,N_34710,N_33312);
and U47916 (N_47916,N_31707,N_35502);
and U47917 (N_47917,N_35567,N_38265);
or U47918 (N_47918,N_34532,N_33033);
xnor U47919 (N_47919,N_31988,N_34356);
xnor U47920 (N_47920,N_34140,N_33538);
xnor U47921 (N_47921,N_36901,N_39647);
and U47922 (N_47922,N_37121,N_36188);
xor U47923 (N_47923,N_30018,N_39097);
and U47924 (N_47924,N_35713,N_32270);
xnor U47925 (N_47925,N_35444,N_32102);
nor U47926 (N_47926,N_34870,N_31358);
nand U47927 (N_47927,N_39387,N_38824);
and U47928 (N_47928,N_34408,N_30179);
nand U47929 (N_47929,N_30920,N_35076);
xor U47930 (N_47930,N_37460,N_32691);
nor U47931 (N_47931,N_30111,N_39417);
and U47932 (N_47932,N_30689,N_36425);
and U47933 (N_47933,N_32382,N_34722);
nand U47934 (N_47934,N_35899,N_30364);
or U47935 (N_47935,N_31040,N_32619);
or U47936 (N_47936,N_39530,N_33256);
nand U47937 (N_47937,N_39984,N_38087);
and U47938 (N_47938,N_31156,N_39255);
nand U47939 (N_47939,N_31361,N_36517);
or U47940 (N_47940,N_33929,N_34631);
or U47941 (N_47941,N_33683,N_36402);
nor U47942 (N_47942,N_37345,N_39230);
nand U47943 (N_47943,N_33638,N_35574);
nor U47944 (N_47944,N_36533,N_38120);
nor U47945 (N_47945,N_36752,N_33746);
nand U47946 (N_47946,N_31864,N_36601);
nand U47947 (N_47947,N_37450,N_33336);
and U47948 (N_47948,N_33116,N_35480);
and U47949 (N_47949,N_39786,N_35152);
nor U47950 (N_47950,N_36190,N_35141);
and U47951 (N_47951,N_31264,N_31501);
and U47952 (N_47952,N_37498,N_32196);
or U47953 (N_47953,N_35199,N_35683);
nand U47954 (N_47954,N_39380,N_30264);
nor U47955 (N_47955,N_36469,N_38040);
and U47956 (N_47956,N_39782,N_35941);
or U47957 (N_47957,N_33897,N_36874);
or U47958 (N_47958,N_38475,N_36454);
and U47959 (N_47959,N_33736,N_38598);
xor U47960 (N_47960,N_39585,N_39891);
nor U47961 (N_47961,N_38615,N_32514);
and U47962 (N_47962,N_39151,N_30010);
and U47963 (N_47963,N_34647,N_37874);
nand U47964 (N_47964,N_30495,N_30672);
nor U47965 (N_47965,N_30575,N_37054);
nand U47966 (N_47966,N_37966,N_39206);
and U47967 (N_47967,N_39543,N_35161);
or U47968 (N_47968,N_39979,N_31571);
or U47969 (N_47969,N_39412,N_33007);
nor U47970 (N_47970,N_31109,N_38520);
nor U47971 (N_47971,N_36005,N_31290);
nor U47972 (N_47972,N_30009,N_38425);
or U47973 (N_47973,N_37309,N_33858);
nand U47974 (N_47974,N_34072,N_32769);
and U47975 (N_47975,N_36305,N_30270);
and U47976 (N_47976,N_30644,N_31469);
or U47977 (N_47977,N_30015,N_33203);
and U47978 (N_47978,N_39323,N_35955);
nand U47979 (N_47979,N_32058,N_39608);
nand U47980 (N_47980,N_30464,N_36339);
xnor U47981 (N_47981,N_39193,N_33101);
nand U47982 (N_47982,N_38956,N_32433);
xor U47983 (N_47983,N_37010,N_31770);
nor U47984 (N_47984,N_33540,N_37322);
or U47985 (N_47985,N_37556,N_37247);
or U47986 (N_47986,N_33495,N_30543);
nand U47987 (N_47987,N_35036,N_34051);
xnor U47988 (N_47988,N_36508,N_32749);
nand U47989 (N_47989,N_31444,N_37078);
nor U47990 (N_47990,N_36050,N_38865);
or U47991 (N_47991,N_36593,N_35096);
or U47992 (N_47992,N_31033,N_39150);
nand U47993 (N_47993,N_36063,N_33875);
and U47994 (N_47994,N_35855,N_36682);
or U47995 (N_47995,N_31583,N_35647);
or U47996 (N_47996,N_38559,N_39505);
nor U47997 (N_47997,N_38440,N_37313);
nor U47998 (N_47998,N_30808,N_34475);
or U47999 (N_47999,N_35933,N_34286);
nor U48000 (N_48000,N_31356,N_34998);
or U48001 (N_48001,N_30298,N_34403);
nand U48002 (N_48002,N_31657,N_38420);
or U48003 (N_48003,N_39954,N_35916);
and U48004 (N_48004,N_33175,N_39918);
or U48005 (N_48005,N_34482,N_38742);
and U48006 (N_48006,N_39760,N_34948);
and U48007 (N_48007,N_35362,N_39507);
xor U48008 (N_48008,N_32759,N_34172);
nor U48009 (N_48009,N_35228,N_34614);
nor U48010 (N_48010,N_38412,N_38500);
nor U48011 (N_48011,N_34675,N_35001);
or U48012 (N_48012,N_39543,N_39273);
xor U48013 (N_48013,N_32143,N_38262);
nand U48014 (N_48014,N_38696,N_37578);
and U48015 (N_48015,N_32391,N_31683);
or U48016 (N_48016,N_37648,N_33387);
nor U48017 (N_48017,N_30411,N_35317);
nand U48018 (N_48018,N_32743,N_38868);
nand U48019 (N_48019,N_32000,N_34267);
and U48020 (N_48020,N_37535,N_36435);
xnor U48021 (N_48021,N_36139,N_39557);
and U48022 (N_48022,N_33046,N_35665);
nor U48023 (N_48023,N_34024,N_31355);
xor U48024 (N_48024,N_31013,N_34313);
nand U48025 (N_48025,N_34987,N_37697);
nand U48026 (N_48026,N_34000,N_38061);
nand U48027 (N_48027,N_35427,N_34113);
and U48028 (N_48028,N_32935,N_34036);
nor U48029 (N_48029,N_30121,N_35192);
nand U48030 (N_48030,N_36604,N_31739);
nor U48031 (N_48031,N_30989,N_35826);
nor U48032 (N_48032,N_38828,N_38784);
nand U48033 (N_48033,N_33970,N_38386);
and U48034 (N_48034,N_33351,N_31328);
and U48035 (N_48035,N_30905,N_31660);
nand U48036 (N_48036,N_37213,N_35167);
nand U48037 (N_48037,N_36009,N_38890);
and U48038 (N_48038,N_33296,N_38331);
or U48039 (N_48039,N_33089,N_33712);
nand U48040 (N_48040,N_34103,N_31722);
nor U48041 (N_48041,N_39191,N_37272);
or U48042 (N_48042,N_38997,N_30970);
or U48043 (N_48043,N_34249,N_32600);
and U48044 (N_48044,N_30243,N_32188);
or U48045 (N_48045,N_34989,N_30794);
nand U48046 (N_48046,N_31379,N_33873);
or U48047 (N_48047,N_33855,N_37751);
or U48048 (N_48048,N_36587,N_36494);
or U48049 (N_48049,N_34060,N_32424);
nor U48050 (N_48050,N_37746,N_34475);
or U48051 (N_48051,N_34913,N_32318);
xor U48052 (N_48052,N_33099,N_36451);
and U48053 (N_48053,N_30916,N_31866);
and U48054 (N_48054,N_33036,N_39528);
nand U48055 (N_48055,N_32170,N_39786);
or U48056 (N_48056,N_38464,N_34552);
and U48057 (N_48057,N_36429,N_37800);
and U48058 (N_48058,N_39726,N_33284);
nor U48059 (N_48059,N_36574,N_35713);
nand U48060 (N_48060,N_34781,N_34058);
nand U48061 (N_48061,N_39466,N_31064);
or U48062 (N_48062,N_32851,N_30441);
nand U48063 (N_48063,N_34818,N_33733);
or U48064 (N_48064,N_30483,N_35568);
xor U48065 (N_48065,N_35176,N_34433);
or U48066 (N_48066,N_32453,N_33949);
nand U48067 (N_48067,N_35957,N_39381);
nor U48068 (N_48068,N_39010,N_35667);
nor U48069 (N_48069,N_32137,N_34254);
nor U48070 (N_48070,N_38400,N_38518);
xor U48071 (N_48071,N_38616,N_35233);
and U48072 (N_48072,N_30865,N_31144);
xor U48073 (N_48073,N_35311,N_32110);
nor U48074 (N_48074,N_36272,N_30335);
or U48075 (N_48075,N_31038,N_32208);
nor U48076 (N_48076,N_39352,N_35952);
or U48077 (N_48077,N_31152,N_35378);
and U48078 (N_48078,N_30041,N_38407);
nor U48079 (N_48079,N_38640,N_37756);
xnor U48080 (N_48080,N_34528,N_36564);
nor U48081 (N_48081,N_34455,N_31561);
nor U48082 (N_48082,N_33127,N_35449);
xor U48083 (N_48083,N_31924,N_33212);
nor U48084 (N_48084,N_37763,N_36416);
nor U48085 (N_48085,N_38866,N_32849);
or U48086 (N_48086,N_31894,N_32702);
and U48087 (N_48087,N_33113,N_39003);
or U48088 (N_48088,N_33288,N_32668);
xnor U48089 (N_48089,N_39278,N_32260);
nor U48090 (N_48090,N_30676,N_30429);
and U48091 (N_48091,N_31911,N_33800);
or U48092 (N_48092,N_34063,N_35408);
nand U48093 (N_48093,N_35359,N_39327);
or U48094 (N_48094,N_37892,N_36354);
nor U48095 (N_48095,N_34096,N_34315);
xnor U48096 (N_48096,N_33757,N_31650);
or U48097 (N_48097,N_30863,N_35050);
nor U48098 (N_48098,N_33323,N_37603);
or U48099 (N_48099,N_35340,N_37850);
or U48100 (N_48100,N_36438,N_39053);
and U48101 (N_48101,N_37174,N_39920);
and U48102 (N_48102,N_34082,N_35792);
nand U48103 (N_48103,N_37780,N_35451);
or U48104 (N_48104,N_31606,N_38905);
or U48105 (N_48105,N_34102,N_32769);
nor U48106 (N_48106,N_32054,N_35619);
or U48107 (N_48107,N_33874,N_39823);
nand U48108 (N_48108,N_33451,N_34305);
nor U48109 (N_48109,N_30804,N_30357);
nand U48110 (N_48110,N_37914,N_30998);
and U48111 (N_48111,N_34617,N_35950);
nor U48112 (N_48112,N_30299,N_36057);
or U48113 (N_48113,N_36847,N_39622);
nor U48114 (N_48114,N_34557,N_36750);
xor U48115 (N_48115,N_36106,N_33688);
nor U48116 (N_48116,N_37279,N_33530);
and U48117 (N_48117,N_30621,N_37278);
and U48118 (N_48118,N_36657,N_31071);
or U48119 (N_48119,N_36425,N_35644);
nand U48120 (N_48120,N_33421,N_37960);
and U48121 (N_48121,N_36303,N_38258);
nor U48122 (N_48122,N_31502,N_32679);
nor U48123 (N_48123,N_33449,N_33226);
nor U48124 (N_48124,N_39208,N_30776);
nand U48125 (N_48125,N_33211,N_34505);
xnor U48126 (N_48126,N_38119,N_34591);
and U48127 (N_48127,N_31188,N_36665);
nor U48128 (N_48128,N_33333,N_34755);
nand U48129 (N_48129,N_37383,N_37003);
or U48130 (N_48130,N_38499,N_31290);
nor U48131 (N_48131,N_30279,N_31179);
and U48132 (N_48132,N_34422,N_34606);
and U48133 (N_48133,N_32715,N_32746);
and U48134 (N_48134,N_37149,N_31234);
or U48135 (N_48135,N_33933,N_37791);
nand U48136 (N_48136,N_37741,N_37366);
nand U48137 (N_48137,N_33231,N_38514);
and U48138 (N_48138,N_31562,N_31898);
nor U48139 (N_48139,N_38649,N_30737);
or U48140 (N_48140,N_31472,N_31466);
nor U48141 (N_48141,N_36398,N_30067);
nand U48142 (N_48142,N_35734,N_35745);
and U48143 (N_48143,N_39690,N_34097);
nor U48144 (N_48144,N_38191,N_30732);
or U48145 (N_48145,N_36154,N_34920);
or U48146 (N_48146,N_39853,N_38763);
or U48147 (N_48147,N_37520,N_39720);
and U48148 (N_48148,N_31267,N_39708);
nand U48149 (N_48149,N_36989,N_33224);
nand U48150 (N_48150,N_34613,N_34762);
nor U48151 (N_48151,N_37679,N_30436);
nand U48152 (N_48152,N_36347,N_35549);
nand U48153 (N_48153,N_39605,N_30134);
nand U48154 (N_48154,N_34584,N_34718);
nor U48155 (N_48155,N_33535,N_36972);
nand U48156 (N_48156,N_36407,N_32112);
nand U48157 (N_48157,N_33400,N_38174);
or U48158 (N_48158,N_31213,N_30481);
nand U48159 (N_48159,N_30882,N_31915);
nand U48160 (N_48160,N_35465,N_38401);
nor U48161 (N_48161,N_30330,N_37946);
or U48162 (N_48162,N_37920,N_38381);
nor U48163 (N_48163,N_39174,N_31093);
or U48164 (N_48164,N_39734,N_33433);
nor U48165 (N_48165,N_34618,N_37006);
nor U48166 (N_48166,N_33730,N_35147);
and U48167 (N_48167,N_31098,N_34188);
nor U48168 (N_48168,N_34807,N_37585);
nand U48169 (N_48169,N_31782,N_36951);
nand U48170 (N_48170,N_36914,N_35295);
xor U48171 (N_48171,N_30491,N_31240);
nand U48172 (N_48172,N_39109,N_39133);
and U48173 (N_48173,N_38474,N_31370);
nand U48174 (N_48174,N_34131,N_39011);
and U48175 (N_48175,N_38740,N_39503);
and U48176 (N_48176,N_32633,N_36629);
or U48177 (N_48177,N_32528,N_38521);
and U48178 (N_48178,N_30084,N_37129);
or U48179 (N_48179,N_36258,N_35822);
nand U48180 (N_48180,N_36782,N_37546);
or U48181 (N_48181,N_36268,N_37073);
and U48182 (N_48182,N_32687,N_38523);
nor U48183 (N_48183,N_34375,N_36676);
nand U48184 (N_48184,N_35862,N_31168);
nand U48185 (N_48185,N_34082,N_38013);
or U48186 (N_48186,N_32343,N_39519);
or U48187 (N_48187,N_38251,N_39392);
nand U48188 (N_48188,N_31325,N_38796);
nand U48189 (N_48189,N_33565,N_36634);
nand U48190 (N_48190,N_39920,N_34580);
nor U48191 (N_48191,N_38083,N_33792);
xor U48192 (N_48192,N_35792,N_30918);
and U48193 (N_48193,N_32752,N_33380);
and U48194 (N_48194,N_38149,N_35922);
nand U48195 (N_48195,N_33721,N_38122);
nand U48196 (N_48196,N_35669,N_37626);
or U48197 (N_48197,N_36346,N_33848);
nand U48198 (N_48198,N_36047,N_33699);
and U48199 (N_48199,N_31340,N_34276);
xor U48200 (N_48200,N_39205,N_32868);
nor U48201 (N_48201,N_32636,N_31650);
xnor U48202 (N_48202,N_34261,N_31287);
nor U48203 (N_48203,N_30093,N_32345);
nand U48204 (N_48204,N_36834,N_32615);
nor U48205 (N_48205,N_30149,N_35688);
or U48206 (N_48206,N_35901,N_37076);
nor U48207 (N_48207,N_38946,N_39027);
nor U48208 (N_48208,N_34991,N_39197);
and U48209 (N_48209,N_36886,N_30121);
nand U48210 (N_48210,N_32657,N_30554);
or U48211 (N_48211,N_32842,N_34018);
nand U48212 (N_48212,N_33519,N_39643);
nor U48213 (N_48213,N_35164,N_30830);
nor U48214 (N_48214,N_35151,N_34267);
or U48215 (N_48215,N_37061,N_32631);
or U48216 (N_48216,N_38641,N_32595);
or U48217 (N_48217,N_38389,N_30393);
nand U48218 (N_48218,N_34654,N_37010);
nand U48219 (N_48219,N_38581,N_34328);
nor U48220 (N_48220,N_38722,N_38301);
nand U48221 (N_48221,N_36653,N_35493);
and U48222 (N_48222,N_32176,N_34914);
and U48223 (N_48223,N_34163,N_32777);
or U48224 (N_48224,N_38615,N_38409);
xnor U48225 (N_48225,N_30137,N_39445);
nor U48226 (N_48226,N_38061,N_38762);
nand U48227 (N_48227,N_32457,N_35317);
and U48228 (N_48228,N_37512,N_30714);
or U48229 (N_48229,N_36316,N_36202);
and U48230 (N_48230,N_30721,N_37633);
and U48231 (N_48231,N_30853,N_34675);
and U48232 (N_48232,N_39201,N_32367);
or U48233 (N_48233,N_38908,N_36433);
and U48234 (N_48234,N_32180,N_35094);
xnor U48235 (N_48235,N_30400,N_37693);
or U48236 (N_48236,N_35856,N_37693);
nor U48237 (N_48237,N_38582,N_35937);
xnor U48238 (N_48238,N_33431,N_32395);
or U48239 (N_48239,N_31052,N_34719);
nor U48240 (N_48240,N_34237,N_34477);
nor U48241 (N_48241,N_30981,N_38694);
nand U48242 (N_48242,N_35714,N_36813);
and U48243 (N_48243,N_33349,N_37599);
nor U48244 (N_48244,N_31660,N_35911);
or U48245 (N_48245,N_31127,N_33510);
nor U48246 (N_48246,N_31788,N_30988);
xor U48247 (N_48247,N_31779,N_35401);
or U48248 (N_48248,N_35990,N_36653);
and U48249 (N_48249,N_31183,N_36615);
or U48250 (N_48250,N_30938,N_36854);
nand U48251 (N_48251,N_30607,N_32255);
nor U48252 (N_48252,N_31195,N_33397);
or U48253 (N_48253,N_37941,N_30278);
and U48254 (N_48254,N_37020,N_36657);
nor U48255 (N_48255,N_35189,N_34105);
nor U48256 (N_48256,N_35203,N_33580);
and U48257 (N_48257,N_31883,N_33926);
nand U48258 (N_48258,N_30038,N_39622);
nand U48259 (N_48259,N_37195,N_36644);
and U48260 (N_48260,N_36257,N_36163);
nor U48261 (N_48261,N_39867,N_37084);
or U48262 (N_48262,N_38157,N_31050);
nand U48263 (N_48263,N_31420,N_39251);
or U48264 (N_48264,N_39610,N_37014);
or U48265 (N_48265,N_36942,N_38709);
or U48266 (N_48266,N_33728,N_30154);
or U48267 (N_48267,N_31720,N_32150);
and U48268 (N_48268,N_39855,N_38402);
and U48269 (N_48269,N_35506,N_35360);
nand U48270 (N_48270,N_37405,N_35331);
or U48271 (N_48271,N_33500,N_34032);
nand U48272 (N_48272,N_39584,N_37277);
nand U48273 (N_48273,N_35865,N_34983);
or U48274 (N_48274,N_35922,N_30637);
xor U48275 (N_48275,N_35367,N_33044);
or U48276 (N_48276,N_39775,N_37314);
and U48277 (N_48277,N_37039,N_32511);
or U48278 (N_48278,N_34083,N_30225);
or U48279 (N_48279,N_33915,N_31831);
and U48280 (N_48280,N_39283,N_39469);
or U48281 (N_48281,N_38404,N_36836);
or U48282 (N_48282,N_35393,N_37998);
nand U48283 (N_48283,N_32956,N_36349);
nor U48284 (N_48284,N_35423,N_38575);
nor U48285 (N_48285,N_33412,N_34713);
nand U48286 (N_48286,N_39085,N_36218);
nor U48287 (N_48287,N_33382,N_30544);
and U48288 (N_48288,N_31052,N_30939);
nor U48289 (N_48289,N_38272,N_37389);
or U48290 (N_48290,N_31199,N_32275);
and U48291 (N_48291,N_37942,N_35078);
and U48292 (N_48292,N_34860,N_39715);
nand U48293 (N_48293,N_31588,N_37741);
and U48294 (N_48294,N_39704,N_38249);
nor U48295 (N_48295,N_39710,N_38857);
or U48296 (N_48296,N_30803,N_33398);
or U48297 (N_48297,N_31455,N_31991);
nand U48298 (N_48298,N_35587,N_37199);
nor U48299 (N_48299,N_31790,N_36908);
or U48300 (N_48300,N_34047,N_39463);
nor U48301 (N_48301,N_31344,N_35689);
and U48302 (N_48302,N_35849,N_34094);
nor U48303 (N_48303,N_32299,N_33175);
or U48304 (N_48304,N_33319,N_32643);
and U48305 (N_48305,N_31548,N_38370);
nor U48306 (N_48306,N_30056,N_32087);
or U48307 (N_48307,N_37794,N_33081);
xor U48308 (N_48308,N_36047,N_35124);
nand U48309 (N_48309,N_31961,N_37410);
nand U48310 (N_48310,N_34469,N_34956);
or U48311 (N_48311,N_36613,N_31395);
and U48312 (N_48312,N_33181,N_35185);
nand U48313 (N_48313,N_31633,N_35723);
or U48314 (N_48314,N_35663,N_34480);
nand U48315 (N_48315,N_36907,N_31446);
nor U48316 (N_48316,N_32154,N_35066);
and U48317 (N_48317,N_38167,N_36246);
and U48318 (N_48318,N_30148,N_38722);
nand U48319 (N_48319,N_34674,N_34046);
or U48320 (N_48320,N_30503,N_30398);
nor U48321 (N_48321,N_36397,N_33812);
nand U48322 (N_48322,N_37421,N_33407);
or U48323 (N_48323,N_35368,N_39558);
nand U48324 (N_48324,N_37807,N_34265);
and U48325 (N_48325,N_30119,N_36266);
and U48326 (N_48326,N_30545,N_34310);
or U48327 (N_48327,N_30738,N_35747);
nor U48328 (N_48328,N_39891,N_38403);
or U48329 (N_48329,N_37065,N_36590);
and U48330 (N_48330,N_33395,N_38516);
nor U48331 (N_48331,N_30333,N_30758);
nand U48332 (N_48332,N_30812,N_34398);
and U48333 (N_48333,N_35122,N_38163);
nand U48334 (N_48334,N_36319,N_32940);
nor U48335 (N_48335,N_38714,N_32665);
and U48336 (N_48336,N_34958,N_30246);
or U48337 (N_48337,N_33663,N_32940);
nand U48338 (N_48338,N_37144,N_39581);
or U48339 (N_48339,N_38013,N_33229);
nor U48340 (N_48340,N_35591,N_38343);
xnor U48341 (N_48341,N_33536,N_37003);
nand U48342 (N_48342,N_37170,N_34680);
or U48343 (N_48343,N_33580,N_39381);
or U48344 (N_48344,N_38924,N_34705);
nand U48345 (N_48345,N_36586,N_31383);
nand U48346 (N_48346,N_31710,N_33140);
or U48347 (N_48347,N_34805,N_34295);
and U48348 (N_48348,N_30608,N_31768);
and U48349 (N_48349,N_35374,N_38704);
nand U48350 (N_48350,N_32897,N_38622);
nor U48351 (N_48351,N_31798,N_34679);
nand U48352 (N_48352,N_37365,N_37389);
or U48353 (N_48353,N_32947,N_35903);
nand U48354 (N_48354,N_34515,N_35290);
nand U48355 (N_48355,N_37879,N_35807);
nor U48356 (N_48356,N_39739,N_35642);
or U48357 (N_48357,N_32269,N_30273);
nand U48358 (N_48358,N_34754,N_31245);
xor U48359 (N_48359,N_31866,N_34769);
and U48360 (N_48360,N_36330,N_34963);
nand U48361 (N_48361,N_37070,N_33120);
and U48362 (N_48362,N_36430,N_32749);
and U48363 (N_48363,N_35092,N_34608);
or U48364 (N_48364,N_31567,N_30322);
and U48365 (N_48365,N_34685,N_36732);
xnor U48366 (N_48366,N_36625,N_37749);
nand U48367 (N_48367,N_36168,N_32316);
xnor U48368 (N_48368,N_38290,N_37783);
nor U48369 (N_48369,N_34270,N_35315);
and U48370 (N_48370,N_30417,N_37081);
nor U48371 (N_48371,N_38586,N_34949);
nor U48372 (N_48372,N_37105,N_33049);
nand U48373 (N_48373,N_35594,N_30096);
nor U48374 (N_48374,N_34530,N_34342);
nand U48375 (N_48375,N_35490,N_38855);
or U48376 (N_48376,N_33861,N_38294);
nand U48377 (N_48377,N_30620,N_38919);
or U48378 (N_48378,N_38525,N_35639);
nand U48379 (N_48379,N_36872,N_34180);
nand U48380 (N_48380,N_32319,N_37631);
or U48381 (N_48381,N_30190,N_38042);
or U48382 (N_48382,N_39470,N_39965);
nand U48383 (N_48383,N_31320,N_32391);
and U48384 (N_48384,N_35260,N_33854);
and U48385 (N_48385,N_39158,N_32314);
nand U48386 (N_48386,N_37503,N_32502);
or U48387 (N_48387,N_37189,N_37250);
nand U48388 (N_48388,N_36542,N_33062);
nand U48389 (N_48389,N_36517,N_37563);
or U48390 (N_48390,N_33537,N_34752);
nand U48391 (N_48391,N_35334,N_35649);
nor U48392 (N_48392,N_38886,N_38985);
nor U48393 (N_48393,N_30815,N_35441);
nand U48394 (N_48394,N_39091,N_37901);
and U48395 (N_48395,N_37341,N_39821);
and U48396 (N_48396,N_36982,N_37688);
and U48397 (N_48397,N_36767,N_30425);
and U48398 (N_48398,N_36991,N_39927);
or U48399 (N_48399,N_35119,N_39309);
nand U48400 (N_48400,N_30819,N_35507);
nand U48401 (N_48401,N_33742,N_35403);
nor U48402 (N_48402,N_31339,N_30421);
and U48403 (N_48403,N_32637,N_30548);
nor U48404 (N_48404,N_35497,N_30456);
or U48405 (N_48405,N_31056,N_34211);
xor U48406 (N_48406,N_33797,N_33277);
and U48407 (N_48407,N_38412,N_37537);
xor U48408 (N_48408,N_36463,N_32397);
nand U48409 (N_48409,N_36165,N_32024);
nand U48410 (N_48410,N_33907,N_35447);
nor U48411 (N_48411,N_37748,N_39571);
and U48412 (N_48412,N_35698,N_39972);
xnor U48413 (N_48413,N_39035,N_31418);
or U48414 (N_48414,N_35274,N_38169);
or U48415 (N_48415,N_34183,N_37227);
nand U48416 (N_48416,N_34500,N_35460);
nor U48417 (N_48417,N_35500,N_38242);
nor U48418 (N_48418,N_33840,N_31477);
nor U48419 (N_48419,N_39097,N_36247);
xor U48420 (N_48420,N_38581,N_33145);
or U48421 (N_48421,N_30702,N_31669);
nor U48422 (N_48422,N_31245,N_34359);
nor U48423 (N_48423,N_36741,N_32221);
and U48424 (N_48424,N_35111,N_37446);
nand U48425 (N_48425,N_36194,N_35739);
nand U48426 (N_48426,N_32126,N_38483);
nand U48427 (N_48427,N_38460,N_30138);
and U48428 (N_48428,N_31893,N_35087);
nand U48429 (N_48429,N_30366,N_36783);
or U48430 (N_48430,N_31695,N_34310);
xor U48431 (N_48431,N_36236,N_33144);
nor U48432 (N_48432,N_31686,N_33143);
or U48433 (N_48433,N_31573,N_32149);
or U48434 (N_48434,N_30283,N_31224);
or U48435 (N_48435,N_33221,N_39161);
or U48436 (N_48436,N_32358,N_38963);
nand U48437 (N_48437,N_38729,N_32503);
or U48438 (N_48438,N_32611,N_30832);
or U48439 (N_48439,N_33153,N_33739);
and U48440 (N_48440,N_39122,N_31735);
nor U48441 (N_48441,N_38767,N_30330);
nor U48442 (N_48442,N_34093,N_38526);
and U48443 (N_48443,N_30235,N_31482);
or U48444 (N_48444,N_30626,N_36913);
or U48445 (N_48445,N_32308,N_33333);
nand U48446 (N_48446,N_34466,N_37522);
nand U48447 (N_48447,N_33210,N_34939);
xor U48448 (N_48448,N_37348,N_33074);
or U48449 (N_48449,N_33318,N_36459);
nand U48450 (N_48450,N_36790,N_38417);
nor U48451 (N_48451,N_33172,N_33167);
nor U48452 (N_48452,N_31572,N_39385);
nand U48453 (N_48453,N_34503,N_31138);
nand U48454 (N_48454,N_37664,N_37332);
and U48455 (N_48455,N_38354,N_33071);
nor U48456 (N_48456,N_38988,N_34602);
nand U48457 (N_48457,N_35611,N_35865);
nand U48458 (N_48458,N_31720,N_30531);
nand U48459 (N_48459,N_39800,N_34415);
and U48460 (N_48460,N_37690,N_30822);
xnor U48461 (N_48461,N_34919,N_30842);
nand U48462 (N_48462,N_34416,N_38700);
nand U48463 (N_48463,N_37765,N_31702);
nand U48464 (N_48464,N_36605,N_32530);
xnor U48465 (N_48465,N_39280,N_33440);
nand U48466 (N_48466,N_32047,N_33661);
nand U48467 (N_48467,N_38364,N_36904);
nand U48468 (N_48468,N_38540,N_38776);
nand U48469 (N_48469,N_32824,N_39817);
nand U48470 (N_48470,N_30924,N_37764);
or U48471 (N_48471,N_39165,N_34523);
nor U48472 (N_48472,N_39636,N_35732);
xor U48473 (N_48473,N_30844,N_31459);
nor U48474 (N_48474,N_35103,N_32295);
nand U48475 (N_48475,N_30976,N_35802);
and U48476 (N_48476,N_33719,N_32831);
and U48477 (N_48477,N_37840,N_35519);
nor U48478 (N_48478,N_31149,N_39723);
or U48479 (N_48479,N_37833,N_35426);
xnor U48480 (N_48480,N_35249,N_31819);
xnor U48481 (N_48481,N_37174,N_36319);
xnor U48482 (N_48482,N_38044,N_38384);
or U48483 (N_48483,N_31339,N_37609);
nand U48484 (N_48484,N_35353,N_33665);
or U48485 (N_48485,N_37344,N_39786);
nand U48486 (N_48486,N_38800,N_31203);
nand U48487 (N_48487,N_34296,N_33078);
nand U48488 (N_48488,N_36776,N_39440);
nor U48489 (N_48489,N_32181,N_37354);
and U48490 (N_48490,N_39090,N_31895);
nor U48491 (N_48491,N_39807,N_39268);
nand U48492 (N_48492,N_38198,N_35457);
and U48493 (N_48493,N_32036,N_34084);
nor U48494 (N_48494,N_32710,N_36833);
xnor U48495 (N_48495,N_31141,N_39379);
nand U48496 (N_48496,N_32888,N_35586);
nor U48497 (N_48497,N_36266,N_33309);
or U48498 (N_48498,N_38378,N_32138);
and U48499 (N_48499,N_30485,N_31843);
or U48500 (N_48500,N_36526,N_37471);
or U48501 (N_48501,N_39760,N_39454);
and U48502 (N_48502,N_38001,N_34199);
or U48503 (N_48503,N_30975,N_34937);
nand U48504 (N_48504,N_33678,N_34484);
nor U48505 (N_48505,N_39015,N_30323);
and U48506 (N_48506,N_30285,N_34841);
or U48507 (N_48507,N_32214,N_39358);
and U48508 (N_48508,N_32965,N_33680);
nand U48509 (N_48509,N_38077,N_30793);
nor U48510 (N_48510,N_31987,N_30378);
or U48511 (N_48511,N_36891,N_34247);
nand U48512 (N_48512,N_30710,N_31479);
nor U48513 (N_48513,N_36763,N_37463);
and U48514 (N_48514,N_39623,N_30085);
nor U48515 (N_48515,N_39402,N_35058);
and U48516 (N_48516,N_39455,N_38214);
and U48517 (N_48517,N_36921,N_37224);
xnor U48518 (N_48518,N_32955,N_30870);
nand U48519 (N_48519,N_30054,N_35211);
and U48520 (N_48520,N_31912,N_35521);
nor U48521 (N_48521,N_31936,N_31409);
xnor U48522 (N_48522,N_33050,N_38586);
nor U48523 (N_48523,N_31771,N_37967);
nand U48524 (N_48524,N_39377,N_39709);
or U48525 (N_48525,N_39105,N_31436);
nor U48526 (N_48526,N_36096,N_34559);
xor U48527 (N_48527,N_37425,N_39973);
nor U48528 (N_48528,N_31256,N_37255);
nand U48529 (N_48529,N_38010,N_37575);
or U48530 (N_48530,N_39799,N_38887);
and U48531 (N_48531,N_32359,N_31741);
or U48532 (N_48532,N_31912,N_36052);
or U48533 (N_48533,N_31991,N_35098);
or U48534 (N_48534,N_39495,N_36072);
nor U48535 (N_48535,N_37201,N_39313);
xnor U48536 (N_48536,N_32535,N_38892);
and U48537 (N_48537,N_33172,N_32251);
or U48538 (N_48538,N_33142,N_38163);
or U48539 (N_48539,N_35246,N_38584);
and U48540 (N_48540,N_38023,N_34622);
and U48541 (N_48541,N_31451,N_38181);
and U48542 (N_48542,N_38861,N_32872);
nand U48543 (N_48543,N_31290,N_38301);
nand U48544 (N_48544,N_36578,N_33700);
and U48545 (N_48545,N_36754,N_33534);
nand U48546 (N_48546,N_33974,N_37785);
and U48547 (N_48547,N_30497,N_37445);
and U48548 (N_48548,N_37488,N_37262);
nand U48549 (N_48549,N_36932,N_39428);
and U48550 (N_48550,N_38205,N_33193);
nor U48551 (N_48551,N_36382,N_32884);
nand U48552 (N_48552,N_38407,N_37591);
nor U48553 (N_48553,N_39301,N_30183);
xnor U48554 (N_48554,N_33928,N_36716);
or U48555 (N_48555,N_34494,N_34591);
nand U48556 (N_48556,N_39845,N_39114);
nor U48557 (N_48557,N_39997,N_35100);
nor U48558 (N_48558,N_33496,N_36069);
nor U48559 (N_48559,N_37296,N_32088);
nand U48560 (N_48560,N_38789,N_36918);
or U48561 (N_48561,N_33624,N_31765);
xor U48562 (N_48562,N_35707,N_38352);
nand U48563 (N_48563,N_34269,N_32046);
or U48564 (N_48564,N_39579,N_30489);
or U48565 (N_48565,N_33502,N_33346);
nand U48566 (N_48566,N_35426,N_39070);
nor U48567 (N_48567,N_37121,N_39997);
or U48568 (N_48568,N_35147,N_32419);
xnor U48569 (N_48569,N_39330,N_34462);
and U48570 (N_48570,N_38184,N_30216);
or U48571 (N_48571,N_37801,N_35525);
nor U48572 (N_48572,N_37041,N_38094);
xor U48573 (N_48573,N_35199,N_32300);
or U48574 (N_48574,N_34890,N_39718);
nor U48575 (N_48575,N_30798,N_34766);
nand U48576 (N_48576,N_35750,N_30514);
and U48577 (N_48577,N_38809,N_35016);
nor U48578 (N_48578,N_38233,N_35993);
nor U48579 (N_48579,N_30214,N_34539);
or U48580 (N_48580,N_31290,N_30065);
nand U48581 (N_48581,N_32288,N_30285);
or U48582 (N_48582,N_34532,N_35566);
and U48583 (N_48583,N_39321,N_30363);
nand U48584 (N_48584,N_36582,N_33024);
xnor U48585 (N_48585,N_30382,N_34953);
and U48586 (N_48586,N_37552,N_34945);
or U48587 (N_48587,N_35489,N_35062);
nand U48588 (N_48588,N_39561,N_30425);
nor U48589 (N_48589,N_38064,N_35751);
and U48590 (N_48590,N_31072,N_31086);
nor U48591 (N_48591,N_35718,N_30380);
xor U48592 (N_48592,N_30354,N_30356);
nand U48593 (N_48593,N_32807,N_35084);
and U48594 (N_48594,N_31275,N_31116);
or U48595 (N_48595,N_32378,N_31925);
nor U48596 (N_48596,N_36868,N_37992);
nand U48597 (N_48597,N_34662,N_30060);
or U48598 (N_48598,N_33340,N_34098);
or U48599 (N_48599,N_31893,N_30358);
nand U48600 (N_48600,N_36576,N_35748);
xnor U48601 (N_48601,N_30922,N_37318);
or U48602 (N_48602,N_39929,N_35510);
or U48603 (N_48603,N_36207,N_33161);
nor U48604 (N_48604,N_33584,N_39425);
xnor U48605 (N_48605,N_34255,N_34557);
and U48606 (N_48606,N_39478,N_31750);
or U48607 (N_48607,N_35821,N_31659);
or U48608 (N_48608,N_30186,N_38274);
nor U48609 (N_48609,N_39040,N_35636);
nor U48610 (N_48610,N_38952,N_37797);
and U48611 (N_48611,N_37807,N_33415);
nand U48612 (N_48612,N_31536,N_30608);
nor U48613 (N_48613,N_32588,N_33595);
nand U48614 (N_48614,N_37593,N_34899);
or U48615 (N_48615,N_32880,N_37540);
nand U48616 (N_48616,N_35707,N_38176);
xor U48617 (N_48617,N_33726,N_31245);
nand U48618 (N_48618,N_35357,N_30375);
and U48619 (N_48619,N_32193,N_36005);
nor U48620 (N_48620,N_31039,N_38055);
nor U48621 (N_48621,N_33057,N_39760);
and U48622 (N_48622,N_34101,N_35383);
nand U48623 (N_48623,N_34932,N_36675);
nor U48624 (N_48624,N_31429,N_34671);
or U48625 (N_48625,N_32879,N_34589);
nand U48626 (N_48626,N_34166,N_30316);
nand U48627 (N_48627,N_36149,N_38738);
and U48628 (N_48628,N_34406,N_34150);
nor U48629 (N_48629,N_36443,N_31090);
and U48630 (N_48630,N_30535,N_31494);
nand U48631 (N_48631,N_39868,N_34652);
xor U48632 (N_48632,N_36228,N_30272);
and U48633 (N_48633,N_34801,N_36881);
or U48634 (N_48634,N_34950,N_36325);
and U48635 (N_48635,N_38085,N_32624);
and U48636 (N_48636,N_32384,N_35079);
xor U48637 (N_48637,N_32954,N_34618);
xnor U48638 (N_48638,N_39881,N_38059);
nand U48639 (N_48639,N_31978,N_35731);
nand U48640 (N_48640,N_37576,N_39990);
nor U48641 (N_48641,N_34548,N_35373);
nor U48642 (N_48642,N_37439,N_32247);
xnor U48643 (N_48643,N_33676,N_30201);
or U48644 (N_48644,N_32147,N_31710);
or U48645 (N_48645,N_34600,N_31338);
or U48646 (N_48646,N_33705,N_35424);
nand U48647 (N_48647,N_35801,N_32090);
xor U48648 (N_48648,N_39910,N_32535);
or U48649 (N_48649,N_34667,N_37751);
and U48650 (N_48650,N_31662,N_35720);
or U48651 (N_48651,N_34161,N_36258);
nor U48652 (N_48652,N_38436,N_39354);
nor U48653 (N_48653,N_36499,N_33273);
xor U48654 (N_48654,N_33326,N_35216);
or U48655 (N_48655,N_35285,N_39876);
and U48656 (N_48656,N_38005,N_31802);
or U48657 (N_48657,N_39942,N_36844);
xor U48658 (N_48658,N_36757,N_32860);
nand U48659 (N_48659,N_36913,N_34150);
or U48660 (N_48660,N_34290,N_34819);
or U48661 (N_48661,N_34369,N_39729);
and U48662 (N_48662,N_30991,N_35630);
or U48663 (N_48663,N_30261,N_37528);
and U48664 (N_48664,N_39762,N_32875);
and U48665 (N_48665,N_33490,N_36076);
nor U48666 (N_48666,N_37988,N_31256);
and U48667 (N_48667,N_33988,N_32217);
or U48668 (N_48668,N_38373,N_34742);
nand U48669 (N_48669,N_35270,N_35622);
and U48670 (N_48670,N_37779,N_36059);
nor U48671 (N_48671,N_38164,N_35546);
or U48672 (N_48672,N_39277,N_35205);
and U48673 (N_48673,N_35430,N_32243);
and U48674 (N_48674,N_36666,N_34303);
nor U48675 (N_48675,N_36542,N_38135);
and U48676 (N_48676,N_33712,N_39503);
nand U48677 (N_48677,N_32919,N_32219);
nor U48678 (N_48678,N_30129,N_37616);
or U48679 (N_48679,N_38392,N_38391);
nand U48680 (N_48680,N_32740,N_35513);
xnor U48681 (N_48681,N_34216,N_39369);
nand U48682 (N_48682,N_38378,N_36210);
nand U48683 (N_48683,N_39389,N_31247);
nand U48684 (N_48684,N_31220,N_31031);
xnor U48685 (N_48685,N_36257,N_38619);
or U48686 (N_48686,N_39835,N_39598);
or U48687 (N_48687,N_37230,N_30362);
and U48688 (N_48688,N_30420,N_34809);
nor U48689 (N_48689,N_36895,N_33028);
and U48690 (N_48690,N_31730,N_39914);
nor U48691 (N_48691,N_38182,N_34897);
nand U48692 (N_48692,N_39191,N_37649);
nand U48693 (N_48693,N_36448,N_33510);
and U48694 (N_48694,N_30499,N_37768);
and U48695 (N_48695,N_37621,N_39546);
or U48696 (N_48696,N_31197,N_36175);
nor U48697 (N_48697,N_31401,N_35567);
and U48698 (N_48698,N_37892,N_38724);
nor U48699 (N_48699,N_35293,N_35284);
xnor U48700 (N_48700,N_34467,N_31350);
or U48701 (N_48701,N_36637,N_33631);
nor U48702 (N_48702,N_34053,N_39025);
nor U48703 (N_48703,N_31572,N_32892);
xor U48704 (N_48704,N_31118,N_33063);
or U48705 (N_48705,N_32691,N_37088);
and U48706 (N_48706,N_31228,N_36458);
xnor U48707 (N_48707,N_33520,N_35644);
and U48708 (N_48708,N_38428,N_35148);
nand U48709 (N_48709,N_32671,N_34859);
xnor U48710 (N_48710,N_31862,N_39370);
nor U48711 (N_48711,N_35793,N_38021);
nor U48712 (N_48712,N_35052,N_33279);
and U48713 (N_48713,N_31828,N_36359);
nor U48714 (N_48714,N_35865,N_31338);
nand U48715 (N_48715,N_34014,N_33123);
and U48716 (N_48716,N_36597,N_37719);
or U48717 (N_48717,N_30545,N_34182);
nor U48718 (N_48718,N_35361,N_39461);
or U48719 (N_48719,N_34497,N_39908);
and U48720 (N_48720,N_36179,N_35876);
nor U48721 (N_48721,N_31602,N_30897);
nand U48722 (N_48722,N_34036,N_39257);
nand U48723 (N_48723,N_36003,N_32445);
nor U48724 (N_48724,N_34715,N_38206);
nor U48725 (N_48725,N_31666,N_36091);
nor U48726 (N_48726,N_34611,N_33063);
nor U48727 (N_48727,N_31833,N_31773);
or U48728 (N_48728,N_37336,N_33418);
nor U48729 (N_48729,N_30946,N_39094);
or U48730 (N_48730,N_38272,N_33456);
and U48731 (N_48731,N_37321,N_35917);
nor U48732 (N_48732,N_31766,N_30888);
nor U48733 (N_48733,N_36316,N_34798);
nor U48734 (N_48734,N_37660,N_30919);
or U48735 (N_48735,N_30745,N_39031);
or U48736 (N_48736,N_33147,N_39322);
nand U48737 (N_48737,N_32148,N_35389);
or U48738 (N_48738,N_39074,N_38518);
nand U48739 (N_48739,N_37020,N_36194);
or U48740 (N_48740,N_39734,N_33657);
or U48741 (N_48741,N_34234,N_34506);
and U48742 (N_48742,N_33316,N_31253);
nand U48743 (N_48743,N_34681,N_34112);
or U48744 (N_48744,N_38354,N_39648);
nor U48745 (N_48745,N_37510,N_34376);
xnor U48746 (N_48746,N_33483,N_34131);
and U48747 (N_48747,N_36439,N_36274);
xor U48748 (N_48748,N_32111,N_38738);
and U48749 (N_48749,N_36476,N_30505);
nor U48750 (N_48750,N_36503,N_36110);
nor U48751 (N_48751,N_35489,N_37024);
nand U48752 (N_48752,N_33323,N_31759);
nand U48753 (N_48753,N_39021,N_34158);
or U48754 (N_48754,N_36555,N_35306);
and U48755 (N_48755,N_31370,N_30025);
nand U48756 (N_48756,N_30089,N_39437);
nand U48757 (N_48757,N_30757,N_31692);
and U48758 (N_48758,N_33560,N_37690);
or U48759 (N_48759,N_37079,N_38042);
xor U48760 (N_48760,N_34427,N_30300);
xnor U48761 (N_48761,N_30488,N_31257);
or U48762 (N_48762,N_39192,N_33403);
nor U48763 (N_48763,N_38580,N_33271);
nand U48764 (N_48764,N_35039,N_31028);
and U48765 (N_48765,N_35877,N_37266);
nor U48766 (N_48766,N_37467,N_36397);
xor U48767 (N_48767,N_32798,N_32660);
nor U48768 (N_48768,N_36473,N_32992);
xnor U48769 (N_48769,N_39439,N_36321);
and U48770 (N_48770,N_38137,N_36989);
or U48771 (N_48771,N_36507,N_34439);
and U48772 (N_48772,N_34340,N_39988);
and U48773 (N_48773,N_31307,N_39422);
or U48774 (N_48774,N_32303,N_37774);
nor U48775 (N_48775,N_36843,N_38537);
xor U48776 (N_48776,N_30146,N_32128);
nand U48777 (N_48777,N_37476,N_30365);
or U48778 (N_48778,N_39484,N_37868);
nor U48779 (N_48779,N_34703,N_33422);
or U48780 (N_48780,N_39909,N_37006);
nand U48781 (N_48781,N_39335,N_34903);
and U48782 (N_48782,N_33726,N_31487);
xnor U48783 (N_48783,N_37247,N_35668);
nand U48784 (N_48784,N_38529,N_34978);
and U48785 (N_48785,N_34632,N_32844);
nor U48786 (N_48786,N_38742,N_32660);
nand U48787 (N_48787,N_30572,N_36163);
xor U48788 (N_48788,N_37429,N_38425);
or U48789 (N_48789,N_33913,N_34675);
nor U48790 (N_48790,N_39952,N_33894);
and U48791 (N_48791,N_36265,N_33589);
or U48792 (N_48792,N_39256,N_32439);
nor U48793 (N_48793,N_33247,N_35039);
or U48794 (N_48794,N_32329,N_37889);
and U48795 (N_48795,N_31791,N_39437);
nand U48796 (N_48796,N_39716,N_37222);
nor U48797 (N_48797,N_35385,N_39564);
xnor U48798 (N_48798,N_34500,N_35484);
nor U48799 (N_48799,N_36235,N_32498);
nand U48800 (N_48800,N_34425,N_31546);
xnor U48801 (N_48801,N_39411,N_30103);
nor U48802 (N_48802,N_30952,N_36918);
nand U48803 (N_48803,N_35732,N_33566);
nand U48804 (N_48804,N_34549,N_34257);
nor U48805 (N_48805,N_34655,N_33762);
or U48806 (N_48806,N_35757,N_36272);
nor U48807 (N_48807,N_31571,N_39623);
nor U48808 (N_48808,N_31144,N_32434);
nand U48809 (N_48809,N_36702,N_31690);
nor U48810 (N_48810,N_36071,N_33534);
nor U48811 (N_48811,N_31194,N_35850);
nand U48812 (N_48812,N_31489,N_34952);
or U48813 (N_48813,N_32281,N_31314);
and U48814 (N_48814,N_30388,N_34786);
or U48815 (N_48815,N_34515,N_34450);
nor U48816 (N_48816,N_36438,N_33805);
and U48817 (N_48817,N_34356,N_30546);
and U48818 (N_48818,N_36059,N_36879);
or U48819 (N_48819,N_37830,N_35363);
nand U48820 (N_48820,N_33816,N_33721);
and U48821 (N_48821,N_32946,N_31807);
nor U48822 (N_48822,N_33952,N_35947);
nand U48823 (N_48823,N_37564,N_30557);
nor U48824 (N_48824,N_33200,N_32521);
xnor U48825 (N_48825,N_31633,N_36364);
or U48826 (N_48826,N_30800,N_32866);
or U48827 (N_48827,N_33933,N_36390);
nand U48828 (N_48828,N_34900,N_30343);
nand U48829 (N_48829,N_34519,N_36118);
nor U48830 (N_48830,N_38406,N_37056);
nor U48831 (N_48831,N_31475,N_33392);
or U48832 (N_48832,N_38290,N_35077);
or U48833 (N_48833,N_30618,N_34096);
nand U48834 (N_48834,N_30516,N_36519);
or U48835 (N_48835,N_31128,N_37416);
or U48836 (N_48836,N_35715,N_33543);
and U48837 (N_48837,N_30291,N_38553);
or U48838 (N_48838,N_35143,N_31925);
xor U48839 (N_48839,N_39880,N_32121);
and U48840 (N_48840,N_31309,N_34324);
nor U48841 (N_48841,N_37428,N_38531);
nor U48842 (N_48842,N_39549,N_30366);
and U48843 (N_48843,N_30519,N_38767);
nand U48844 (N_48844,N_34074,N_36092);
or U48845 (N_48845,N_35441,N_38004);
nand U48846 (N_48846,N_38373,N_32529);
nor U48847 (N_48847,N_34427,N_37276);
or U48848 (N_48848,N_36845,N_33078);
nor U48849 (N_48849,N_36191,N_34578);
and U48850 (N_48850,N_39686,N_38358);
or U48851 (N_48851,N_37971,N_39417);
or U48852 (N_48852,N_32615,N_32789);
nor U48853 (N_48853,N_35826,N_35348);
nor U48854 (N_48854,N_38808,N_39330);
nor U48855 (N_48855,N_39977,N_32059);
nor U48856 (N_48856,N_30232,N_31122);
or U48857 (N_48857,N_37349,N_39073);
nor U48858 (N_48858,N_34267,N_38257);
xor U48859 (N_48859,N_38057,N_30530);
nor U48860 (N_48860,N_39789,N_31111);
or U48861 (N_48861,N_32041,N_36891);
or U48862 (N_48862,N_34670,N_37732);
and U48863 (N_48863,N_35295,N_30990);
nand U48864 (N_48864,N_39986,N_35369);
nor U48865 (N_48865,N_31429,N_31125);
nand U48866 (N_48866,N_32396,N_33912);
or U48867 (N_48867,N_37496,N_38582);
nor U48868 (N_48868,N_33985,N_32465);
xnor U48869 (N_48869,N_30355,N_36397);
nor U48870 (N_48870,N_36491,N_30219);
or U48871 (N_48871,N_36986,N_32686);
nand U48872 (N_48872,N_35628,N_32360);
xor U48873 (N_48873,N_32139,N_32772);
or U48874 (N_48874,N_36906,N_35724);
nand U48875 (N_48875,N_34325,N_38647);
or U48876 (N_48876,N_30290,N_30568);
nand U48877 (N_48877,N_31548,N_34459);
nand U48878 (N_48878,N_38012,N_36737);
xor U48879 (N_48879,N_36426,N_36946);
and U48880 (N_48880,N_34870,N_36257);
nor U48881 (N_48881,N_38665,N_39666);
nand U48882 (N_48882,N_34706,N_32716);
nor U48883 (N_48883,N_32852,N_33637);
nor U48884 (N_48884,N_37764,N_34160);
nor U48885 (N_48885,N_32412,N_38166);
nand U48886 (N_48886,N_38482,N_33786);
xnor U48887 (N_48887,N_30162,N_35172);
and U48888 (N_48888,N_39682,N_33075);
or U48889 (N_48889,N_36358,N_35797);
nand U48890 (N_48890,N_36794,N_32048);
nand U48891 (N_48891,N_36754,N_30837);
nand U48892 (N_48892,N_30995,N_31948);
nand U48893 (N_48893,N_34667,N_31020);
nand U48894 (N_48894,N_32862,N_36488);
or U48895 (N_48895,N_36655,N_37201);
or U48896 (N_48896,N_31385,N_33629);
nor U48897 (N_48897,N_33995,N_32066);
and U48898 (N_48898,N_31569,N_36656);
and U48899 (N_48899,N_32190,N_39755);
and U48900 (N_48900,N_35251,N_38435);
nor U48901 (N_48901,N_37698,N_35195);
and U48902 (N_48902,N_36546,N_32826);
and U48903 (N_48903,N_39336,N_31040);
nor U48904 (N_48904,N_32189,N_32038);
nor U48905 (N_48905,N_30014,N_37413);
or U48906 (N_48906,N_31052,N_34475);
or U48907 (N_48907,N_32373,N_39400);
nand U48908 (N_48908,N_32143,N_32338);
or U48909 (N_48909,N_37558,N_37559);
nand U48910 (N_48910,N_31543,N_36337);
xor U48911 (N_48911,N_34416,N_30522);
or U48912 (N_48912,N_30338,N_32461);
nand U48913 (N_48913,N_36167,N_37272);
nor U48914 (N_48914,N_36110,N_34364);
and U48915 (N_48915,N_39562,N_32994);
xor U48916 (N_48916,N_35236,N_32070);
xor U48917 (N_48917,N_36489,N_36446);
or U48918 (N_48918,N_35981,N_32445);
or U48919 (N_48919,N_32780,N_38759);
nand U48920 (N_48920,N_37600,N_38594);
nor U48921 (N_48921,N_31977,N_31868);
or U48922 (N_48922,N_37450,N_38135);
or U48923 (N_48923,N_34909,N_30846);
or U48924 (N_48924,N_31958,N_30065);
nand U48925 (N_48925,N_36363,N_34814);
or U48926 (N_48926,N_39664,N_34499);
xnor U48927 (N_48927,N_31645,N_37236);
nand U48928 (N_48928,N_38328,N_33386);
nand U48929 (N_48929,N_30434,N_34841);
nand U48930 (N_48930,N_39818,N_33776);
and U48931 (N_48931,N_30530,N_34588);
and U48932 (N_48932,N_35996,N_35279);
and U48933 (N_48933,N_31378,N_32570);
nor U48934 (N_48934,N_36870,N_30278);
nor U48935 (N_48935,N_36470,N_30765);
and U48936 (N_48936,N_36611,N_31849);
xnor U48937 (N_48937,N_39814,N_37316);
nor U48938 (N_48938,N_36025,N_30538);
nor U48939 (N_48939,N_37231,N_30932);
nor U48940 (N_48940,N_30942,N_36969);
nand U48941 (N_48941,N_37265,N_30055);
and U48942 (N_48942,N_31987,N_30326);
nand U48943 (N_48943,N_30156,N_37508);
or U48944 (N_48944,N_35345,N_38318);
xor U48945 (N_48945,N_36853,N_35778);
and U48946 (N_48946,N_30049,N_35370);
or U48947 (N_48947,N_39334,N_37177);
nor U48948 (N_48948,N_33460,N_30208);
nand U48949 (N_48949,N_35376,N_39251);
nor U48950 (N_48950,N_31160,N_31973);
and U48951 (N_48951,N_38647,N_31029);
nor U48952 (N_48952,N_33280,N_37732);
or U48953 (N_48953,N_38271,N_34194);
nor U48954 (N_48954,N_36567,N_30440);
or U48955 (N_48955,N_33535,N_36043);
or U48956 (N_48956,N_39969,N_33991);
or U48957 (N_48957,N_32220,N_38665);
and U48958 (N_48958,N_30723,N_33407);
xor U48959 (N_48959,N_35472,N_39891);
and U48960 (N_48960,N_34368,N_30303);
nand U48961 (N_48961,N_38687,N_36475);
xor U48962 (N_48962,N_39534,N_32966);
nor U48963 (N_48963,N_39400,N_34327);
nor U48964 (N_48964,N_34252,N_35405);
nand U48965 (N_48965,N_37626,N_32213);
and U48966 (N_48966,N_32511,N_33188);
or U48967 (N_48967,N_36437,N_32902);
nor U48968 (N_48968,N_33773,N_39207);
or U48969 (N_48969,N_32643,N_32944);
nand U48970 (N_48970,N_34251,N_32434);
and U48971 (N_48971,N_34349,N_37733);
or U48972 (N_48972,N_37058,N_38248);
and U48973 (N_48973,N_31636,N_38108);
nand U48974 (N_48974,N_38985,N_36658);
nand U48975 (N_48975,N_33025,N_30247);
nor U48976 (N_48976,N_36991,N_33540);
nor U48977 (N_48977,N_37946,N_38318);
or U48978 (N_48978,N_37781,N_30569);
nor U48979 (N_48979,N_37886,N_34909);
and U48980 (N_48980,N_37648,N_31242);
or U48981 (N_48981,N_34459,N_37735);
nand U48982 (N_48982,N_37854,N_37889);
nand U48983 (N_48983,N_30190,N_37494);
nand U48984 (N_48984,N_34736,N_39860);
or U48985 (N_48985,N_38677,N_31968);
xnor U48986 (N_48986,N_33921,N_34593);
nor U48987 (N_48987,N_33343,N_31623);
nor U48988 (N_48988,N_33890,N_34672);
nor U48989 (N_48989,N_33403,N_34272);
or U48990 (N_48990,N_32847,N_32111);
nor U48991 (N_48991,N_39847,N_33782);
or U48992 (N_48992,N_30190,N_35696);
or U48993 (N_48993,N_34625,N_39821);
nor U48994 (N_48994,N_37790,N_32503);
nand U48995 (N_48995,N_36638,N_37258);
nor U48996 (N_48996,N_30502,N_39792);
nor U48997 (N_48997,N_36919,N_38038);
and U48998 (N_48998,N_36014,N_31673);
nor U48999 (N_48999,N_30764,N_32795);
nor U49000 (N_49000,N_39985,N_35642);
nand U49001 (N_49001,N_33705,N_39776);
and U49002 (N_49002,N_30275,N_38208);
and U49003 (N_49003,N_39311,N_36828);
and U49004 (N_49004,N_39098,N_34872);
nor U49005 (N_49005,N_39702,N_38195);
or U49006 (N_49006,N_31261,N_36990);
nor U49007 (N_49007,N_39378,N_39873);
and U49008 (N_49008,N_39771,N_38488);
nor U49009 (N_49009,N_32831,N_33556);
or U49010 (N_49010,N_31578,N_32268);
or U49011 (N_49011,N_35923,N_38155);
or U49012 (N_49012,N_36770,N_33457);
nand U49013 (N_49013,N_30298,N_34586);
and U49014 (N_49014,N_35772,N_33310);
nand U49015 (N_49015,N_38319,N_38467);
and U49016 (N_49016,N_32740,N_33068);
nand U49017 (N_49017,N_32929,N_39686);
and U49018 (N_49018,N_30967,N_33793);
nor U49019 (N_49019,N_37112,N_33917);
nor U49020 (N_49020,N_39948,N_36719);
and U49021 (N_49021,N_35891,N_38856);
and U49022 (N_49022,N_36194,N_33559);
nor U49023 (N_49023,N_37671,N_30122);
nand U49024 (N_49024,N_35139,N_31436);
nor U49025 (N_49025,N_39062,N_31674);
or U49026 (N_49026,N_39095,N_39177);
and U49027 (N_49027,N_35332,N_39640);
or U49028 (N_49028,N_37715,N_34439);
nand U49029 (N_49029,N_30143,N_37663);
nor U49030 (N_49030,N_32889,N_37905);
nand U49031 (N_49031,N_38904,N_35529);
and U49032 (N_49032,N_38130,N_32557);
or U49033 (N_49033,N_36505,N_37697);
nand U49034 (N_49034,N_30530,N_34263);
nand U49035 (N_49035,N_38676,N_35427);
and U49036 (N_49036,N_38775,N_38534);
and U49037 (N_49037,N_36086,N_31216);
or U49038 (N_49038,N_36885,N_35964);
nand U49039 (N_49039,N_34600,N_33740);
or U49040 (N_49040,N_31778,N_39364);
nand U49041 (N_49041,N_33243,N_33506);
and U49042 (N_49042,N_38904,N_37985);
nor U49043 (N_49043,N_39880,N_32902);
and U49044 (N_49044,N_34634,N_33186);
or U49045 (N_49045,N_34934,N_36887);
nor U49046 (N_49046,N_36791,N_38103);
or U49047 (N_49047,N_31866,N_39142);
nor U49048 (N_49048,N_34637,N_31137);
nor U49049 (N_49049,N_38556,N_35771);
nand U49050 (N_49050,N_39034,N_30532);
nor U49051 (N_49051,N_39860,N_34761);
nor U49052 (N_49052,N_33918,N_39041);
or U49053 (N_49053,N_30698,N_38146);
and U49054 (N_49054,N_31472,N_39721);
or U49055 (N_49055,N_38029,N_30625);
and U49056 (N_49056,N_37282,N_34880);
xnor U49057 (N_49057,N_35636,N_36496);
nand U49058 (N_49058,N_35107,N_38396);
nand U49059 (N_49059,N_35505,N_30861);
and U49060 (N_49060,N_33892,N_37016);
xor U49061 (N_49061,N_36448,N_37978);
or U49062 (N_49062,N_38546,N_32844);
nand U49063 (N_49063,N_36572,N_39907);
and U49064 (N_49064,N_38062,N_39894);
nand U49065 (N_49065,N_39816,N_33146);
nor U49066 (N_49066,N_35170,N_32239);
xnor U49067 (N_49067,N_30002,N_30218);
or U49068 (N_49068,N_34546,N_31902);
or U49069 (N_49069,N_35061,N_34969);
and U49070 (N_49070,N_36083,N_33958);
or U49071 (N_49071,N_37052,N_33468);
xnor U49072 (N_49072,N_39357,N_35569);
and U49073 (N_49073,N_34845,N_32994);
and U49074 (N_49074,N_37328,N_34411);
or U49075 (N_49075,N_34856,N_36075);
or U49076 (N_49076,N_36681,N_32715);
nor U49077 (N_49077,N_31559,N_33143);
nor U49078 (N_49078,N_31485,N_38788);
and U49079 (N_49079,N_37078,N_30313);
nor U49080 (N_49080,N_33130,N_38217);
and U49081 (N_49081,N_39029,N_32507);
nand U49082 (N_49082,N_31865,N_33735);
and U49083 (N_49083,N_30543,N_36197);
nand U49084 (N_49084,N_32631,N_36623);
xor U49085 (N_49085,N_33956,N_34890);
and U49086 (N_49086,N_30955,N_36431);
nand U49087 (N_49087,N_36604,N_34866);
and U49088 (N_49088,N_34904,N_35292);
nor U49089 (N_49089,N_35920,N_35065);
nand U49090 (N_49090,N_36970,N_32709);
nand U49091 (N_49091,N_35682,N_31029);
and U49092 (N_49092,N_35591,N_33621);
nor U49093 (N_49093,N_33948,N_37895);
nand U49094 (N_49094,N_32371,N_32502);
nor U49095 (N_49095,N_33509,N_36440);
or U49096 (N_49096,N_35968,N_39045);
xor U49097 (N_49097,N_37878,N_35214);
nand U49098 (N_49098,N_38727,N_37141);
and U49099 (N_49099,N_37794,N_31080);
or U49100 (N_49100,N_33792,N_30854);
nand U49101 (N_49101,N_34996,N_32590);
xnor U49102 (N_49102,N_39113,N_30952);
or U49103 (N_49103,N_32321,N_33528);
or U49104 (N_49104,N_35673,N_35181);
nor U49105 (N_49105,N_35917,N_38293);
or U49106 (N_49106,N_36917,N_37054);
nor U49107 (N_49107,N_35530,N_36825);
nor U49108 (N_49108,N_30344,N_31293);
xor U49109 (N_49109,N_32946,N_38072);
nor U49110 (N_49110,N_37401,N_33843);
nand U49111 (N_49111,N_33922,N_39103);
or U49112 (N_49112,N_31483,N_38630);
nor U49113 (N_49113,N_39378,N_33843);
and U49114 (N_49114,N_30941,N_38151);
or U49115 (N_49115,N_33634,N_30650);
and U49116 (N_49116,N_34447,N_33356);
nand U49117 (N_49117,N_39665,N_35916);
nor U49118 (N_49118,N_37659,N_33451);
or U49119 (N_49119,N_39122,N_38012);
or U49120 (N_49120,N_36949,N_35661);
or U49121 (N_49121,N_38088,N_32729);
xor U49122 (N_49122,N_31610,N_36233);
nand U49123 (N_49123,N_35953,N_39857);
or U49124 (N_49124,N_31842,N_31010);
or U49125 (N_49125,N_37772,N_34645);
nor U49126 (N_49126,N_38587,N_39666);
nand U49127 (N_49127,N_33251,N_34470);
xor U49128 (N_49128,N_35519,N_35448);
nor U49129 (N_49129,N_38623,N_36566);
or U49130 (N_49130,N_31910,N_36606);
nand U49131 (N_49131,N_31371,N_30680);
nand U49132 (N_49132,N_31496,N_31478);
nand U49133 (N_49133,N_36563,N_37799);
nor U49134 (N_49134,N_35048,N_33812);
nand U49135 (N_49135,N_33813,N_30569);
xor U49136 (N_49136,N_35500,N_34582);
nor U49137 (N_49137,N_30853,N_35173);
nor U49138 (N_49138,N_39091,N_32914);
nor U49139 (N_49139,N_33418,N_35386);
or U49140 (N_49140,N_34940,N_38780);
or U49141 (N_49141,N_33848,N_38266);
nand U49142 (N_49142,N_37748,N_32175);
and U49143 (N_49143,N_39705,N_38606);
xor U49144 (N_49144,N_38862,N_38773);
and U49145 (N_49145,N_31480,N_31819);
nand U49146 (N_49146,N_30641,N_34755);
and U49147 (N_49147,N_39680,N_35742);
and U49148 (N_49148,N_32487,N_36032);
xor U49149 (N_49149,N_34332,N_38118);
and U49150 (N_49150,N_32951,N_39991);
and U49151 (N_49151,N_35507,N_39865);
and U49152 (N_49152,N_33219,N_33362);
nor U49153 (N_49153,N_37162,N_31673);
xor U49154 (N_49154,N_34420,N_30278);
and U49155 (N_49155,N_32617,N_39501);
xnor U49156 (N_49156,N_34592,N_33246);
and U49157 (N_49157,N_33210,N_34325);
nand U49158 (N_49158,N_39470,N_30662);
nor U49159 (N_49159,N_39787,N_30411);
and U49160 (N_49160,N_35180,N_32690);
or U49161 (N_49161,N_37130,N_37746);
nor U49162 (N_49162,N_37442,N_30711);
nor U49163 (N_49163,N_33016,N_36466);
nand U49164 (N_49164,N_37482,N_31926);
nand U49165 (N_49165,N_33668,N_36535);
and U49166 (N_49166,N_31600,N_33709);
nor U49167 (N_49167,N_31237,N_36235);
or U49168 (N_49168,N_34944,N_35655);
xnor U49169 (N_49169,N_38171,N_37604);
or U49170 (N_49170,N_30069,N_38281);
nor U49171 (N_49171,N_31891,N_37084);
xnor U49172 (N_49172,N_31192,N_36342);
and U49173 (N_49173,N_32977,N_39569);
or U49174 (N_49174,N_38545,N_36947);
and U49175 (N_49175,N_39687,N_31904);
or U49176 (N_49176,N_34465,N_37963);
or U49177 (N_49177,N_32932,N_32365);
or U49178 (N_49178,N_31673,N_31625);
xnor U49179 (N_49179,N_39048,N_30299);
and U49180 (N_49180,N_35652,N_38701);
and U49181 (N_49181,N_36170,N_37204);
and U49182 (N_49182,N_38245,N_37803);
or U49183 (N_49183,N_30617,N_38331);
nand U49184 (N_49184,N_36805,N_37427);
and U49185 (N_49185,N_31503,N_36509);
nor U49186 (N_49186,N_33503,N_39276);
and U49187 (N_49187,N_31167,N_37803);
nand U49188 (N_49188,N_37912,N_33477);
xor U49189 (N_49189,N_35583,N_36937);
nor U49190 (N_49190,N_34191,N_35391);
and U49191 (N_49191,N_31166,N_37123);
nand U49192 (N_49192,N_30970,N_34815);
nand U49193 (N_49193,N_39154,N_39632);
nor U49194 (N_49194,N_30716,N_31692);
nand U49195 (N_49195,N_37166,N_36774);
xor U49196 (N_49196,N_36233,N_38803);
nor U49197 (N_49197,N_39107,N_38354);
nor U49198 (N_49198,N_37121,N_38340);
nand U49199 (N_49199,N_31988,N_31002);
or U49200 (N_49200,N_33114,N_38082);
nor U49201 (N_49201,N_38975,N_34650);
and U49202 (N_49202,N_34455,N_34581);
or U49203 (N_49203,N_38296,N_35082);
xor U49204 (N_49204,N_34208,N_36076);
nand U49205 (N_49205,N_34314,N_39671);
nand U49206 (N_49206,N_38086,N_37783);
and U49207 (N_49207,N_34374,N_39742);
nand U49208 (N_49208,N_36006,N_34597);
nor U49209 (N_49209,N_39467,N_31514);
nor U49210 (N_49210,N_33751,N_39318);
nand U49211 (N_49211,N_35515,N_34097);
nand U49212 (N_49212,N_35347,N_33710);
and U49213 (N_49213,N_34602,N_35603);
nor U49214 (N_49214,N_39782,N_31315);
and U49215 (N_49215,N_32351,N_30744);
and U49216 (N_49216,N_32534,N_39244);
and U49217 (N_49217,N_30605,N_31680);
and U49218 (N_49218,N_34298,N_33771);
nand U49219 (N_49219,N_35412,N_36565);
and U49220 (N_49220,N_32770,N_30349);
or U49221 (N_49221,N_31761,N_36508);
or U49222 (N_49222,N_34006,N_39759);
and U49223 (N_49223,N_31718,N_36944);
nand U49224 (N_49224,N_34962,N_38529);
nand U49225 (N_49225,N_31337,N_35788);
nor U49226 (N_49226,N_33682,N_30293);
or U49227 (N_49227,N_37922,N_33800);
or U49228 (N_49228,N_33261,N_32780);
or U49229 (N_49229,N_36094,N_33293);
xor U49230 (N_49230,N_36139,N_32404);
or U49231 (N_49231,N_39518,N_30892);
or U49232 (N_49232,N_32234,N_39858);
nor U49233 (N_49233,N_39230,N_37433);
nand U49234 (N_49234,N_37545,N_34902);
nor U49235 (N_49235,N_36542,N_33779);
nor U49236 (N_49236,N_30157,N_36485);
nand U49237 (N_49237,N_35165,N_38410);
nor U49238 (N_49238,N_30422,N_35000);
and U49239 (N_49239,N_38623,N_32802);
nand U49240 (N_49240,N_30515,N_31578);
and U49241 (N_49241,N_30583,N_38785);
nor U49242 (N_49242,N_36056,N_36207);
and U49243 (N_49243,N_36579,N_34640);
xor U49244 (N_49244,N_34184,N_33770);
or U49245 (N_49245,N_36343,N_38671);
xor U49246 (N_49246,N_31882,N_34580);
nor U49247 (N_49247,N_34870,N_35708);
nand U49248 (N_49248,N_36606,N_37042);
or U49249 (N_49249,N_31006,N_37253);
or U49250 (N_49250,N_30194,N_37511);
and U49251 (N_49251,N_39033,N_37875);
nor U49252 (N_49252,N_37009,N_36011);
nor U49253 (N_49253,N_32586,N_36306);
or U49254 (N_49254,N_34049,N_33170);
and U49255 (N_49255,N_34199,N_32796);
nand U49256 (N_49256,N_35523,N_39481);
nand U49257 (N_49257,N_33913,N_38435);
or U49258 (N_49258,N_31420,N_32631);
and U49259 (N_49259,N_30077,N_37701);
nor U49260 (N_49260,N_34711,N_33182);
nand U49261 (N_49261,N_30192,N_34953);
or U49262 (N_49262,N_30007,N_34413);
or U49263 (N_49263,N_35078,N_30445);
xor U49264 (N_49264,N_30658,N_36815);
nand U49265 (N_49265,N_34639,N_35417);
xnor U49266 (N_49266,N_39801,N_30548);
and U49267 (N_49267,N_36834,N_38551);
and U49268 (N_49268,N_35973,N_33949);
nor U49269 (N_49269,N_35236,N_37607);
nand U49270 (N_49270,N_31729,N_30145);
nor U49271 (N_49271,N_32256,N_31849);
nand U49272 (N_49272,N_33062,N_35913);
and U49273 (N_49273,N_36944,N_32208);
and U49274 (N_49274,N_36130,N_32276);
or U49275 (N_49275,N_38415,N_39498);
xnor U49276 (N_49276,N_32581,N_36830);
xor U49277 (N_49277,N_39534,N_31598);
and U49278 (N_49278,N_37695,N_37221);
nor U49279 (N_49279,N_39743,N_33890);
or U49280 (N_49280,N_32836,N_39617);
or U49281 (N_49281,N_36540,N_32467);
nand U49282 (N_49282,N_39722,N_38418);
nand U49283 (N_49283,N_34421,N_32998);
nand U49284 (N_49284,N_37511,N_31120);
nor U49285 (N_49285,N_31418,N_30541);
or U49286 (N_49286,N_33522,N_36975);
or U49287 (N_49287,N_39185,N_36456);
or U49288 (N_49288,N_38782,N_30029);
or U49289 (N_49289,N_35545,N_39627);
and U49290 (N_49290,N_30240,N_30010);
nor U49291 (N_49291,N_31527,N_36684);
nand U49292 (N_49292,N_38114,N_39394);
and U49293 (N_49293,N_37385,N_31739);
xnor U49294 (N_49294,N_39017,N_31634);
and U49295 (N_49295,N_34954,N_33032);
nand U49296 (N_49296,N_34618,N_39373);
nand U49297 (N_49297,N_37896,N_38110);
nand U49298 (N_49298,N_39081,N_31177);
xnor U49299 (N_49299,N_31774,N_33541);
nor U49300 (N_49300,N_30837,N_35893);
xor U49301 (N_49301,N_35086,N_32233);
nor U49302 (N_49302,N_33940,N_38554);
and U49303 (N_49303,N_39110,N_35361);
or U49304 (N_49304,N_34819,N_36449);
and U49305 (N_49305,N_37583,N_30331);
xnor U49306 (N_49306,N_39460,N_39709);
and U49307 (N_49307,N_36702,N_30342);
nand U49308 (N_49308,N_30156,N_33839);
or U49309 (N_49309,N_35376,N_34333);
and U49310 (N_49310,N_31842,N_32756);
nor U49311 (N_49311,N_38584,N_33362);
nand U49312 (N_49312,N_35640,N_33266);
nand U49313 (N_49313,N_35104,N_32037);
nor U49314 (N_49314,N_39549,N_34544);
nor U49315 (N_49315,N_35312,N_31564);
or U49316 (N_49316,N_32975,N_35686);
nor U49317 (N_49317,N_36115,N_34436);
xnor U49318 (N_49318,N_38353,N_31555);
nor U49319 (N_49319,N_32248,N_36071);
xor U49320 (N_49320,N_37201,N_34701);
and U49321 (N_49321,N_35681,N_35178);
xnor U49322 (N_49322,N_34129,N_32004);
nor U49323 (N_49323,N_32943,N_32871);
and U49324 (N_49324,N_33168,N_30331);
and U49325 (N_49325,N_37968,N_39407);
nand U49326 (N_49326,N_33104,N_35888);
nor U49327 (N_49327,N_37381,N_32697);
and U49328 (N_49328,N_30889,N_35796);
or U49329 (N_49329,N_34578,N_34959);
and U49330 (N_49330,N_36954,N_36219);
xor U49331 (N_49331,N_31240,N_39853);
xnor U49332 (N_49332,N_37480,N_37215);
or U49333 (N_49333,N_35977,N_33765);
or U49334 (N_49334,N_36697,N_33278);
nand U49335 (N_49335,N_37567,N_30594);
nand U49336 (N_49336,N_32064,N_36992);
nand U49337 (N_49337,N_36778,N_36145);
nand U49338 (N_49338,N_31677,N_39841);
nor U49339 (N_49339,N_34944,N_37679);
and U49340 (N_49340,N_36482,N_36674);
and U49341 (N_49341,N_38518,N_37762);
or U49342 (N_49342,N_30001,N_31885);
nand U49343 (N_49343,N_31206,N_37504);
or U49344 (N_49344,N_34229,N_33388);
nor U49345 (N_49345,N_36394,N_38559);
nor U49346 (N_49346,N_33447,N_39307);
xor U49347 (N_49347,N_30062,N_35667);
nor U49348 (N_49348,N_32827,N_31030);
nor U49349 (N_49349,N_33925,N_34102);
xor U49350 (N_49350,N_36755,N_35302);
and U49351 (N_49351,N_33238,N_32064);
nor U49352 (N_49352,N_31253,N_37602);
or U49353 (N_49353,N_32376,N_31585);
nor U49354 (N_49354,N_38895,N_35601);
or U49355 (N_49355,N_34673,N_30034);
nand U49356 (N_49356,N_36884,N_37836);
or U49357 (N_49357,N_35542,N_31283);
or U49358 (N_49358,N_38838,N_36986);
xor U49359 (N_49359,N_30847,N_35798);
nand U49360 (N_49360,N_32475,N_32763);
nor U49361 (N_49361,N_39358,N_30499);
nand U49362 (N_49362,N_36456,N_35094);
or U49363 (N_49363,N_31461,N_30941);
and U49364 (N_49364,N_35033,N_37228);
and U49365 (N_49365,N_35787,N_33888);
xor U49366 (N_49366,N_34010,N_39007);
nor U49367 (N_49367,N_35185,N_30657);
or U49368 (N_49368,N_35765,N_33577);
and U49369 (N_49369,N_37498,N_34132);
nand U49370 (N_49370,N_39627,N_37014);
nor U49371 (N_49371,N_37383,N_33126);
nand U49372 (N_49372,N_30618,N_30805);
nand U49373 (N_49373,N_38805,N_39556);
or U49374 (N_49374,N_31262,N_34295);
nand U49375 (N_49375,N_37313,N_31077);
nand U49376 (N_49376,N_31736,N_38231);
nor U49377 (N_49377,N_39903,N_32689);
xor U49378 (N_49378,N_39933,N_30235);
or U49379 (N_49379,N_37975,N_39419);
nand U49380 (N_49380,N_31565,N_37642);
and U49381 (N_49381,N_31684,N_33230);
nand U49382 (N_49382,N_39390,N_38754);
and U49383 (N_49383,N_33551,N_37377);
and U49384 (N_49384,N_38105,N_33927);
nand U49385 (N_49385,N_30816,N_39006);
or U49386 (N_49386,N_34248,N_38753);
and U49387 (N_49387,N_38698,N_34381);
nand U49388 (N_49388,N_33862,N_37092);
and U49389 (N_49389,N_31186,N_37908);
and U49390 (N_49390,N_32247,N_36950);
and U49391 (N_49391,N_36002,N_33066);
and U49392 (N_49392,N_30619,N_31647);
or U49393 (N_49393,N_34530,N_32695);
nand U49394 (N_49394,N_35430,N_35872);
or U49395 (N_49395,N_38889,N_37495);
and U49396 (N_49396,N_36709,N_30676);
xnor U49397 (N_49397,N_36864,N_39310);
or U49398 (N_49398,N_39130,N_31757);
and U49399 (N_49399,N_37103,N_37545);
or U49400 (N_49400,N_34109,N_35202);
or U49401 (N_49401,N_32878,N_31461);
and U49402 (N_49402,N_35051,N_38105);
nor U49403 (N_49403,N_37486,N_39340);
or U49404 (N_49404,N_37314,N_34788);
nor U49405 (N_49405,N_30408,N_32034);
nand U49406 (N_49406,N_37127,N_37308);
and U49407 (N_49407,N_33588,N_34766);
xnor U49408 (N_49408,N_37724,N_39821);
or U49409 (N_49409,N_37153,N_31857);
nor U49410 (N_49410,N_30455,N_37790);
and U49411 (N_49411,N_32321,N_37751);
nand U49412 (N_49412,N_39844,N_36057);
or U49413 (N_49413,N_39647,N_34745);
or U49414 (N_49414,N_30273,N_33015);
or U49415 (N_49415,N_30421,N_38130);
xor U49416 (N_49416,N_38488,N_36391);
nor U49417 (N_49417,N_36030,N_38632);
nor U49418 (N_49418,N_34440,N_39802);
and U49419 (N_49419,N_39589,N_34423);
nor U49420 (N_49420,N_38179,N_36570);
or U49421 (N_49421,N_34098,N_36674);
nor U49422 (N_49422,N_34370,N_34309);
nand U49423 (N_49423,N_31274,N_32172);
nand U49424 (N_49424,N_31128,N_38606);
and U49425 (N_49425,N_39635,N_33671);
nand U49426 (N_49426,N_38728,N_31668);
xor U49427 (N_49427,N_39138,N_38621);
nand U49428 (N_49428,N_32311,N_31544);
or U49429 (N_49429,N_38935,N_33706);
nand U49430 (N_49430,N_35543,N_38942);
nand U49431 (N_49431,N_33774,N_36544);
xor U49432 (N_49432,N_34250,N_35109);
or U49433 (N_49433,N_34255,N_37355);
nand U49434 (N_49434,N_32333,N_30273);
nor U49435 (N_49435,N_36297,N_39728);
nand U49436 (N_49436,N_33884,N_30161);
or U49437 (N_49437,N_38376,N_35056);
nand U49438 (N_49438,N_32786,N_34124);
and U49439 (N_49439,N_35079,N_34075);
or U49440 (N_49440,N_30317,N_34920);
xor U49441 (N_49441,N_37291,N_38797);
nand U49442 (N_49442,N_30601,N_37244);
and U49443 (N_49443,N_34216,N_37466);
and U49444 (N_49444,N_35061,N_38476);
nor U49445 (N_49445,N_30466,N_38366);
or U49446 (N_49446,N_33590,N_34968);
xor U49447 (N_49447,N_38534,N_31359);
and U49448 (N_49448,N_31425,N_39985);
or U49449 (N_49449,N_32455,N_37165);
or U49450 (N_49450,N_36811,N_38481);
or U49451 (N_49451,N_37682,N_35211);
nand U49452 (N_49452,N_31148,N_31818);
nand U49453 (N_49453,N_33736,N_35606);
or U49454 (N_49454,N_36831,N_35810);
xnor U49455 (N_49455,N_37058,N_39922);
nor U49456 (N_49456,N_39921,N_31039);
and U49457 (N_49457,N_35112,N_37270);
nand U49458 (N_49458,N_36233,N_36421);
nor U49459 (N_49459,N_37086,N_34748);
and U49460 (N_49460,N_36860,N_31271);
nor U49461 (N_49461,N_39312,N_37639);
nor U49462 (N_49462,N_38603,N_39467);
nand U49463 (N_49463,N_33233,N_31132);
and U49464 (N_49464,N_30142,N_33950);
and U49465 (N_49465,N_34294,N_30840);
nor U49466 (N_49466,N_30248,N_33779);
nand U49467 (N_49467,N_33959,N_30300);
nand U49468 (N_49468,N_32842,N_39719);
nor U49469 (N_49469,N_36296,N_37216);
or U49470 (N_49470,N_36343,N_31595);
and U49471 (N_49471,N_36912,N_34750);
nor U49472 (N_49472,N_39563,N_35152);
or U49473 (N_49473,N_30491,N_32886);
or U49474 (N_49474,N_38627,N_30427);
or U49475 (N_49475,N_36523,N_30223);
or U49476 (N_49476,N_30396,N_38103);
xnor U49477 (N_49477,N_35310,N_34683);
or U49478 (N_49478,N_33535,N_37550);
xor U49479 (N_49479,N_30156,N_39224);
or U49480 (N_49480,N_33517,N_32630);
or U49481 (N_49481,N_36977,N_35647);
nor U49482 (N_49482,N_39645,N_32175);
nor U49483 (N_49483,N_33676,N_37650);
or U49484 (N_49484,N_34942,N_36573);
nand U49485 (N_49485,N_33192,N_30742);
xor U49486 (N_49486,N_30727,N_39494);
nand U49487 (N_49487,N_37409,N_32150);
nor U49488 (N_49488,N_37584,N_39404);
nand U49489 (N_49489,N_31003,N_37228);
nand U49490 (N_49490,N_33131,N_34349);
nand U49491 (N_49491,N_31326,N_38677);
or U49492 (N_49492,N_31548,N_30839);
or U49493 (N_49493,N_36482,N_33852);
and U49494 (N_49494,N_38820,N_33293);
or U49495 (N_49495,N_34322,N_39814);
or U49496 (N_49496,N_38000,N_33474);
or U49497 (N_49497,N_34346,N_39922);
or U49498 (N_49498,N_38096,N_39285);
and U49499 (N_49499,N_30488,N_38062);
nand U49500 (N_49500,N_32408,N_33285);
xor U49501 (N_49501,N_35788,N_39975);
or U49502 (N_49502,N_37721,N_34581);
and U49503 (N_49503,N_30663,N_32446);
nor U49504 (N_49504,N_30606,N_38169);
nand U49505 (N_49505,N_31284,N_31135);
nor U49506 (N_49506,N_39128,N_33612);
and U49507 (N_49507,N_36861,N_32399);
nor U49508 (N_49508,N_31092,N_31199);
or U49509 (N_49509,N_38237,N_35340);
nand U49510 (N_49510,N_38667,N_30629);
nor U49511 (N_49511,N_32907,N_35084);
and U49512 (N_49512,N_33863,N_35049);
or U49513 (N_49513,N_31478,N_32553);
xnor U49514 (N_49514,N_35451,N_38892);
xor U49515 (N_49515,N_37172,N_31387);
nand U49516 (N_49516,N_30473,N_34391);
or U49517 (N_49517,N_38387,N_39799);
xnor U49518 (N_49518,N_37361,N_32576);
nor U49519 (N_49519,N_34950,N_33861);
nor U49520 (N_49520,N_34996,N_34282);
and U49521 (N_49521,N_30618,N_36239);
or U49522 (N_49522,N_34829,N_31117);
or U49523 (N_49523,N_38364,N_37198);
or U49524 (N_49524,N_36022,N_34876);
and U49525 (N_49525,N_32871,N_31721);
nor U49526 (N_49526,N_33139,N_34000);
nor U49527 (N_49527,N_30211,N_34191);
nand U49528 (N_49528,N_35342,N_37936);
or U49529 (N_49529,N_38557,N_35390);
nor U49530 (N_49530,N_34501,N_39355);
nand U49531 (N_49531,N_31457,N_35452);
xor U49532 (N_49532,N_39374,N_38109);
and U49533 (N_49533,N_36093,N_38438);
or U49534 (N_49534,N_39209,N_30005);
or U49535 (N_49535,N_35853,N_30360);
and U49536 (N_49536,N_30054,N_33252);
nor U49537 (N_49537,N_39639,N_30735);
and U49538 (N_49538,N_30448,N_39562);
and U49539 (N_49539,N_32776,N_31569);
and U49540 (N_49540,N_33409,N_38552);
nand U49541 (N_49541,N_32416,N_34609);
and U49542 (N_49542,N_39288,N_30064);
nand U49543 (N_49543,N_32772,N_34478);
nor U49544 (N_49544,N_31059,N_34678);
or U49545 (N_49545,N_38957,N_39583);
or U49546 (N_49546,N_31321,N_35048);
and U49547 (N_49547,N_35933,N_33469);
and U49548 (N_49548,N_33209,N_31716);
or U49549 (N_49549,N_34525,N_34002);
nor U49550 (N_49550,N_38253,N_38056);
or U49551 (N_49551,N_34713,N_37753);
nor U49552 (N_49552,N_36322,N_38110);
nor U49553 (N_49553,N_35381,N_32873);
and U49554 (N_49554,N_37130,N_31476);
or U49555 (N_49555,N_31495,N_30240);
nand U49556 (N_49556,N_37256,N_38830);
nor U49557 (N_49557,N_32897,N_30710);
and U49558 (N_49558,N_31601,N_37810);
and U49559 (N_49559,N_39298,N_37859);
nor U49560 (N_49560,N_35351,N_37081);
and U49561 (N_49561,N_30121,N_33210);
nor U49562 (N_49562,N_39721,N_35189);
and U49563 (N_49563,N_38790,N_33071);
nand U49564 (N_49564,N_34953,N_33867);
nor U49565 (N_49565,N_31236,N_32003);
and U49566 (N_49566,N_34141,N_32318);
nand U49567 (N_49567,N_34958,N_33736);
nand U49568 (N_49568,N_30655,N_31882);
nand U49569 (N_49569,N_33550,N_34925);
or U49570 (N_49570,N_31320,N_34502);
and U49571 (N_49571,N_30193,N_30867);
xnor U49572 (N_49572,N_30861,N_39420);
nor U49573 (N_49573,N_36409,N_34972);
nand U49574 (N_49574,N_33300,N_34686);
nor U49575 (N_49575,N_30939,N_33188);
or U49576 (N_49576,N_31663,N_31921);
nor U49577 (N_49577,N_32766,N_34441);
nand U49578 (N_49578,N_36366,N_35917);
xnor U49579 (N_49579,N_39183,N_30818);
nor U49580 (N_49580,N_34722,N_32261);
xor U49581 (N_49581,N_30107,N_30166);
and U49582 (N_49582,N_33728,N_36640);
or U49583 (N_49583,N_39617,N_36949);
and U49584 (N_49584,N_30985,N_30763);
nand U49585 (N_49585,N_34913,N_34196);
and U49586 (N_49586,N_39588,N_35103);
nand U49587 (N_49587,N_34469,N_37062);
or U49588 (N_49588,N_31650,N_39761);
nand U49589 (N_49589,N_31535,N_31293);
xor U49590 (N_49590,N_32477,N_36180);
and U49591 (N_49591,N_30013,N_31966);
xnor U49592 (N_49592,N_32763,N_35692);
nand U49593 (N_49593,N_34572,N_34233);
nand U49594 (N_49594,N_31744,N_33306);
and U49595 (N_49595,N_31085,N_37410);
nor U49596 (N_49596,N_39633,N_35770);
nand U49597 (N_49597,N_32630,N_39982);
or U49598 (N_49598,N_34950,N_32874);
nor U49599 (N_49599,N_30755,N_33877);
or U49600 (N_49600,N_34023,N_37345);
nor U49601 (N_49601,N_39042,N_39744);
or U49602 (N_49602,N_34649,N_35899);
nand U49603 (N_49603,N_32259,N_30050);
and U49604 (N_49604,N_38168,N_34739);
or U49605 (N_49605,N_36304,N_31823);
and U49606 (N_49606,N_31043,N_37788);
or U49607 (N_49607,N_32976,N_31828);
and U49608 (N_49608,N_34132,N_34288);
nor U49609 (N_49609,N_34607,N_36241);
nor U49610 (N_49610,N_36015,N_34319);
xor U49611 (N_49611,N_35872,N_36960);
xor U49612 (N_49612,N_35575,N_38513);
nor U49613 (N_49613,N_39784,N_34807);
and U49614 (N_49614,N_32685,N_34600);
and U49615 (N_49615,N_35683,N_37438);
or U49616 (N_49616,N_35170,N_39931);
and U49617 (N_49617,N_38938,N_37740);
nor U49618 (N_49618,N_34156,N_31743);
nand U49619 (N_49619,N_37463,N_32943);
nand U49620 (N_49620,N_37349,N_38836);
nand U49621 (N_49621,N_32715,N_38097);
nand U49622 (N_49622,N_34435,N_33722);
nand U49623 (N_49623,N_39989,N_38550);
nor U49624 (N_49624,N_30116,N_34039);
xnor U49625 (N_49625,N_39937,N_37300);
xor U49626 (N_49626,N_35082,N_33545);
and U49627 (N_49627,N_35932,N_31890);
nor U49628 (N_49628,N_34237,N_33379);
nor U49629 (N_49629,N_33152,N_37947);
nor U49630 (N_49630,N_36573,N_31028);
xor U49631 (N_49631,N_32677,N_30086);
nor U49632 (N_49632,N_36726,N_30999);
nor U49633 (N_49633,N_31709,N_31101);
nand U49634 (N_49634,N_34721,N_36989);
and U49635 (N_49635,N_33980,N_32528);
nor U49636 (N_49636,N_36334,N_38675);
nand U49637 (N_49637,N_36324,N_30416);
nor U49638 (N_49638,N_31256,N_36495);
and U49639 (N_49639,N_34624,N_37155);
nor U49640 (N_49640,N_32672,N_39806);
nand U49641 (N_49641,N_37134,N_38858);
nand U49642 (N_49642,N_32596,N_30075);
and U49643 (N_49643,N_38487,N_35549);
nor U49644 (N_49644,N_39606,N_32635);
xor U49645 (N_49645,N_38010,N_30759);
and U49646 (N_49646,N_30768,N_34075);
and U49647 (N_49647,N_38767,N_37501);
nand U49648 (N_49648,N_34766,N_34207);
nand U49649 (N_49649,N_33691,N_39937);
xnor U49650 (N_49650,N_39948,N_31592);
or U49651 (N_49651,N_31091,N_33046);
nand U49652 (N_49652,N_37345,N_35935);
and U49653 (N_49653,N_36250,N_31096);
and U49654 (N_49654,N_35184,N_39212);
nand U49655 (N_49655,N_33102,N_37357);
nand U49656 (N_49656,N_30944,N_37313);
and U49657 (N_49657,N_35001,N_30278);
and U49658 (N_49658,N_31719,N_31527);
or U49659 (N_49659,N_37728,N_33493);
xnor U49660 (N_49660,N_31463,N_33590);
nor U49661 (N_49661,N_35568,N_36174);
xnor U49662 (N_49662,N_32814,N_31743);
nand U49663 (N_49663,N_32430,N_38541);
or U49664 (N_49664,N_39235,N_35123);
and U49665 (N_49665,N_30335,N_33126);
or U49666 (N_49666,N_35011,N_36901);
and U49667 (N_49667,N_32408,N_34616);
nand U49668 (N_49668,N_36825,N_30201);
or U49669 (N_49669,N_31738,N_32730);
or U49670 (N_49670,N_31435,N_34961);
nand U49671 (N_49671,N_35584,N_39533);
nor U49672 (N_49672,N_34151,N_33261);
xor U49673 (N_49673,N_31683,N_37372);
nor U49674 (N_49674,N_31654,N_35940);
or U49675 (N_49675,N_36621,N_36680);
nand U49676 (N_49676,N_35419,N_32903);
nor U49677 (N_49677,N_37971,N_33652);
nor U49678 (N_49678,N_35642,N_30798);
nand U49679 (N_49679,N_38907,N_35698);
nand U49680 (N_49680,N_37629,N_37283);
nor U49681 (N_49681,N_37874,N_31942);
nand U49682 (N_49682,N_37655,N_36037);
nand U49683 (N_49683,N_39658,N_30177);
nor U49684 (N_49684,N_38480,N_30452);
xor U49685 (N_49685,N_34453,N_37222);
and U49686 (N_49686,N_34873,N_30743);
or U49687 (N_49687,N_33392,N_35303);
xor U49688 (N_49688,N_34870,N_35452);
nand U49689 (N_49689,N_39198,N_35935);
and U49690 (N_49690,N_32827,N_37845);
nand U49691 (N_49691,N_36054,N_32667);
or U49692 (N_49692,N_32107,N_33120);
or U49693 (N_49693,N_38537,N_36770);
and U49694 (N_49694,N_35614,N_35244);
and U49695 (N_49695,N_30653,N_32219);
and U49696 (N_49696,N_38540,N_31236);
and U49697 (N_49697,N_32338,N_38102);
or U49698 (N_49698,N_37897,N_32422);
or U49699 (N_49699,N_32250,N_34881);
nand U49700 (N_49700,N_38905,N_37415);
or U49701 (N_49701,N_30409,N_38049);
or U49702 (N_49702,N_38771,N_39705);
nor U49703 (N_49703,N_30823,N_32089);
xor U49704 (N_49704,N_36322,N_36939);
xor U49705 (N_49705,N_38462,N_39685);
or U49706 (N_49706,N_38210,N_30178);
nand U49707 (N_49707,N_34671,N_37764);
nand U49708 (N_49708,N_31906,N_30443);
or U49709 (N_49709,N_38193,N_36830);
nand U49710 (N_49710,N_32878,N_39783);
and U49711 (N_49711,N_30498,N_32650);
nor U49712 (N_49712,N_37169,N_35038);
and U49713 (N_49713,N_31583,N_36937);
nor U49714 (N_49714,N_30517,N_36885);
and U49715 (N_49715,N_37433,N_37268);
and U49716 (N_49716,N_39545,N_32890);
nand U49717 (N_49717,N_35998,N_33935);
and U49718 (N_49718,N_31120,N_30249);
nor U49719 (N_49719,N_31534,N_34867);
or U49720 (N_49720,N_31065,N_31531);
nor U49721 (N_49721,N_32348,N_33707);
and U49722 (N_49722,N_39702,N_32016);
and U49723 (N_49723,N_30281,N_30991);
nand U49724 (N_49724,N_37449,N_32425);
or U49725 (N_49725,N_30438,N_37007);
nand U49726 (N_49726,N_34015,N_35778);
nand U49727 (N_49727,N_31280,N_30053);
nand U49728 (N_49728,N_37680,N_33791);
or U49729 (N_49729,N_31357,N_37973);
nand U49730 (N_49730,N_39930,N_38490);
nand U49731 (N_49731,N_38909,N_30297);
and U49732 (N_49732,N_34104,N_32282);
or U49733 (N_49733,N_37218,N_39812);
and U49734 (N_49734,N_35355,N_39411);
xor U49735 (N_49735,N_33017,N_33316);
nand U49736 (N_49736,N_30258,N_38667);
nand U49737 (N_49737,N_36526,N_33668);
or U49738 (N_49738,N_30499,N_32012);
nor U49739 (N_49739,N_35963,N_35792);
or U49740 (N_49740,N_36181,N_39322);
and U49741 (N_49741,N_31590,N_34814);
nand U49742 (N_49742,N_35327,N_39243);
nand U49743 (N_49743,N_35687,N_35212);
nand U49744 (N_49744,N_38705,N_39001);
nand U49745 (N_49745,N_34848,N_39728);
or U49746 (N_49746,N_35354,N_35613);
and U49747 (N_49747,N_39628,N_37315);
and U49748 (N_49748,N_31437,N_30230);
or U49749 (N_49749,N_33068,N_34440);
nand U49750 (N_49750,N_33752,N_37405);
nor U49751 (N_49751,N_37893,N_36088);
nor U49752 (N_49752,N_39006,N_32059);
nor U49753 (N_49753,N_37569,N_36280);
xnor U49754 (N_49754,N_30934,N_38033);
nand U49755 (N_49755,N_39495,N_32940);
and U49756 (N_49756,N_33657,N_36236);
or U49757 (N_49757,N_31170,N_34792);
nor U49758 (N_49758,N_35846,N_36051);
xnor U49759 (N_49759,N_36389,N_35892);
nand U49760 (N_49760,N_37123,N_35718);
nor U49761 (N_49761,N_33066,N_36238);
nand U49762 (N_49762,N_35349,N_30969);
nor U49763 (N_49763,N_36438,N_36026);
and U49764 (N_49764,N_36683,N_32704);
nor U49765 (N_49765,N_36273,N_37668);
xor U49766 (N_49766,N_36012,N_34061);
and U49767 (N_49767,N_39757,N_37362);
nor U49768 (N_49768,N_33810,N_36852);
nor U49769 (N_49769,N_35301,N_34463);
xor U49770 (N_49770,N_36277,N_33271);
and U49771 (N_49771,N_38360,N_38962);
nand U49772 (N_49772,N_35743,N_33918);
or U49773 (N_49773,N_32547,N_39403);
xnor U49774 (N_49774,N_35205,N_34321);
or U49775 (N_49775,N_35490,N_37970);
nor U49776 (N_49776,N_39323,N_36982);
or U49777 (N_49777,N_33121,N_34375);
or U49778 (N_49778,N_32761,N_37084);
nor U49779 (N_49779,N_30622,N_32750);
or U49780 (N_49780,N_34844,N_30124);
or U49781 (N_49781,N_37889,N_31079);
nand U49782 (N_49782,N_35815,N_37139);
nand U49783 (N_49783,N_39946,N_35324);
and U49784 (N_49784,N_32585,N_36978);
nor U49785 (N_49785,N_33310,N_32398);
nand U49786 (N_49786,N_38564,N_30415);
or U49787 (N_49787,N_38415,N_38424);
xor U49788 (N_49788,N_36820,N_33562);
nor U49789 (N_49789,N_37072,N_37071);
or U49790 (N_49790,N_34091,N_34547);
and U49791 (N_49791,N_32237,N_37077);
and U49792 (N_49792,N_32802,N_35809);
and U49793 (N_49793,N_37626,N_38334);
and U49794 (N_49794,N_34820,N_34120);
and U49795 (N_49795,N_33339,N_38790);
nor U49796 (N_49796,N_33759,N_36494);
nand U49797 (N_49797,N_36553,N_34256);
or U49798 (N_49798,N_38939,N_34622);
and U49799 (N_49799,N_37868,N_31871);
and U49800 (N_49800,N_34036,N_35455);
and U49801 (N_49801,N_33230,N_35886);
and U49802 (N_49802,N_35090,N_30097);
nand U49803 (N_49803,N_39475,N_33705);
nand U49804 (N_49804,N_34329,N_32547);
nor U49805 (N_49805,N_30053,N_38814);
nor U49806 (N_49806,N_37882,N_32115);
or U49807 (N_49807,N_38865,N_37793);
or U49808 (N_49808,N_38503,N_35923);
nor U49809 (N_49809,N_36689,N_36202);
xnor U49810 (N_49810,N_38365,N_37127);
nand U49811 (N_49811,N_34563,N_39649);
and U49812 (N_49812,N_38201,N_31387);
and U49813 (N_49813,N_31375,N_36990);
nor U49814 (N_49814,N_33653,N_37539);
nand U49815 (N_49815,N_32975,N_32598);
nor U49816 (N_49816,N_38006,N_38820);
nor U49817 (N_49817,N_34001,N_39532);
and U49818 (N_49818,N_34203,N_30055);
nand U49819 (N_49819,N_38429,N_39748);
nand U49820 (N_49820,N_32198,N_38062);
nand U49821 (N_49821,N_39541,N_32210);
nand U49822 (N_49822,N_31983,N_39254);
xor U49823 (N_49823,N_38796,N_30568);
and U49824 (N_49824,N_35200,N_37744);
or U49825 (N_49825,N_35736,N_31435);
or U49826 (N_49826,N_35070,N_30791);
xnor U49827 (N_49827,N_30544,N_33024);
nand U49828 (N_49828,N_35363,N_31394);
nand U49829 (N_49829,N_38828,N_30031);
and U49830 (N_49830,N_37529,N_37091);
and U49831 (N_49831,N_39318,N_33171);
nand U49832 (N_49832,N_31153,N_39960);
and U49833 (N_49833,N_31033,N_31920);
or U49834 (N_49834,N_32043,N_38039);
or U49835 (N_49835,N_38728,N_32645);
nor U49836 (N_49836,N_34504,N_33816);
and U49837 (N_49837,N_31353,N_36349);
and U49838 (N_49838,N_38537,N_34129);
and U49839 (N_49839,N_34756,N_32249);
or U49840 (N_49840,N_39648,N_38015);
or U49841 (N_49841,N_35766,N_31534);
nand U49842 (N_49842,N_32660,N_38166);
or U49843 (N_49843,N_32372,N_30267);
or U49844 (N_49844,N_34453,N_30661);
nor U49845 (N_49845,N_38289,N_33988);
and U49846 (N_49846,N_39588,N_32989);
nand U49847 (N_49847,N_38771,N_36580);
or U49848 (N_49848,N_30947,N_36556);
nand U49849 (N_49849,N_39325,N_37393);
nor U49850 (N_49850,N_36250,N_38167);
nand U49851 (N_49851,N_35093,N_38595);
nand U49852 (N_49852,N_36481,N_30458);
nand U49853 (N_49853,N_31326,N_35102);
and U49854 (N_49854,N_35170,N_31535);
and U49855 (N_49855,N_35189,N_36448);
and U49856 (N_49856,N_39880,N_33060);
and U49857 (N_49857,N_33813,N_37212);
nor U49858 (N_49858,N_33420,N_38887);
xnor U49859 (N_49859,N_30436,N_37298);
nor U49860 (N_49860,N_33825,N_33989);
nand U49861 (N_49861,N_38568,N_31367);
or U49862 (N_49862,N_38864,N_37820);
and U49863 (N_49863,N_37502,N_34964);
nor U49864 (N_49864,N_31319,N_37397);
and U49865 (N_49865,N_31741,N_36286);
xor U49866 (N_49866,N_38278,N_39273);
or U49867 (N_49867,N_37307,N_34307);
nor U49868 (N_49868,N_33928,N_31021);
or U49869 (N_49869,N_32227,N_31058);
nand U49870 (N_49870,N_36970,N_39393);
or U49871 (N_49871,N_34182,N_30171);
nor U49872 (N_49872,N_38189,N_31445);
or U49873 (N_49873,N_31573,N_34095);
nor U49874 (N_49874,N_36130,N_38854);
and U49875 (N_49875,N_32559,N_30058);
nor U49876 (N_49876,N_34284,N_32504);
and U49877 (N_49877,N_33995,N_38948);
nand U49878 (N_49878,N_32775,N_33984);
xnor U49879 (N_49879,N_37973,N_37781);
nand U49880 (N_49880,N_35946,N_36827);
nor U49881 (N_49881,N_33038,N_38731);
and U49882 (N_49882,N_36039,N_39382);
and U49883 (N_49883,N_36230,N_34046);
or U49884 (N_49884,N_37800,N_32970);
or U49885 (N_49885,N_37896,N_32648);
nor U49886 (N_49886,N_39264,N_39820);
and U49887 (N_49887,N_39367,N_30470);
and U49888 (N_49888,N_35380,N_36855);
or U49889 (N_49889,N_32536,N_33033);
nor U49890 (N_49890,N_35097,N_37628);
or U49891 (N_49891,N_36049,N_34634);
or U49892 (N_49892,N_35772,N_34247);
nand U49893 (N_49893,N_36970,N_32813);
nor U49894 (N_49894,N_37631,N_36980);
and U49895 (N_49895,N_32500,N_35140);
or U49896 (N_49896,N_34978,N_36982);
nand U49897 (N_49897,N_32215,N_30364);
nor U49898 (N_49898,N_39572,N_32494);
nor U49899 (N_49899,N_36839,N_39519);
nor U49900 (N_49900,N_35546,N_33383);
xnor U49901 (N_49901,N_30804,N_36847);
nor U49902 (N_49902,N_33472,N_33154);
or U49903 (N_49903,N_36113,N_36044);
nor U49904 (N_49904,N_34133,N_35700);
xor U49905 (N_49905,N_32206,N_37430);
nor U49906 (N_49906,N_33121,N_30358);
nand U49907 (N_49907,N_31921,N_32628);
or U49908 (N_49908,N_39401,N_37102);
nand U49909 (N_49909,N_38993,N_34817);
xor U49910 (N_49910,N_37356,N_34251);
nand U49911 (N_49911,N_32693,N_31174);
and U49912 (N_49912,N_38597,N_38816);
xor U49913 (N_49913,N_33051,N_34700);
nand U49914 (N_49914,N_35145,N_34400);
nor U49915 (N_49915,N_36637,N_37034);
or U49916 (N_49916,N_36239,N_35339);
xor U49917 (N_49917,N_33969,N_35556);
nor U49918 (N_49918,N_30209,N_35212);
nor U49919 (N_49919,N_36313,N_31639);
nor U49920 (N_49920,N_39156,N_33975);
nand U49921 (N_49921,N_32434,N_37230);
nand U49922 (N_49922,N_36197,N_35878);
nand U49923 (N_49923,N_39949,N_34577);
nand U49924 (N_49924,N_30465,N_38888);
or U49925 (N_49925,N_37558,N_38806);
nand U49926 (N_49926,N_36502,N_31089);
and U49927 (N_49927,N_35403,N_36997);
nand U49928 (N_49928,N_36774,N_33083);
nor U49929 (N_49929,N_32516,N_32713);
and U49930 (N_49930,N_32398,N_30015);
or U49931 (N_49931,N_34474,N_31827);
or U49932 (N_49932,N_34061,N_34193);
or U49933 (N_49933,N_33217,N_30419);
nand U49934 (N_49934,N_39021,N_38382);
and U49935 (N_49935,N_35561,N_39881);
nor U49936 (N_49936,N_33547,N_33261);
and U49937 (N_49937,N_31269,N_39246);
nor U49938 (N_49938,N_30314,N_37843);
xnor U49939 (N_49939,N_32176,N_33422);
or U49940 (N_49940,N_36915,N_38094);
nor U49941 (N_49941,N_33128,N_34177);
nor U49942 (N_49942,N_36258,N_30660);
xnor U49943 (N_49943,N_38985,N_30769);
or U49944 (N_49944,N_36863,N_35399);
or U49945 (N_49945,N_36722,N_34120);
and U49946 (N_49946,N_33347,N_32001);
nor U49947 (N_49947,N_33759,N_30176);
or U49948 (N_49948,N_33341,N_32030);
and U49949 (N_49949,N_35926,N_36919);
nor U49950 (N_49950,N_38252,N_35538);
nand U49951 (N_49951,N_31564,N_37684);
and U49952 (N_49952,N_36767,N_30094);
or U49953 (N_49953,N_37689,N_35264);
nor U49954 (N_49954,N_35984,N_33855);
and U49955 (N_49955,N_32041,N_31751);
and U49956 (N_49956,N_37923,N_36528);
or U49957 (N_49957,N_39121,N_32333);
and U49958 (N_49958,N_30109,N_33413);
and U49959 (N_49959,N_32213,N_34158);
nor U49960 (N_49960,N_30630,N_39542);
xor U49961 (N_49961,N_30786,N_38995);
or U49962 (N_49962,N_34030,N_39818);
and U49963 (N_49963,N_34504,N_30621);
nor U49964 (N_49964,N_35615,N_36547);
or U49965 (N_49965,N_32045,N_34994);
and U49966 (N_49966,N_32417,N_39638);
and U49967 (N_49967,N_37573,N_32074);
and U49968 (N_49968,N_39156,N_36724);
nor U49969 (N_49969,N_39084,N_34969);
and U49970 (N_49970,N_33195,N_39061);
xnor U49971 (N_49971,N_38081,N_35803);
nor U49972 (N_49972,N_39013,N_37102);
nand U49973 (N_49973,N_38941,N_34534);
xor U49974 (N_49974,N_36555,N_30744);
nand U49975 (N_49975,N_35608,N_36710);
nor U49976 (N_49976,N_31984,N_30680);
or U49977 (N_49977,N_34430,N_30762);
nor U49978 (N_49978,N_39181,N_39884);
nand U49979 (N_49979,N_39840,N_34243);
and U49980 (N_49980,N_34111,N_36376);
and U49981 (N_49981,N_33967,N_32212);
xor U49982 (N_49982,N_35529,N_34918);
and U49983 (N_49983,N_36986,N_36509);
xor U49984 (N_49984,N_31298,N_34117);
nor U49985 (N_49985,N_32616,N_35902);
or U49986 (N_49986,N_32492,N_36441);
or U49987 (N_49987,N_36636,N_38044);
xnor U49988 (N_49988,N_32962,N_35689);
or U49989 (N_49989,N_38895,N_37713);
and U49990 (N_49990,N_35203,N_37409);
nand U49991 (N_49991,N_32945,N_38000);
nor U49992 (N_49992,N_32733,N_34353);
or U49993 (N_49993,N_33897,N_39640);
nor U49994 (N_49994,N_32615,N_39414);
nand U49995 (N_49995,N_34723,N_35355);
or U49996 (N_49996,N_31977,N_35687);
and U49997 (N_49997,N_37163,N_38168);
nand U49998 (N_49998,N_34874,N_31030);
xnor U49999 (N_49999,N_32516,N_35675);
or UO_0 (O_0,N_42380,N_42939);
nand UO_1 (O_1,N_48567,N_49426);
and UO_2 (O_2,N_44049,N_45369);
or UO_3 (O_3,N_46745,N_43027);
and UO_4 (O_4,N_43742,N_40909);
xnor UO_5 (O_5,N_47984,N_41703);
nor UO_6 (O_6,N_46155,N_48647);
and UO_7 (O_7,N_47427,N_47360);
or UO_8 (O_8,N_46975,N_42463);
nor UO_9 (O_9,N_40875,N_45840);
or UO_10 (O_10,N_49210,N_41353);
xnor UO_11 (O_11,N_43262,N_48862);
or UO_12 (O_12,N_47246,N_46293);
xnor UO_13 (O_13,N_44123,N_40734);
or UO_14 (O_14,N_43031,N_42815);
nor UO_15 (O_15,N_41616,N_43875);
or UO_16 (O_16,N_48933,N_49552);
nor UO_17 (O_17,N_48217,N_49508);
nand UO_18 (O_18,N_41959,N_41964);
nand UO_19 (O_19,N_48074,N_45480);
or UO_20 (O_20,N_46238,N_40673);
nor UO_21 (O_21,N_45180,N_42529);
xor UO_22 (O_22,N_45416,N_46043);
nand UO_23 (O_23,N_42956,N_48974);
and UO_24 (O_24,N_43663,N_48125);
and UO_25 (O_25,N_42114,N_46270);
nand UO_26 (O_26,N_46440,N_41183);
nand UO_27 (O_27,N_44252,N_48696);
nand UO_28 (O_28,N_49966,N_41386);
nand UO_29 (O_29,N_44198,N_44546);
or UO_30 (O_30,N_47341,N_44143);
or UO_31 (O_31,N_40610,N_46590);
nor UO_32 (O_32,N_43273,N_40419);
nand UO_33 (O_33,N_41016,N_45805);
nor UO_34 (O_34,N_46256,N_40376);
nor UO_35 (O_35,N_48656,N_41018);
and UO_36 (O_36,N_49217,N_47198);
nand UO_37 (O_37,N_49884,N_45919);
and UO_38 (O_38,N_46338,N_49303);
and UO_39 (O_39,N_46508,N_42216);
nand UO_40 (O_40,N_45932,N_42084);
nor UO_41 (O_41,N_40936,N_45496);
and UO_42 (O_42,N_42474,N_46767);
and UO_43 (O_43,N_48912,N_40753);
and UO_44 (O_44,N_44615,N_48820);
nor UO_45 (O_45,N_43548,N_45136);
nand UO_46 (O_46,N_42763,N_47499);
xnor UO_47 (O_47,N_44483,N_49047);
and UO_48 (O_48,N_44011,N_42963);
xnor UO_49 (O_49,N_47437,N_47339);
nand UO_50 (O_50,N_44171,N_41865);
or UO_51 (O_51,N_43820,N_46237);
and UO_52 (O_52,N_43084,N_48456);
nand UO_53 (O_53,N_49161,N_45109);
nor UO_54 (O_54,N_45551,N_48192);
xnor UO_55 (O_55,N_47089,N_42108);
or UO_56 (O_56,N_40067,N_45084);
nor UO_57 (O_57,N_47058,N_41645);
or UO_58 (O_58,N_40732,N_43142);
and UO_59 (O_59,N_47564,N_46273);
and UO_60 (O_60,N_49469,N_42879);
and UO_61 (O_61,N_43796,N_49227);
and UO_62 (O_62,N_44758,N_41780);
xor UO_63 (O_63,N_44312,N_44187);
or UO_64 (O_64,N_42133,N_40184);
and UO_65 (O_65,N_42777,N_41818);
xor UO_66 (O_66,N_43741,N_40560);
xor UO_67 (O_67,N_40629,N_42661);
nor UO_68 (O_68,N_40624,N_45568);
xnor UO_69 (O_69,N_47624,N_45954);
nand UO_70 (O_70,N_43572,N_46481);
nand UO_71 (O_71,N_44807,N_41311);
nand UO_72 (O_72,N_49898,N_48551);
or UO_73 (O_73,N_40090,N_41144);
and UO_74 (O_74,N_46373,N_43402);
nand UO_75 (O_75,N_45926,N_43994);
and UO_76 (O_76,N_47962,N_48495);
xor UO_77 (O_77,N_47705,N_40145);
nor UO_78 (O_78,N_43594,N_42030);
xnor UO_79 (O_79,N_40522,N_48538);
nand UO_80 (O_80,N_45029,N_41702);
nor UO_81 (O_81,N_42220,N_45090);
nor UO_82 (O_82,N_41833,N_40821);
or UO_83 (O_83,N_45765,N_44728);
and UO_84 (O_84,N_48597,N_42495);
or UO_85 (O_85,N_47155,N_49954);
nor UO_86 (O_86,N_48154,N_47830);
nand UO_87 (O_87,N_48478,N_46396);
nor UO_88 (O_88,N_42425,N_45392);
or UO_89 (O_89,N_40994,N_47486);
and UO_90 (O_90,N_48208,N_42271);
nand UO_91 (O_91,N_47207,N_44401);
and UO_92 (O_92,N_47033,N_44754);
nand UO_93 (O_93,N_40105,N_46452);
nor UO_94 (O_94,N_43393,N_42910);
and UO_95 (O_95,N_40437,N_43394);
nand UO_96 (O_96,N_48520,N_49211);
nor UO_97 (O_97,N_49914,N_47225);
and UO_98 (O_98,N_49710,N_45096);
or UO_99 (O_99,N_44033,N_46777);
nand UO_100 (O_100,N_42979,N_40187);
nor UO_101 (O_101,N_43154,N_45962);
nand UO_102 (O_102,N_44492,N_49176);
and UO_103 (O_103,N_41003,N_43133);
nor UO_104 (O_104,N_47647,N_49031);
or UO_105 (O_105,N_48831,N_46902);
nand UO_106 (O_106,N_48642,N_47684);
or UO_107 (O_107,N_40160,N_43264);
and UO_108 (O_108,N_47036,N_47555);
nand UO_109 (O_109,N_40772,N_46500);
and UO_110 (O_110,N_40574,N_49216);
or UO_111 (O_111,N_41303,N_47409);
and UO_112 (O_112,N_44950,N_40243);
and UO_113 (O_113,N_41807,N_41285);
or UO_114 (O_114,N_45708,N_45667);
xnor UO_115 (O_115,N_42081,N_43693);
and UO_116 (O_116,N_49802,N_43595);
nor UO_117 (O_117,N_46750,N_47854);
xor UO_118 (O_118,N_42546,N_40873);
nand UO_119 (O_119,N_40444,N_40965);
nor UO_120 (O_120,N_46161,N_43275);
nor UO_121 (O_121,N_49281,N_47343);
or UO_122 (O_122,N_49196,N_46300);
nand UO_123 (O_123,N_49055,N_40702);
or UO_124 (O_124,N_40967,N_40795);
nor UO_125 (O_125,N_49475,N_44451);
nor UO_126 (O_126,N_47773,N_45344);
and UO_127 (O_127,N_44679,N_48124);
nor UO_128 (O_128,N_41592,N_47590);
nor UO_129 (O_129,N_49715,N_48499);
nor UO_130 (O_130,N_46025,N_44172);
or UO_131 (O_131,N_42078,N_44732);
nand UO_132 (O_132,N_49647,N_43202);
and UO_133 (O_133,N_45356,N_43854);
xnor UO_134 (O_134,N_43819,N_46790);
xor UO_135 (O_135,N_49910,N_42427);
or UO_136 (O_136,N_44605,N_46067);
xor UO_137 (O_137,N_44381,N_46091);
nand UO_138 (O_138,N_47806,N_49698);
nor UO_139 (O_139,N_40670,N_40338);
and UO_140 (O_140,N_42395,N_40694);
nand UO_141 (O_141,N_41613,N_42276);
nor UO_142 (O_142,N_43690,N_49493);
nor UO_143 (O_143,N_44391,N_41727);
nor UO_144 (O_144,N_46261,N_44870);
nand UO_145 (O_145,N_47826,N_45968);
or UO_146 (O_146,N_40023,N_47132);
or UO_147 (O_147,N_45066,N_43459);
or UO_148 (O_148,N_41165,N_43258);
nor UO_149 (O_149,N_41894,N_47292);
and UO_150 (O_150,N_49976,N_49583);
nand UO_151 (O_151,N_46847,N_41086);
nor UO_152 (O_152,N_46857,N_41880);
nor UO_153 (O_153,N_41571,N_45106);
nand UO_154 (O_154,N_40827,N_47235);
or UO_155 (O_155,N_47559,N_41141);
nor UO_156 (O_156,N_44278,N_47012);
nor UO_157 (O_157,N_43589,N_47181);
or UO_158 (O_158,N_46395,N_48368);
nor UO_159 (O_159,N_47189,N_44894);
or UO_160 (O_160,N_45536,N_49120);
xor UO_161 (O_161,N_46428,N_41939);
xor UO_162 (O_162,N_42522,N_41428);
and UO_163 (O_163,N_49347,N_49791);
and UO_164 (O_164,N_46220,N_42695);
nor UO_165 (O_165,N_43059,N_48754);
or UO_166 (O_166,N_41798,N_49795);
and UO_167 (O_167,N_47999,N_44439);
nand UO_168 (O_168,N_43921,N_46687);
xor UO_169 (O_169,N_43051,N_45347);
nor UO_170 (O_170,N_44181,N_45266);
nor UO_171 (O_171,N_49341,N_40495);
and UO_172 (O_172,N_46712,N_46641);
or UO_173 (O_173,N_42420,N_48510);
and UO_174 (O_174,N_43998,N_47395);
or UO_175 (O_175,N_48859,N_49456);
and UO_176 (O_176,N_43178,N_48362);
nand UO_177 (O_177,N_41387,N_44408);
xor UO_178 (O_178,N_40575,N_41301);
nand UO_179 (O_179,N_44458,N_43032);
xor UO_180 (O_180,N_42561,N_45380);
and UO_181 (O_181,N_46927,N_42547);
or UO_182 (O_182,N_47160,N_49402);
or UO_183 (O_183,N_49010,N_45905);
nor UO_184 (O_184,N_47669,N_40234);
nor UO_185 (O_185,N_43138,N_41279);
nand UO_186 (O_186,N_46855,N_40481);
nor UO_187 (O_187,N_46805,N_43426);
nor UO_188 (O_188,N_44477,N_41815);
or UO_189 (O_189,N_40616,N_43509);
nand UO_190 (O_190,N_46680,N_46168);
or UO_191 (O_191,N_46032,N_44395);
or UO_192 (O_192,N_43917,N_46706);
and UO_193 (O_193,N_40484,N_48320);
nor UO_194 (O_194,N_44529,N_48359);
nand UO_195 (O_195,N_40406,N_46719);
xnor UO_196 (O_196,N_41671,N_42778);
and UO_197 (O_197,N_48643,N_49250);
nand UO_198 (O_198,N_42850,N_45238);
nand UO_199 (O_199,N_47878,N_41034);
nand UO_200 (O_200,N_48190,N_46808);
nand UO_201 (O_201,N_48824,N_46662);
or UO_202 (O_202,N_48562,N_41942);
nor UO_203 (O_203,N_47286,N_48527);
nand UO_204 (O_204,N_40354,N_47986);
and UO_205 (O_205,N_44199,N_45607);
nor UO_206 (O_206,N_49973,N_46118);
and UO_207 (O_207,N_40297,N_47828);
nand UO_208 (O_208,N_45538,N_40845);
and UO_209 (O_209,N_49495,N_40622);
nor UO_210 (O_210,N_43408,N_47776);
nand UO_211 (O_211,N_40810,N_48171);
nor UO_212 (O_212,N_46848,N_49332);
nand UO_213 (O_213,N_46145,N_49145);
and UO_214 (O_214,N_48336,N_41364);
nor UO_215 (O_215,N_41922,N_45047);
or UO_216 (O_216,N_46498,N_43360);
nand UO_217 (O_217,N_42229,N_44032);
nor UO_218 (O_218,N_44229,N_49205);
nor UO_219 (O_219,N_49713,N_42486);
or UO_220 (O_220,N_44261,N_45375);
or UO_221 (O_221,N_46289,N_45437);
and UO_222 (O_222,N_41973,N_48429);
or UO_223 (O_223,N_48428,N_47903);
nand UO_224 (O_224,N_46983,N_43017);
and UO_225 (O_225,N_43267,N_40887);
nor UO_226 (O_226,N_42072,N_41039);
and UO_227 (O_227,N_44518,N_41210);
nor UO_228 (O_228,N_48826,N_44791);
xnor UO_229 (O_229,N_45974,N_41219);
and UO_230 (O_230,N_42239,N_45807);
xnor UO_231 (O_231,N_40508,N_40278);
and UO_232 (O_232,N_49178,N_45717);
or UO_233 (O_233,N_46497,N_48835);
or UO_234 (O_234,N_41581,N_44989);
and UO_235 (O_235,N_42365,N_41770);
nor UO_236 (O_236,N_49126,N_49989);
nor UO_237 (O_237,N_41501,N_41935);
or UO_238 (O_238,N_47600,N_45633);
and UO_239 (O_239,N_46593,N_44760);
nor UO_240 (O_240,N_47754,N_47054);
or UO_241 (O_241,N_49536,N_45918);
or UO_242 (O_242,N_42281,N_40153);
nor UO_243 (O_243,N_42351,N_49461);
and UO_244 (O_244,N_44089,N_42165);
and UO_245 (O_245,N_47118,N_44410);
nand UO_246 (O_246,N_47083,N_49311);
and UO_247 (O_247,N_43941,N_45198);
nor UO_248 (O_248,N_43907,N_49735);
or UO_249 (O_249,N_45652,N_49768);
nor UO_250 (O_250,N_48674,N_48852);
nand UO_251 (O_251,N_44836,N_48945);
nand UO_252 (O_252,N_40775,N_40170);
nor UO_253 (O_253,N_42241,N_47127);
and UO_254 (O_254,N_41468,N_49784);
or UO_255 (O_255,N_42368,N_45020);
nand UO_256 (O_256,N_41845,N_41157);
nor UO_257 (O_257,N_45235,N_47011);
nand UO_258 (O_258,N_45834,N_49357);
nor UO_259 (O_259,N_42137,N_41225);
nand UO_260 (O_260,N_46066,N_45600);
and UO_261 (O_261,N_44079,N_44887);
nand UO_262 (O_262,N_43783,N_48389);
and UO_263 (O_263,N_41600,N_49744);
or UO_264 (O_264,N_44498,N_40139);
nor UO_265 (O_265,N_45202,N_45139);
nor UO_266 (O_266,N_43168,N_45639);
and UO_267 (O_267,N_47656,N_45014);
nor UO_268 (O_268,N_45851,N_45979);
nand UO_269 (O_269,N_42119,N_48247);
nor UO_270 (O_270,N_46909,N_48929);
and UO_271 (O_271,N_44924,N_42525);
nand UO_272 (O_272,N_45604,N_44224);
and UO_273 (O_273,N_44030,N_41675);
xnor UO_274 (O_274,N_46194,N_43828);
or UO_275 (O_275,N_43158,N_47197);
nor UO_276 (O_276,N_45690,N_45646);
or UO_277 (O_277,N_40364,N_43518);
xor UO_278 (O_278,N_41680,N_42617);
nor UO_279 (O_279,N_42584,N_45204);
or UO_280 (O_280,N_47163,N_47631);
nor UO_281 (O_281,N_46501,N_47263);
or UO_282 (O_282,N_42987,N_45352);
nand UO_283 (O_283,N_48166,N_44660);
nand UO_284 (O_284,N_46341,N_42443);
or UO_285 (O_285,N_45439,N_48179);
and UO_286 (O_286,N_48895,N_45177);
xor UO_287 (O_287,N_42378,N_43952);
nand UO_288 (O_288,N_41649,N_44276);
nand UO_289 (O_289,N_45850,N_45613);
nand UO_290 (O_290,N_45371,N_40631);
and UO_291 (O_291,N_43339,N_47652);
or UO_292 (O_292,N_44179,N_45981);
or UO_293 (O_293,N_45809,N_48507);
xor UO_294 (O_294,N_41133,N_43901);
nand UO_295 (O_295,N_47508,N_41902);
nand UO_296 (O_296,N_48480,N_48170);
and UO_297 (O_297,N_41478,N_47980);
xor UO_298 (O_298,N_45476,N_48356);
nand UO_299 (O_299,N_49361,N_43553);
nand UO_300 (O_300,N_48329,N_48786);
nor UO_301 (O_301,N_46477,N_47834);
xnor UO_302 (O_302,N_49248,N_48063);
nand UO_303 (O_303,N_42475,N_46409);
xor UO_304 (O_304,N_42779,N_42382);
nand UO_305 (O_305,N_45944,N_40615);
and UO_306 (O_306,N_47412,N_49068);
and UO_307 (O_307,N_41456,N_41374);
nand UO_308 (O_308,N_45363,N_40202);
and UO_309 (O_309,N_46153,N_46647);
xor UO_310 (O_310,N_42934,N_43809);
and UO_311 (O_311,N_48689,N_44644);
nor UO_312 (O_312,N_40877,N_47137);
nor UO_313 (O_313,N_46587,N_47825);
and UO_314 (O_314,N_42790,N_48644);
nand UO_315 (O_315,N_41921,N_49353);
or UO_316 (O_316,N_48203,N_41615);
and UO_317 (O_317,N_42549,N_41860);
nand UO_318 (O_318,N_49520,N_47688);
or UO_319 (O_319,N_46491,N_46350);
and UO_320 (O_320,N_45407,N_40547);
and UO_321 (O_321,N_43764,N_41677);
or UO_322 (O_322,N_48901,N_48746);
or UO_323 (O_323,N_41669,N_40712);
or UO_324 (O_324,N_44251,N_48846);
or UO_325 (O_325,N_43358,N_44453);
nor UO_326 (O_326,N_48244,N_44610);
xor UO_327 (O_327,N_44675,N_42406);
nor UO_328 (O_328,N_42265,N_45195);
nor UO_329 (O_329,N_49669,N_46627);
nand UO_330 (O_330,N_46417,N_46512);
nor UO_331 (O_331,N_48012,N_40774);
nand UO_332 (O_332,N_43855,N_41074);
xor UO_333 (O_333,N_47406,N_40523);
nand UO_334 (O_334,N_42446,N_43460);
nand UO_335 (O_335,N_40533,N_45804);
nor UO_336 (O_336,N_42295,N_47781);
nand UO_337 (O_337,N_43386,N_48013);
or UO_338 (O_338,N_43463,N_44023);
and UO_339 (O_339,N_40796,N_41495);
or UO_340 (O_340,N_44250,N_43420);
or UO_341 (O_341,N_42951,N_45854);
and UO_342 (O_342,N_43385,N_46112);
nor UO_343 (O_343,N_42997,N_45355);
nand UO_344 (O_344,N_46208,N_47212);
nand UO_345 (O_345,N_42578,N_41631);
or UO_346 (O_346,N_48789,N_45304);
nor UO_347 (O_347,N_48543,N_46765);
nand UO_348 (O_348,N_47203,N_41442);
nor UO_349 (O_349,N_48361,N_48314);
nor UO_350 (O_350,N_49567,N_48489);
nand UO_351 (O_351,N_47757,N_41608);
and UO_352 (O_352,N_46158,N_42393);
and UO_353 (O_353,N_47269,N_49575);
xor UO_354 (O_354,N_44690,N_40907);
nor UO_355 (O_355,N_42319,N_44722);
and UO_356 (O_356,N_47604,N_48873);
nand UO_357 (O_357,N_43419,N_42678);
nor UO_358 (O_358,N_41232,N_47226);
and UO_359 (O_359,N_44674,N_40480);
nor UO_360 (O_360,N_40841,N_45389);
nor UO_361 (O_361,N_49832,N_43269);
and UO_362 (O_362,N_41812,N_47112);
or UO_363 (O_363,N_43771,N_44471);
or UO_364 (O_364,N_41842,N_41890);
or UO_365 (O_365,N_46223,N_43644);
and UO_366 (O_366,N_49002,N_41978);
xor UO_367 (O_367,N_42297,N_47231);
nor UO_368 (O_368,N_42776,N_46252);
nand UO_369 (O_369,N_45626,N_49220);
or UO_370 (O_370,N_45822,N_46799);
and UO_371 (O_371,N_40687,N_46316);
nand UO_372 (O_372,N_43152,N_46495);
and UO_373 (O_373,N_44954,N_42655);
or UO_374 (O_374,N_44371,N_41981);
or UO_375 (O_375,N_49501,N_41548);
nand UO_376 (O_376,N_49027,N_43316);
nor UO_377 (O_377,N_47432,N_47971);
nor UO_378 (O_378,N_40749,N_49035);
or UO_379 (O_379,N_42189,N_44227);
and UO_380 (O_380,N_43612,N_48875);
or UO_381 (O_381,N_41874,N_48571);
nor UO_382 (O_382,N_49607,N_47446);
or UO_383 (O_383,N_45346,N_40174);
and UO_384 (O_384,N_48781,N_44621);
or UO_385 (O_385,N_44648,N_48164);
nand UO_386 (O_386,N_49075,N_48467);
or UO_387 (O_387,N_49807,N_44053);
nand UO_388 (O_388,N_44988,N_46020);
nor UO_389 (O_389,N_48686,N_42709);
nand UO_390 (O_390,N_48815,N_48816);
and UO_391 (O_391,N_44632,N_41660);
or UO_392 (O_392,N_42723,N_48558);
nand UO_393 (O_393,N_49844,N_47420);
or UO_394 (O_394,N_43411,N_48632);
nor UO_395 (O_395,N_46478,N_42006);
xor UO_396 (O_396,N_49690,N_45887);
or UO_397 (O_397,N_45008,N_40498);
or UO_398 (O_398,N_48313,N_40422);
nor UO_399 (O_399,N_49252,N_44963);
or UO_400 (O_400,N_42478,N_49565);
and UO_401 (O_401,N_41469,N_40564);
and UO_402 (O_402,N_40445,N_45296);
or UO_403 (O_403,N_48959,N_41075);
xnor UO_404 (O_404,N_46663,N_41797);
nor UO_405 (O_405,N_49907,N_48080);
nand UO_406 (O_406,N_40750,N_48157);
or UO_407 (O_407,N_48800,N_46071);
and UO_408 (O_408,N_43815,N_45628);
xnor UO_409 (O_409,N_49457,N_48923);
nor UO_410 (O_410,N_41603,N_45274);
nand UO_411 (O_411,N_46146,N_47362);
xor UO_412 (O_412,N_42759,N_49112);
xor UO_413 (O_413,N_48505,N_40960);
and UO_414 (O_414,N_41828,N_49429);
nor UO_415 (O_415,N_43655,N_46311);
xnor UO_416 (O_416,N_47029,N_44971);
nand UO_417 (O_417,N_44406,N_45171);
nand UO_418 (O_418,N_46258,N_47314);
and UO_419 (O_419,N_48617,N_40843);
nand UO_420 (O_420,N_47936,N_49694);
nand UO_421 (O_421,N_43638,N_46424);
nor UO_422 (O_422,N_43222,N_41763);
and UO_423 (O_423,N_48782,N_45327);
xnor UO_424 (O_424,N_41782,N_42038);
and UO_425 (O_425,N_44488,N_43097);
nor UO_426 (O_426,N_45410,N_49162);
or UO_427 (O_427,N_48328,N_45669);
or UO_428 (O_428,N_47535,N_45243);
and UO_429 (O_429,N_46450,N_41861);
nand UO_430 (O_430,N_47037,N_41796);
nand UO_431 (O_431,N_43148,N_43825);
nand UO_432 (O_432,N_40016,N_42955);
nor UO_433 (O_433,N_40721,N_46953);
or UO_434 (O_434,N_49854,N_45806);
nand UO_435 (O_435,N_43469,N_46901);
and UO_436 (O_436,N_42774,N_45126);
and UO_437 (O_437,N_43713,N_48107);
and UO_438 (O_438,N_41775,N_48196);
and UO_439 (O_439,N_45566,N_44098);
nor UO_440 (O_440,N_49174,N_43444);
nor UO_441 (O_441,N_48834,N_47227);
and UO_442 (O_442,N_40627,N_42719);
nand UO_443 (O_443,N_45693,N_42052);
and UO_444 (O_444,N_45435,N_41586);
nor UO_445 (O_445,N_44910,N_47682);
or UO_446 (O_446,N_43060,N_44581);
nor UO_447 (O_447,N_43403,N_48837);
nor UO_448 (O_448,N_40066,N_41424);
and UO_449 (O_449,N_41988,N_49719);
nor UO_450 (O_450,N_46462,N_43132);
or UO_451 (O_451,N_44221,N_45398);
nor UO_452 (O_452,N_43192,N_42316);
or UO_453 (O_453,N_44829,N_45577);
and UO_454 (O_454,N_42911,N_49249);
nand UO_455 (O_455,N_45452,N_40193);
nand UO_456 (O_456,N_46057,N_45993);
or UO_457 (O_457,N_41834,N_48370);
nor UO_458 (O_458,N_43942,N_43197);
nand UO_459 (O_459,N_41244,N_43954);
or UO_460 (O_460,N_46921,N_47172);
or UO_461 (O_461,N_40691,N_45221);
nor UO_462 (O_462,N_41102,N_45741);
or UO_463 (O_463,N_40349,N_43581);
and UO_464 (O_464,N_44263,N_42410);
nand UO_465 (O_465,N_41674,N_48713);
nor UO_466 (O_466,N_41111,N_46367);
and UO_467 (O_467,N_49298,N_44995);
and UO_468 (O_468,N_42277,N_49280);
nand UO_469 (O_469,N_45419,N_43407);
and UO_470 (O_470,N_48084,N_47312);
nand UO_471 (O_471,N_41863,N_45225);
nand UO_472 (O_472,N_48832,N_40018);
xor UO_473 (O_473,N_41646,N_41593);
and UO_474 (O_474,N_45283,N_40428);
or UO_475 (O_475,N_47009,N_42880);
nor UO_476 (O_476,N_44268,N_41426);
nor UO_477 (O_477,N_46014,N_47790);
nor UO_478 (O_478,N_46055,N_47620);
nand UO_479 (O_479,N_49494,N_40925);
nor UO_480 (O_480,N_45220,N_48606);
nand UO_481 (O_481,N_46916,N_40356);
nor UO_482 (O_482,N_42208,N_49411);
nand UO_483 (O_483,N_42002,N_47018);
nor UO_484 (O_484,N_49776,N_45616);
or UO_485 (O_485,N_45552,N_41378);
and UO_486 (O_486,N_49105,N_42353);
nand UO_487 (O_487,N_49093,N_48673);
and UO_488 (O_488,N_43867,N_43353);
nor UO_489 (O_489,N_42775,N_43786);
or UO_490 (O_490,N_40207,N_43226);
and UO_491 (O_491,N_44375,N_44780);
nand UO_492 (O_492,N_43071,N_46693);
nor UO_493 (O_493,N_45839,N_42315);
nor UO_494 (O_494,N_45390,N_45555);
or UO_495 (O_495,N_47487,N_46290);
or UO_496 (O_496,N_49579,N_45168);
xor UO_497 (O_497,N_43272,N_46410);
nand UO_498 (O_498,N_44222,N_46127);
or UO_499 (O_499,N_45027,N_42913);
xor UO_500 (O_500,N_49337,N_48349);
nand UO_501 (O_501,N_49645,N_41015);
nand UO_502 (O_502,N_48075,N_43255);
or UO_503 (O_503,N_46271,N_42235);
nor UO_504 (O_504,N_45543,N_41135);
nand UO_505 (O_505,N_47328,N_47618);
and UO_506 (O_506,N_44782,N_44638);
or UO_507 (O_507,N_46580,N_43800);
and UO_508 (O_508,N_47094,N_48133);
nor UO_509 (O_509,N_40520,N_46147);
and UO_510 (O_510,N_42825,N_46733);
nand UO_511 (O_511,N_44151,N_43897);
xor UO_512 (O_512,N_43150,N_46700);
nand UO_513 (O_513,N_46298,N_46439);
and UO_514 (O_514,N_42715,N_47043);
nor UO_515 (O_515,N_48939,N_40502);
nand UO_516 (O_516,N_41622,N_41350);
nand UO_517 (O_517,N_44220,N_44326);
nand UO_518 (O_518,N_41661,N_42817);
xnor UO_519 (O_519,N_49521,N_45559);
nand UO_520 (O_520,N_47295,N_44243);
nand UO_521 (O_521,N_45780,N_49338);
nor UO_522 (O_522,N_43038,N_47431);
nor UO_523 (O_523,N_42550,N_45963);
and UO_524 (O_524,N_43557,N_46074);
xnor UO_525 (O_525,N_41897,N_49870);
and UO_526 (O_526,N_49608,N_46454);
nor UO_527 (O_527,N_46636,N_44163);
or UO_528 (O_528,N_48321,N_46374);
and UO_529 (O_529,N_48081,N_40307);
nand UO_530 (O_530,N_46917,N_45069);
nand UO_531 (O_531,N_49225,N_44486);
nand UO_532 (O_532,N_45362,N_44456);
and UO_533 (O_533,N_42167,N_47002);
or UO_534 (O_534,N_46747,N_42482);
nor UO_535 (O_535,N_49177,N_40779);
nor UO_536 (O_536,N_45192,N_42656);
and UO_537 (O_537,N_40743,N_43758);
nand UO_538 (O_538,N_41938,N_41314);
nor UO_539 (O_539,N_44866,N_49664);
and UO_540 (O_540,N_47958,N_48736);
nor UO_541 (O_541,N_49169,N_40300);
xnor UO_542 (O_542,N_48770,N_48760);
or UO_543 (O_543,N_49388,N_41151);
or UO_544 (O_544,N_42557,N_47305);
and UO_545 (O_545,N_44819,N_48180);
and UO_546 (O_546,N_44811,N_44515);
nor UO_547 (O_547,N_42632,N_47567);
nand UO_548 (O_548,N_44235,N_49066);
and UO_549 (O_549,N_45964,N_40555);
xor UO_550 (O_550,N_44154,N_44478);
and UO_551 (O_551,N_47115,N_40390);
nor UO_552 (O_552,N_46758,N_42519);
nand UO_553 (O_553,N_49449,N_46292);
nor UO_554 (O_554,N_47281,N_40776);
nand UO_555 (O_555,N_48682,N_47007);
nor UO_556 (O_556,N_44082,N_43153);
nor UO_557 (O_557,N_41373,N_42390);
and UO_558 (O_558,N_46685,N_43956);
nand UO_559 (O_559,N_41968,N_43030);
xnor UO_560 (O_560,N_47642,N_46039);
and UO_561 (O_561,N_46376,N_44715);
or UO_562 (O_562,N_44302,N_49228);
and UO_563 (O_563,N_41835,N_49135);
nor UO_564 (O_564,N_48324,N_47883);
or UO_565 (O_565,N_40259,N_40602);
or UO_566 (O_566,N_48739,N_46570);
and UO_567 (O_567,N_43043,N_42197);
nand UO_568 (O_568,N_48550,N_42718);
nor UO_569 (O_569,N_41509,N_49692);
or UO_570 (O_570,N_42730,N_45461);
or UO_571 (O_571,N_49840,N_46553);
xor UO_572 (O_572,N_42364,N_42140);
nand UO_573 (O_573,N_47498,N_41492);
xor UO_574 (O_574,N_44568,N_49492);
nand UO_575 (O_575,N_42240,N_44986);
xnor UO_576 (O_576,N_44669,N_46726);
nand UO_577 (O_577,N_47939,N_43253);
or UO_578 (O_578,N_46274,N_42083);
nand UO_579 (O_579,N_49741,N_44232);
and UO_580 (O_580,N_46965,N_48535);
or UO_581 (O_581,N_47477,N_41092);
nand UO_582 (O_582,N_48791,N_49464);
nand UO_583 (O_583,N_45294,N_42049);
or UO_584 (O_584,N_48762,N_42574);
nor UO_585 (O_585,N_40138,N_40266);
and UO_586 (O_586,N_41920,N_48511);
nor UO_587 (O_587,N_49371,N_46937);
nor UO_588 (O_588,N_46922,N_48657);
and UO_589 (O_589,N_43996,N_41830);
nand UO_590 (O_590,N_42325,N_48172);
nor UO_591 (O_591,N_44781,N_44024);
nor UO_592 (O_592,N_47119,N_45895);
xor UO_593 (O_593,N_41783,N_40131);
nor UO_594 (O_594,N_46761,N_43863);
or UO_595 (O_595,N_42448,N_48973);
nand UO_596 (O_596,N_43837,N_45128);
and UO_597 (O_597,N_49283,N_45697);
nor UO_598 (O_598,N_48430,N_42492);
nor UO_599 (O_599,N_42321,N_47074);
and UO_600 (O_600,N_47660,N_40137);
nand UO_601 (O_601,N_48009,N_47404);
or UO_602 (O_602,N_47614,N_42826);
or UO_603 (O_603,N_46048,N_47324);
or UO_604 (O_604,N_41717,N_48473);
nor UO_605 (O_605,N_41460,N_49825);
xnor UO_606 (O_606,N_41427,N_44670);
or UO_607 (O_607,N_48195,N_47670);
nor UO_608 (O_608,N_49486,N_49133);
and UO_609 (O_609,N_44919,N_44572);
and UO_610 (O_610,N_48002,N_40835);
nor UO_611 (O_611,N_41741,N_48156);
and UO_612 (O_612,N_43035,N_47873);
and UO_613 (O_613,N_41766,N_48741);
nor UO_614 (O_614,N_46612,N_40014);
nand UO_615 (O_615,N_45466,N_45070);
nor UO_616 (O_616,N_42717,N_42476);
nand UO_617 (O_617,N_47460,N_43821);
xnor UO_618 (O_618,N_43895,N_47373);
or UO_619 (O_619,N_47177,N_49515);
or UO_620 (O_620,N_47640,N_47838);
nor UO_621 (O_621,N_40370,N_42021);
nand UO_622 (O_622,N_43946,N_42286);
or UO_623 (O_623,N_47174,N_47028);
or UO_624 (O_624,N_45892,N_44752);
nor UO_625 (O_625,N_46502,N_42349);
xor UO_626 (O_626,N_43686,N_43932);
nor UO_627 (O_627,N_44176,N_41246);
and UO_628 (O_628,N_47753,N_45024);
or UO_629 (O_629,N_43458,N_43209);
or UO_630 (O_630,N_40728,N_45773);
and UO_631 (O_631,N_40189,N_47617);
nor UO_632 (O_632,N_46277,N_46725);
nand UO_633 (O_633,N_48141,N_48677);
or UO_634 (O_634,N_49241,N_48386);
and UO_635 (O_635,N_49095,N_43291);
and UO_636 (O_636,N_48981,N_40769);
nand UO_637 (O_637,N_40968,N_40217);
or UO_638 (O_638,N_40975,N_45351);
and UO_639 (O_639,N_44128,N_41691);
nor UO_640 (O_640,N_45510,N_49782);
and UO_641 (O_641,N_47287,N_43603);
and UO_642 (O_642,N_44569,N_40630);
xor UO_643 (O_643,N_40915,N_44380);
or UO_644 (O_644,N_48792,N_42401);
or UO_645 (O_645,N_47441,N_45517);
or UO_646 (O_646,N_40597,N_45876);
nand UO_647 (O_647,N_48825,N_43338);
nor UO_648 (O_648,N_47357,N_45808);
nor UO_649 (O_649,N_41223,N_40948);
nor UO_650 (O_650,N_43004,N_43474);
and UO_651 (O_651,N_41021,N_41068);
or UO_652 (O_652,N_40336,N_41673);
and UO_653 (O_653,N_46272,N_43293);
or UO_654 (O_654,N_48201,N_41987);
xnor UO_655 (O_655,N_46442,N_49476);
nor UO_656 (O_656,N_40468,N_40250);
or UO_657 (O_657,N_45323,N_41853);
nand UO_658 (O_658,N_45370,N_41925);
nand UO_659 (O_659,N_47200,N_40452);
or UO_660 (O_660,N_42441,N_40707);
or UO_661 (O_661,N_41330,N_49394);
and UO_662 (O_662,N_42346,N_49650);
nor UO_663 (O_663,N_43963,N_40716);
or UO_664 (O_664,N_47955,N_46667);
nor UO_665 (O_665,N_42128,N_42658);
nand UO_666 (O_666,N_47022,N_44551);
or UO_667 (O_667,N_45771,N_45978);
nand UO_668 (O_668,N_47008,N_41536);
nor UO_669 (O_669,N_43743,N_43120);
and UO_670 (O_670,N_45700,N_48054);
nand UO_671 (O_671,N_41278,N_42702);
nor UO_672 (O_672,N_45300,N_42821);
and UO_673 (O_673,N_41192,N_43040);
or UO_674 (O_674,N_49004,N_40270);
nor UO_675 (O_675,N_45845,N_45455);
and UO_676 (O_676,N_45411,N_49599);
nor UO_677 (O_677,N_40692,N_41816);
and UO_678 (O_678,N_46468,N_45713);
or UO_679 (O_679,N_46562,N_43427);
nand UO_680 (O_680,N_49305,N_42568);
nor UO_681 (O_681,N_49224,N_42577);
nor UO_682 (O_682,N_47003,N_42231);
and UO_683 (O_683,N_40335,N_49988);
xor UO_684 (O_684,N_41899,N_42185);
or UO_685 (O_685,N_41936,N_45431);
nor UO_686 (O_686,N_47731,N_44856);
nor UO_687 (O_687,N_44206,N_48580);
and UO_688 (O_688,N_46392,N_42660);
and UO_689 (O_689,N_43528,N_47976);
nor UO_690 (O_690,N_43781,N_48425);
nor UO_691 (O_691,N_43072,N_42690);
and UO_692 (O_692,N_41665,N_49355);
nand UO_693 (O_693,N_43566,N_42263);
and UO_694 (O_694,N_43696,N_48263);
or UO_695 (O_695,N_44597,N_41785);
and UO_696 (O_696,N_40046,N_47667);
nand UO_697 (O_697,N_46757,N_41802);
or UO_698 (O_698,N_40544,N_43928);
nor UO_699 (O_699,N_48759,N_44764);
nor UO_700 (O_700,N_47388,N_48024);
nor UO_701 (O_701,N_40087,N_45540);
xnor UO_702 (O_702,N_49287,N_45190);
or UO_703 (O_703,N_42835,N_47595);
or UO_704 (O_704,N_40304,N_41035);
nor UO_705 (O_705,N_46132,N_47923);
or UO_706 (O_706,N_46156,N_43111);
or UO_707 (O_707,N_42290,N_46370);
nor UO_708 (O_708,N_44443,N_47717);
nand UO_709 (O_709,N_49505,N_41559);
and UO_710 (O_710,N_49991,N_44394);
nor UO_711 (O_711,N_43962,N_40007);
or UO_712 (O_712,N_49172,N_41042);
nor UO_713 (O_713,N_47998,N_48943);
and UO_714 (O_714,N_49945,N_49566);
nand UO_715 (O_715,N_40147,N_46475);
and UO_716 (O_716,N_41367,N_44992);
and UO_717 (O_717,N_44591,N_46538);
nand UO_718 (O_718,N_47538,N_49693);
or UO_719 (O_719,N_40123,N_48145);
nand UO_720 (O_720,N_41821,N_48864);
nand UO_721 (O_721,N_40181,N_42404);
and UO_722 (O_722,N_41462,N_43960);
and UO_723 (O_723,N_40279,N_43090);
nor UO_724 (O_724,N_49580,N_44685);
or UO_725 (O_725,N_47194,N_40874);
or UO_726 (O_726,N_40085,N_48604);
and UO_727 (O_727,N_49632,N_49522);
nor UO_728 (O_728,N_47741,N_49401);
nand UO_729 (O_729,N_42771,N_46383);
nand UO_730 (O_730,N_46385,N_40267);
nand UO_731 (O_731,N_48518,N_48611);
nand UO_732 (O_732,N_41013,N_42092);
nor UO_733 (O_733,N_44810,N_46697);
nor UO_734 (O_734,N_45801,N_42536);
nor UO_735 (O_735,N_45367,N_40075);
and UO_736 (O_736,N_40177,N_46876);
nand UO_737 (O_737,N_46264,N_44305);
nand UO_738 (O_738,N_44000,N_49413);
nor UO_739 (O_739,N_40314,N_44502);
and UO_740 (O_740,N_49187,N_45869);
nand UO_741 (O_741,N_44667,N_40321);
or UO_742 (O_742,N_48587,N_42169);
or UO_743 (O_743,N_47952,N_47641);
and UO_744 (O_744,N_44666,N_48576);
and UO_745 (O_745,N_45870,N_49555);
and UO_746 (O_746,N_41728,N_42885);
nand UO_747 (O_747,N_43343,N_48339);
or UO_748 (O_748,N_40558,N_40666);
or UO_749 (O_749,N_44871,N_41610);
nor UO_750 (O_750,N_48049,N_49670);
and UO_751 (O_751,N_43347,N_47644);
nand UO_752 (O_752,N_49705,N_47361);
nor UO_753 (O_753,N_41927,N_49503);
nor UO_754 (O_754,N_46188,N_41143);
or UO_755 (O_755,N_41479,N_47592);
xnor UO_756 (O_756,N_48162,N_42653);
xnor UO_757 (O_757,N_40609,N_41142);
or UO_758 (O_758,N_40158,N_46851);
and UO_759 (O_759,N_45514,N_44279);
nor UO_760 (O_760,N_43325,N_45092);
nor UO_761 (O_761,N_41377,N_42634);
nor UO_762 (O_762,N_45890,N_44987);
and UO_763 (O_763,N_44822,N_43813);
or UO_764 (O_764,N_43823,N_45306);
xnor UO_765 (O_765,N_48985,N_47734);
and UO_766 (O_766,N_43715,N_45695);
nor UO_767 (O_767,N_47428,N_48836);
nand UO_768 (O_768,N_41576,N_47013);
and UO_769 (O_769,N_41535,N_43337);
nor UO_770 (O_770,N_41422,N_47425);
and UO_771 (O_771,N_41838,N_43480);
and UO_772 (O_772,N_45387,N_47601);
or UO_773 (O_773,N_49767,N_40901);
or UO_774 (O_774,N_43359,N_49707);
nand UO_775 (O_775,N_44343,N_49375);
and UO_776 (O_776,N_41362,N_45681);
xnor UO_777 (O_777,N_49076,N_46554);
xnor UO_778 (O_778,N_46734,N_48986);
or UO_779 (O_779,N_40120,N_44411);
nand UO_780 (O_780,N_45293,N_42958);
or UO_781 (O_781,N_41642,N_41837);
or UO_782 (O_782,N_40253,N_44712);
nor UO_783 (O_783,N_45917,N_47101);
nor UO_784 (O_784,N_47476,N_46138);
nand UO_785 (O_785,N_45038,N_43439);
nand UO_786 (O_786,N_41844,N_46176);
or UO_787 (O_787,N_47308,N_48398);
or UO_788 (O_788,N_43164,N_46509);
nor UO_789 (O_789,N_40474,N_47786);
or UO_790 (O_790,N_40343,N_43634);
and UO_791 (O_791,N_47161,N_40410);
or UO_792 (O_792,N_42429,N_49867);
or UO_793 (O_793,N_48783,N_47398);
xor UO_794 (O_794,N_47243,N_41187);
nand UO_795 (O_795,N_42982,N_47363);
nor UO_796 (O_796,N_47580,N_46720);
nor UO_797 (O_797,N_48549,N_46072);
or UO_798 (O_798,N_43180,N_42819);
and UO_799 (O_799,N_45992,N_40019);
or UO_800 (O_800,N_48325,N_45163);
or UO_801 (O_801,N_46963,N_45430);
or UO_802 (O_802,N_46897,N_49800);
nor UO_803 (O_803,N_41061,N_49638);
and UO_804 (O_804,N_41738,N_47714);
and UO_805 (O_805,N_47451,N_48879);
or UO_806 (O_806,N_47895,N_44170);
and UO_807 (O_807,N_43472,N_41259);
nand UO_808 (O_808,N_41748,N_43128);
and UO_809 (O_809,N_44937,N_47509);
or UO_810 (O_810,N_40487,N_43559);
or UO_811 (O_811,N_49984,N_44281);
nor UO_812 (O_812,N_48501,N_42412);
or UO_813 (O_813,N_41626,N_44364);
or UO_814 (O_814,N_42750,N_46488);
nand UO_815 (O_815,N_46567,N_49318);
nand UO_816 (O_816,N_43574,N_44113);
xnor UO_817 (O_817,N_46211,N_48284);
nand UO_818 (O_818,N_40262,N_44070);
nor UO_819 (O_819,N_49130,N_42969);
and UO_820 (O_820,N_40392,N_48521);
nor UO_821 (O_821,N_47130,N_42729);
nand UO_822 (O_822,N_40990,N_46620);
or UO_823 (O_823,N_48109,N_44109);
and UO_824 (O_824,N_41849,N_43113);
or UO_825 (O_825,N_40519,N_44040);
or UO_826 (O_826,N_43131,N_47823);
nor UO_827 (O_827,N_49736,N_49900);
and UO_828 (O_828,N_45188,N_46024);
or UO_829 (O_829,N_44012,N_47309);
nor UO_830 (O_830,N_46569,N_47400);
or UO_831 (O_831,N_47024,N_44622);
nor UO_832 (O_832,N_42394,N_40509);
or UO_833 (O_833,N_49805,N_46243);
or UO_834 (O_834,N_42339,N_41032);
nand UO_835 (O_835,N_44702,N_43840);
and UO_836 (O_836,N_47915,N_46122);
or UO_837 (O_837,N_41166,N_49820);
and UO_838 (O_838,N_44264,N_41282);
nand UO_839 (O_839,N_41699,N_44628);
and UO_840 (O_840,N_42905,N_49787);
nand UO_841 (O_841,N_46007,N_43521);
nand UO_842 (O_842,N_40911,N_40175);
or UO_843 (O_843,N_48413,N_49339);
and UO_844 (O_844,N_46579,N_43401);
and UO_845 (O_845,N_43471,N_45907);
or UO_846 (O_846,N_43326,N_46416);
and UO_847 (O_847,N_42517,N_42094);
xor UO_848 (O_848,N_49259,N_46840);
nand UO_849 (O_849,N_48322,N_43282);
and UO_850 (O_850,N_46918,N_40108);
and UO_851 (O_851,N_43723,N_43081);
and UO_852 (O_852,N_47778,N_45880);
or UO_853 (O_853,N_40503,N_41886);
or UO_854 (O_854,N_49550,N_49553);
nor UO_855 (O_855,N_44306,N_45742);
and UO_856 (O_856,N_46482,N_41212);
nand UO_857 (O_857,N_44895,N_47702);
or UO_858 (O_858,N_48962,N_43462);
nand UO_859 (O_859,N_41088,N_43248);
and UO_860 (O_860,N_42555,N_49621);
nor UO_861 (O_861,N_41506,N_43047);
nor UO_862 (O_862,N_46728,N_45058);
nor UO_863 (O_863,N_46351,N_47218);
nand UO_864 (O_864,N_47353,N_47598);
nand UO_865 (O_865,N_47569,N_45673);
nor UO_866 (O_866,N_49185,N_44291);
nand UO_867 (O_867,N_48833,N_41087);
nand UO_868 (O_868,N_46459,N_45815);
nand UO_869 (O_869,N_49823,N_41277);
and UO_870 (O_870,N_48136,N_46170);
nand UO_871 (O_871,N_45977,N_49728);
nand UO_872 (O_872,N_49153,N_40870);
nor UO_873 (O_873,N_45000,N_49458);
nor UO_874 (O_874,N_44697,N_48420);
nor UO_875 (O_875,N_48942,N_43641);
nand UO_876 (O_876,N_40413,N_45988);
xnor UO_877 (O_877,N_41900,N_44071);
and UO_878 (O_878,N_48579,N_41575);
and UO_879 (O_879,N_44850,N_46601);
nor UO_880 (O_880,N_46534,N_42122);
and UO_881 (O_881,N_42836,N_40438);
or UO_882 (O_882,N_46988,N_49261);
or UO_883 (O_883,N_47888,N_46204);
or UO_884 (O_884,N_41369,N_41155);
nor UO_885 (O_885,N_47072,N_48984);
and UO_886 (O_886,N_44372,N_46051);
nor UO_887 (O_887,N_48991,N_49761);
or UO_888 (O_888,N_48144,N_44528);
or UO_889 (O_889,N_41708,N_41910);
or UO_890 (O_890,N_49725,N_42136);
and UO_891 (O_891,N_40805,N_42221);
xor UO_892 (O_892,N_44396,N_49641);
nand UO_893 (O_893,N_44861,N_47077);
nor UO_894 (O_894,N_47989,N_47438);
or UO_895 (O_895,N_41119,N_44898);
nand UO_896 (O_896,N_48855,N_48821);
xor UO_897 (O_897,N_48953,N_47851);
and UO_898 (O_898,N_48993,N_44905);
or UO_899 (O_899,N_48462,N_40918);
or UO_900 (O_900,N_40840,N_48874);
and UO_901 (O_901,N_44437,N_49648);
or UO_902 (O_902,N_41097,N_49972);
nor UO_903 (O_903,N_49278,N_45074);
nor UO_904 (O_904,N_46499,N_43894);
and UO_905 (O_905,N_47672,N_44504);
xnor UO_906 (O_906,N_42087,N_47298);
nand UO_907 (O_907,N_44671,N_45159);
and UO_908 (O_908,N_46191,N_40471);
and UO_909 (O_909,N_45191,N_43838);
and UO_910 (O_910,N_44792,N_46263);
nand UO_911 (O_911,N_45064,N_40476);
and UO_912 (O_912,N_42090,N_45194);
nor UO_913 (O_913,N_49140,N_45976);
or UO_914 (O_914,N_48183,N_40328);
and UO_915 (O_915,N_43449,N_46031);
or UO_916 (O_916,N_40639,N_43582);
or UO_917 (O_917,N_42754,N_47145);
or UO_918 (O_918,N_45874,N_40924);
nand UO_919 (O_919,N_42409,N_41656);
and UO_920 (O_920,N_41025,N_40675);
nor UO_921 (O_921,N_43699,N_49340);
and UO_922 (O_922,N_40064,N_47972);
nand UO_923 (O_923,N_45497,N_46827);
nand UO_924 (O_924,N_48351,N_47148);
or UO_925 (O_925,N_49792,N_43177);
nand UO_926 (O_926,N_46883,N_40851);
xnor UO_927 (O_927,N_42289,N_41001);
or UO_928 (O_928,N_48936,N_42228);
nand UO_929 (O_929,N_41697,N_49941);
nor UO_930 (O_930,N_44403,N_43776);
nor UO_931 (O_931,N_41312,N_40643);
nor UO_932 (O_932,N_42838,N_43519);
or UO_933 (O_933,N_49063,N_43627);
nand UO_934 (O_934,N_48883,N_42533);
and UO_935 (O_935,N_46483,N_49917);
and UO_936 (O_936,N_42161,N_47758);
nor UO_937 (O_937,N_48234,N_49680);
and UO_938 (O_938,N_41134,N_47706);
or UO_939 (O_939,N_46287,N_41023);
or UO_940 (O_940,N_42740,N_43331);
nand UO_941 (O_941,N_48406,N_48046);
nor UO_942 (O_942,N_40762,N_48950);
nor UO_943 (O_943,N_43187,N_44014);
and UO_944 (O_944,N_41541,N_43524);
or UO_945 (O_945,N_42465,N_48707);
or UO_946 (O_946,N_47168,N_44190);
and UO_947 (O_947,N_49688,N_43846);
and UO_948 (O_948,N_48934,N_41474);
nand UO_949 (O_949,N_40327,N_49998);
and UO_950 (O_950,N_47658,N_41895);
or UO_951 (O_951,N_47524,N_40185);
nor UO_952 (O_952,N_47216,N_49268);
nor UO_953 (O_953,N_42326,N_42456);
nor UO_954 (O_954,N_49158,N_40096);
and UO_955 (O_955,N_49359,N_41182);
nand UO_956 (O_956,N_49069,N_41043);
and UO_957 (O_957,N_49186,N_49969);
or UO_958 (O_958,N_47108,N_41048);
nor UO_959 (O_959,N_40715,N_45671);
nand UO_960 (O_960,N_42244,N_42024);
or UO_961 (O_961,N_49056,N_47455);
or UO_962 (O_962,N_46826,N_41662);
nand UO_963 (O_963,N_47964,N_42046);
or UO_964 (O_964,N_43501,N_45826);
nor UO_965 (O_965,N_40849,N_43378);
or UO_966 (O_966,N_43205,N_46336);
xor UO_967 (O_967,N_48542,N_45288);
nor UO_968 (O_968,N_43558,N_49663);
xor UO_969 (O_969,N_45758,N_47820);
and UO_970 (O_970,N_43700,N_44629);
nand UO_971 (O_971,N_40341,N_48704);
or UO_972 (O_972,N_40977,N_42562);
nor UO_973 (O_973,N_45023,N_43841);
or UO_974 (O_974,N_49689,N_46253);
nor UO_975 (O_975,N_45825,N_49939);
nand UO_976 (O_976,N_45746,N_41970);
nor UO_977 (O_977,N_40302,N_47144);
xor UO_978 (O_978,N_47922,N_49060);
and UO_979 (O_979,N_46674,N_49279);
nor UO_980 (O_980,N_41247,N_41389);
and UO_981 (O_981,N_43899,N_48401);
nand UO_982 (O_982,N_40912,N_43600);
nor UO_983 (O_983,N_42596,N_44923);
nand UO_984 (O_984,N_42981,N_44441);
xor UO_985 (O_985,N_46731,N_40801);
or UO_986 (O_986,N_42812,N_44313);
or UO_987 (O_987,N_43502,N_46437);
nand UO_988 (O_988,N_43050,N_40449);
nor UO_989 (O_989,N_47926,N_41383);
nor UO_990 (O_990,N_45061,N_49835);
or UO_991 (O_991,N_46193,N_48392);
and UO_992 (O_992,N_41470,N_42909);
and UO_993 (O_993,N_41952,N_41806);
nand UO_994 (O_994,N_42945,N_43300);
and UO_995 (O_995,N_43436,N_46541);
and UO_996 (O_996,N_40248,N_46582);
nor UO_997 (O_997,N_41937,N_41238);
xnor UO_998 (O_998,N_45428,N_49384);
nand UO_999 (O_999,N_45733,N_46305);
nor UO_1000 (O_1000,N_47805,N_44370);
nor UO_1001 (O_1001,N_49231,N_42246);
xor UO_1002 (O_1002,N_46241,N_44523);
nor UO_1003 (O_1003,N_46645,N_44323);
and UO_1004 (O_1004,N_49011,N_49350);
and UO_1005 (O_1005,N_42903,N_44260);
and UO_1006 (O_1006,N_40755,N_41635);
nor UO_1007 (O_1007,N_47071,N_46828);
and UO_1008 (O_1008,N_43787,N_47056);
nand UO_1009 (O_1009,N_44104,N_48334);
and UO_1010 (O_1010,N_43387,N_47374);
or UO_1011 (O_1011,N_41496,N_45587);
xnor UO_1012 (O_1012,N_43630,N_45910);
nor UO_1013 (O_1013,N_49786,N_42728);
and UO_1014 (O_1014,N_49937,N_40567);
or UO_1015 (O_1015,N_44327,N_40678);
nor UO_1016 (O_1016,N_42142,N_45388);
nand UO_1017 (O_1017,N_49813,N_45262);
nor UO_1018 (O_1018,N_43818,N_48132);
nor UO_1019 (O_1019,N_41788,N_49277);
nor UO_1020 (O_1020,N_43802,N_46823);
nand UO_1021 (O_1021,N_41547,N_41319);
or UO_1022 (O_1022,N_45789,N_40040);
or UO_1023 (O_1023,N_49974,N_43049);
or UO_1024 (O_1024,N_45558,N_49574);
and UO_1025 (O_1025,N_43737,N_45494);
and UO_1026 (O_1026,N_44977,N_40326);
nand UO_1027 (O_1027,N_44676,N_47176);
or UO_1028 (O_1028,N_43231,N_43311);
xor UO_1029 (O_1029,N_48488,N_48225);
xnor UO_1030 (O_1030,N_44228,N_40939);
nand UO_1031 (O_1031,N_49275,N_46792);
nand UO_1032 (O_1032,N_40617,N_43259);
or UO_1033 (O_1033,N_41118,N_44795);
xor UO_1034 (O_1034,N_48422,N_46236);
or UO_1035 (O_1035,N_46708,N_40736);
and UO_1036 (O_1036,N_41218,N_43792);
nor UO_1037 (O_1037,N_46406,N_49273);
nor UO_1038 (O_1038,N_47140,N_40797);
xor UO_1039 (O_1039,N_48938,N_44876);
and UO_1040 (O_1040,N_49528,N_47128);
and UO_1041 (O_1041,N_49198,N_45384);
and UO_1042 (O_1042,N_42348,N_49766);
xnor UO_1043 (O_1043,N_46389,N_41947);
nand UO_1044 (O_1044,N_48178,N_45827);
or UO_1045 (O_1045,N_44688,N_42129);
xnor UO_1046 (O_1046,N_47991,N_45941);
and UO_1047 (O_1047,N_44998,N_47102);
nor UO_1048 (O_1048,N_41209,N_49390);
and UO_1049 (O_1049,N_47152,N_41060);
or UO_1050 (O_1050,N_44500,N_40985);
or UO_1051 (O_1051,N_44862,N_48288);
or UO_1052 (O_1052,N_45244,N_41400);
or UO_1053 (O_1053,N_43010,N_42654);
nand UO_1054 (O_1054,N_40580,N_46976);
nand UO_1055 (O_1055,N_43380,N_43423);
nand UO_1056 (O_1056,N_42607,N_49438);
and UO_1057 (O_1057,N_48778,N_41694);
and UO_1058 (O_1058,N_46739,N_46420);
and UO_1059 (O_1059,N_40178,N_48448);
nand UO_1060 (O_1060,N_46992,N_47222);
nand UO_1061 (O_1061,N_46487,N_49896);
or UO_1062 (O_1062,N_43418,N_40618);
or UO_1063 (O_1063,N_43112,N_44161);
and UO_1064 (O_1064,N_43490,N_46784);
or UO_1065 (O_1065,N_47560,N_48152);
and UO_1066 (O_1066,N_48001,N_45542);
and UO_1067 (O_1067,N_45151,N_43976);
or UO_1068 (O_1068,N_41787,N_43965);
nor UO_1069 (O_1069,N_49346,N_43544);
or UO_1070 (O_1070,N_49415,N_49637);
nand UO_1071 (O_1071,N_42580,N_48271);
nor UO_1072 (O_1072,N_44854,N_40880);
nand UO_1073 (O_1073,N_46796,N_47045);
xor UO_1074 (O_1074,N_47832,N_47978);
or UO_1075 (O_1075,N_41204,N_41879);
xor UO_1076 (O_1076,N_49387,N_41822);
nand UO_1077 (O_1077,N_40155,N_41394);
nand UO_1078 (O_1078,N_40587,N_44541);
nand UO_1079 (O_1079,N_49488,N_40176);
and UO_1080 (O_1080,N_40917,N_48954);
xnor UO_1081 (O_1081,N_42855,N_45663);
nand UO_1082 (O_1082,N_41342,N_42932);
or UO_1083 (O_1083,N_47039,N_49349);
and UO_1084 (O_1084,N_45287,N_41258);
nand UO_1085 (O_1085,N_44028,N_42716);
nand UO_1086 (O_1086,N_49878,N_45036);
nor UO_1087 (O_1087,N_40394,N_46038);
or UO_1088 (O_1088,N_44997,N_49499);
nand UO_1089 (O_1089,N_47856,N_48570);
nor UO_1090 (O_1090,N_41887,N_42889);
nor UO_1091 (O_1091,N_41288,N_48857);
nor UO_1092 (O_1092,N_40059,N_48635);
and UO_1093 (O_1093,N_49316,N_45471);
and UO_1094 (O_1094,N_40073,N_44783);
nor UO_1095 (O_1095,N_45467,N_48999);
or UO_1096 (O_1096,N_45579,N_46033);
and UO_1097 (O_1097,N_46882,N_43689);
or UO_1098 (O_1098,N_44140,N_45961);
or UO_1099 (O_1099,N_41059,N_49631);
and UO_1100 (O_1100,N_44330,N_41653);
nand UO_1101 (O_1101,N_44029,N_45672);
and UO_1102 (O_1102,N_48931,N_44720);
and UO_1103 (O_1103,N_49986,N_42015);
or UO_1104 (O_1104,N_48969,N_49569);
nor UO_1105 (O_1105,N_43826,N_45508);
nand UO_1106 (O_1106,N_44059,N_45739);
and UO_1107 (O_1107,N_44393,N_45463);
and UO_1108 (O_1108,N_49956,N_47782);
or UO_1109 (O_1109,N_47117,N_43950);
and UO_1110 (O_1110,N_43563,N_45752);
or UO_1111 (O_1111,N_43585,N_49364);
xor UO_1112 (O_1112,N_49405,N_41370);
and UO_1113 (O_1113,N_42473,N_44449);
nand UO_1114 (O_1114,N_46791,N_42116);
nor UO_1115 (O_1115,N_42765,N_43384);
xnor UO_1116 (O_1116,N_49310,N_42840);
nor UO_1117 (O_1117,N_42629,N_47435);
nand UO_1118 (O_1118,N_45864,N_42032);
nand UO_1119 (O_1119,N_41846,N_45810);
or UO_1120 (O_1120,N_49229,N_43003);
nor UO_1121 (O_1121,N_41000,N_47151);
xnor UO_1122 (O_1122,N_42662,N_44606);
nor UO_1123 (O_1123,N_40970,N_41640);
and UO_1124 (O_1124,N_44407,N_49873);
and UO_1125 (O_1125,N_49890,N_45853);
nand UO_1126 (O_1126,N_47170,N_49958);
nand UO_1127 (O_1127,N_44843,N_41056);
or UO_1128 (O_1128,N_49810,N_41093);
and UO_1129 (O_1129,N_41189,N_46089);
and UO_1130 (O_1130,N_43785,N_40199);
nor UO_1131 (O_1131,N_41291,N_47973);
nand UO_1132 (O_1132,N_47091,N_49313);
or UO_1133 (O_1133,N_43271,N_46471);
and UO_1134 (O_1134,N_40448,N_40667);
nor UO_1135 (O_1135,N_46754,N_44242);
nor UO_1136 (O_1136,N_41323,N_49197);
or UO_1137 (O_1137,N_44426,N_40109);
and UO_1138 (O_1138,N_49436,N_42058);
nand UO_1139 (O_1139,N_46930,N_43005);
and UO_1140 (O_1140,N_45324,N_41856);
and UO_1141 (O_1141,N_46952,N_44786);
nor UO_1142 (O_1142,N_46912,N_49821);
nor UO_1143 (O_1143,N_47889,N_40577);
or UO_1144 (O_1144,N_41692,N_49617);
or UO_1145 (O_1145,N_47848,N_47333);
and UO_1146 (O_1146,N_47804,N_41533);
or UO_1147 (O_1147,N_42878,N_46908);
xor UO_1148 (O_1148,N_40647,N_47573);
or UO_1149 (O_1149,N_48526,N_47985);
nand UO_1150 (O_1150,N_41611,N_42583);
or UO_1151 (O_1151,N_48131,N_41073);
nand UO_1152 (O_1152,N_46044,N_48065);
nand UO_1153 (O_1153,N_46576,N_47996);
or UO_1154 (O_1154,N_41672,N_41024);
or UO_1155 (O_1155,N_41110,N_49380);
nor UO_1156 (O_1156,N_41931,N_40499);
nor UO_1157 (O_1157,N_46288,N_47220);
or UO_1158 (O_1158,N_45627,N_47515);
nor UO_1159 (O_1159,N_49215,N_45473);
nand UO_1160 (O_1160,N_41053,N_41002);
and UO_1161 (O_1161,N_40881,N_41368);
and UO_1162 (O_1162,N_42166,N_45153);
nand UO_1163 (O_1163,N_42756,N_44867);
and UO_1164 (O_1164,N_43473,N_47545);
xor UO_1165 (O_1165,N_43613,N_44460);
xnor UO_1166 (O_1166,N_48299,N_40674);
or UO_1167 (O_1167,N_45142,N_43424);
nor UO_1168 (O_1168,N_40899,N_48691);
and UO_1169 (O_1169,N_47901,N_43236);
nand UO_1170 (O_1170,N_41131,N_47244);
or UO_1171 (O_1171,N_49203,N_42942);
nand UO_1172 (O_1172,N_48891,N_42616);
and UO_1173 (O_1173,N_49594,N_41250);
and UO_1174 (O_1174,N_41503,N_49116);
nand UO_1175 (O_1175,N_46692,N_48056);
nand UO_1176 (O_1176,N_45987,N_47630);
or UO_1177 (O_1177,N_49826,N_45261);
nor UO_1178 (O_1178,N_45557,N_46322);
and UO_1179 (O_1179,N_42809,N_41153);
and UO_1180 (O_1180,N_41081,N_49930);
nor UO_1181 (O_1181,N_42031,N_41396);
nor UO_1182 (O_1182,N_47429,N_45541);
xor UO_1183 (O_1183,N_48886,N_40946);
nor UO_1184 (O_1184,N_44435,N_40355);
nand UO_1185 (O_1185,N_49949,N_40458);
nand UO_1186 (O_1186,N_48699,N_41554);
or UO_1187 (O_1187,N_43445,N_44149);
xor UO_1188 (O_1188,N_44938,N_41986);
or UO_1189 (O_1189,N_47021,N_47689);
nor UO_1190 (O_1190,N_44789,N_46804);
nand UO_1191 (O_1191,N_49755,N_45691);
nand UO_1192 (O_1192,N_46951,N_42706);
nand UO_1193 (O_1193,N_46785,N_41275);
or UO_1194 (O_1194,N_43268,N_47995);
or UO_1195 (O_1195,N_46137,N_46560);
or UO_1196 (O_1196,N_43107,N_44316);
xor UO_1197 (O_1197,N_43692,N_48844);
nor UO_1198 (O_1198,N_48213,N_47407);
nor UO_1199 (O_1199,N_40042,N_44322);
or UO_1200 (O_1200,N_44489,N_41491);
and UO_1201 (O_1201,N_46382,N_40565);
nor UO_1202 (O_1202,N_41688,N_48910);
nor UO_1203 (O_1203,N_40477,N_45820);
xnor UO_1204 (O_1204,N_42828,N_40563);
nor UO_1205 (O_1205,N_41359,N_46323);
nor UO_1206 (O_1206,N_46229,N_41704);
or UO_1207 (O_1207,N_44708,N_48250);
or UO_1208 (O_1208,N_42342,N_48393);
xor UO_1209 (O_1209,N_40894,N_49365);
nand UO_1210 (O_1210,N_47966,N_48390);
nand UO_1211 (O_1211,N_43513,N_43302);
or UO_1212 (O_1212,N_46318,N_42317);
nor UO_1213 (O_1213,N_40002,N_44665);
or UO_1214 (O_1214,N_46763,N_44402);
nor UO_1215 (O_1215,N_49053,N_42106);
xnor UO_1216 (O_1216,N_46076,N_40269);
and UO_1217 (O_1217,N_44160,N_49863);
xnor UO_1218 (O_1218,N_41969,N_44016);
and UO_1219 (O_1219,N_47100,N_43567);
or UO_1220 (O_1220,N_43640,N_40790);
or UO_1221 (O_1221,N_41851,N_43221);
xnor UO_1222 (O_1222,N_40568,N_46240);
or UO_1223 (O_1223,N_41990,N_47695);
nor UO_1224 (O_1224,N_48814,N_49370);
nand UO_1225 (O_1225,N_41271,N_49233);
nor UO_1226 (O_1226,N_45490,N_46545);
or UO_1227 (O_1227,N_40106,N_49788);
xnor UO_1228 (O_1228,N_48496,N_45155);
and UO_1229 (O_1229,N_49490,N_47745);
nand UO_1230 (O_1230,N_46163,N_47632);
nand UO_1231 (O_1231,N_48082,N_45830);
and UO_1232 (O_1232,N_41095,N_47042);
xor UO_1233 (O_1233,N_44299,N_45483);
nor UO_1234 (O_1234,N_42983,N_47184);
nand UO_1235 (O_1235,N_42832,N_47494);
nor UO_1236 (O_1236,N_46345,N_40312);
nand UO_1237 (O_1237,N_45226,N_42977);
and UO_1238 (O_1238,N_41188,N_41534);
or UO_1239 (O_1239,N_48071,N_45718);
xor UO_1240 (O_1240,N_45386,N_41108);
nand UO_1241 (O_1241,N_40895,N_42642);
or UO_1242 (O_1242,N_48665,N_44328);
and UO_1243 (O_1243,N_44607,N_49881);
nand UO_1244 (O_1244,N_42245,N_47245);
nor UO_1245 (O_1245,N_48738,N_46356);
and UO_1246 (O_1246,N_46445,N_45045);
nand UO_1247 (O_1247,N_41193,N_40169);
or UO_1248 (O_1248,N_49221,N_43643);
or UO_1249 (O_1249,N_45044,N_41563);
nor UO_1250 (O_1250,N_43716,N_44068);
or UO_1251 (O_1251,N_46919,N_46461);
nand UO_1252 (O_1252,N_43964,N_47057);
xnor UO_1253 (O_1253,N_43375,N_47916);
nor UO_1254 (O_1254,N_48276,N_45469);
and UO_1255 (O_1255,N_41129,N_49119);
nand UO_1256 (O_1256,N_41621,N_40161);
or UO_1257 (O_1257,N_41639,N_40763);
nor UO_1258 (O_1258,N_40159,N_47886);
nor UO_1259 (O_1259,N_40127,N_43514);
nand UO_1260 (O_1260,N_45133,N_47928);
or UO_1261 (O_1261,N_42975,N_46332);
and UO_1262 (O_1262,N_45254,N_49644);
xnor UO_1263 (O_1263,N_41531,N_43760);
nor UO_1264 (O_1264,N_46111,N_43276);
xor UO_1265 (O_1265,N_47771,N_47942);
and UO_1266 (O_1266,N_43650,N_43681);
or UO_1267 (O_1267,N_42929,N_44935);
and UO_1268 (O_1268,N_42123,N_44209);
nor UO_1269 (O_1269,N_47505,N_44167);
and UO_1270 (O_1270,N_49164,N_45424);
or UO_1271 (O_1271,N_43538,N_41208);
or UO_1272 (O_1272,N_41678,N_42649);
or UO_1273 (O_1273,N_42787,N_40436);
or UO_1274 (O_1274,N_49348,N_41726);
and UO_1275 (O_1275,N_42920,N_45871);
and UO_1276 (O_1276,N_47068,N_48502);
nand UO_1277 (O_1277,N_46259,N_46493);
and UO_1278 (O_1278,N_40429,N_42954);
nor UO_1279 (O_1279,N_45878,N_43569);
nand UO_1280 (O_1280,N_46511,N_47365);
or UO_1281 (O_1281,N_48088,N_40826);
or UO_1282 (O_1282,N_43766,N_46633);
or UO_1283 (O_1283,N_46753,N_47802);
nand UO_1284 (O_1284,N_46313,N_45500);
or UO_1285 (O_1285,N_44054,N_49636);
or UO_1286 (O_1286,N_46436,N_47141);
or UO_1287 (O_1287,N_44691,N_41033);
nor UO_1288 (O_1288,N_43995,N_44122);
xor UO_1289 (O_1289,N_46353,N_49619);
nand UO_1290 (O_1290,N_45156,N_41416);
nor UO_1291 (O_1291,N_46821,N_44112);
xor UO_1292 (O_1292,N_45049,N_48650);
nand UO_1293 (O_1293,N_44826,N_47974);
nand UO_1294 (O_1294,N_45930,N_48252);
nor UO_1295 (O_1295,N_41248,N_46523);
and UO_1296 (O_1296,N_42102,N_41761);
xnor UO_1297 (O_1297,N_42048,N_43982);
and UO_1298 (O_1298,N_49382,N_44668);
nand UO_1299 (O_1299,N_46426,N_40703);
nor UO_1300 (O_1300,N_41017,N_45172);
xor UO_1301 (O_1301,N_47034,N_42236);
and UO_1302 (O_1302,N_49125,N_48135);
nand UO_1303 (O_1303,N_45852,N_46853);
and UO_1304 (O_1304,N_47044,N_41776);
nor UO_1305 (O_1305,N_47625,N_49014);
and UO_1306 (O_1306,N_47483,N_42487);
nor UO_1307 (O_1307,N_42866,N_48122);
nor UO_1308 (O_1308,N_45303,N_48522);
nor UO_1309 (O_1309,N_40773,N_42460);
nor UO_1310 (O_1310,N_45122,N_41349);
and UO_1311 (O_1311,N_42207,N_40395);
nor UO_1312 (O_1312,N_47792,N_49894);
nor UO_1313 (O_1313,N_45239,N_43493);
or UO_1314 (O_1314,N_47105,N_45784);
or UO_1315 (O_1315,N_43379,N_42891);
nor UO_1316 (O_1316,N_46585,N_48927);
xor UO_1317 (O_1317,N_49603,N_41146);
or UO_1318 (O_1318,N_40179,N_47378);
nor UO_1319 (O_1319,N_46173,N_46617);
nor UO_1320 (O_1320,N_42376,N_42294);
nand UO_1321 (O_1321,N_49817,N_41296);
and UO_1322 (O_1322,N_46812,N_48417);
or UO_1323 (O_1323,N_46354,N_44886);
or UO_1324 (O_1324,N_48416,N_42152);
nor UO_1325 (O_1325,N_47844,N_49082);
nor UO_1326 (O_1326,N_44329,N_44207);
and UO_1327 (O_1327,N_46041,N_40905);
or UO_1328 (O_1328,N_40830,N_49999);
or UO_1329 (O_1329,N_47504,N_45209);
xnor UO_1330 (O_1330,N_41245,N_48992);
and UO_1331 (O_1331,N_41755,N_42665);
nor UO_1332 (O_1332,N_40249,N_46099);
or UO_1333 (O_1333,N_45865,N_42900);
or UO_1334 (O_1334,N_41664,N_41732);
nand UO_1335 (O_1335,N_47272,N_47389);
nand UO_1336 (O_1336,N_46415,N_43156);
nand UO_1337 (O_1337,N_42215,N_42922);
nor UO_1338 (O_1338,N_42450,N_45144);
and UO_1339 (O_1339,N_47415,N_42633);
nand UO_1340 (O_1340,N_43747,N_40913);
nor UO_1341 (O_1341,N_45137,N_47143);
and UO_1342 (O_1342,N_40681,N_49942);
nor UO_1343 (O_1343,N_46097,N_45213);
or UO_1344 (O_1344,N_49025,N_48968);
and UO_1345 (O_1345,N_40758,N_41385);
and UO_1346 (O_1346,N_47426,N_45754);
and UO_1347 (O_1347,N_48695,N_40163);
nand UO_1348 (O_1348,N_43611,N_41300);
or UO_1349 (O_1349,N_40291,N_40540);
and UO_1350 (O_1350,N_42397,N_45597);
nand UO_1351 (O_1351,N_45307,N_45684);
nor UO_1352 (O_1352,N_41455,N_40151);
nor UO_1353 (O_1353,N_46698,N_42823);
nor UO_1354 (O_1354,N_45040,N_42369);
and UO_1355 (O_1355,N_48055,N_43430);
nand UO_1356 (O_1356,N_49328,N_43816);
nor UO_1357 (O_1357,N_40237,N_42614);
and UO_1358 (O_1358,N_46034,N_42937);
nand UO_1359 (O_1359,N_48474,N_47230);
xnor UO_1360 (O_1360,N_46126,N_47594);
or UO_1361 (O_1361,N_45863,N_44376);
and UO_1362 (O_1362,N_41527,N_42543);
or UO_1363 (O_1363,N_45114,N_44902);
and UO_1364 (O_1364,N_41028,N_42959);
nor UO_1365 (O_1365,N_42044,N_44927);
nand UO_1366 (O_1366,N_42747,N_46166);
nand UO_1367 (O_1367,N_43200,N_46842);
or UO_1368 (O_1368,N_41313,N_45636);
nor UO_1369 (O_1369,N_46485,N_44397);
or UO_1370 (O_1370,N_41126,N_48486);
nor UO_1371 (O_1371,N_40226,N_49437);
nand UO_1372 (O_1372,N_47523,N_45844);
or UO_1373 (O_1373,N_45610,N_41594);
nand UO_1374 (O_1374,N_48982,N_43765);
nand UO_1375 (O_1375,N_40357,N_48871);
or UO_1376 (O_1376,N_42887,N_41184);
nor UO_1377 (O_1377,N_49668,N_49598);
nor UO_1378 (O_1378,N_40714,N_42488);
and UO_1379 (O_1379,N_48684,N_49590);
xnor UO_1380 (O_1380,N_45731,N_47860);
or UO_1381 (O_1381,N_42001,N_46845);
nand UO_1382 (O_1382,N_45354,N_49345);
and UO_1383 (O_1383,N_46028,N_46279);
or UO_1384 (O_1384,N_47949,N_45095);
xnor UO_1385 (O_1385,N_43476,N_45894);
or UO_1386 (O_1386,N_48797,N_45129);
nand UO_1387 (O_1387,N_49141,N_42359);
xor UO_1388 (O_1388,N_47685,N_41229);
nand UO_1389 (O_1389,N_42917,N_48724);
nor UO_1390 (O_1390,N_43206,N_42175);
and UO_1391 (O_1391,N_48315,N_40943);
nor UO_1392 (O_1392,N_42847,N_47738);
and UO_1393 (O_1393,N_43217,N_45951);
or UO_1394 (O_1394,N_40551,N_43013);
nor UO_1395 (O_1395,N_46551,N_41701);
and UO_1396 (O_1396,N_48671,N_48388);
or UO_1397 (O_1397,N_45685,N_45756);
nor UO_1398 (O_1398,N_46589,N_43312);
and UO_1399 (O_1399,N_43654,N_49267);
nand UO_1400 (O_1400,N_44538,N_40554);
nand UO_1401 (O_1401,N_43376,N_44178);
nor UO_1402 (O_1402,N_49961,N_48709);
nand UO_1403 (O_1403,N_44966,N_44574);
nor UO_1404 (O_1404,N_46971,N_45453);
or UO_1405 (O_1405,N_44262,N_42292);
xnor UO_1406 (O_1406,N_41764,N_41163);
xnor UO_1407 (O_1407,N_48142,N_48265);
nor UO_1408 (O_1408,N_41233,N_40128);
nor UO_1409 (O_1409,N_42182,N_45409);
or UO_1410 (O_1410,N_41029,N_46375);
or UO_1411 (O_1411,N_44102,N_46715);
and UO_1412 (O_1412,N_45924,N_49200);
nor UO_1413 (O_1413,N_49478,N_47777);
nand UO_1414 (O_1414,N_40688,N_48553);
or UO_1415 (O_1415,N_48688,N_46065);
or UO_1416 (O_1416,N_46079,N_44073);
or UO_1417 (O_1417,N_42203,N_46816);
xnor UO_1418 (O_1418,N_41794,N_46212);
and UO_1419 (O_1419,N_45942,N_45292);
nor UO_1420 (O_1420,N_40908,N_45747);
nor UO_1421 (O_1421,N_43052,N_42712);
or UO_1422 (O_1422,N_42449,N_47863);
xnor UO_1423 (O_1423,N_48008,N_42639);
nand UO_1424 (O_1424,N_40272,N_47063);
or UO_1425 (O_1425,N_40407,N_48355);
nand UO_1426 (O_1426,N_48727,N_44423);
or UO_1427 (O_1427,N_47501,N_44197);
xor UO_1428 (O_1428,N_45567,N_47959);
xor UO_1429 (O_1429,N_44308,N_49519);
nor UO_1430 (O_1430,N_49356,N_42643);
nand UO_1431 (O_1431,N_43239,N_44964);
and UO_1432 (O_1432,N_41050,N_44110);
nor UO_1433 (O_1433,N_46565,N_48036);
nand UO_1434 (O_1434,N_45665,N_48994);
and UO_1435 (O_1435,N_46907,N_40111);
and UO_1436 (O_1436,N_48326,N_44787);
nor UO_1437 (O_1437,N_45744,N_44004);
or UO_1438 (O_1438,N_46594,N_44418);
and UO_1439 (O_1439,N_48182,N_42873);
and UO_1440 (O_1440,N_40676,N_46027);
or UO_1441 (O_1441,N_48123,N_43182);
or UO_1442 (O_1442,N_40621,N_43884);
nor UO_1443 (O_1443,N_47142,N_40579);
nand UO_1444 (O_1444,N_42338,N_48545);
or UO_1445 (O_1445,N_42586,N_41709);
or UO_1446 (O_1446,N_46997,N_42332);
or UO_1447 (O_1447,N_45640,N_44647);
or UO_1448 (O_1448,N_47469,N_46874);
or UO_1449 (O_1449,N_43008,N_47852);
nand UO_1450 (O_1450,N_49849,N_43454);
nand UO_1451 (O_1451,N_48761,N_46262);
nor UO_1452 (O_1452,N_48051,N_41644);
nor UO_1453 (O_1453,N_46378,N_44374);
nor UO_1454 (O_1454,N_45725,N_42680);
xnor UO_1455 (O_1455,N_41919,N_42035);
xor UO_1456 (O_1456,N_42868,N_40697);
and UO_1457 (O_1457,N_46340,N_41476);
and UO_1458 (O_1458,N_47795,N_49602);
nand UO_1459 (O_1459,N_45678,N_45152);
nand UO_1460 (O_1460,N_42335,N_42206);
nor UO_1461 (O_1461,N_43879,N_48705);
nor UO_1462 (O_1462,N_48779,N_46646);
nor UO_1463 (O_1463,N_47377,N_49084);
nand UO_1464 (O_1464,N_43726,N_40466);
or UO_1465 (O_1465,N_40930,N_48771);
nor UO_1466 (O_1466,N_47744,N_42079);
xor UO_1467 (O_1467,N_49128,N_45837);
or UO_1468 (O_1468,N_41347,N_48989);
or UO_1469 (O_1469,N_40365,N_45520);
nor UO_1470 (O_1470,N_45333,N_44155);
and UO_1471 (O_1471,N_44036,N_43833);
and UO_1472 (O_1472,N_41620,N_40048);
nor UO_1473 (O_1473,N_48896,N_46895);
nand UO_1474 (O_1474,N_44450,N_49885);
nand UO_1475 (O_1475,N_40696,N_45119);
and UO_1476 (O_1476,N_40559,N_41328);
or UO_1477 (O_1477,N_45131,N_45051);
nand UO_1478 (O_1478,N_42947,N_48949);
nor UO_1479 (O_1479,N_46189,N_47673);
nand UO_1480 (O_1480,N_40434,N_45281);
nor UO_1481 (O_1481,N_45117,N_41200);
or UO_1482 (O_1482,N_42990,N_45107);
nand UO_1483 (O_1483,N_44424,N_45482);
nor UO_1484 (O_1484,N_47885,N_42033);
xnor UO_1485 (O_1485,N_43265,N_47073);
and UO_1486 (O_1486,N_41502,N_41528);
nor UO_1487 (O_1487,N_41843,N_47103);
nor UO_1488 (O_1488,N_43020,N_48274);
and UO_1489 (O_1489,N_45757,N_48530);
and UO_1490 (O_1490,N_40399,N_40592);
and UO_1491 (O_1491,N_44446,N_45632);
nand UO_1492 (O_1492,N_48435,N_41605);
nor UO_1493 (O_1493,N_46104,N_41112);
nand UO_1494 (O_1494,N_43886,N_40834);
and UO_1495 (O_1495,N_47938,N_45675);
or UO_1496 (O_1496,N_49981,N_48487);
nand UO_1497 (O_1497,N_46820,N_48649);
and UO_1498 (O_1498,N_48033,N_44050);
nor UO_1499 (O_1499,N_44332,N_45057);
or UO_1500 (O_1500,N_44303,N_46556);
nor UO_1501 (O_1501,N_40657,N_46190);
nand UO_1502 (O_1502,N_40529,N_43985);
nor UO_1503 (O_1503,N_42451,N_40112);
nand UO_1504 (O_1504,N_42876,N_47394);
and UO_1505 (O_1505,N_45085,N_46722);
or UO_1506 (O_1506,N_48255,N_42258);
or UO_1507 (O_1507,N_44091,N_40680);
or UO_1508 (O_1508,N_41953,N_42986);
or UO_1509 (O_1509,N_40748,N_40264);
or UO_1510 (O_1510,N_43199,N_45609);
and UO_1511 (O_1511,N_44983,N_41911);
and UO_1512 (O_1512,N_40497,N_49809);
or UO_1513 (O_1513,N_41270,N_41966);
or UO_1514 (O_1514,N_43811,N_42389);
nand UO_1515 (O_1515,N_40196,N_44433);
nand UO_1516 (O_1516,N_47214,N_46358);
nand UO_1517 (O_1517,N_45624,N_43904);
nand UO_1518 (O_1518,N_46732,N_46865);
xor UO_1519 (O_1519,N_47544,N_48672);
nand UO_1520 (O_1520,N_45374,N_42303);
nor UO_1521 (O_1521,N_40117,N_42720);
and UO_1522 (O_1522,N_49462,N_47260);
nand UO_1523 (O_1523,N_45715,N_41420);
and UO_1524 (O_1524,N_41659,N_44645);
nor UO_1525 (O_1525,N_48711,N_43146);
nor UO_1526 (O_1526,N_47743,N_43489);
nand UO_1527 (O_1527,N_41145,N_49166);
or UO_1528 (O_1528,N_43596,N_40594);
or UO_1529 (O_1529,N_41363,N_45990);
xor UO_1530 (O_1530,N_43892,N_47540);
nor UO_1531 (O_1531,N_46225,N_46547);
and UO_1532 (O_1532,N_44018,N_40689);
and UO_1533 (O_1533,N_43735,N_42158);
and UO_1534 (O_1534,N_41873,N_42931);
nand UO_1535 (O_1535,N_49381,N_41080);
and UO_1536 (O_1536,N_47240,N_46544);
nand UO_1537 (O_1537,N_43250,N_41601);
xnor UO_1538 (O_1538,N_48863,N_44618);
nor UO_1539 (O_1539,N_48605,N_44440);
and UO_1540 (O_1540,N_44852,N_43719);
or UO_1541 (O_1541,N_49049,N_40890);
xor UO_1542 (O_1542,N_43349,N_45289);
xnor UO_1543 (O_1543,N_44210,N_49606);
xnor UO_1544 (O_1544,N_43374,N_46666);
and UO_1545 (O_1545,N_41217,N_41765);
nor UO_1546 (O_1546,N_43980,N_42520);
or UO_1547 (O_1547,N_46301,N_46516);
nor UO_1548 (O_1548,N_48687,N_42933);
nand UO_1549 (O_1549,N_49622,N_40556);
xor UO_1550 (O_1550,N_49026,N_46584);
and UO_1551 (O_1551,N_40380,N_45399);
nor UO_1552 (O_1552,N_46085,N_40274);
and UO_1553 (O_1553,N_47086,N_42831);
nand UO_1554 (O_1554,N_41561,N_41713);
nor UO_1555 (O_1555,N_43256,N_44721);
nand UO_1556 (O_1556,N_47084,N_45799);
nand UO_1557 (O_1557,N_43675,N_44186);
and UO_1558 (O_1558,N_43229,N_49541);
and UO_1559 (O_1559,N_41346,N_46363);
or UO_1560 (O_1560,N_44096,N_42222);
and UO_1561 (O_1561,N_44507,N_40787);
or UO_1562 (O_1562,N_44942,N_45611);
and UO_1563 (O_1563,N_41354,N_47351);
and UO_1564 (O_1564,N_42356,N_46718);
or UO_1565 (O_1565,N_43483,N_42118);
nand UO_1566 (O_1566,N_40800,N_47338);
nor UO_1567 (O_1567,N_44133,N_45265);
or UO_1568 (O_1568,N_44769,N_41588);
and UO_1569 (O_1569,N_42795,N_43487);
and UO_1570 (O_1570,N_40035,N_42155);
or UO_1571 (O_1571,N_47283,N_44743);
and UO_1572 (O_1572,N_46418,N_49561);
and UO_1573 (O_1573,N_49468,N_40060);
nor UO_1574 (O_1574,N_45427,N_40315);
and UO_1575 (O_1575,N_41555,N_45544);
or UO_1576 (O_1576,N_46181,N_41768);
nor UO_1577 (O_1577,N_44959,N_45991);
or UO_1578 (O_1578,N_49721,N_47816);
xnor UO_1579 (O_1579,N_41063,N_49420);
nand UO_1580 (O_1580,N_43512,N_43211);
nor UO_1581 (O_1581,N_40612,N_41810);
or UO_1582 (O_1582,N_47981,N_48753);
xnor UO_1583 (O_1583,N_48763,N_48218);
xor UO_1584 (O_1584,N_48161,N_48126);
and UO_1585 (O_1585,N_42752,N_42700);
nor UO_1586 (O_1586,N_44723,N_48513);
and UO_1587 (O_1587,N_48777,N_44755);
nand UO_1588 (O_1588,N_48098,N_47847);
and UO_1589 (O_1589,N_40792,N_42531);
nand UO_1590 (O_1590,N_41685,N_44619);
or UO_1591 (O_1591,N_42219,N_44640);
or UO_1592 (O_1592,N_49459,N_43653);
and UO_1593 (O_1593,N_45193,N_49085);
and UO_1594 (O_1594,N_45982,N_49466);
nand UO_1595 (O_1595,N_46949,N_48531);
or UO_1596 (O_1596,N_47422,N_48563);
or UO_1597 (O_1597,N_41585,N_43061);
nor UO_1598 (O_1598,N_45679,N_41877);
nor UO_1599 (O_1599,N_40803,N_49175);
and UO_1600 (O_1600,N_48742,N_47692);
nor UO_1601 (O_1601,N_47157,N_48935);
xor UO_1602 (O_1602,N_49058,N_41747);
nand UO_1603 (O_1603,N_43754,N_45608);
nor UO_1604 (O_1604,N_42385,N_46771);
nand UO_1605 (O_1605,N_40604,N_47934);
or UO_1606 (O_1606,N_40974,N_42422);
or UO_1607 (O_1607,N_44392,N_47124);
or UO_1608 (O_1608,N_49218,N_47456);
and UO_1609 (O_1609,N_40699,N_48806);
nor UO_1610 (O_1610,N_45174,N_42505);
nor UO_1611 (O_1611,N_47440,N_46755);
and UO_1612 (O_1612,N_43806,N_47211);
or UO_1613 (O_1613,N_45495,N_43831);
nor UO_1614 (O_1614,N_49526,N_49798);
xor UO_1615 (O_1615,N_42895,N_43442);
and UO_1616 (O_1616,N_45071,N_48561);
nor UO_1617 (O_1617,N_44200,N_45258);
or UO_1618 (O_1618,N_48285,N_49525);
nand UO_1619 (O_1619,N_49255,N_40020);
or UO_1620 (O_1620,N_48111,N_45264);
nor UO_1621 (O_1621,N_46694,N_41508);
or UO_1622 (O_1622,N_43797,N_49460);
nand UO_1623 (O_1623,N_48937,N_45087);
or UO_1624 (O_1624,N_43185,N_41627);
nand UO_1625 (O_1625,N_40638,N_47683);
nor UO_1626 (O_1626,N_45836,N_47829);
or UO_1627 (O_1627,N_41156,N_41722);
nor UO_1628 (O_1628,N_45447,N_40143);
or UO_1629 (O_1629,N_40103,N_43468);
xor UO_1630 (O_1630,N_42970,N_43845);
xor UO_1631 (O_1631,N_46809,N_40284);
nor UO_1632 (O_1632,N_41714,N_44827);
or UO_1633 (O_1633,N_42017,N_41289);
and UO_1634 (O_1634,N_47831,N_43972);
nand UO_1635 (O_1635,N_42331,N_48970);
and UO_1636 (O_1636,N_46119,N_49023);
or UO_1637 (O_1637,N_48515,N_40642);
xnor UO_1638 (O_1638,N_40799,N_41399);
nor UO_1639 (O_1639,N_45945,N_46337);
and UO_1640 (O_1640,N_48948,N_42992);
xnor UO_1641 (O_1641,N_49173,N_47461);
or UO_1642 (O_1642,N_41847,N_41679);
or UO_1643 (O_1643,N_49861,N_43041);
and UO_1644 (O_1644,N_49769,N_47154);
and UO_1645 (O_1645,N_44765,N_48685);
and UO_1646 (O_1646,N_45394,N_44587);
or UO_1647 (O_1647,N_47615,N_43711);
nor UO_1648 (O_1648,N_44277,N_47262);
nand UO_1649 (O_1649,N_45798,N_40816);
or UO_1650 (O_1650,N_41595,N_45868);
and UO_1651 (O_1651,N_40628,N_46011);
nor UO_1652 (O_1652,N_47940,N_40473);
and UO_1653 (O_1653,N_47606,N_44432);
or UO_1654 (O_1654,N_44216,N_47562);
or UO_1655 (O_1655,N_45176,N_40319);
nor UO_1656 (O_1656,N_43062,N_41687);
or UO_1657 (O_1657,N_40044,N_40934);
nor UO_1658 (O_1658,N_43587,N_47202);
or UO_1659 (O_1659,N_49077,N_42237);
and UO_1660 (O_1660,N_46640,N_40280);
nor UO_1661 (O_1661,N_40034,N_48880);
nand UO_1662 (O_1662,N_44304,N_49020);
nor UO_1663 (O_1663,N_44926,N_47158);
nand UO_1664 (O_1664,N_40663,N_48536);
xor UO_1665 (O_1665,N_45623,N_42154);
xor UO_1666 (O_1666,N_48402,N_46696);
and UO_1667 (O_1667,N_40332,N_42858);
and UO_1668 (O_1668,N_44553,N_49134);
nand UO_1669 (O_1669,N_41779,N_48764);
xor UO_1670 (O_1670,N_43190,N_45111);
or UO_1671 (O_1671,N_46429,N_46335);
nand UO_1672 (O_1672,N_48678,N_42247);
nand UO_1673 (O_1673,N_43320,N_48264);
or UO_1674 (O_1674,N_42553,N_46387);
and UO_1675 (O_1675,N_48978,N_44585);
nand UO_1676 (O_1676,N_42650,N_47237);
and UO_1677 (O_1677,N_45358,N_42509);
and UO_1678 (O_1678,N_44776,N_43057);
nor UO_1679 (O_1679,N_44095,N_45330);
nor UO_1680 (O_1680,N_48645,N_44641);
nor UO_1681 (O_1681,N_45549,N_44980);
or UO_1682 (O_1682,N_40342,N_43074);
or UO_1683 (O_1683,N_43577,N_45727);
nor UO_1684 (O_1684,N_44512,N_45664);
and UO_1685 (O_1685,N_44378,N_40833);
or UO_1686 (O_1686,N_44890,N_45298);
nor UO_1687 (O_1687,N_49061,N_47608);
nand UO_1688 (O_1688,N_46492,N_45879);
nand UO_1689 (O_1689,N_43238,N_45630);
and UO_1690 (O_1690,N_46994,N_47712);
or UO_1691 (O_1691,N_43920,N_42403);
xnor UO_1692 (O_1692,N_46113,N_49451);
and UO_1693 (O_1693,N_47933,N_46944);
and UO_1694 (O_1694,N_45162,N_49307);
or UO_1695 (O_1695,N_48023,N_44280);
or UO_1696 (O_1696,N_40525,N_49427);
nand UO_1697 (O_1697,N_47992,N_49103);
xnor UO_1698 (O_1698,N_40510,N_42057);
or UO_1699 (O_1699,N_42151,N_46615);
xnor UO_1700 (O_1700,N_43801,N_46810);
nand UO_1701 (O_1701,N_44808,N_46344);
or UO_1702 (O_1702,N_47271,N_45775);
or UO_1703 (O_1703,N_40162,N_42445);
and UO_1704 (O_1704,N_42162,N_49804);
nor UO_1705 (O_1705,N_49723,N_44021);
and UO_1706 (O_1706,N_46017,N_42904);
nand UO_1707 (O_1707,N_42813,N_44839);
and UO_1708 (O_1708,N_43637,N_41800);
and UO_1709 (O_1709,N_42461,N_46596);
nor UO_1710 (O_1710,N_42559,N_45273);
nand UO_1711 (O_1711,N_44903,N_41769);
nor UO_1712 (O_1712,N_48745,N_45353);
nor UO_1713 (O_1713,N_42935,N_43488);
nand UO_1714 (O_1714,N_43435,N_47693);
nor UO_1715 (O_1715,N_43865,N_48372);
nand UO_1716 (O_1716,N_41107,N_45813);
xor UO_1717 (O_1717,N_44468,N_48528);
xnor UO_1718 (O_1718,N_44265,N_49080);
and UO_1719 (O_1719,N_44353,N_42485);
xor UO_1720 (O_1720,N_42582,N_45769);
xnor UO_1721 (O_1721,N_46435,N_49857);
and UO_1722 (O_1722,N_49875,N_47720);
nor UO_1723 (O_1723,N_45873,N_43234);
nor UO_1724 (O_1724,N_41715,N_43999);
xnor UO_1725 (O_1725,N_42099,N_45996);
nand UO_1726 (O_1726,N_43397,N_42386);
nand UO_1727 (O_1727,N_43701,N_47659);
or UO_1728 (O_1728,N_48860,N_41590);
and UO_1729 (O_1729,N_41085,N_43872);
nor UO_1730 (O_1730,N_40398,N_43421);
xnor UO_1731 (O_1731,N_48459,N_48540);
nor UO_1732 (O_1732,N_45637,N_49336);
nand UO_1733 (O_1733,N_48149,N_44350);
nor UO_1734 (O_1734,N_42737,N_46928);
nor UO_1735 (O_1735,N_44153,N_43207);
and UO_1736 (O_1736,N_47550,N_44425);
nand UO_1737 (O_1737,N_40611,N_46080);
or UO_1738 (O_1738,N_43916,N_40527);
or UO_1739 (O_1739,N_44052,N_43042);
xnor UO_1740 (O_1740,N_43278,N_42532);
xor UO_1741 (O_1741,N_43731,N_49088);
nand UO_1742 (O_1742,N_44900,N_43115);
nand UO_1743 (O_1743,N_42496,N_43054);
nand UO_1744 (O_1744,N_43870,N_49089);
nand UO_1745 (O_1745,N_48068,N_49383);
or UO_1746 (O_1746,N_45585,N_48552);
or UO_1747 (O_1747,N_47284,N_48061);
and UO_1748 (O_1748,N_49704,N_40649);
nand UO_1749 (O_1749,N_48668,N_46319);
nor UO_1750 (O_1750,N_46974,N_40718);
nand UO_1751 (O_1751,N_48679,N_49874);
nand UO_1752 (O_1752,N_46955,N_42641);
nand UO_1753 (O_1753,N_43216,N_47444);
nand UO_1754 (O_1754,N_43866,N_46202);
nor UO_1755 (O_1755,N_40526,N_42884);
or UO_1756 (O_1756,N_42785,N_40896);
nor UO_1757 (O_1757,N_41497,N_46035);
nand UO_1758 (O_1758,N_43849,N_40677);
or UO_1759 (O_1759,N_42157,N_43887);
nand UO_1760 (O_1760,N_45285,N_43181);
nor UO_1761 (O_1761,N_49147,N_45573);
or UO_1762 (O_1762,N_45793,N_42054);
xnor UO_1763 (O_1763,N_43324,N_41808);
nand UO_1764 (O_1764,N_41538,N_43718);
nor UO_1765 (O_1765,N_45884,N_41140);
and UO_1766 (O_1766,N_46084,N_47653);
or UO_1767 (O_1767,N_44740,N_46672);
and UO_1768 (O_1768,N_42480,N_42405);
nand UO_1769 (O_1769,N_49902,N_48708);
xor UO_1770 (O_1770,N_40212,N_49562);
and UO_1771 (O_1771,N_47561,N_49613);
and UO_1772 (O_1772,N_49911,N_47195);
and UO_1773 (O_1773,N_40222,N_49094);
and UO_1774 (O_1774,N_44901,N_46443);
or UO_1775 (O_1775,N_46709,N_49171);
or UO_1776 (O_1776,N_42799,N_46231);
or UO_1777 (O_1777,N_41795,N_44745);
or UO_1778 (O_1778,N_46180,N_45946);
xor UO_1779 (O_1779,N_49306,N_44289);
xor UO_1780 (O_1780,N_47761,N_46197);
nand UO_1781 (O_1781,N_47051,N_49568);
nand UO_1782 (O_1782,N_40524,N_44696);
or UO_1783 (O_1783,N_48904,N_44703);
or UO_1784 (O_1784,N_44409,N_47066);
or UO_1785 (O_1785,N_44695,N_47179);
nand UO_1786 (O_1786,N_42408,N_48600);
and UO_1787 (O_1787,N_46954,N_42732);
xor UO_1788 (O_1788,N_47247,N_42447);
xnor UO_1789 (O_1789,N_40283,N_47236);
and UO_1790 (O_1790,N_47473,N_44351);
or UO_1791 (O_1791,N_45501,N_44993);
nand UO_1792 (O_1792,N_43092,N_45893);
or UO_1793 (O_1793,N_44194,N_41552);
nor UO_1794 (O_1794,N_47756,N_41859);
nor UO_1795 (O_1795,N_40097,N_49040);
nor UO_1796 (O_1796,N_42923,N_44673);
xnor UO_1797 (O_1797,N_49737,N_40847);
xor UO_1798 (O_1798,N_47085,N_45580);
and UO_1799 (O_1799,N_40235,N_44842);
nor UO_1800 (O_1800,N_48205,N_45732);
or UO_1801 (O_1801,N_42145,N_42560);
nand UO_1802 (O_1802,N_43619,N_42803);
and UO_1803 (O_1803,N_46172,N_49822);
or UO_1804 (O_1804,N_42187,N_48269);
xor UO_1805 (O_1805,N_42901,N_43116);
or UO_1806 (O_1806,N_48773,N_46527);
and UO_1807 (O_1807,N_47414,N_43977);
nor UO_1808 (O_1808,N_41893,N_46203);
nand UO_1809 (O_1809,N_42489,N_47392);
nor UO_1810 (O_1810,N_47408,N_49376);
nor UO_1811 (O_1811,N_40378,N_42402);
nand UO_1812 (O_1812,N_43677,N_47131);
or UO_1813 (O_1813,N_40987,N_48767);
xnor UO_1814 (O_1814,N_41683,N_48503);
or UO_1815 (O_1815,N_44077,N_47334);
or UO_1816 (O_1816,N_48584,N_44062);
and UO_1817 (O_1817,N_48630,N_45875);
and UO_1818 (O_1818,N_49924,N_40275);
or UO_1819 (O_1819,N_40494,N_45028);
or UO_1820 (O_1820,N_43966,N_48366);
xnor UO_1821 (O_1821,N_49232,N_47858);
or UO_1822 (O_1822,N_40132,N_48437);
xor UO_1823 (O_1823,N_41274,N_45418);
nand UO_1824 (O_1824,N_46433,N_48403);
and UO_1825 (O_1825,N_45312,N_40050);
nand UO_1826 (O_1826,N_44939,N_44816);
nor UO_1827 (O_1827,N_47493,N_44193);
xor UO_1828 (O_1828,N_42439,N_44796);
nand UO_1829 (O_1829,N_47965,N_42093);
nand UO_1830 (O_1830,N_41871,N_42113);
nand UO_1831 (O_1831,N_40922,N_43274);
nor UO_1832 (O_1832,N_45444,N_48090);
or UO_1833 (O_1833,N_43541,N_41123);
and UO_1834 (O_1834,N_41337,N_45039);
nand UO_1835 (O_1835,N_44586,N_47530);
nor UO_1836 (O_1836,N_41276,N_42552);
nand UO_1837 (O_1837,N_41130,N_44556);
nor UO_1838 (O_1838,N_45383,N_40133);
or UO_1839 (O_1839,N_48534,N_48199);
nor UO_1840 (O_1840,N_42538,N_45564);
nor UO_1841 (O_1841,N_45229,N_42677);
nand UO_1842 (O_1842,N_48245,N_48249);
nor UO_1843 (O_1843,N_44255,N_44309);
nand UO_1844 (O_1844,N_40001,N_42149);
xor UO_1845 (O_1845,N_47921,N_45019);
xnor UO_1846 (O_1846,N_40501,N_40028);
or UO_1847 (O_1847,N_46128,N_43212);
nor UO_1848 (O_1848,N_44837,N_47742);
nand UO_1849 (O_1849,N_48383,N_46019);
nor UO_1850 (O_1850,N_47050,N_45319);
and UO_1851 (O_1851,N_47527,N_41266);
and UO_1852 (O_1852,N_44230,N_43280);
nor UO_1853 (O_1853,N_40489,N_43305);
or UO_1854 (O_1854,N_41943,N_44779);
nand UO_1855 (O_1855,N_40731,N_47582);
nand UO_1856 (O_1856,N_41309,N_43022);
or UO_1857 (O_1857,N_45458,N_40658);
nor UO_1858 (O_1858,N_46216,N_44635);
xnor UO_1859 (O_1859,N_42060,N_49005);
or UO_1860 (O_1860,N_43323,N_46657);
xor UO_1861 (O_1861,N_42340,N_45211);
and UO_1862 (O_1862,N_40424,N_43628);
nand UO_1863 (O_1863,N_44067,N_49258);
or UO_1864 (O_1864,N_44258,N_49300);
nor UO_1865 (O_1865,N_47185,N_41724);
or UO_1866 (O_1866,N_45359,N_48693);
nor UO_1867 (O_1867,N_41195,N_42384);
nor UO_1868 (O_1868,N_44714,N_49016);
xor UO_1869 (O_1869,N_40933,N_46444);
nor UO_1870 (O_1870,N_44969,N_48337);
nand UO_1871 (O_1871,N_49904,N_41523);
nand UO_1872 (O_1872,N_47924,N_47563);
nor UO_1873 (O_1873,N_44537,N_43651);
and UO_1874 (O_1874,N_47371,N_43902);
or UO_1875 (O_1875,N_42734,N_45689);
or UO_1876 (O_1876,N_43618,N_42193);
nand UO_1877 (O_1877,N_44464,N_46105);
nand UO_1878 (O_1878,N_43608,N_49042);
and UO_1879 (O_1879,N_43365,N_43063);
nand UO_1880 (O_1880,N_40999,N_48582);
nor UO_1881 (O_1881,N_48585,N_47822);
nand UO_1882 (O_1882,N_45751,N_44256);
and UO_1883 (O_1883,N_41214,N_46548);
and UO_1884 (O_1884,N_49554,N_44233);
nor UO_1885 (O_1885,N_43366,N_49948);
nand UO_1886 (O_1886,N_45912,N_42457);
or UO_1887 (O_1887,N_46366,N_47120);
nand UO_1888 (O_1888,N_44363,N_48020);
nand UO_1889 (O_1889,N_43687,N_46749);
xor UO_1890 (O_1890,N_41290,N_46160);
and UO_1891 (O_1891,N_46724,N_44911);
nor UO_1892 (O_1892,N_44341,N_42587);
nand UO_1893 (O_1893,N_40710,N_41757);
or UO_1894 (O_1894,N_41099,N_42147);
nor UO_1895 (O_1895,N_49957,N_49748);
nor UO_1896 (O_1896,N_46782,N_44931);
nand UO_1897 (O_1897,N_46779,N_40904);
nor UO_1898 (O_1898,N_49977,N_48286);
or UO_1899 (O_1899,N_43939,N_44738);
nor UO_1900 (O_1900,N_43171,N_48287);
xnor UO_1901 (O_1901,N_43377,N_45295);
nor UO_1902 (O_1902,N_41065,N_48750);
nand UO_1903 (O_1903,N_48802,N_46269);
nand UO_1904 (O_1904,N_49915,N_48772);
nand UO_1905 (O_1905,N_47868,N_42268);
nor UO_1906 (O_1906,N_40457,N_40557);
xnor UO_1907 (O_1907,N_45764,N_49839);
nand UO_1908 (O_1908,N_46807,N_46571);
nand UO_1909 (O_1909,N_42864,N_48560);
nor UO_1910 (O_1910,N_45301,N_40921);
or UO_1911 (O_1911,N_46858,N_47581);
and UO_1912 (O_1912,N_44726,N_40277);
nand UO_1913 (O_1913,N_48493,N_44804);
xnor UO_1914 (O_1914,N_47772,N_45112);
nor UO_1915 (O_1915,N_47839,N_45308);
nor UO_1916 (O_1916,N_42890,N_43767);
nor UO_1917 (O_1917,N_45824,N_49477);
nor UO_1918 (O_1918,N_47070,N_44236);
xnor UO_1919 (O_1919,N_49276,N_41602);
nor UO_1920 (O_1920,N_41382,N_40811);
and UO_1921 (O_1921,N_40047,N_43371);
nand UO_1922 (O_1922,N_41137,N_40192);
or UO_1923 (O_1923,N_45120,N_41784);
nor UO_1924 (O_1924,N_40427,N_41958);
nor UO_1925 (O_1925,N_42279,N_47350);
nand UO_1926 (O_1926,N_49107,N_47988);
nor UO_1927 (O_1927,N_40417,N_49796);
or UO_1928 (O_1928,N_43912,N_40372);
nor UO_1929 (O_1929,N_48726,N_40944);
and UO_1930 (O_1930,N_40823,N_43218);
nor UO_1931 (O_1931,N_45270,N_45189);
nor UO_1932 (O_1932,N_45755,N_46329);
or UO_1933 (O_1933,N_48610,N_49391);
nor UO_1934 (O_1934,N_49219,N_41648);
or UO_1935 (O_1935,N_40391,N_45762);
and UO_1936 (O_1936,N_46684,N_49073);
nor UO_1937 (O_1937,N_43450,N_45146);
nor UO_1938 (O_1938,N_47911,N_44162);
or UO_1939 (O_1939,N_49090,N_44658);
nand UO_1940 (O_1940,N_42800,N_47241);
nor UO_1941 (O_1941,N_43135,N_45975);
nor UO_1942 (O_1942,N_43243,N_42419);
nor UO_1943 (O_1943,N_49202,N_42980);
or UO_1944 (O_1944,N_43822,N_40652);
xnor UO_1945 (O_1945,N_46182,N_45249);
nor UO_1946 (O_1946,N_49630,N_42592);
or UO_1947 (O_1947,N_48464,N_49441);
and UO_1948 (O_1948,N_44951,N_42960);
and UO_1949 (O_1949,N_40634,N_42938);
nor UO_1950 (O_1950,N_49570,N_48718);
nand UO_1951 (O_1951,N_42314,N_45524);
or UO_1952 (O_1952,N_43301,N_49487);
nand UO_1953 (O_1953,N_44948,N_47447);
or UO_1954 (O_1954,N_49291,N_41231);
or UO_1955 (O_1955,N_44146,N_43546);
nor UO_1956 (O_1956,N_43086,N_42609);
or UO_1957 (O_1957,N_41974,N_47584);
nor UO_1958 (O_1958,N_43346,N_46047);
xor UO_1959 (O_1959,N_42518,N_42783);
or UO_1960 (O_1960,N_48227,N_45602);
nand UO_1961 (O_1961,N_49419,N_45927);
nand UO_1962 (O_1962,N_42966,N_49074);
nor UO_1963 (O_1963,N_48168,N_49324);
nand UO_1964 (O_1964,N_44858,N_45257);
nor UO_1965 (O_1965,N_45442,N_49757);
xnor UO_1966 (O_1966,N_43688,N_46053);
or UO_1967 (O_1967,N_44943,N_49952);
or UO_1968 (O_1968,N_42352,N_48346);
xnor UO_1969 (O_1969,N_43992,N_40415);
nor UO_1970 (O_1970,N_48296,N_47019);
nor UO_1971 (O_1971,N_41607,N_43913);
and UO_1972 (O_1972,N_44377,N_47280);
or UO_1973 (O_1973,N_42088,N_49659);
nor UO_1974 (O_1974,N_43286,N_40980);
nand UO_1975 (O_1975,N_41490,N_42898);
nor UO_1976 (O_1976,N_46349,N_48432);
nand UO_1977 (O_1977,N_40070,N_42844);
nor UO_1978 (O_1978,N_47510,N_40411);
and UO_1979 (O_1979,N_43232,N_49333);
or UO_1980 (O_1980,N_46789,N_40317);
xnor UO_1981 (O_1981,N_46157,N_46302);
nor UO_1982 (O_1982,N_44088,N_42693);
nor UO_1983 (O_1983,N_47175,N_48348);
nor UO_1984 (O_1984,N_40541,N_40375);
or UO_1985 (O_1985,N_45795,N_44319);
xnor UO_1986 (O_1986,N_43125,N_48089);
or UO_1987 (O_1987,N_49811,N_44817);
or UO_1988 (O_1988,N_46458,N_48623);
nand UO_1989 (O_1989,N_46940,N_47464);
and UO_1990 (O_1990,N_45928,N_44976);
xor UO_1991 (O_1991,N_45545,N_44417);
nor UO_1992 (O_1992,N_46108,N_42143);
nand UO_1993 (O_1993,N_44214,N_47579);
nor UO_1994 (O_1994,N_45788,N_47390);
nand UO_1995 (O_1995,N_49106,N_46425);
nand UO_1996 (O_1996,N_46629,N_47090);
xor UO_1997 (O_1997,N_45816,N_46265);
or UO_1998 (O_1998,N_48847,N_46131);
or UO_1999 (O_1999,N_49633,N_45877);
and UO_2000 (O_2000,N_43431,N_44085);
nand UO_2001 (O_2001,N_40722,N_47961);
nand UO_2002 (O_2002,N_40882,N_49052);
and UO_2003 (O_2003,N_47136,N_42132);
nor UO_2004 (O_2004,N_40136,N_47945);
nor UO_2005 (O_2005,N_42608,N_46434);
xnor UO_2006 (O_2006,N_40337,N_47433);
nor UO_2007 (O_2007,N_48599,N_40115);
and UO_2008 (O_2008,N_40983,N_40751);
nand UO_2009 (O_2009,N_49916,N_48058);
xor UO_2010 (O_2010,N_43091,N_41854);
nand UO_2011 (O_2011,N_47811,N_42444);
or UO_2012 (O_2012,N_46268,N_41892);
nand UO_2013 (O_2013,N_40684,N_41658);
or UO_2014 (O_2014,N_41069,N_41263);
xor UO_2015 (O_2015,N_42604,N_44025);
and UO_2016 (O_2016,N_48928,N_42534);
nor UO_2017 (O_2017,N_41809,N_43763);
and UO_2018 (O_2018,N_49136,N_48343);
or UO_2019 (O_2019,N_42985,N_43666);
nand UO_2020 (O_2020,N_49747,N_44010);
nand UO_2021 (O_2021,N_40771,N_43087);
xor UO_2022 (O_2022,N_47801,N_45841);
nor UO_2023 (O_2023,N_41811,N_44583);
or UO_2024 (O_2024,N_41941,N_41539);
and UO_2025 (O_2025,N_45446,N_49081);
nand UO_2026 (O_2026,N_48817,N_47419);
or UO_2027 (O_2027,N_49584,N_49846);
or UO_2028 (O_2028,N_47718,N_41062);
and UO_2029 (O_2029,N_45631,N_45737);
nand UO_2030 (O_2030,N_45846,N_45819);
and UO_2031 (O_2031,N_46473,N_42606);
and UO_2032 (O_2032,N_45916,N_47953);
or UO_2033 (O_2033,N_40004,N_44226);
or UO_2034 (O_2034,N_41431,N_43793);
and UO_2035 (O_2035,N_42121,N_44653);
or UO_2036 (O_2036,N_49558,N_45236);
nor UO_2037 (O_2037,N_40246,N_42195);
nand UO_2038 (O_2038,N_42183,N_40668);
or UO_2039 (O_2039,N_42978,N_42845);
xnor UO_2040 (O_2040,N_46530,N_49799);
nand UO_2041 (O_2041,N_48150,N_46304);
or UO_2042 (O_2042,N_44881,N_48902);
nor UO_2043 (O_2043,N_46005,N_46945);
and UO_2044 (O_2044,N_48660,N_40808);
or UO_2045 (O_2045,N_46179,N_49434);
or UO_2046 (O_2046,N_43284,N_41011);
and UO_2047 (O_2047,N_46081,N_43947);
xnor UO_2048 (O_2048,N_48318,N_41261);
nor UO_2049 (O_2049,N_45753,N_47032);
or UO_2050 (O_2050,N_49514,N_41415);
nand UO_2051 (O_2051,N_48583,N_46201);
nand UO_2052 (O_2052,N_49117,N_43551);
and UO_2053 (O_2053,N_41957,N_48624);
or UO_2054 (O_2054,N_49071,N_49270);
or UO_2055 (O_2055,N_44620,N_48394);
nand UO_2056 (O_2056,N_41161,N_47759);
and UO_2057 (O_2057,N_42009,N_41875);
nand UO_2058 (O_2058,N_45583,N_47865);
or UO_2059 (O_2059,N_46000,N_49160);
nor UO_2060 (O_2060,N_42400,N_40958);
nand UO_2061 (O_2061,N_40991,N_46599);
and UO_2062 (O_2062,N_41260,N_42301);
or UO_2063 (O_2063,N_42366,N_41745);
nand UO_2064 (O_2064,N_47799,N_45674);
or UO_2065 (O_2065,N_43707,N_46910);
and UO_2066 (O_2066,N_47944,N_40383);
nand UO_2067 (O_2067,N_44491,N_49484);
nor UO_2068 (O_2068,N_47668,N_43327);
nand UO_2069 (O_2069,N_44897,N_44762);
and UO_2070 (O_2070,N_42426,N_45206);
nand UO_2071 (O_2071,N_46139,N_46446);
nor UO_2072 (O_2072,N_40242,N_43245);
nor UO_2073 (O_2073,N_46605,N_43105);
and UO_2074 (O_2074,N_42924,N_47466);
xor UO_2075 (O_2075,N_45728,N_43591);
nand UO_2076 (O_2076,N_42766,N_40416);
nor UO_2077 (O_2077,N_48371,N_46148);
and UO_2078 (O_2078,N_43345,N_49531);
or UO_2079 (O_2079,N_45721,N_43441);
nor UO_2080 (O_2080,N_46925,N_41084);
nand UO_2081 (O_2081,N_49990,N_48087);
xnor UO_2082 (O_2082,N_49834,N_44045);
and UO_2083 (O_2083,N_43464,N_45657);
and UO_2084 (O_2084,N_40387,N_44929);
nand UO_2085 (O_2085,N_43632,N_43145);
nor UO_2086 (O_2086,N_45263,N_48365);
nor UO_2087 (O_2087,N_48060,N_45761);
and UO_2088 (O_2088,N_42283,N_49836);
xor UO_2089 (O_2089,N_49687,N_43428);
nor UO_2090 (O_2090,N_43079,N_49471);
nor UO_2091 (O_2091,N_41564,N_49330);
xnor UO_2092 (O_2092,N_43318,N_41956);
xnor UO_2093 (O_2093,N_47282,N_49086);
nand UO_2094 (O_2094,N_40071,N_49872);
xor UO_2095 (O_2095,N_45886,N_48965);
nor UO_2096 (O_2096,N_40459,N_41196);
or UO_2097 (O_2097,N_47703,N_42273);
and UO_2098 (O_2098,N_49078,N_45680);
nor UO_2099 (O_2099,N_41475,N_44550);
and UO_2100 (O_2100,N_46334,N_46464);
nor UO_2101 (O_2101,N_42593,N_46449);
xor UO_2102 (O_2102,N_49749,N_48946);
or UO_2103 (O_2103,N_44849,N_43096);
xnor UO_2104 (O_2104,N_49292,N_47099);
and UO_2105 (O_2105,N_44564,N_44382);
or UO_2106 (O_2106,N_46911,N_40295);
and UO_2107 (O_2107,N_49428,N_44156);
and UO_2108 (O_2108,N_47234,N_40462);
or UO_2109 (O_2109,N_40713,N_45983);
nand UO_2110 (O_2110,N_41681,N_45462);
or UO_2111 (O_2111,N_43510,N_43048);
and UO_2112 (O_2112,N_40570,N_47511);
or UO_2113 (O_2113,N_49170,N_47503);
or UO_2114 (O_2114,N_41524,N_41464);
and UO_2115 (O_2115,N_47654,N_45565);
nor UO_2116 (O_2116,N_48038,N_44061);
nor UO_2117 (O_2117,N_48484,N_47397);
or UO_2118 (O_2118,N_44636,N_45457);
and UO_2119 (O_2119,N_45067,N_49323);
or UO_2120 (O_2120,N_40804,N_45349);
nor UO_2121 (O_2121,N_41190,N_42272);
and UO_2122 (O_2122,N_43937,N_40984);
nand UO_2123 (O_2123,N_47107,N_43543);
or UO_2124 (O_2124,N_43101,N_41557);
nor UO_2125 (O_2125,N_44692,N_41624);
nand UO_2126 (O_2126,N_46705,N_45676);
and UO_2127 (O_2127,N_46096,N_43909);
or UO_2128 (O_2128,N_41518,N_45115);
nand UO_2129 (O_2129,N_47968,N_45026);
nand UO_2130 (O_2130,N_42177,N_43157);
or UO_2131 (O_2131,N_41630,N_40324);
nand UO_2132 (O_2132,N_47814,N_44882);
and UO_2133 (O_2133,N_42896,N_47445);
xnor UO_2134 (O_2134,N_40121,N_49444);
and UO_2135 (O_2135,N_46359,N_49576);
xor UO_2136 (O_2136,N_44841,N_49373);
or UO_2137 (O_2137,N_48241,N_46938);
or UO_2138 (O_2138,N_41625,N_42014);
or UO_2139 (O_2139,N_42004,N_42537);
and UO_2140 (O_2140,N_49319,N_47516);
and UO_2141 (O_2141,N_42865,N_48588);
xor UO_2142 (O_2142,N_49504,N_43299);
and UO_2143 (O_2143,N_45433,N_45958);
nand UO_2144 (O_2144,N_40124,N_49389);
nand UO_2145 (O_2145,N_42710,N_48774);
nor UO_2146 (O_2146,N_43943,N_46775);
nor UO_2147 (O_2147,N_40806,N_42308);
and UO_2148 (O_2148,N_44705,N_49403);
nor UO_2149 (O_2149,N_40822,N_41945);
nor UO_2150 (O_2150,N_40856,N_43001);
or UO_2151 (O_2151,N_45505,N_44559);
or UO_2152 (O_2152,N_43406,N_47349);
xnor UO_2153 (O_2153,N_43710,N_47352);
nor UO_2154 (O_2154,N_40362,N_45537);
nand UO_2155 (O_2155,N_42071,N_47914);
or UO_2156 (O_2156,N_45621,N_46015);
and UO_2157 (O_2157,N_40058,N_42095);
nor UO_2158 (O_2158,N_44912,N_48655);
or UO_2159 (O_2159,N_44241,N_44009);
nor UO_2160 (O_2160,N_46140,N_43364);
or UO_2161 (O_2161,N_47927,N_45938);
nand UO_2162 (O_2162,N_41872,N_46068);
or UO_2163 (O_2163,N_40493,N_43119);
nand UO_2164 (O_2164,N_41178,N_46257);
or UO_2165 (O_2165,N_43382,N_49480);
and UO_2166 (O_2166,N_41055,N_44960);
xnor UO_2167 (O_2167,N_41158,N_48319);
and UO_2168 (O_2168,N_47929,N_46503);
and UO_2169 (O_2169,N_45645,N_40768);
and UO_2170 (O_2170,N_40435,N_41358);
and UO_2171 (O_2171,N_45848,N_45724);
and UO_2172 (O_2172,N_45943,N_43289);
or UO_2173 (O_2173,N_43694,N_49703);
nand UO_2174 (O_2174,N_48768,N_41045);
nor UO_2175 (O_2175,N_43568,N_48556);
nand UO_2176 (O_2176,N_44932,N_46234);
nand UO_2177 (O_2177,N_43590,N_48957);
nand UO_2178 (O_2178,N_41778,N_42761);
nor UO_2179 (O_2179,N_41553,N_42464);
or UO_2180 (O_2180,N_41930,N_48451);
nor UO_2181 (O_2181,N_40778,N_45282);
nand UO_2182 (O_2182,N_47104,N_42638);
nor UO_2183 (O_2183,N_43779,N_46465);
and UO_2184 (O_2184,N_43933,N_49246);
nor UO_2185 (O_2185,N_46677,N_45033);
and UO_2186 (O_2186,N_43586,N_43565);
xor UO_2187 (O_2187,N_41739,N_49304);
nor UO_2188 (O_2188,N_47951,N_47719);
nand UO_2189 (O_2189,N_42696,N_46688);
or UO_2190 (O_2190,N_47344,N_42760);
or UO_2191 (O_2191,N_44436,N_48031);
nor UO_2192 (O_2192,N_45404,N_47728);
nand UO_2193 (O_2193,N_42324,N_44682);
and UO_2194 (O_2194,N_47930,N_49155);
xor UO_2195 (O_2195,N_49271,N_40294);
and UO_2196 (O_2196,N_42640,N_48581);
nand UO_2197 (O_2197,N_47897,N_40962);
or UO_2198 (O_2198,N_49070,N_42780);
nand UO_2199 (O_2199,N_47208,N_47791);
xnor UO_2200 (O_2200,N_44566,N_42284);
xnor UO_2201 (O_2201,N_47522,N_45511);
nand UO_2202 (O_2202,N_45169,N_49604);
or UO_2203 (O_2203,N_47678,N_41989);
nand UO_2204 (O_2204,N_43448,N_42681);
nand UO_2205 (O_2205,N_45025,N_48261);
nand UO_2206 (O_2206,N_44487,N_46989);
or UO_2207 (O_2207,N_46678,N_41124);
nor UO_2208 (O_2208,N_48177,N_44598);
nor UO_2209 (O_2209,N_48532,N_43356);
and UO_2210 (O_2210,N_47205,N_49592);
xor UO_2211 (O_2211,N_40443,N_45617);
nor UO_2212 (O_2212,N_42647,N_47943);
and UO_2213 (O_2213,N_47320,N_42953);
and UO_2214 (O_2214,N_46716,N_46427);
or UO_2215 (O_2215,N_44573,N_49137);
or UO_2216 (O_2216,N_45554,N_41197);
and UO_2217 (O_2217,N_40401,N_48409);
or UO_2218 (O_2218,N_43134,N_43333);
nand UO_2219 (O_2219,N_44833,N_44915);
nand UO_2220 (O_2220,N_47960,N_42357);
nand UO_2221 (O_2221,N_42034,N_41707);
nand UO_2222 (O_2222,N_41414,N_45196);
nor UO_2223 (O_2223,N_44342,N_46609);
or UO_2224 (O_2224,N_44934,N_46561);
or UO_2225 (O_2225,N_44962,N_47701);
or UO_2226 (O_2226,N_45464,N_46914);
or UO_2227 (O_2227,N_49801,N_41820);
and UO_2228 (O_2228,N_45939,N_46867);
nor UO_2229 (O_2229,N_46894,N_49167);
nand UO_2230 (O_2230,N_44930,N_47874);
nor UO_2231 (O_2231,N_43093,N_49691);
or UO_2232 (O_2232,N_45007,N_46564);
and UO_2233 (O_2233,N_43409,N_40454);
or UO_2234 (O_2234,N_44175,N_45786);
and UO_2235 (O_2235,N_49282,N_40812);
nor UO_2236 (O_2236,N_40733,N_42688);
nand UO_2237 (O_2237,N_43507,N_43593);
or UO_2238 (O_2238,N_43893,N_44592);
or UO_2239 (O_2239,N_48415,N_44039);
and UO_2240 (O_2240,N_47348,N_48352);
and UO_2241 (O_2241,N_47794,N_44953);
nand UO_2242 (O_2242,N_47591,N_43780);
nand UO_2243 (O_2243,N_49109,N_48967);
and UO_2244 (O_2244,N_44516,N_44092);
and UO_2245 (O_2245,N_46230,N_41104);
xor UO_2246 (O_2246,N_43103,N_41228);
and UO_2247 (O_2247,N_43434,N_46998);
nand UO_2248 (O_2248,N_49138,N_46742);
nand UO_2249 (O_2249,N_49679,N_46555);
nand UO_2250 (O_2250,N_44686,N_42260);
nand UO_2251 (O_2251,N_49168,N_47347);
xnor UO_2252 (O_2252,N_47014,N_41302);
or UO_2253 (O_2253,N_42925,N_44991);
and UO_2254 (O_2254,N_49667,N_45643);
nand UO_2255 (O_2255,N_41799,N_43888);
or UO_2256 (O_2256,N_41031,N_43322);
nor UO_2257 (O_2257,N_43633,N_45134);
and UO_2258 (O_2258,N_43294,N_42870);
nand UO_2259 (O_2259,N_40465,N_44825);
nor UO_2260 (O_2260,N_47517,N_46169);
nand UO_2261 (O_2261,N_43317,N_45449);
nand UO_2262 (O_2262,N_49573,N_41128);
nor UO_2263 (O_2263,N_43861,N_48661);
and UO_2264 (O_2264,N_41461,N_48884);
and UO_2265 (O_2265,N_47030,N_43605);
or UO_2266 (O_2266,N_47321,N_40552);
and UO_2267 (O_2267,N_47691,N_43242);
and UO_2268 (O_2268,N_43170,N_40233);
nand UO_2269 (O_2269,N_42068,N_49556);
and UO_2270 (O_2270,N_48544,N_42579);
xor UO_2271 (O_2271,N_45561,N_42788);
and UO_2272 (O_2272,N_44150,N_47626);
nand UO_2273 (O_2273,N_44956,N_45184);
xor UO_2274 (O_2274,N_41227,N_48494);
nor UO_2275 (O_2275,N_43805,N_47891);
nand UO_2276 (O_2276,N_41743,N_49946);
and UO_2277 (O_2277,N_41411,N_41591);
nand UO_2278 (O_2278,N_46936,N_42861);
or UO_2279 (O_2279,N_48175,N_44718);
xor UO_2280 (O_2280,N_41749,N_40490);
or UO_2281 (O_2281,N_46558,N_41735);
and UO_2282 (O_2282,N_43114,N_45434);
nand UO_2283 (O_2283,N_42184,N_48476);
nor UO_2284 (O_2284,N_49326,N_49101);
nand UO_2285 (O_2285,N_48418,N_47798);
nand UO_2286 (O_2286,N_47570,N_49842);
nor UO_2287 (O_2287,N_48698,N_43626);
xnor UO_2288 (O_2288,N_44965,N_40397);
and UO_2289 (O_2289,N_42670,N_42089);
and UO_2290 (O_2290,N_41676,N_46069);
nand UO_2291 (O_2291,N_45104,N_49422);
xor UO_2292 (O_2292,N_40061,N_46474);
or UO_2293 (O_2293,N_42421,N_46834);
and UO_2294 (O_2294,N_41762,N_46419);
nor UO_2295 (O_2295,N_42069,N_40231);
or UO_2296 (O_2296,N_46432,N_44820);
nor UO_2297 (O_2297,N_49352,N_42059);
nand UO_2298 (O_2298,N_46117,N_45796);
and UO_2299 (O_2299,N_45402,N_49289);
or UO_2300 (O_2300,N_42563,N_48045);
or UO_2301 (O_2301,N_42542,N_42595);
nor UO_2302 (O_2302,N_48143,N_45659);
xnor UO_2303 (O_2303,N_49423,N_48357);
nor UO_2304 (O_2304,N_49740,N_49947);
or UO_2305 (O_2305,N_48176,N_45578);
nand UO_2306 (O_2306,N_43669,N_41357);
xor UO_2307 (O_2307,N_41825,N_40738);
nor UO_2308 (O_2308,N_42278,N_48885);
nor UO_2309 (O_2309,N_40126,N_43971);
or UO_2310 (O_2310,N_47520,N_41734);
and UO_2311 (O_2311,N_49421,N_44737);
and UO_2312 (O_2312,N_49143,N_48574);
nor UO_2313 (O_2313,N_41267,N_49092);
nand UO_2314 (O_2314,N_49322,N_45256);
and UO_2315 (O_2315,N_40208,N_42988);
nand UO_2316 (O_2316,N_47979,N_46086);
or UO_2317 (O_2317,N_40043,N_45531);
xnor UO_2318 (O_2318,N_44558,N_42820);
nand UO_2319 (O_2319,N_41340,N_49674);
and UO_2320 (O_2320,N_47291,N_41179);
or UO_2321 (O_2321,N_47532,N_43703);
nor UO_2322 (O_2322,N_47049,N_43842);
or UO_2323 (O_2323,N_43404,N_47857);
xnor UO_2324 (O_2324,N_41160,N_40488);
nand UO_2325 (O_2325,N_41351,N_48341);
nand UO_2326 (O_2326,N_47300,N_46421);
and UO_2327 (O_2327,N_41604,N_43733);
and UO_2328 (O_2328,N_46573,N_48104);
nand UO_2329 (O_2329,N_45847,N_40385);
nand UO_2330 (O_2330,N_42056,N_42360);
and UO_2331 (O_2331,N_43749,N_40402);
and UO_2332 (O_2332,N_44473,N_49780);
or UO_2333 (O_2333,N_45278,N_48628);
nor UO_2334 (O_2334,N_43935,N_48011);
and UO_2335 (O_2335,N_45422,N_41792);
nor UO_2336 (O_2336,N_41933,N_48301);
nor UO_2337 (O_2337,N_46956,N_47767);
or UO_2338 (O_2338,N_46218,N_48976);
xor UO_2339 (O_2339,N_49510,N_44974);
or UO_2340 (O_2340,N_46380,N_41273);
and UO_2341 (O_2341,N_42941,N_40897);
xor UO_2342 (O_2342,N_44589,N_42230);
nand UO_2343 (O_2343,N_42350,N_49847);
nor UO_2344 (O_2344,N_40964,N_42469);
xnor UO_2345 (O_2345,N_46494,N_43026);
nor UO_2346 (O_2346,N_41481,N_40172);
and UO_2347 (O_2347,N_41971,N_48793);
xor UO_2348 (O_2348,N_43915,N_46695);
and UO_2349 (O_2349,N_47649,N_47116);
nand UO_2350 (O_2350,N_40068,N_44115);
nand UO_2351 (O_2351,N_49111,N_47098);
and UO_2352 (O_2352,N_43437,N_48554);
nand UO_2353 (O_2353,N_49722,N_46691);
nand UO_2354 (O_2354,N_40464,N_45921);
nor UO_2355 (O_2355,N_40135,N_46308);
nand UO_2356 (O_2356,N_47025,N_46546);
xor UO_2357 (O_2357,N_47436,N_49841);
nand UO_2358 (O_2358,N_42860,N_43208);
xor UO_2359 (O_2359,N_46841,N_48323);
or UO_2360 (O_2360,N_41395,N_41652);
nor UO_2361 (O_2361,N_47607,N_42794);
nand UO_2362 (O_2362,N_46892,N_40784);
nor UO_2363 (O_2363,N_43983,N_41352);
and UO_2364 (O_2364,N_45113,N_41985);
or UO_2365 (O_2365,N_49009,N_49657);
nand UO_2366 (O_2366,N_41198,N_49683);
nor UO_2367 (O_2367,N_48787,N_45272);
nor UO_2368 (O_2368,N_44815,N_48729);
or UO_2369 (O_2369,N_49743,N_41499);
or UO_2370 (O_2370,N_43891,N_48461);
xor UO_2371 (O_2371,N_41453,N_41690);
nor UO_2372 (O_2372,N_43160,N_44920);
or UO_2373 (O_2373,N_42020,N_42683);
and UO_2374 (O_2374,N_45376,N_40039);
xor UO_2375 (O_2375,N_44346,N_43381);
or UO_2376 (O_2376,N_42666,N_45425);
nor UO_2377 (O_2377,N_45653,N_43410);
or UO_2378 (O_2378,N_47627,N_49410);
or UO_2379 (O_2379,N_43990,N_47356);
and UO_2380 (O_2380,N_48776,N_48706);
nand UO_2381 (O_2381,N_49851,N_46177);
and UO_2382 (O_2382,N_46595,N_48027);
and UO_2383 (O_2383,N_41381,N_46934);
or UO_2384 (O_2384,N_41147,N_40700);
nand UO_2385 (O_2385,N_49266,N_43646);
nand UO_2386 (O_2386,N_49182,N_48725);
nor UO_2387 (O_2387,N_49378,N_47557);
or UO_2388 (O_2388,N_40286,N_49918);
and UO_2389 (O_2389,N_47434,N_48204);
and UO_2390 (O_2390,N_40220,N_48015);
or UO_2391 (O_2391,N_41777,N_49649);
and UO_2392 (O_2392,N_44742,N_40122);
nand UO_2393 (O_2393,N_49104,N_40450);
or UO_2394 (O_2394,N_43089,N_48830);
nand UO_2395 (O_2395,N_44845,N_46036);
and UO_2396 (O_2396,N_40973,N_44860);
and UO_2397 (O_2397,N_43578,N_47946);
nor UO_2398 (O_2398,N_46795,N_42135);
xor UO_2399 (O_2399,N_47732,N_45499);
nor UO_2400 (O_2400,N_49970,N_41465);
nand UO_2401 (O_2401,N_44582,N_47297);
and UO_2402 (O_2402,N_46794,N_46008);
and UO_2403 (O_2403,N_47997,N_48191);
nor UO_2404 (O_2404,N_49448,N_42179);
nand UO_2405 (O_2405,N_44480,N_46981);
nand UO_2406 (O_2406,N_42300,N_42407);
nor UO_2407 (O_2407,N_44560,N_48658);
nor UO_2408 (O_2408,N_49830,N_43529);
and UO_2409 (O_2409,N_40809,N_40585);
nand UO_2410 (O_2410,N_40206,N_49491);
nand UO_2411 (O_2411,N_40764,N_47537);
nand UO_2412 (O_2412,N_47666,N_44008);
or UO_2413 (O_2413,N_49781,N_41999);
or UO_2414 (O_2414,N_41477,N_49517);
and UO_2415 (O_2415,N_44314,N_45714);
nor UO_2416 (O_2416,N_49585,N_43025);
or UO_2417 (O_2417,N_45186,N_48810);
and UO_2418 (O_2418,N_48813,N_44577);
xnor UO_2419 (O_2419,N_45933,N_41946);
nand UO_2420 (O_2420,N_43979,N_47840);
nand UO_2421 (O_2421,N_45922,N_43625);
and UO_2422 (O_2422,N_45147,N_46669);
and UO_2423 (O_2423,N_49778,N_48165);
or UO_2424 (O_2424,N_45574,N_46377);
nand UO_2425 (O_2425,N_49548,N_40625);
or UO_2426 (O_2426,N_47646,N_46815);
nor UO_2427 (O_2427,N_46762,N_40793);
nor UO_2428 (O_2428,N_48850,N_45575);
and UO_2429 (O_2429,N_43570,N_44481);
nor UO_2430 (O_2430,N_41100,N_42362);
and UO_2431 (O_2431,N_48445,N_43725);
or UO_2432 (O_2432,N_45772,N_41742);
nand UO_2433 (O_2433,N_43532,N_40504);
or UO_2434 (O_2434,N_45097,N_44563);
and UO_2435 (O_2435,N_40228,N_49708);
nor UO_2436 (O_2436,N_41457,N_45556);
nor UO_2437 (O_2437,N_40094,N_49965);
or UO_2438 (O_2438,N_47268,N_45286);
or UO_2439 (O_2439,N_48380,N_48005);
nor UO_2440 (O_2440,N_40076,N_46639);
and UO_2441 (O_2441,N_44106,N_45638);
and UO_2442 (O_2442,N_46995,N_40837);
nor UO_2443 (O_2443,N_44118,N_42416);
or UO_2444 (O_2444,N_47525,N_46018);
and UO_2445 (O_2445,N_44790,N_45103);
nand UO_2446 (O_2446,N_41234,N_40386);
and UO_2447 (O_2447,N_46150,N_41666);
or UO_2448 (O_2448,N_46730,N_40013);
or UO_2449 (O_2449,N_48097,N_42051);
nand UO_2450 (O_2450,N_49537,N_46896);
nor UO_2451 (O_2451,N_43015,N_40350);
and UO_2452 (O_2452,N_48347,N_46978);
and UO_2453 (O_2453,N_49363,N_41638);
and UO_2454 (O_2454,N_49897,N_46803);
and UO_2455 (O_2455,N_47850,N_40012);
or UO_2456 (O_2456,N_41505,N_49544);
nor UO_2457 (O_2457,N_43500,N_49560);
nor UO_2458 (O_2458,N_42996,N_42139);
and UO_2459 (O_2459,N_42344,N_47610);
nor UO_2460 (O_2460,N_44595,N_49655);
nor UO_2461 (O_2461,N_45041,N_42383);
nor UO_2462 (O_2462,N_43991,N_40027);
nor UO_2463 (O_2463,N_49062,N_43314);
nor UO_2464 (O_2464,N_48909,N_48622);
and UO_2465 (O_2465,N_40209,N_48851);
nand UO_2466 (O_2466,N_47628,N_41408);
nor UO_2467 (O_2467,N_47481,N_47768);
and UO_2468 (O_2468,N_44751,N_43537);
and UO_2469 (O_2469,N_41473,N_46506);
and UO_2470 (O_2470,N_47006,N_46199);
nor UO_2471 (O_2471,N_43470,N_48733);
nor UO_2472 (O_2472,N_42435,N_47789);
nand UO_2473 (O_2473,N_41866,N_42571);
or UO_2474 (O_2474,N_41655,N_42347);
or UO_2475 (O_2475,N_49642,N_42566);
or UO_2476 (O_2476,N_41912,N_40288);
xor UO_2477 (O_2477,N_42829,N_41801);
nand UO_2478 (O_2478,N_44063,N_45068);
or UO_2479 (O_2479,N_48210,N_49045);
nor UO_2480 (O_2480,N_46759,N_45723);
or UO_2481 (O_2481,N_47565,N_48812);
nand UO_2482 (O_2482,N_41700,N_45089);
or UO_2483 (O_2483,N_41733,N_46423);
or UO_2484 (O_2484,N_45148,N_42358);
nor UO_2485 (O_2485,N_44223,N_48780);
and UO_2486 (O_2486,N_48128,N_44524);
nand UO_2487 (O_2487,N_43329,N_47345);
nor UO_2488 (O_2488,N_45997,N_48514);
nand UO_2489 (O_2489,N_40780,N_42731);
or UO_2490 (O_2490,N_42168,N_42144);
nand UO_2491 (O_2491,N_48052,N_41516);
nor UO_2492 (O_2492,N_42466,N_44813);
or UO_2493 (O_2493,N_40650,N_45227);
nor UO_2494 (O_2494,N_49386,N_49843);
or UO_2495 (O_2495,N_48073,N_44476);
and UO_2496 (O_2496,N_43191,N_49577);
nand UO_2497 (O_2497,N_46115,N_48452);
nand UO_2498 (O_2498,N_47866,N_41082);
nand UO_2499 (O_2499,N_46676,N_46404);
and UO_2500 (O_2500,N_40798,N_46864);
nand UO_2501 (O_2501,N_40623,N_48616);
xnor UO_2502 (O_2502,N_45438,N_48694);
xor UO_2503 (O_2503,N_42572,N_47881);
nor UO_2504 (O_2504,N_41774,N_44231);
or UO_2505 (O_2505,N_41429,N_40216);
nand UO_2506 (O_2506,N_41175,N_41840);
and UO_2507 (O_2507,N_41405,N_41360);
nand UO_2508 (O_2508,N_40794,N_49931);
nor UO_2509 (O_2509,N_40305,N_43934);
nor UO_2510 (O_2510,N_40296,N_41174);
nor UO_2511 (O_2511,N_42818,N_47876);
nand UO_2512 (O_2512,N_43465,N_45707);
or UO_2513 (O_2513,N_44865,N_43520);
nor UO_2514 (O_2514,N_49226,N_45127);
nor UO_2515 (O_2515,N_49808,N_49706);
or UO_2516 (O_2516,N_44134,N_44459);
or UO_2517 (O_2517,N_47067,N_42636);
or UO_2518 (O_2518,N_45381,N_46642);
and UO_2519 (O_2519,N_49646,N_44219);
or UO_2520 (O_2520,N_46221,N_42738);
xnor UO_2521 (O_2521,N_40735,N_44001);
xnor UO_2522 (O_2522,N_49880,N_41454);
or UO_2523 (O_2523,N_40008,N_41243);
nand UO_2524 (O_2524,N_44284,N_42971);
nor UO_2525 (O_2525,N_42707,N_42257);
and UO_2526 (O_2526,N_47849,N_44152);
and UO_2527 (O_2527,N_49926,N_48338);
nand UO_2528 (O_2528,N_45984,N_48291);
nor UO_2529 (O_2529,N_42918,N_49610);
nand UO_2530 (O_2530,N_45688,N_45042);
and UO_2531 (O_2531,N_48040,N_46013);
nor UO_2532 (O_2532,N_43108,N_44687);
nor UO_2533 (O_2533,N_46889,N_41542);
nand UO_2534 (O_2534,N_43997,N_44933);
nor UO_2535 (O_2535,N_40024,N_40353);
and UO_2536 (O_2536,N_41379,N_42626);
and UO_2537 (O_2537,N_48477,N_42218);
and UO_2538 (O_2538,N_48796,N_45778);
nand UO_2539 (O_2539,N_46093,N_41452);
and UO_2540 (O_2540,N_46164,N_45232);
or UO_2541 (O_2541,N_49206,N_43803);
nor UO_2542 (O_2542,N_40855,N_45479);
and UO_2543 (O_2543,N_45118,N_47905);
xor UO_2544 (O_2544,N_48602,N_47275);
nand UO_2545 (O_2545,N_48426,N_43485);
or UO_2546 (O_2546,N_45534,N_48353);
nor UO_2547 (O_2547,N_49358,N_42679);
and UO_2548 (O_2548,N_40239,N_45814);
or UO_2549 (O_2549,N_40368,N_44205);
and UO_2550 (O_2550,N_40950,N_47896);
nor UO_2551 (O_2551,N_47583,N_45960);
xnor UO_2552 (O_2552,N_48996,N_40451);
nor UO_2553 (O_2553,N_41546,N_42470);
or UO_2554 (O_2554,N_40104,N_45341);
or UO_2555 (O_2555,N_48460,N_46135);
and UO_2556 (O_2556,N_43009,N_42211);
nand UO_2557 (O_2557,N_44213,N_47430);
or UO_2558 (O_2558,N_40846,N_43219);
or UO_2559 (O_2559,N_46817,N_40561);
nor UO_2560 (O_2560,N_43099,N_49317);
and UO_2561 (O_2561,N_45787,N_44530);
or UO_2562 (O_2562,N_44741,N_42170);
nand UO_2563 (O_2563,N_44921,N_48639);
and UO_2564 (O_2564,N_41230,N_42512);
xnor UO_2565 (O_2565,N_49699,N_42062);
nand UO_2566 (O_2566,N_41116,N_48997);
nor UO_2567 (O_2567,N_40593,N_43457);
and UO_2568 (O_2568,N_49240,N_43285);
xor UO_2569 (O_2569,N_46400,N_41338);
and UO_2570 (O_2570,N_45166,N_42527);
and UO_2571 (O_2571,N_40982,N_41316);
and UO_2572 (O_2572,N_44405,N_47123);
nor UO_2573 (O_2573,N_41173,N_46307);
and UO_2574 (O_2574,N_47199,N_48454);
or UO_2575 (O_2575,N_42733,N_42849);
and UO_2576 (O_2576,N_41540,N_47005);
and UO_2577 (O_2577,N_45995,N_48216);
or UO_2578 (O_2578,N_49714,N_45197);
xor UO_2579 (O_2579,N_40583,N_45649);
and UO_2580 (O_2580,N_46597,N_41047);
or UO_2581 (O_2581,N_41298,N_43244);
and UO_2582 (O_2582,N_44601,N_45797);
nor UO_2583 (O_2583,N_42615,N_42459);
nand UO_2584 (O_2584,N_49483,N_43610);
or UO_2585 (O_2585,N_47173,N_43034);
nand UO_2586 (O_2586,N_49726,N_40157);
nand UO_2587 (O_2587,N_42510,N_43927);
and UO_2588 (O_2588,N_40549,N_49724);
or UO_2589 (O_2589,N_49325,N_48138);
nand UO_2590 (O_2590,N_49507,N_47821);
nor UO_2591 (O_2591,N_47596,N_45644);
or UO_2592 (O_2592,N_48303,N_45734);
xnor UO_2593 (O_2593,N_49745,N_40282);
nor UO_2594 (O_2594,N_46887,N_47817);
and UO_2595 (O_2595,N_46947,N_47906);
xor UO_2596 (O_2596,N_46625,N_49295);
or UO_2597 (O_2597,N_49589,N_45173);
or UO_2598 (O_2598,N_44875,N_47696);
and UO_2599 (O_2599,N_49605,N_44968);
nor UO_2600 (O_2600,N_47957,N_45770);
and UO_2601 (O_2601,N_41565,N_41867);
or UO_2602 (O_2602,N_43019,N_42875);
xor UO_2603 (O_2603,N_45906,N_44794);
and UO_2604 (O_2604,N_40920,N_47713);
and UO_2605 (O_2605,N_49315,N_45956);
and UO_2606 (O_2606,N_49819,N_41589);
nor UO_2607 (O_2607,N_42096,N_42894);
nand UO_2608 (O_2608,N_42430,N_47909);
or UO_2609 (O_2609,N_41530,N_47514);
nor UO_2610 (O_2610,N_49732,N_41598);
or UO_2611 (O_2611,N_45950,N_48524);
or UO_2612 (O_2612,N_45654,N_45081);
nor UO_2613 (O_2613,N_49597,N_45937);
nand UO_2614 (O_2614,N_46029,N_48103);
and UO_2615 (O_2615,N_44646,N_45260);
xnor UO_2616 (O_2616,N_46987,N_49189);
nand UO_2617 (O_2617,N_48198,N_45006);
nor UO_2618 (O_2618,N_41511,N_45903);
and UO_2619 (O_2619,N_40110,N_49975);
and UO_2620 (O_2620,N_44493,N_41826);
or UO_2621 (O_2621,N_44496,N_45412);
or UO_2622 (O_2622,N_48667,N_42764);
or UO_2623 (O_2623,N_49913,N_42452);
nor UO_2624 (O_2624,N_48720,N_43315);
and UO_2625 (O_2625,N_41221,N_43078);
xor UO_2626 (O_2626,N_48775,N_41882);
or UO_2627 (O_2627,N_44273,N_40021);
nor UO_2628 (O_2628,N_48664,N_40581);
and UO_2629 (O_2629,N_49412,N_43953);
nand UO_2630 (O_2630,N_41759,N_47729);
nand UO_2631 (O_2631,N_45591,N_46786);
or UO_2632 (O_2632,N_43416,N_41525);
or UO_2633 (O_2633,N_41537,N_46630);
nand UO_2634 (O_2634,N_40759,N_45606);
nor UO_2635 (O_2635,N_43494,N_40813);
xnor UO_2636 (O_2636,N_49572,N_45791);
xnor UO_2637 (O_2637,N_48900,N_45361);
and UO_2638 (O_2638,N_44352,N_46738);
nand UO_2639 (O_2639,N_44121,N_49201);
nor UO_2640 (O_2640,N_45948,N_45043);
nand UO_2641 (O_2641,N_40923,N_49595);
and UO_2642 (O_2642,N_48559,N_42689);
nand UO_2643 (O_2643,N_42164,N_46054);
nand UO_2644 (O_2644,N_47551,N_40589);
or UO_2645 (O_2645,N_40334,N_42309);
nand UO_2646 (O_2646,N_45321,N_40929);
or UO_2647 (O_2647,N_45102,N_43184);
nor UO_2648 (O_2648,N_43330,N_45280);
and UO_2649 (O_2649,N_40857,N_43900);
and UO_2650 (O_2650,N_46242,N_43306);
and UO_2651 (O_2651,N_45325,N_42601);
and UO_2652 (O_2652,N_42994,N_46870);
nand UO_2653 (O_2653,N_46200,N_41331);
xor UO_2654 (O_2654,N_42886,N_49955);
nor UO_2655 (O_2655,N_45242,N_42504);
and UO_2656 (O_2656,N_47296,N_40301);
or UO_2657 (O_2657,N_47069,N_44578);
nand UO_2658 (O_2658,N_47330,N_40469);
and UO_2659 (O_2659,N_44340,N_45989);
nand UO_2660 (O_2660,N_44562,N_45246);
nor UO_2661 (O_2661,N_41994,N_41651);
xor UO_2662 (O_2662,N_48396,N_43341);
nand UO_2663 (O_2663,N_46061,N_41181);
or UO_2664 (O_2664,N_47187,N_46326);
nor UO_2665 (O_2665,N_41695,N_43220);
nand UO_2666 (O_2666,N_46297,N_40989);
or UO_2667 (O_2667,N_47497,N_45474);
and UO_2668 (O_2668,N_45178,N_43658);
and UO_2669 (O_2669,N_47699,N_41010);
and UO_2670 (O_2670,N_40754,N_46964);
nor UO_2671 (O_2671,N_48533,N_46267);
nand UO_2672 (O_2672,N_41186,N_42345);
or UO_2673 (O_2673,N_48565,N_46030);
nor UO_2674 (O_2674,N_49654,N_48595);
or UO_2675 (O_2675,N_48019,N_44166);
nand UO_2676 (O_2676,N_45108,N_40906);
nor UO_2677 (O_2677,N_45050,N_47871);
nand UO_2678 (O_2678,N_44590,N_43662);
xnor UO_2679 (O_2679,N_44246,N_43685);
or UO_2680 (O_2680,N_44269,N_46854);
and UO_2681 (O_2681,N_43002,N_42789);
or UO_2682 (O_2682,N_43678,N_48758);
xor UO_2683 (O_2683,N_43531,N_48730);
or UO_2684 (O_2684,N_48547,N_42011);
nand UO_2685 (O_2685,N_40951,N_43067);
or UO_2686 (O_2686,N_48752,N_46299);
or UO_2687 (O_2687,N_42883,N_44188);
or UO_2688 (O_2688,N_48298,N_44840);
xnor UO_2689 (O_2689,N_40928,N_46224);
and UO_2690 (O_2690,N_41940,N_47454);
and UO_2691 (O_2691,N_42973,N_44196);
nand UO_2692 (O_2692,N_46844,N_42944);
nand UO_2693 (O_2693,N_48856,N_49879);
nor UO_2694 (O_2694,N_44828,N_45034);
or UO_2695 (O_2695,N_48340,N_45001);
and UO_2696 (O_2696,N_42805,N_43930);
nor UO_2697 (O_2697,N_46144,N_45305);
nor UO_2698 (O_2698,N_48333,N_40654);
nor UO_2699 (O_2699,N_47253,N_43303);
xor UO_2700 (O_2700,N_42399,N_47380);
nand UO_2701 (O_2701,N_49374,N_48497);
and UO_2702 (O_2702,N_42086,N_46390);
nor UO_2703 (O_2703,N_44064,N_45443);
and UO_2704 (O_2704,N_44047,N_44812);
nand UO_2705 (O_2705,N_43748,N_46711);
and UO_2706 (O_2706,N_42687,N_45413);
nand UO_2707 (O_2707,N_41437,N_44659);
nor UO_2708 (O_2708,N_44623,N_49485);
or UO_2709 (O_2709,N_40935,N_42171);
and UO_2710 (O_2710,N_43391,N_48256);
or UO_2711 (O_2711,N_41120,N_49435);
nor UO_2712 (O_2712,N_41657,N_40051);
or UO_2713 (O_2713,N_44909,N_46552);
and UO_2714 (O_2714,N_42103,N_49022);
or UO_2715 (O_2715,N_45766,N_41754);
nand UO_2716 (O_2716,N_47869,N_40590);
nor UO_2717 (O_2717,N_46661,N_43224);
nand UO_2718 (O_2718,N_49019,N_44238);
and UO_2719 (O_2719,N_44164,N_44318);
nor UO_2720 (O_2720,N_47775,N_43321);
nor UO_2721 (O_2721,N_43389,N_44129);
and UO_2722 (O_2722,N_42881,N_47690);
nand UO_2723 (O_2723,N_49718,N_47462);
nand UO_2724 (O_2724,N_44099,N_42943);
nor UO_2725 (O_2725,N_40701,N_47122);
xor UO_2726 (O_2726,N_43744,N_45021);
xnor UO_2727 (O_2727,N_44832,N_42212);
and UO_2728 (O_2728,N_41744,N_49453);
or UO_2729 (O_2729,N_45091,N_44183);
nor UO_2730 (O_2730,N_41614,N_48246);
and UO_2731 (O_2731,N_43225,N_42091);
nand UO_2732 (O_2732,N_42146,N_42117);
and UO_2733 (O_2733,N_47546,N_42254);
nand UO_2734 (O_2734,N_48721,N_46333);
nor UO_2735 (O_2735,N_47810,N_41402);
nand UO_2736 (O_2736,N_47381,N_40258);
or UO_2737 (O_2737,N_43056,N_40727);
or UO_2738 (O_2738,N_49099,N_45035);
nor UO_2739 (O_2739,N_41049,N_42926);
and UO_2740 (O_2740,N_48908,N_46970);
or UO_2741 (O_2741,N_40256,N_41855);
or UO_2742 (O_2742,N_48267,N_43313);
nand UO_2743 (O_2743,N_48930,N_40957);
or UO_2744 (O_2744,N_48412,N_42045);
nor UO_2745 (O_2745,N_47576,N_48827);
nor UO_2746 (O_2746,N_44043,N_40339);
nand UO_2747 (O_2747,N_40323,N_43824);
nand UO_2748 (O_2748,N_46557,N_42502);
nand UO_2749 (O_2749,N_48134,N_47285);
or UO_2750 (O_2750,N_40745,N_45228);
and UO_2751 (O_2751,N_40453,N_49673);
or UO_2752 (O_2752,N_48714,N_44941);
xor UO_2753 (O_2753,N_42280,N_49559);
xnor UO_2754 (O_2754,N_40229,N_41365);
nand UO_2755 (O_2755,N_43073,N_41169);
or UO_2756 (O_2756,N_46394,N_44717);
nor UO_2757 (O_2757,N_40726,N_43332);
nand UO_2758 (O_2758,N_45110,N_48100);
xor UO_2759 (O_2759,N_47894,N_40003);
nand UO_2760 (O_2760,N_47213,N_41991);
or UO_2761 (O_2761,N_48345,N_44027);
xor UO_2762 (O_2762,N_49869,N_45175);
nand UO_2763 (O_2763,N_40514,N_48050);
xnor UO_2764 (O_2764,N_47730,N_46702);
nor UO_2765 (O_2765,N_47887,N_40995);
nor UO_2766 (O_2766,N_42627,N_48609);
nor UO_2767 (O_2767,N_42714,N_43862);
or UO_2768 (O_2768,N_47884,N_48958);
or UO_2769 (O_2769,N_49195,N_44855);
nand UO_2770 (O_2770,N_46850,N_47609);
nand UO_2771 (O_2771,N_49922,N_44652);
or UO_2772 (O_2772,N_44532,N_45130);
nand UO_2773 (O_2773,N_40089,N_42630);
or UO_2774 (O_2774,N_41199,N_44985);
xnor UO_2775 (O_2775,N_47096,N_47450);
xnor UO_2776 (O_2776,N_40475,N_43695);
nor UO_2777 (O_2777,N_43007,N_40467);
or UO_2778 (O_2778,N_46455,N_46856);
or UO_2779 (O_2779,N_47387,N_41566);
nor UO_2780 (O_2780,N_48095,N_41494);
or UO_2781 (O_2781,N_44748,N_44434);
xor UO_2782 (O_2782,N_40872,N_43672);
nand UO_2783 (O_2783,N_45250,N_49547);
nand UO_2784 (O_2784,N_42837,N_40767);
nand UO_2785 (O_2785,N_46214,N_42085);
xnor UO_2786 (O_2786,N_40791,N_40430);
nand UO_2787 (O_2787,N_49445,N_49686);
and UO_2788 (O_2788,N_46505,N_48809);
nand UO_2789 (O_2789,N_48254,N_43298);
nand UO_2790 (O_2790,N_41406,N_44527);
and UO_2791 (O_2791,N_40868,N_49758);
nand UO_2792 (O_2792,N_44539,N_44248);
or UO_2793 (O_2793,N_40534,N_42882);
and UO_2794 (O_2794,N_44108,N_47449);
and UO_2795 (O_2795,N_45150,N_41864);
or UO_2796 (O_2796,N_45441,N_45904);
nand UO_2797 (O_2797,N_41596,N_46592);
nand UO_2798 (O_2798,N_48956,N_45116);
nand UO_2799 (O_2799,N_46217,N_48163);
xor UO_2800 (O_2800,N_44557,N_44387);
nor UO_2801 (O_2801,N_48765,N_41904);
nand UO_2802 (O_2802,N_44657,N_43847);
nand UO_2803 (O_2803,N_46371,N_43484);
nor UO_2804 (O_2804,N_46228,N_43334);
or UO_2805 (O_2805,N_43757,N_45581);
nand UO_2806 (O_2806,N_40690,N_43756);
and UO_2807 (O_2807,N_44947,N_43583);
and UO_2808 (O_2808,N_49204,N_42635);
nand UO_2809 (O_2809,N_47833,N_47507);
xnor UO_2810 (O_2810,N_48564,N_44245);
nor UO_2811 (O_2811,N_47183,N_40244);
nand UO_2812 (O_2812,N_41380,N_49110);
nor UO_2813 (O_2813,N_42269,N_49262);
or UO_2814 (O_2814,N_49772,N_44247);
and UO_2815 (O_2815,N_46355,N_41550);
xor UO_2816 (O_2816,N_42198,N_49293);
and UO_2817 (O_2817,N_41896,N_43014);
or UO_2818 (O_2818,N_46125,N_40348);
and UO_2819 (O_2819,N_49150,N_48466);
nor UO_2820 (O_2820,N_42976,N_45855);
or UO_2821 (O_2821,N_44768,N_46050);
nand UO_2822 (O_2822,N_40142,N_48840);
or UO_2823 (O_2823,N_45357,N_48598);
nand UO_2824 (O_2824,N_47645,N_46198);
or UO_2825 (O_2825,N_40891,N_46778);
nand UO_2826 (O_2826,N_44144,N_43684);
xnor UO_2827 (O_2827,N_48822,N_41848);
nor UO_2828 (O_2828,N_46165,N_43110);
or UO_2829 (O_2829,N_46891,N_42436);
and UO_2830 (O_2830,N_44979,N_46878);
and UO_2831 (O_2831,N_48275,N_43196);
nor UO_2832 (O_2832,N_40945,N_47643);
or UO_2833 (O_2833,N_46448,N_43873);
xor UO_2834 (O_2834,N_48053,N_43088);
xor UO_2835 (O_2835,N_43908,N_40026);
nand UO_2836 (O_2836,N_44847,N_49238);
or UO_2837 (O_2837,N_44631,N_46783);
nor UO_2838 (O_2838,N_47676,N_41070);
xor UO_2839 (O_2839,N_43413,N_46681);
nand UO_2840 (O_2840,N_45299,N_49190);
or UO_2841 (O_2841,N_49037,N_46748);
nor UO_2842 (O_2842,N_45726,N_48378);
and UO_2843 (O_2843,N_43136,N_48231);
and UO_2844 (O_2844,N_48239,N_45205);
and UO_2845 (O_2845,N_43213,N_41521);
nor UO_2846 (O_2846,N_48843,N_42275);
nand UO_2847 (O_2847,N_42307,N_46413);
nand UO_2848 (O_2848,N_44240,N_48805);
and UO_2849 (O_2849,N_42355,N_49612);
nand UO_2850 (O_2850,N_44389,N_48876);
nor UO_2851 (O_2851,N_47293,N_40409);
and UO_2852 (O_2852,N_40240,N_41609);
nor UO_2853 (O_2853,N_49399,N_41443);
or UO_2854 (O_2854,N_42833,N_43782);
or UO_2855 (O_2855,N_41928,N_40396);
xor UO_2856 (O_2856,N_48117,N_48728);
and UO_2857 (O_2857,N_49889,N_41078);
nor UO_2858 (O_2858,N_47541,N_43118);
or UO_2859 (O_2859,N_43352,N_40693);
or UO_2860 (O_2860,N_46957,N_40961);
or UO_2861 (O_2861,N_43340,N_42417);
nand UO_2862 (O_2862,N_45396,N_46574);
and UO_2863 (O_2863,N_43251,N_43053);
nor UO_2864 (O_2864,N_44838,N_43649);
and UO_2865 (O_2865,N_48666,N_43761);
nor UO_2866 (O_2866,N_46282,N_47159);
and UO_2867 (O_2867,N_49746,N_49342);
and UO_2868 (O_2868,N_46572,N_46447);
or UO_2869 (O_2869,N_43773,N_49237);
xnor UO_2870 (O_2870,N_47411,N_48443);
and UO_2871 (O_2871,N_49265,N_47401);
nor UO_2872 (O_2872,N_43925,N_41252);
nand UO_2873 (O_2873,N_43290,N_45507);
or UO_2874 (O_2874,N_42252,N_48129);
nand UO_2875 (O_2875,N_45079,N_41888);
or UO_2876 (O_2876,N_42539,N_44315);
nand UO_2877 (O_2877,N_48592,N_46766);
or UO_2878 (O_2878,N_43247,N_48439);
or UO_2879 (O_2879,N_41485,N_49760);
and UO_2880 (O_2880,N_46330,N_48188);
and UO_2881 (O_2881,N_44535,N_40766);
nor UO_2882 (O_2882,N_43673,N_40605);
nor UO_2883 (O_2883,N_49463,N_41072);
and UO_2884 (O_2884,N_42701,N_45315);
nand UO_2885 (O_2885,N_41577,N_46075);
and UO_2886 (O_2886,N_43835,N_44536);
and UO_2887 (O_2887,N_45472,N_44616);
and UO_2888 (O_2888,N_47950,N_48232);
xnor UO_2889 (O_2889,N_46219,N_46134);
nand UO_2890 (O_2890,N_41917,N_43495);
and UO_2891 (O_2891,N_44761,N_49244);
nand UO_2892 (O_2892,N_42867,N_41239);
nor UO_2893 (O_2893,N_48151,N_42782);
xnor UO_2894 (O_2894,N_42341,N_44006);
or UO_2895 (O_2895,N_46095,N_43279);
or UO_2896 (O_2896,N_43790,N_43505);
xnor UO_2897 (O_2897,N_47774,N_44286);
xor UO_2898 (O_2898,N_47399,N_49586);
and UO_2899 (O_2899,N_47875,N_40869);
nand UO_2900 (O_2900,N_45620,N_40433);
or UO_2901 (O_2901,N_41079,N_40084);
and UO_2902 (O_2902,N_45504,N_43140);
nand UO_2903 (O_2903,N_40251,N_40069);
and UO_2904 (O_2904,N_44325,N_46361);
and UO_2905 (O_2905,N_45082,N_42767);
or UO_2906 (O_2906,N_44844,N_49886);
and UO_2907 (O_2907,N_40655,N_46746);
or UO_2908 (O_2908,N_40053,N_42558);
nand UO_2909 (O_2909,N_46275,N_45720);
xor UO_2910 (O_2910,N_41532,N_44534);
nand UO_2911 (O_2911,N_46581,N_48589);
or UO_2912 (O_2912,N_45160,N_47121);
nor UO_2913 (O_2913,N_45181,N_40214);
or UO_2914 (O_2914,N_49043,N_47078);
xor UO_2915 (O_2915,N_44642,N_40389);
nor UO_2916 (O_2916,N_46532,N_41827);
nand UO_2917 (O_2917,N_41543,N_43287);
nand UO_2918 (O_2918,N_48159,N_44711);
or UO_2919 (O_2919,N_43124,N_49181);
nand UO_2920 (O_2920,N_42310,N_43388);
nor UO_2921 (O_2921,N_44100,N_45509);
xnor UO_2922 (O_2922,N_46958,N_47188);
xnor UO_2923 (O_2923,N_46403,N_40518);
or UO_2924 (O_2924,N_48971,N_41152);
nand UO_2925 (O_2925,N_42950,N_41723);
or UO_2926 (O_2926,N_49571,N_49247);
and UO_2927 (O_2927,N_41926,N_40359);
nor UO_2928 (O_2928,N_45415,N_49015);
nor UO_2929 (O_2929,N_47528,N_45073);
nor UO_2930 (O_2930,N_49753,N_49848);
and UO_2931 (O_2931,N_40091,N_47238);
and UO_2932 (O_2932,N_48481,N_43919);
or UO_2933 (O_2933,N_41203,N_44914);
and UO_2934 (O_2934,N_49409,N_47000);
nand UO_2935 (O_2935,N_40737,N_46690);
nor UO_2936 (O_2936,N_44680,N_40055);
nor UO_2937 (O_2937,N_45170,N_46634);
nor UO_2938 (O_2938,N_44510,N_42659);
or UO_2939 (O_2939,N_40988,N_42304);
nand UO_2940 (O_2940,N_44362,N_47531);
nor UO_2941 (O_2941,N_48676,N_40505);
or UO_2942 (O_2942,N_48498,N_40582);
or UO_2943 (O_2943,N_40152,N_45792);
and UO_2944 (O_2944,N_45010,N_45277);
nor UO_2945 (O_2945,N_42110,N_47547);
xor UO_2946 (O_2946,N_44031,N_46246);
and UO_2947 (O_2947,N_49450,N_42554);
nand UO_2948 (O_2948,N_46689,N_47812);
nor UO_2949 (O_2949,N_40648,N_43194);
and UO_2950 (O_2950,N_48491,N_43357);
xnor UO_2951 (O_2951,N_46102,N_45302);
xor UO_2952 (O_2952,N_46744,N_44354);
and UO_2953 (O_2953,N_40854,N_44087);
nand UO_2954 (O_2954,N_45183,N_48951);
nand UO_2955 (O_2955,N_49455,N_40218);
or UO_2956 (O_2956,N_44716,N_41172);
nor UO_2957 (O_2957,N_43629,N_43497);
xnor UO_2958 (O_2958,N_42722,N_41514);
nand UO_2959 (O_2959,N_49731,N_46519);
nor UO_2960 (O_2960,N_40535,N_42007);
or UO_2961 (O_2961,N_45535,N_42851);
nor UO_2962 (O_2962,N_43398,N_46578);
nor UO_2963 (O_2963,N_44522,N_48455);
nor UO_2964 (O_2964,N_49702,N_47877);
nand UO_2965 (O_2965,N_41654,N_45571);
or UO_2966 (O_2966,N_43759,N_47274);
xnor UO_2967 (O_2967,N_47619,N_46699);
xnor UO_2968 (O_2968,N_41150,N_45310);
nor UO_2969 (O_2969,N_49653,N_47150);
nand UO_2970 (O_2970,N_46133,N_46070);
nand UO_2971 (O_2971,N_40303,N_47393);
nand UO_2972 (O_2972,N_45716,N_44570);
nand UO_2973 (O_2973,N_43918,N_49858);
or UO_2974 (O_2974,N_46339,N_40952);
nand UO_2975 (O_2975,N_40099,N_44184);
xor UO_2976 (O_2976,N_45309,N_46972);
nor UO_2977 (O_2977,N_47708,N_49516);
nor UO_2978 (O_2978,N_40431,N_47458);
and UO_2979 (O_2979,N_47114,N_44639);
or UO_2980 (O_2980,N_47765,N_48197);
or UO_2981 (O_2981,N_43068,N_41979);
and UO_2982 (O_2982,N_48932,N_49284);
nand UO_2983 (O_2983,N_45030,N_42293);
or UO_2984 (O_2984,N_48941,N_41915);
and UO_2985 (O_2985,N_43461,N_46656);
nor UO_2986 (O_2986,N_44107,N_43183);
nand UO_2987 (O_2987,N_42261,N_43885);
nand UO_2988 (O_2988,N_47153,N_42361);
nand UO_2989 (O_2989,N_40914,N_43098);
and UO_2990 (O_2990,N_42160,N_45776);
nor UO_2991 (O_2991,N_49803,N_41758);
and UO_2992 (O_2992,N_49297,N_42138);
or UO_2993 (O_2993,N_41336,N_43525);
and UO_2994 (O_2994,N_41308,N_49344);
nor UO_2995 (O_2995,N_41730,N_49392);
nor UO_2996 (O_2996,N_49696,N_43350);
and UO_2997 (O_2997,N_43527,N_46438);
or UO_2998 (O_2998,N_43635,N_44169);
nand UO_2999 (O_2999,N_45687,N_46929);
nor UO_3000 (O_3000,N_47650,N_42336);
or UO_3001 (O_3001,N_44431,N_48305);
nor UO_3002 (O_3002,N_41862,N_40197);
or UO_3003 (O_3003,N_42210,N_43355);
and UO_3004 (O_3004,N_41255,N_40367);
or UO_3005 (O_3005,N_45589,N_40719);
and UO_3006 (O_3006,N_46515,N_43535);
nor UO_3007 (O_3007,N_42377,N_40513);
or UO_3008 (O_3008,N_47385,N_44588);
nor UO_3009 (O_3009,N_41459,N_48014);
and UO_3010 (O_3010,N_46517,N_44225);
nand UO_3011 (O_3011,N_46839,N_47956);
xnor UO_3012 (O_3012,N_41562,N_44359);
xnor UO_3013 (O_3013,N_40065,N_45491);
nor UO_3014 (O_3014,N_42266,N_44174);
nand UO_3015 (O_3015,N_48849,N_42112);
nand UO_3016 (O_3016,N_43012,N_46010);
nor UO_3017 (O_3017,N_46245,N_48869);
nand UO_3018 (O_3018,N_41520,N_47475);
or UO_3019 (O_3019,N_47323,N_47215);
xor UO_3020 (O_3020,N_45368,N_44879);
and UO_3021 (O_3021,N_40308,N_40144);
and UO_3022 (O_3022,N_47715,N_47941);
nor UO_3023 (O_3023,N_41629,N_48035);
or UO_3024 (O_3024,N_40320,N_47266);
nand UO_3025 (O_3025,N_49962,N_41641);
and UO_3026 (O_3026,N_47633,N_41526);
or UO_3027 (O_3027,N_46463,N_49272);
nor UO_3028 (O_3028,N_42256,N_46362);
and UO_3029 (O_3029,N_42892,N_47059);
or UO_3030 (O_3030,N_43881,N_49763);
nor UO_3031 (O_3031,N_49765,N_45397);
nand UO_3032 (O_3032,N_42327,N_41580);
nor UO_3033 (O_3033,N_42107,N_46619);
xnor UO_3034 (O_3034,N_43974,N_49360);
nor UO_3035 (O_3035,N_45539,N_47722);
nand UO_3036 (O_3036,N_49950,N_44945);
nand UO_3037 (O_3037,N_49139,N_45214);
xnor UO_3038 (O_3038,N_48683,N_46904);
nor UO_3039 (O_3039,N_47813,N_46836);
and UO_3040 (O_3040,N_42961,N_42070);
nor UO_3041 (O_3041,N_41322,N_47307);
nor UO_3042 (O_3042,N_46244,N_41294);
nor UO_3043 (O_3043,N_40098,N_43957);
or UO_3044 (O_3044,N_48801,N_44355);
nand UO_3045 (O_3045,N_41823,N_49993);
or UO_3046 (O_3046,N_47663,N_47982);
nor UO_3047 (O_3047,N_48652,N_49006);
nor UO_3048 (O_3048,N_43584,N_40255);
or UO_3049 (O_3049,N_42010,N_43829);
and UO_3050 (O_3050,N_46109,N_45601);
xnor UO_3051 (O_3051,N_46431,N_47593);
nor UO_3052 (O_3052,N_40057,N_47842);
xnor UO_3053 (O_3053,N_46583,N_49179);
nand UO_3054 (O_3054,N_48140,N_47146);
nand UO_3055 (O_3055,N_46968,N_47342);
or UO_3056 (O_3056,N_44967,N_41384);
or UO_3057 (O_3057,N_45379,N_47824);
xnor UO_3058 (O_3058,N_47335,N_47815);
or UO_3059 (O_3059,N_40850,N_46802);
nand UO_3060 (O_3060,N_44189,N_41517);
xnor UO_3061 (O_3061,N_48961,N_43223);
xor UO_3062 (O_3062,N_43708,N_43082);
or UO_3063 (O_3063,N_40938,N_48044);
xnor UO_3064 (O_3064,N_42039,N_41215);
and UO_3065 (O_3065,N_48047,N_40045);
nor UO_3066 (O_3066,N_49903,N_44936);
and UO_3067 (O_3067,N_47880,N_48578);
or UO_3068 (O_3068,N_44602,N_48964);
nor UO_3069 (O_3069,N_47639,N_41361);
and UO_3070 (O_3070,N_40165,N_42824);
nand UO_3071 (O_3071,N_42952,N_42735);
xor UO_3072 (O_3072,N_48363,N_41009);
and UO_3073 (O_3073,N_48209,N_44744);
nand UO_3074 (O_3074,N_42927,N_42109);
or UO_3075 (O_3075,N_46966,N_49700);
and UO_3076 (O_3076,N_41280,N_47553);
nand UO_3077 (O_3077,N_47488,N_44484);
or UO_3078 (O_3078,N_49030,N_42725);
and UO_3079 (O_3079,N_45077,N_40600);
nor UO_3080 (O_3080,N_40819,N_47721);
nand UO_3081 (O_3081,N_48215,N_42854);
nor UO_3082 (O_3082,N_49235,N_44414);
nand UO_3083 (O_3083,N_41870,N_46846);
nor UO_3084 (O_3084,N_48034,N_44630);
or UO_3085 (O_3085,N_47079,N_47472);
or UO_3086 (O_3086,N_47336,N_47126);
nor UO_3087 (O_3087,N_40442,N_49943);
and UO_3088 (O_3088,N_43429,N_40955);
or UO_3089 (O_3089,N_41814,N_49865);
nand UO_3090 (O_3090,N_40997,N_44889);
nand UO_3091 (O_3091,N_44599,N_46457);
xnor UO_3092 (O_3092,N_47572,N_45241);
or UO_3093 (O_3093,N_47841,N_41623);
nand UO_3094 (O_3094,N_49021,N_40005);
and UO_3095 (O_3095,N_44609,N_49512);
nor UO_3096 (O_3096,N_40030,N_46710);
and UO_3097 (O_3097,N_40744,N_43906);
nor UO_3098 (O_3098,N_41515,N_46280);
nor UO_3099 (O_3099,N_48327,N_47315);
and UO_3100 (O_3100,N_45247,N_44422);
nor UO_3101 (O_3101,N_40725,N_44499);
nor UO_3102 (O_3102,N_45923,N_40761);
nand UO_3103 (O_3103,N_47191,N_42621);
and UO_3104 (O_3104,N_46183,N_46250);
nand UO_3105 (O_3105,N_45365,N_49756);
or UO_3106 (O_3106,N_43948,N_44613);
nor UO_3107 (O_3107,N_44907,N_46232);
xnor UO_3108 (O_3108,N_47845,N_43417);
xor UO_3109 (O_3109,N_46654,N_41052);
nor UO_3110 (O_3110,N_47661,N_44017);
or UO_3111 (O_3111,N_45199,N_48861);
or UO_3112 (O_3112,N_45857,N_45533);
nand UO_3113 (O_3113,N_49677,N_41251);
nand UO_3114 (O_3114,N_48384,N_44485);
nand UO_3115 (O_3115,N_40223,N_49905);
and UO_3116 (O_3116,N_48310,N_45527);
and UO_3117 (O_3117,N_44399,N_44874);
and UO_3118 (O_3118,N_45629,N_46776);
nor UO_3119 (O_3119,N_44211,N_45485);
nor UO_3120 (O_3120,N_47835,N_45908);
or UO_3121 (O_3121,N_48710,N_41211);
nand UO_3122 (O_3122,N_45872,N_44584);
nand UO_3123 (O_3123,N_48017,N_46982);
and UO_3124 (O_3124,N_47827,N_43123);
nand UO_3125 (O_3125,N_43104,N_49299);
nand UO_3126 (O_3126,N_46717,N_49783);
or UO_3127 (O_3127,N_48899,N_46624);
and UO_3128 (O_3128,N_43179,N_49794);
nor UO_3129 (O_3129,N_43412,N_44126);
nor UO_3130 (O_3130,N_44955,N_42388);
or UO_3131 (O_3131,N_42125,N_42745);
nand UO_3132 (O_3132,N_46315,N_43491);
and UO_3133 (O_3133,N_48092,N_41836);
or UO_3134 (O_3134,N_43143,N_48397);
nand UO_3135 (O_3135,N_44626,N_49433);
or UO_3136 (O_3136,N_47337,N_48206);
nand UO_3137 (O_3137,N_40408,N_43161);
and UO_3138 (O_3138,N_40403,N_43100);
and UO_3139 (O_3139,N_48253,N_40664);
nand UO_3140 (O_3140,N_47196,N_43712);
or UO_3141 (O_3141,N_43770,N_43832);
and UO_3142 (O_3142,N_42067,N_40369);
nand UO_3143 (O_3143,N_44767,N_43975);
or UO_3144 (O_3144,N_40976,N_41998);
xnor UO_3145 (O_3145,N_48748,N_46818);
nand UO_3146 (O_3146,N_44801,N_41106);
xnor UO_3147 (O_3147,N_48458,N_46001);
or UO_3148 (O_3148,N_46206,N_49497);
nor UO_3149 (O_3149,N_43659,N_43598);
or UO_3150 (O_3150,N_48297,N_40287);
and UO_3151 (O_3151,N_41441,N_42874);
or UO_3152 (O_3152,N_40993,N_47796);
nand UO_3153 (O_3153,N_47948,N_42440);
and UO_3154 (O_3154,N_40377,N_45269);
and UO_3155 (O_3155,N_43817,N_46735);
nand UO_3156 (O_3156,N_42330,N_44730);
nor UO_3157 (O_3157,N_46984,N_44799);
or UO_3158 (O_3158,N_48716,N_44131);
and UO_3159 (O_3159,N_42251,N_49354);
nor UO_3160 (O_3160,N_47180,N_49148);
or UO_3161 (O_3161,N_42570,N_46467);
or UO_3162 (O_3162,N_49430,N_49593);
nor UO_3163 (O_3163,N_42075,N_49833);
xnor UO_3164 (O_3164,N_42494,N_42637);
or UO_3165 (O_3165,N_44735,N_48222);
nand UO_3166 (O_3166,N_44494,N_41869);
and UO_3167 (O_3167,N_41551,N_42991);
nand UO_3168 (O_3168,N_44994,N_44442);
and UO_3169 (O_3169,N_48749,N_48983);
or UO_3170 (O_3170,N_48732,N_47861);
or UO_3171 (O_3171,N_44124,N_43664);
and UO_3172 (O_3172,N_48391,N_41858);
nor UO_3173 (O_3173,N_47016,N_48889);
nor UO_3174 (O_3174,N_49032,N_45522);
nor UO_3175 (O_3175,N_44834,N_40665);
and UO_3176 (O_3176,N_43717,N_43967);
or UO_3177 (O_3177,N_45003,N_42311);
nand UO_3178 (O_3178,N_41458,N_43083);
nand UO_3179 (O_3179,N_44454,N_41030);
or UO_3180 (O_3180,N_41569,N_42047);
or UO_3181 (O_3181,N_49041,N_46088);
nor UO_3182 (O_3182,N_48032,N_48919);
xor UO_3183 (O_3183,N_42514,N_40194);
nor UO_3184 (O_3184,N_44878,N_48572);
nand UO_3185 (O_3185,N_42846,N_45668);
and UO_3186 (O_3186,N_45658,N_44145);
and UO_3187 (O_3187,N_41634,N_40232);
and UO_3188 (O_3188,N_47221,N_44379);
and UO_3189 (O_3189,N_40972,N_43545);
nor UO_3190 (O_3190,N_45271,N_48308);
and UO_3191 (O_3191,N_48903,N_41617);
and UO_3192 (O_3192,N_40082,N_49711);
nor UO_3193 (O_3193,N_46946,N_40926);
or UO_3194 (O_3194,N_48447,N_40672);
nand UO_3195 (O_3195,N_42181,N_49533);
nand UO_3196 (O_3196,N_43309,N_41091);
and UO_3197 (O_3197,N_40404,N_48734);
or UO_3198 (O_3198,N_49978,N_40669);
nor UO_3199 (O_3199,N_49829,N_47574);
and UO_3200 (O_3200,N_44805,N_47521);
xor UO_3201 (O_3201,N_49257,N_40491);
or UO_3202 (O_3202,N_42073,N_44831);
xor UO_3203 (O_3203,N_49368,N_45526);
and UO_3204 (O_3204,N_46563,N_40276);
and UO_3205 (O_3205,N_42025,N_45703);
and UO_3206 (O_3206,N_48119,N_45488);
nand UO_3207 (O_3207,N_49734,N_44249);
and UO_3208 (O_3208,N_49008,N_40483);
xnor UO_3209 (O_3209,N_42148,N_41829);
nor UO_3210 (O_3210,N_49611,N_46235);
and UO_3211 (O_3211,N_41549,N_49129);
nor UO_3212 (O_3212,N_49087,N_42501);
or UO_3213 (O_3213,N_48788,N_41884);
nor UO_3214 (O_3214,N_40942,N_46898);
xor UO_3215 (O_3215,N_45838,N_40482);
nand UO_3216 (O_3216,N_48517,N_43016);
nand UO_3217 (O_3217,N_40959,N_47223);
nand UO_3218 (O_3218,N_49929,N_44678);
and UO_3219 (O_3219,N_41841,N_47784);
nor UO_3220 (O_3220,N_48048,N_47621);
and UO_3221 (O_3221,N_49440,N_43722);
xnor UO_3222 (O_3222,N_47459,N_47391);
or UO_3223 (O_3223,N_44293,N_47662);
nor UO_3224 (O_3224,N_45615,N_42598);
or UO_3225 (O_3225,N_43215,N_44797);
and UO_3226 (O_3226,N_47279,N_44614);
xnor UO_3227 (O_3227,N_46022,N_43775);
nand UO_3228 (O_3228,N_45121,N_45200);
nor UO_3229 (O_3229,N_47106,N_44390);
nor UO_3230 (O_3230,N_48808,N_48947);
nand UO_3231 (O_3231,N_49079,N_43774);
xor UO_3232 (O_3232,N_46602,N_46456);
nor UO_3233 (O_3233,N_47182,N_47062);
or UO_3234 (O_3234,N_45423,N_45666);
nor UO_3235 (O_3235,N_47366,N_47242);
and UO_3236 (O_3236,N_40191,N_44042);
nor UO_3237 (O_3237,N_48411,N_43859);
nor UO_3238 (O_3238,N_48913,N_42312);
nor UO_3239 (O_3239,N_46046,N_49048);
nor UO_3240 (O_3240,N_45179,N_44990);
nand UO_3241 (O_3241,N_44065,N_42458);
and UO_3242 (O_3242,N_42746,N_48354);
and UO_3243 (O_3243,N_43798,N_41348);
nor UO_3244 (O_3244,N_43853,N_44360);
or UO_3245 (O_3245,N_47088,N_47048);
or UO_3246 (O_3246,N_43882,N_43599);
xnor UO_3247 (O_3247,N_45867,N_47470);
nand UO_3248 (O_3248,N_47740,N_46852);
nand UO_3249 (O_3249,N_45326,N_49938);
or UO_3250 (O_3250,N_41929,N_42605);
or UO_3251 (O_3251,N_42432,N_47229);
or UO_3252 (O_3252,N_47113,N_46296);
nand UO_3253 (O_3253,N_42742,N_47634);
nand UO_3254 (O_3254,N_45694,N_46550);
or UO_3255 (O_3255,N_48057,N_47750);
and UO_3256 (O_3256,N_41071,N_48158);
nor UO_3257 (O_3257,N_45738,N_46083);
nand UO_3258 (O_3258,N_41813,N_47490);
nand UO_3259 (O_3259,N_40888,N_49524);
and UO_3260 (O_3260,N_46479,N_43498);
and UO_3261 (O_3261,N_41560,N_43175);
xor UO_3262 (O_3262,N_40739,N_46635);
xor UO_3263 (O_3263,N_44288,N_45934);
nor UO_3264 (O_3264,N_48546,N_46513);
nand UO_3265 (O_3265,N_45915,N_43058);
or UO_3266 (O_3266,N_49675,N_42565);
and UO_3267 (O_3267,N_48110,N_45331);
or UO_3268 (O_3268,N_42131,N_43814);
nand UO_3269 (O_3269,N_41012,N_45861);
nand UO_3270 (O_3270,N_46616,N_48408);
and UO_3271 (O_3271,N_48987,N_48076);
or UO_3272 (O_3272,N_42363,N_47311);
or UO_3273 (O_3273,N_40500,N_44681);
nand UO_3274 (O_3274,N_40056,N_46798);
nand UO_3275 (O_3275,N_44802,N_45957);
nand UO_3276 (O_3276,N_40129,N_46073);
and UO_3277 (O_3277,N_43745,N_48083);
xor UO_3278 (O_3278,N_43938,N_40325);
nand UO_3279 (O_3279,N_42691,N_49876);
and UO_3280 (O_3280,N_49987,N_43044);
or UO_3281 (O_3281,N_48169,N_48638);
xnor UO_3282 (O_3282,N_40545,N_45366);
nand UO_3283 (O_3283,N_41793,N_48385);
nand UO_3284 (O_3284,N_47442,N_48769);
nand UO_3285 (O_3285,N_41663,N_46357);
or UO_3286 (O_3286,N_44412,N_41132);
or UO_3287 (O_3287,N_46638,N_44975);
or UO_3288 (O_3288,N_48621,N_45124);
nand UO_3289 (O_3289,N_44482,N_42255);
nand UO_3290 (O_3290,N_44384,N_49072);
nor UO_3291 (O_3291,N_45562,N_44952);
or UO_3292 (O_3292,N_49982,N_46248);
nand UO_3293 (O_3293,N_48030,N_46933);
nor UO_3294 (O_3294,N_42624,N_43167);
nor UO_3295 (O_3295,N_45952,N_49296);
nor UO_3296 (O_3296,N_49932,N_45832);
nand UO_3297 (O_3297,N_47918,N_49828);
nand UO_3298 (O_3298,N_44212,N_40760);
nand UO_3299 (O_3299,N_44385,N_49831);
nor UO_3300 (O_3300,N_44611,N_47267);
and UO_3301 (O_3301,N_45222,N_47549);
or UO_3302 (O_3302,N_47534,N_45525);
nand UO_3303 (O_3303,N_44366,N_40292);
and UO_3304 (O_3304,N_49893,N_46942);
nand UO_3305 (O_3305,N_46327,N_46186);
and UO_3306 (O_3306,N_45748,N_44774);
and UO_3307 (O_3307,N_40521,N_44713);
xnor UO_3308 (O_3308,N_40245,N_44180);
or UO_3309 (O_3309,N_42524,N_40536);
or UO_3310 (O_3310,N_46484,N_47111);
or UO_3311 (O_3311,N_40885,N_46489);
nand UO_3312 (O_3312,N_46129,N_45972);
and UO_3313 (O_3313,N_48977,N_46507);
nor UO_3314 (O_3314,N_43959,N_44864);
or UO_3315 (O_3315,N_40273,N_44335);
or UO_3316 (O_3316,N_44141,N_41366);
xnor UO_3317 (O_3317,N_43369,N_42603);
and UO_3318 (O_3318,N_40783,N_43109);
nand UO_3319 (O_3319,N_45712,N_41125);
or UO_3320 (O_3320,N_40290,N_40038);
or UO_3321 (O_3321,N_48219,N_42141);
nand UO_3322 (O_3322,N_41176,N_40898);
nor UO_3323 (O_3323,N_40293,N_43137);
and UO_3324 (O_3324,N_45860,N_43661);
or UO_3325 (O_3325,N_45053,N_40405);
nand UO_3326 (O_3326,N_49530,N_47053);
nand UO_3327 (O_3327,N_40824,N_47638);
or UO_3328 (O_3328,N_42946,N_47920);
nand UO_3329 (O_3329,N_49396,N_40682);
and UO_3330 (O_3330,N_48243,N_41619);
or UO_3331 (O_3331,N_45268,N_43812);
and UO_3332 (O_3332,N_49557,N_47027);
nor UO_3333 (O_3333,N_41819,N_49417);
nor UO_3334 (O_3334,N_40825,N_46707);
nor UO_3335 (O_3335,N_47489,N_48890);
or UO_3336 (O_3336,N_44883,N_44973);
xor UO_3337 (O_3337,N_46106,N_40204);
or UO_3338 (O_3338,N_45132,N_40333);
nand UO_3339 (O_3339,N_49639,N_43522);
or UO_3340 (O_3340,N_45401,N_41167);
xnor UO_3341 (O_3341,N_45216,N_40268);
nand UO_3342 (O_3342,N_43011,N_48273);
and UO_3343 (O_3343,N_44913,N_45429);
xor UO_3344 (O_3344,N_40516,N_47686);
nand UO_3345 (O_3345,N_48228,N_45650);
nor UO_3346 (O_3346,N_48342,N_46671);
nor UO_3347 (O_3347,N_42202,N_45516);
or UO_3348 (O_3348,N_43266,N_45518);
nand UO_3349 (O_3349,N_40746,N_46653);
and UO_3350 (O_3350,N_44074,N_48975);
xnor UO_3351 (O_3351,N_45618,N_42610);
nor UO_3352 (O_3352,N_44349,N_45885);
and UO_3353 (O_3353,N_48293,N_45037);
nor UO_3354 (O_3354,N_41647,N_46618);
and UO_3355 (O_3355,N_43631,N_40439);
or UO_3356 (O_3356,N_45167,N_45400);
nand UO_3357 (O_3357,N_40271,N_40910);
nor UO_3358 (O_3358,N_40828,N_41752);
nand UO_3359 (O_3359,N_41014,N_44643);
nor UO_3360 (O_3360,N_44157,N_45596);
nand UO_3361 (O_3361,N_45276,N_42016);
and UO_3362 (O_3362,N_49770,N_43186);
nand UO_3363 (O_3363,N_41005,N_44357);
and UO_3364 (O_3364,N_48500,N_46107);
nor UO_3365 (O_3365,N_48853,N_42037);
nor UO_3366 (O_3366,N_49624,N_43858);
nor UO_3367 (O_3367,N_43149,N_49039);
nor UO_3368 (O_3368,N_48828,N_46835);
nor UO_3369 (O_3369,N_42333,N_42748);
or UO_3370 (O_3370,N_49207,N_43029);
or UO_3371 (O_3371,N_46060,N_45935);
or UO_3372 (O_3372,N_45101,N_42540);
or UO_3373 (O_3373,N_44117,N_42066);
nor UO_3374 (O_3374,N_41268,N_48952);
or UO_3375 (O_3375,N_45492,N_43195);
or UO_3376 (O_3376,N_41574,N_42962);
or UO_3377 (O_3377,N_43077,N_49532);
or UO_3378 (O_3378,N_43203,N_48200);
or UO_3379 (O_3379,N_46868,N_43753);
nand UO_3380 (O_3380,N_40646,N_46875);
or UO_3381 (O_3381,N_40752,N_47135);
nor UO_3382 (O_3382,N_46167,N_46016);
xnor UO_3383 (O_3383,N_46453,N_42704);
or UO_3384 (O_3384,N_40963,N_46764);
nor UO_3385 (O_3385,N_44093,N_45223);
nand UO_3386 (O_3386,N_41310,N_44747);
nor UO_3387 (O_3387,N_49909,N_46607);
xnor UO_3388 (O_3388,N_40515,N_43987);
nand UO_3389 (O_3389,N_47026,N_45595);
or UO_3390 (O_3390,N_49024,N_43367);
nand UO_3391 (O_3391,N_42150,N_43466);
nor UO_3392 (O_3392,N_49123,N_48173);
or UO_3393 (O_3393,N_42483,N_46303);
nor UO_3394 (O_3394,N_47319,N_43981);
and UO_3395 (O_3395,N_40842,N_42967);
or UO_3396 (O_3396,N_47276,N_41643);
and UO_3397 (O_3397,N_45677,N_41410);
and UO_3398 (O_3398,N_45529,N_48662);
nor UO_3399 (O_3399,N_40329,N_45605);
nand UO_3400 (O_3400,N_48586,N_46829);
nor UO_3401 (O_3401,N_41103,N_46306);
or UO_3402 (O_3402,N_44076,N_40031);
and UO_3403 (O_3403,N_42798,N_40671);
nor UO_3404 (O_3404,N_47664,N_47655);
or UO_3405 (O_3405,N_41901,N_42853);
or UO_3406 (O_3406,N_49695,N_42126);
nand UO_3407 (O_3407,N_44041,N_45800);
xor UO_3408 (O_3408,N_46830,N_48757);
and UO_3409 (O_3409,N_42773,N_48094);
nand UO_3410 (O_3410,N_49256,N_45165);
nor UO_3411 (O_3411,N_46514,N_49269);
nor UO_3412 (O_3412,N_40656,N_47166);
xnor UO_3413 (O_3413,N_44324,N_40572);
and UO_3414 (O_3414,N_43969,N_41868);
nor UO_3415 (O_3415,N_48160,N_44337);
nand UO_3416 (O_3416,N_40709,N_46650);
or UO_3417 (O_3417,N_42373,N_45929);
nor UO_3418 (O_3418,N_46568,N_45576);
and UO_3419 (O_3419,N_45502,N_41407);
nand UO_3420 (O_3420,N_40361,N_49546);
or UO_3421 (O_3421,N_40507,N_46879);
or UO_3422 (O_3422,N_45343,N_45279);
or UO_3423 (O_3423,N_46736,N_44908);
nor UO_3424 (O_3424,N_44637,N_45417);
nor UO_3425 (O_3425,N_44552,N_45290);
or UO_3426 (O_3426,N_49033,N_43453);
or UO_3427 (O_3427,N_41114,N_48784);
and UO_3428 (O_3428,N_46837,N_49465);
nand UO_3429 (O_3429,N_40661,N_49660);
xor UO_3430 (O_3430,N_49790,N_46284);
or UO_3431 (O_3431,N_46890,N_46999);
and UO_3432 (O_3432,N_49236,N_42848);
nor UO_3433 (O_3433,N_48212,N_40588);
xor UO_3434 (O_3434,N_42827,N_47304);
nor UO_3435 (O_3435,N_46320,N_46522);
nor UO_3436 (O_3436,N_48062,N_43455);
nand UO_3437 (O_3437,N_42194,N_45831);
and UO_3438 (O_3438,N_43363,N_41696);
nor UO_3439 (O_3439,N_48277,N_46116);
nand UO_3440 (O_3440,N_42291,N_49243);
and UO_3441 (O_3441,N_44347,N_47859);
or UO_3442 (O_3442,N_44925,N_49651);
nand UO_3443 (O_3443,N_48640,N_45598);
and UO_3444 (O_3444,N_43508,N_46703);
or UO_3445 (O_3445,N_43940,N_47892);
and UO_3446 (O_3446,N_49163,N_43456);
and UO_3447 (O_3447,N_49098,N_44447);
nand UO_3448 (O_3448,N_45454,N_40418);
or UO_3449 (O_3449,N_49506,N_48114);
and UO_3450 (O_3450,N_43237,N_47749);
and UO_3451 (O_3451,N_40171,N_45284);
or UO_3452 (O_3452,N_46052,N_46611);
and UO_3453 (O_3453,N_40979,N_44617);
nor UO_3454 (O_3454,N_41578,N_48653);
and UO_3455 (O_3455,N_40100,N_47837);
and UO_3456 (O_3456,N_41019,N_43249);
or UO_3457 (O_3457,N_41344,N_45660);
nor UO_3458 (O_3458,N_48280,N_47769);
or UO_3459 (O_3459,N_42318,N_42548);
nand UO_3460 (O_3460,N_42498,N_40820);
xnor UO_3461 (O_3461,N_47797,N_40645);
or UO_3462 (O_3462,N_46398,N_49581);
nand UO_3463 (O_3463,N_40757,N_43777);
nand UO_3464 (O_3464,N_49616,N_49234);
or UO_3465 (O_3465,N_48358,N_46679);
or UO_3466 (O_3466,N_43989,N_48712);
or UO_3467 (O_3467,N_45054,N_42497);
nor UO_3468 (O_3468,N_41831,N_40817);
nand UO_3469 (O_3469,N_41889,N_41284);
or UO_3470 (O_3470,N_43993,N_45018);
xnor UO_3471 (O_3471,N_40186,N_44823);
nor UO_3472 (O_3472,N_47622,N_49871);
nand UO_3473 (O_3473,N_48492,N_42664);
or UO_3474 (O_3474,N_42646,N_48268);
or UO_3475 (O_3475,N_44814,N_40079);
and UO_3476 (O_3476,N_42298,N_47506);
nand UO_3477 (O_3477,N_48043,N_47255);
nand UO_3478 (O_3478,N_41484,N_48990);
or UO_3479 (O_3479,N_46422,N_46899);
nor UO_3480 (O_3480,N_45883,N_49983);
nand UO_3481 (O_3481,N_46213,N_41612);
or UO_3482 (O_3482,N_44531,N_40717);
nor UO_3483 (O_3483,N_42711,N_46348);
nand UO_3484 (O_3484,N_44051,N_45318);
nand UO_3485 (O_3485,N_40340,N_47937);
nand UO_3486 (O_3486,N_45477,N_48260);
nor UO_3487 (O_3487,N_47081,N_42585);
xnor UO_3488 (O_3488,N_40814,N_45790);
xnor UO_3489 (O_3489,N_48108,N_46401);
or UO_3490 (O_3490,N_43166,N_47138);
nand UO_3491 (O_3491,N_41883,N_49114);
nor UO_3492 (O_3492,N_45395,N_45445);
nand UO_3493 (O_3493,N_42415,N_41636);
and UO_3494 (O_3494,N_45704,N_43961);
nor UO_3495 (O_3495,N_42120,N_48702);
nand UO_3496 (O_3496,N_42115,N_41881);
nand UO_3497 (O_3497,N_46249,N_45641);
nand UO_3498 (O_3498,N_47484,N_43890);
or UO_3499 (O_3499,N_45481,N_41283);
and UO_3500 (O_3500,N_49666,N_49959);
nor UO_3501 (O_3501,N_47217,N_49779);
nand UO_3502 (O_3502,N_46100,N_45889);
and UO_3503 (O_3503,N_45750,N_47383);
or UO_3504 (O_3504,N_49142,N_49083);
nor UO_3505 (O_3505,N_41004,N_48670);
or UO_3506 (O_3506,N_40550,N_46814);
nand UO_3507 (O_3507,N_43151,N_40224);
xor UO_3508 (O_3508,N_47355,N_49294);
nand UO_3509 (O_3509,N_43539,N_41992);
nand UO_3510 (O_3510,N_48442,N_43530);
xnor UO_3511 (O_3511,N_41891,N_41224);
nand UO_3512 (O_3512,N_46369,N_41057);
or UO_3513 (O_3513,N_49054,N_40478);
nand UO_3514 (O_3514,N_48059,N_40485);
or UO_3515 (O_3515,N_49542,N_49738);
xnor UO_3516 (O_3516,N_46365,N_48944);
or UO_3517 (O_3517,N_43526,N_42190);
or UO_3518 (O_3518,N_48003,N_47597);
nor UO_3519 (O_3519,N_46977,N_42499);
nor UO_3520 (O_3520,N_45622,N_40022);
nand UO_3521 (O_3521,N_44706,N_47474);
xnor UO_3522 (O_3522,N_46414,N_40200);
nor UO_3523 (O_3523,N_44922,N_46797);
and UO_3524 (O_3524,N_42428,N_44416);
and UO_3525 (O_3525,N_41718,N_49274);
and UO_3526 (O_3526,N_40782,N_47665);
and UO_3527 (O_3527,N_44661,N_48841);
or UO_3528 (O_3528,N_41257,N_41716);
nand UO_3529 (O_3529,N_47807,N_46286);
or UO_3530 (O_3530,N_43351,N_44533);
nand UO_3531 (O_3531,N_48893,N_41618);
xnor UO_3532 (O_3532,N_42786,N_40660);
xnor UO_3533 (O_3533,N_43874,N_40025);
nand UO_3534 (O_3534,N_49393,N_40636);
nor UO_3535 (O_3535,N_43810,N_41026);
or UO_3536 (O_3536,N_48907,N_43193);
and UO_3537 (O_3537,N_44548,N_41022);
or UO_3538 (O_3538,N_43075,N_49334);
nand UO_3539 (O_3539,N_40037,N_47413);
nand UO_3540 (O_3540,N_42708,N_45802);
nand UO_3541 (O_3541,N_42625,N_48619);
nor UO_3542 (O_3542,N_46162,N_45219);
nand UO_3543 (O_3543,N_47954,N_45203);
nor UO_3544 (O_3544,N_43295,N_45651);
nor UO_3545 (O_3545,N_47675,N_42753);
nor UO_3546 (O_3546,N_44333,N_46913);
nand UO_3547 (O_3547,N_49121,N_40331);
nor UO_3548 (O_3548,N_45230,N_43440);
nor UO_3549 (O_3549,N_41264,N_49551);
or UO_3550 (O_3550,N_46658,N_49223);
nor UO_3551 (O_3551,N_44259,N_41498);
and UO_3552 (O_3552,N_45135,N_49290);
nand UO_3553 (O_3553,N_48877,N_41307);
nand UO_3554 (O_3554,N_47599,N_45342);
or UO_3555 (O_3555,N_43036,N_42995);
nor UO_3556 (O_3556,N_48463,N_43174);
or UO_3557 (O_3557,N_45320,N_44116);
and UO_3558 (O_3558,N_44627,N_40049);
nand UO_3559 (O_3559,N_42209,N_45584);
nor UO_3560 (O_3560,N_49720,N_41790);
and UO_3561 (O_3561,N_43665,N_47423);
or UO_3562 (O_3562,N_41751,N_41404);
nor UO_3563 (O_3563,N_44356,N_47698);
xor UO_3564 (O_3564,N_46026,N_46040);
or UO_3565 (O_3565,N_45967,N_49439);
nand UO_3566 (O_3566,N_41397,N_45440);
and UO_3567 (O_3567,N_44338,N_47612);
or UO_3568 (O_3568,N_43102,N_49716);
nor UO_3569 (O_3569,N_43515,N_48421);
nor UO_3570 (O_3570,N_41885,N_45317);
or UO_3571 (O_3571,N_47492,N_48307);
or UO_3572 (O_3572,N_47376,N_47061);
nand UO_3573 (O_3573,N_47566,N_48423);
and UO_3574 (O_3574,N_40781,N_49245);
and UO_3575 (O_3575,N_46151,N_41791);
nand UO_3576 (O_3576,N_49131,N_43122);
nand UO_3577 (O_3577,N_45056,N_42784);
and UO_3578 (O_3578,N_41299,N_48367);
nand UO_3579 (O_3579,N_49587,N_46399);
nand UO_3580 (O_3580,N_43922,N_42396);
or UO_3581 (O_3581,N_45891,N_43970);
nand UO_3582 (O_3582,N_41324,N_48627);
or UO_3583 (O_3583,N_40148,N_49351);
or UO_3584 (O_3584,N_41432,N_40310);
nand UO_3585 (O_3585,N_44884,N_40118);
xor UO_3586 (O_3586,N_44072,N_46788);
and UO_3587 (O_3587,N_46960,N_44125);
or UO_3588 (O_3588,N_45818,N_44873);
and UO_3589 (O_3589,N_48295,N_46673);
nor UO_3590 (O_3590,N_45642,N_45185);
nand UO_3591 (O_3591,N_47872,N_48882);
or UO_3592 (O_3592,N_47368,N_47568);
or UO_3593 (O_3593,N_47064,N_41007);
and UO_3594 (O_3594,N_44505,N_40366);
and UO_3595 (O_3595,N_45821,N_41236);
or UO_3596 (O_3596,N_47359,N_46543);
and UO_3597 (O_3597,N_40141,N_44296);
nand UO_3598 (O_3598,N_48229,N_42238);
nand UO_3599 (O_3599,N_42224,N_44663);
nand UO_3600 (O_3600,N_44982,N_46822);
nand UO_3601 (O_3601,N_45648,N_40532);
and UO_3602 (O_3602,N_46524,N_43045);
nand UO_3603 (O_3603,N_48419,N_47290);
or UO_3604 (O_3604,N_49529,N_49146);
or UO_3605 (O_3605,N_43263,N_40953);
or UO_3606 (O_3606,N_46476,N_47687);
or UO_3607 (O_3607,N_43478,N_44283);
nand UO_3608 (O_3608,N_47935,N_44571);
nand UO_3609 (O_3609,N_44139,N_46811);
nor UO_3610 (O_3610,N_42264,N_41471);
nand UO_3611 (O_3611,N_42619,N_42468);
nor UO_3612 (O_3612,N_42023,N_49513);
or UO_3613 (O_3613,N_42180,N_46098);
nand UO_3614 (O_3614,N_43736,N_41293);
nor UO_3615 (O_3615,N_42322,N_42652);
xor UO_3616 (O_3616,N_44147,N_41824);
and UO_3617 (O_3617,N_47780,N_49582);
or UO_3618 (O_3618,N_42907,N_46675);
xnor UO_3619 (O_3619,N_41036,N_40903);
and UO_3620 (O_3620,N_47264,N_49301);
and UO_3621 (O_3621,N_44818,N_40802);
and UO_3622 (O_3622,N_43383,N_41916);
and UO_3623 (O_3623,N_48381,N_45603);
nand UO_3624 (O_3624,N_46393,N_44239);
xor UO_3625 (O_3625,N_44101,N_43503);
nor UO_3626 (O_3626,N_48914,N_41686);
xnor UO_3627 (O_3627,N_49527,N_49253);
nand UO_3628 (O_3628,N_42050,N_45767);
and UO_3629 (O_3629,N_41430,N_40167);
nor UO_3630 (O_3630,N_41329,N_42100);
or UO_3631 (O_3631,N_42442,N_49482);
nand UO_3632 (O_3632,N_44857,N_45382);
nor UO_3633 (O_3633,N_40006,N_46769);
or UO_3634 (O_3634,N_44798,N_44672);
and UO_3635 (O_3635,N_43028,N_47248);
nand UO_3636 (O_3636,N_47252,N_46407);
nor UO_3637 (O_3637,N_43724,N_40054);
xor UO_3638 (O_3638,N_40421,N_47372);
and UO_3639 (O_3639,N_46152,N_48282);
and UO_3640 (O_3640,N_43542,N_46787);
and UO_3641 (O_3641,N_46121,N_43534);
and UO_3642 (O_3642,N_46460,N_42080);
and UO_3643 (O_3643,N_43911,N_41789);
or UO_3644 (O_3644,N_45322,N_47331);
or UO_3645 (O_3645,N_47536,N_43451);
and UO_3646 (O_3646,N_42196,N_41265);
and UO_3647 (O_3647,N_42082,N_41467);
nand UO_3648 (O_3648,N_45015,N_49314);
nor UO_3649 (O_3649,N_49793,N_44026);
nor UO_3650 (O_3650,N_41567,N_42041);
and UO_3651 (O_3651,N_43549,N_43739);
nor UO_3652 (O_3652,N_43869,N_41164);
xor UO_3653 (O_3653,N_44274,N_48066);
nand UO_3654 (O_3654,N_40423,N_46187);
nor UO_3655 (O_3655,N_46178,N_43228);
nor UO_3656 (O_3656,N_47636,N_46408);
nand UO_3657 (O_3657,N_43252,N_49406);
and UO_3658 (O_3658,N_46087,N_48819);
or UO_3659 (O_3659,N_42957,N_41286);
nand UO_3660 (O_3660,N_44700,N_41507);
nand UO_3661 (O_3661,N_46185,N_49578);
nand UO_3662 (O_3662,N_49588,N_46613);
and UO_3663 (O_3663,N_41960,N_40659);
nand UO_3664 (O_3664,N_48251,N_42491);
nor UO_3665 (O_3665,N_46598,N_47603);
and UO_3666 (O_3666,N_46082,N_48620);
nor UO_3667 (O_3667,N_48955,N_42055);
nor UO_3668 (O_3668,N_44851,N_45785);
nand UO_3669 (O_3669,N_48960,N_46002);
or UO_3670 (O_3670,N_46184,N_47931);
xor UO_3671 (O_3671,N_44298,N_45328);
or UO_3672 (O_3672,N_44899,N_42213);
nand UO_3673 (O_3673,N_40932,N_40134);
or UO_3674 (O_3674,N_49980,N_42930);
and UO_3675 (O_3675,N_40956,N_47902);
nand UO_3676 (O_3676,N_47167,N_46768);
nor UO_3677 (O_3677,N_47418,N_42914);
nor UO_3678 (O_3678,N_41439,N_46869);
nor UO_3679 (O_3679,N_45009,N_49919);
or UO_3680 (O_3680,N_47250,N_46801);
and UO_3681 (O_3681,N_46831,N_41972);
nand UO_3682 (O_3682,N_45823,N_45925);
xor UO_3683 (O_3683,N_44877,N_40083);
nor UO_3684 (O_3684,N_40859,N_43728);
or UO_3685 (O_3685,N_47882,N_49944);
or UO_3686 (O_3686,N_42792,N_42437);
or UO_3687 (O_3687,N_45478,N_40322);
xor UO_3688 (O_3688,N_41803,N_40456);
and UO_3689 (O_3689,N_49920,N_48042);
nor UO_3690 (O_3690,N_42462,N_46159);
and UO_3691 (O_3691,N_44848,N_44731);
nor UO_3692 (O_3692,N_41109,N_49838);
or UO_3693 (O_3693,N_44777,N_47277);
or UO_3694 (O_3694,N_40211,N_42594);
and UO_3695 (O_3695,N_47109,N_43697);
or UO_3696 (O_3696,N_47818,N_47867);
and UO_3697 (O_3697,N_43189,N_42993);
and UO_3698 (O_3698,N_40313,N_46588);
and UO_3699 (O_3699,N_42061,N_43372);
nand UO_3700 (O_3700,N_48569,N_45233);
nor UO_3701 (O_3701,N_46062,N_41185);
or UO_3702 (O_3702,N_44208,N_46472);
or UO_3703 (O_3703,N_43839,N_46324);
xnor UO_3704 (O_3704,N_45408,N_46529);
nand UO_3705 (O_3705,N_40382,N_48377);
or UO_3706 (O_3706,N_48506,N_49850);
or UO_3707 (O_3707,N_49100,N_49789);
xnor UO_3708 (O_3708,N_42172,N_44561);
and UO_3709 (O_3709,N_45338,N_49500);
nand UO_3710 (O_3710,N_46683,N_48079);
nand UO_3711 (O_3711,N_48010,N_41006);
and UO_3712 (O_3712,N_40815,N_48603);
or UO_3713 (O_3713,N_42431,N_49672);
or UO_3714 (O_3714,N_40447,N_42074);
or UO_3715 (O_3715,N_47908,N_40263);
nand UO_3716 (O_3716,N_42830,N_49489);
or UO_3717 (O_3717,N_49367,N_46985);
and UO_3718 (O_3718,N_42467,N_48637);
xnor UO_3719 (O_3719,N_42974,N_43165);
nand UO_3720 (O_3720,N_48659,N_47055);
or UO_3721 (O_3721,N_42005,N_47386);
nand UO_3722 (O_3722,N_44015,N_49395);
nor UO_3723 (O_3723,N_49933,N_44103);
nand UO_3724 (O_3724,N_43499,N_47539);
and UO_3725 (O_3725,N_44600,N_43868);
nand UO_3726 (O_3726,N_43852,N_42387);
nor UO_3727 (O_3727,N_46860,N_48469);
and UO_3728 (O_3728,N_48625,N_45940);
or UO_3729 (O_3729,N_42674,N_45255);
nor UO_3730 (O_3730,N_45335,N_47310);
nor UO_3731 (O_3731,N_41923,N_43335);
nor UO_3732 (O_3732,N_48922,N_40538);
xor UO_3733 (O_3733,N_42188,N_49369);
nand UO_3734 (O_3734,N_49113,N_48731);
and UO_3735 (O_3735,N_46384,N_48651);
or UO_3736 (O_3736,N_47912,N_49628);
nand UO_3737 (O_3737,N_46090,N_48335);
nor UO_3738 (O_3738,N_47468,N_41805);
or UO_3739 (O_3739,N_49963,N_40644);
or UO_3740 (O_3740,N_40770,N_44724);
nand UO_3741 (O_3741,N_45393,N_44310);
nor UO_3742 (O_3742,N_45920,N_45224);
or UO_3743 (O_3743,N_40360,N_40511);
or UO_3744 (O_3744,N_48294,N_41409);
and UO_3745 (O_3745,N_47616,N_44311);
or UO_3746 (O_3746,N_42644,N_42770);
nor UO_3747 (O_3747,N_40807,N_46347);
nand UO_3748 (O_3748,N_40998,N_48703);
nand UO_3749 (O_3749,N_48407,N_41961);
and UO_3750 (O_3750,N_42130,N_40981);
nor UO_3751 (O_3751,N_48697,N_45297);
nor UO_3752 (O_3752,N_43988,N_41332);
and UO_3753 (O_3753,N_46606,N_42989);
nand UO_3754 (O_3754,N_48387,N_42233);
or UO_3755 (O_3755,N_42672,N_45914);
nor UO_3756 (O_3756,N_46701,N_44508);
nand UO_3757 (O_3757,N_47326,N_47917);
nor UO_3758 (O_3758,N_44750,N_48479);
nand UO_3759 (O_3759,N_40595,N_43808);
or UO_3760 (O_3760,N_42972,N_47093);
nand UO_3761 (O_3761,N_44514,N_48614);
and UO_3762 (O_3762,N_45859,N_48636);
or UO_3763 (O_3763,N_45065,N_41320);
and UO_3764 (O_3764,N_49543,N_46741);
nand UO_3765 (O_3765,N_42968,N_49816);
or UO_3766 (O_3766,N_43709,N_42757);
nand UO_3767 (O_3767,N_44612,N_44770);
nor UO_3768 (O_3768,N_43438,N_47762);
nor UO_3769 (O_3769,N_47156,N_44159);
and UO_3770 (O_3770,N_47329,N_47004);
nor UO_3771 (O_3771,N_46045,N_41772);
xnor UO_3772 (O_3772,N_40213,N_47733);
nor UO_3773 (O_3773,N_44944,N_44331);
nand UO_3774 (O_3774,N_41914,N_49928);
nor UO_3775 (O_3775,N_43033,N_48085);
nor UO_3776 (O_3776,N_48186,N_48744);
nor UO_3777 (O_3777,N_49860,N_46504);
and UO_3778 (O_3778,N_40653,N_49697);
nor UO_3779 (O_3779,N_40916,N_49678);
and UO_3780 (O_3780,N_40088,N_42176);
and UO_3781 (O_3781,N_49003,N_43679);
nand UO_3782 (O_3782,N_47605,N_45829);
nand UO_3783 (O_3783,N_41435,N_45612);
and UO_3784 (O_3784,N_43555,N_49091);
nand UO_3785 (O_3785,N_46866,N_43414);
nand UO_3786 (O_3786,N_44094,N_41325);
and UO_3787 (O_3787,N_48523,N_41326);
or UO_3788 (O_3788,N_46309,N_49108);
nand UO_3789 (O_3789,N_44729,N_40306);
and UO_3790 (O_3790,N_47206,N_44651);
and UO_3791 (O_3791,N_41201,N_46686);
nand UO_3792 (O_3792,N_42173,N_42053);
nor UO_3793 (O_3793,N_45141,N_43750);
xnor UO_3794 (O_3794,N_45022,N_48449);
xnor UO_3795 (O_3795,N_44463,N_46621);
and UO_3796 (O_3796,N_43296,N_44201);
nand UO_3797 (O_3797,N_46533,N_49591);
and UO_3798 (O_3798,N_42411,N_46528);
nand UO_3799 (O_3799,N_47679,N_49329);
or UO_3800 (O_3800,N_49431,N_41804);
and UO_3801 (O_3801,N_48369,N_40400);
nand UO_3802 (O_3802,N_42859,N_46660);
nor UO_3803 (O_3803,N_40363,N_48593);
nand UO_3804 (O_3804,N_44455,N_41712);
nand UO_3805 (O_3805,N_47586,N_49007);
and UO_3806 (O_3806,N_45528,N_45161);
or UO_3807 (O_3807,N_43348,N_45965);
or UO_3808 (O_3808,N_45563,N_47097);
nand UO_3809 (O_3809,N_44701,N_47316);
and UO_3810 (O_3810,N_47201,N_45016);
nor UO_3811 (O_3811,N_48858,N_45182);
or UO_3812 (O_3812,N_43482,N_46536);
and UO_3813 (O_3813,N_46729,N_43475);
nand UO_3814 (O_3814,N_43304,N_45060);
nand UO_3815 (O_3815,N_48304,N_43172);
nand UO_3816 (O_3816,N_49891,N_42806);
nor UO_3817 (O_3817,N_40886,N_40704);
and UO_3818 (O_3818,N_41667,N_44771);
nand UO_3819 (O_3819,N_40578,N_42697);
nor UO_3820 (O_3820,N_49951,N_41240);
and UO_3821 (O_3821,N_47169,N_43523);
or UO_3822 (O_3822,N_40150,N_48803);
xnor UO_3823 (O_3823,N_42249,N_42225);
xnor UO_3824 (O_3824,N_49656,N_41982);
nor UO_3825 (O_3825,N_40765,N_46077);
xor UO_3826 (O_3826,N_48690,N_43807);
nor UO_3827 (O_3827,N_46905,N_46510);
nor UO_3828 (O_3828,N_42857,N_41413);
or UO_3829 (O_3829,N_42516,N_43467);
or UO_3830 (O_3830,N_46990,N_40927);
or UO_3831 (O_3831,N_46780,N_45986);
xnor UO_3832 (O_3832,N_45350,N_44766);
nand UO_3833 (O_3833,N_46649,N_47724);
or UO_3834 (O_3834,N_49034,N_41076);
xnor UO_3835 (O_3835,N_44501,N_41194);
and UO_3836 (O_3836,N_46880,N_40015);
or UO_3837 (O_3837,N_44287,N_49447);
and UO_3838 (O_3838,N_46637,N_45017);
nor UO_3839 (O_3839,N_45590,N_41556);
and UO_3840 (O_3840,N_42802,N_49038);
nor UO_3841 (O_3841,N_43080,N_40706);
and UO_3842 (O_3842,N_45012,N_47322);
and UO_3843 (O_3843,N_41162,N_40662);
xnor UO_3844 (O_3844,N_43621,N_46626);
nand UO_3845 (O_3845,N_40092,N_40969);
nor UO_3846 (O_3846,N_43843,N_49327);
and UO_3847 (O_3847,N_45532,N_48436);
nor UO_3848 (O_3848,N_42713,N_42839);
nand UO_3849 (O_3849,N_48106,N_47301);
or UO_3850 (O_3850,N_49286,N_49824);
or UO_3851 (O_3851,N_44785,N_40584);
nand UO_3852 (O_3852,N_49967,N_43447);
and UO_3853 (O_3853,N_45487,N_47421);
or UO_3854 (O_3854,N_41689,N_40201);
xnor UO_3855 (O_3855,N_44853,N_46486);
and UO_3856 (O_3856,N_43936,N_41113);
nand UO_3857 (O_3857,N_41786,N_42302);
or UO_3858 (O_3858,N_44057,N_42077);
nor UO_3859 (O_3859,N_47249,N_47299);
nor UO_3860 (O_3860,N_41544,N_43261);
or UO_3861 (O_3861,N_45759,N_47228);
or UO_3862 (O_3862,N_48037,N_45011);
nand UO_3863 (O_3863,N_40971,N_49180);
nand UO_3864 (O_3864,N_41682,N_46372);
and UO_3865 (O_3865,N_40562,N_48509);
or UO_3866 (O_3866,N_44545,N_40902);
nor UO_3867 (O_3867,N_42843,N_47060);
or UO_3868 (O_3868,N_43624,N_47529);
and UO_3869 (O_3869,N_49868,N_46143);
and UO_3870 (O_3870,N_47500,N_43579);
and UO_3871 (O_3871,N_48167,N_44254);
xnor UO_3872 (O_3872,N_48331,N_40330);
nor UO_3873 (O_3873,N_46466,N_47803);
xnor UO_3874 (O_3874,N_45218,N_46364);
nand UO_3875 (O_3875,N_43169,N_44709);
or UO_3876 (O_3876,N_41737,N_40346);
nor UO_3877 (O_3877,N_44060,N_44565);
nand UO_3878 (O_3878,N_40463,N_43623);
nand UO_3879 (O_3879,N_41321,N_41339);
nand UO_3880 (O_3880,N_45842,N_41584);
and UO_3881 (O_3881,N_45811,N_40640);
nand UO_3882 (O_3882,N_41529,N_47899);
nor UO_3883 (O_3883,N_45486,N_40388);
or UO_3884 (O_3884,N_45031,N_40316);
nor UO_3885 (O_3885,N_40236,N_43734);
nand UO_3886 (O_3886,N_43425,N_49194);
and UO_3887 (O_3887,N_45625,N_41375);
nand UO_3888 (O_3888,N_45456,N_43147);
nor UO_3889 (O_3889,N_49545,N_47766);
nand UO_3890 (O_3890,N_43636,N_44345);
nor UO_3891 (O_3891,N_48112,N_45086);
nand UO_3892 (O_3892,N_47035,N_43984);
nand UO_3893 (O_3893,N_47526,N_43443);
nand UO_3894 (O_3894,N_45729,N_42721);
nor UO_3895 (O_3895,N_48740,N_44707);
or UO_3896 (O_3896,N_48118,N_47637);
or UO_3897 (O_3897,N_41725,N_45709);
or UO_3898 (O_3898,N_49855,N_42511);
nand UO_3899 (O_3899,N_49385,N_46873);
and UO_3900 (O_3900,N_42915,N_46441);
and UO_3901 (O_3901,N_40586,N_42768);
nand UO_3902 (O_3902,N_49424,N_48539);
nor UO_3903 (O_3903,N_45696,N_46521);
or UO_3904 (O_3904,N_49260,N_42551);
nand UO_3905 (O_3905,N_49096,N_49968);
nor UO_3906 (O_3906,N_41371,N_44470);
nand UO_3907 (O_3907,N_40140,N_43064);
nand UO_3908 (O_3908,N_40358,N_48865);
xnor UO_3909 (O_3909,N_49183,N_46542);
nand UO_3910 (O_3910,N_47259,N_48137);
nor UO_3911 (O_3911,N_42201,N_47737);
nand UO_3912 (O_3912,N_46751,N_41949);
or UO_3913 (O_3913,N_40543,N_47354);
xnor UO_3914 (O_3914,N_40986,N_48434);
nor UO_3915 (O_3915,N_42724,N_47723);
and UO_3916 (O_3916,N_43319,N_40517);
and UO_3917 (O_3917,N_45515,N_46490);
nand UO_3918 (O_3918,N_48490,N_47403);
nor UO_3919 (O_3919,N_42008,N_46727);
nand UO_3920 (O_3920,N_49017,N_45519);
nor UO_3921 (O_3921,N_46379,N_49064);
nor UO_3922 (O_3922,N_46331,N_46520);
and UO_3923 (O_3923,N_43592,N_48238);
or UO_3924 (O_3924,N_44368,N_42513);
and UO_3925 (O_3925,N_41372,N_47747);
and UO_3926 (O_3926,N_43667,N_41832);
or UO_3927 (O_3927,N_49764,N_42098);
or UO_3928 (O_3928,N_43752,N_40041);
nor UO_3929 (O_3929,N_40009,N_47589);
or UO_3930 (O_3930,N_40711,N_48202);
and UO_3931 (O_3931,N_40113,N_44892);
nor UO_3932 (O_3932,N_49044,N_43945);
or UO_3933 (O_3933,N_49213,N_45736);
nor UO_3934 (O_3934,N_44019,N_47265);
nand UO_3935 (O_3935,N_44267,N_47171);
nand UO_3936 (O_3936,N_41281,N_43310);
or UO_3937 (O_3937,N_44002,N_42299);
nor UO_3938 (O_3938,N_44244,N_43037);
nor UO_3939 (O_3939,N_43564,N_45275);
or UO_3940 (O_3940,N_47471,N_48972);
or UO_3941 (O_3941,N_42841,N_48427);
or UO_3942 (O_3942,N_48475,N_45592);
nand UO_3943 (O_3943,N_45138,N_46773);
nand UO_3944 (O_3944,N_49681,N_45985);
nand UO_3945 (O_3945,N_46078,N_44137);
nor UO_3946 (O_3946,N_48279,N_40599);
or UO_3947 (O_3947,N_44339,N_42156);
and UO_3948 (O_3948,N_44317,N_45157);
nor UO_3949 (O_3949,N_45745,N_42526);
or UO_3950 (O_3950,N_48548,N_46740);
nand UO_3951 (O_3951,N_42434,N_49888);
nor UO_3952 (O_3952,N_46266,N_45493);
and UO_3953 (O_3953,N_43400,N_44893);
nor UO_3954 (O_3954,N_44388,N_46932);
and UO_3955 (O_3955,N_43486,N_49473);
nand UO_3956 (O_3956,N_42438,N_46962);
nand UO_3957 (O_3957,N_44022,N_48465);
and UO_3958 (O_3958,N_44270,N_46806);
nand UO_3959 (O_3959,N_47270,N_40183);
nand UO_3960 (O_3960,N_48568,N_42521);
or UO_3961 (O_3961,N_41955,N_46979);
nand UO_3962 (O_3962,N_42591,N_42192);
nor UO_3963 (O_3963,N_46381,N_45898);
xnor UO_3964 (O_3964,N_43671,N_42205);
nand UO_3965 (O_3965,N_44429,N_43477);
or UO_3966 (O_3966,N_43607,N_40683);
nand UO_3967 (O_3967,N_41750,N_48634);
nand UO_3968 (O_3968,N_41154,N_44906);
xnor UO_3969 (O_3969,N_40492,N_40838);
nor UO_3970 (O_3970,N_47087,N_47020);
nand UO_3971 (O_3971,N_44369,N_43674);
xnor UO_3972 (O_3972,N_48350,N_48715);
or UO_3973 (O_3973,N_42104,N_43606);
and UO_3974 (O_3974,N_40078,N_47346);
nand UO_3975 (O_3975,N_47779,N_45682);
or UO_3976 (O_3976,N_49242,N_44957);
or UO_3977 (O_3977,N_44090,N_49729);
nand UO_3978 (O_3978,N_49157,N_45470);
and UO_3979 (O_3979,N_44168,N_41341);
and UO_3980 (O_3980,N_47808,N_42040);
and UO_3981 (O_3981,N_40747,N_47015);
nor UO_3982 (O_3982,N_41438,N_46325);
and UO_3983 (O_3983,N_41237,N_41287);
and UO_3984 (O_3984,N_45971,N_49308);
or UO_3985 (O_3985,N_43328,N_42477);
or UO_3986 (O_3986,N_40862,N_48236);
nand UO_3987 (O_3987,N_42684,N_48120);
nand UO_3988 (O_3988,N_41493,N_49563);
or UO_3989 (O_3989,N_46136,N_40831);
nor UO_3990 (O_3990,N_41876,N_43188);
and UO_3991 (O_3991,N_48607,N_47977);
or UO_3992 (O_3992,N_41583,N_42320);
nand UO_3993 (O_3993,N_47251,N_49193);
and UO_3994 (O_3994,N_43704,N_47047);
or UO_3995 (O_3995,N_40858,N_44037);
nand UO_3996 (O_3996,N_48468,N_43354);
nand UO_3997 (O_3997,N_45856,N_45560);
and UO_3998 (O_3998,N_45099,N_42808);
nand UO_3999 (O_3999,N_42217,N_44506);
and UO_4000 (O_4000,N_42726,N_41096);
or UO_4001 (O_4001,N_40740,N_41434);
nor UO_4002 (O_4002,N_45032,N_41907);
nand UO_4003 (O_4003,N_44521,N_48867);
and UO_4004 (O_4004,N_40892,N_49730);
nor UO_4005 (O_4005,N_41993,N_41206);
and UO_4006 (O_4006,N_48375,N_48747);
nand UO_4007 (O_4007,N_45421,N_45337);
and UO_4008 (O_4008,N_45460,N_43844);
nand UO_4009 (O_4009,N_48400,N_42762);
or UO_4010 (O_4010,N_45888,N_46525);
and UO_4011 (O_4011,N_47233,N_47748);
or UO_4012 (O_4012,N_47787,N_43127);
nor UO_4013 (O_4013,N_41472,N_43738);
or UO_4014 (O_4014,N_48646,N_44056);
nand UO_4015 (O_4015,N_48737,N_43944);
xor UO_4016 (O_4016,N_44136,N_42744);
nand UO_4017 (O_4017,N_47623,N_43405);
xor UO_4018 (O_4018,N_44733,N_46959);
nand UO_4019 (O_4019,N_42682,N_44869);
and UO_4020 (O_4020,N_44757,N_46781);
and UO_4021 (O_4021,N_43533,N_42064);
or UO_4022 (O_4022,N_42699,N_46310);
or UO_4023 (O_4023,N_48259,N_44336);
or UO_4024 (O_4024,N_46648,N_45372);
and UO_4025 (O_4025,N_43830,N_49906);
nand UO_4026 (O_4026,N_46935,N_48963);
xor UO_4027 (O_4027,N_45953,N_48512);
nand UO_4028 (O_4028,N_48756,N_48483);
nand UO_4029 (O_4029,N_46283,N_42781);
xnor UO_4030 (O_4030,N_40931,N_42288);
nand UO_4031 (O_4031,N_43848,N_47680);
nand UO_4032 (O_4032,N_48555,N_44005);
xnor UO_4033 (O_4033,N_40542,N_42602);
or UO_4034 (O_4034,N_44148,N_48194);
nand UO_4035 (O_4035,N_46655,N_43889);
nor UO_4036 (O_4036,N_48818,N_48248);
nor UO_4037 (O_4037,N_41482,N_46714);
and UO_4038 (O_4038,N_43588,N_44075);
or UO_4039 (O_4039,N_46222,N_40344);
and UO_4040 (O_4040,N_40708,N_44608);
nor UO_4041 (O_4041,N_46861,N_42667);
or UO_4042 (O_4042,N_41090,N_43283);
nor UO_4043 (O_4043,N_44650,N_41177);
and UO_4044 (O_4044,N_42253,N_40241);
xor UO_4045 (O_4045,N_44365,N_49302);
or UO_4046 (O_4046,N_44105,N_43121);
or UO_4047 (O_4047,N_46496,N_45055);
nor UO_4048 (O_4048,N_45339,N_41305);
nor UO_4049 (O_4049,N_41767,N_40072);
nand UO_4050 (O_4050,N_41343,N_40530);
or UO_4051 (O_4051,N_45403,N_46659);
nand UO_4052 (O_4052,N_47375,N_43144);
xnor UO_4053 (O_4053,N_48026,N_42611);
and UO_4054 (O_4054,N_44044,N_45391);
nand UO_4055 (O_4055,N_41105,N_41083);
nand UO_4056 (O_4056,N_46575,N_49866);
or UO_4057 (O_4057,N_48525,N_44182);
nor UO_4058 (O_4058,N_44916,N_43517);
nand UO_4059 (O_4059,N_41450,N_49372);
xor UO_4060 (O_4060,N_40635,N_46643);
xor UO_4061 (O_4061,N_43778,N_40878);
nand UO_4062 (O_4062,N_49614,N_44253);
and UO_4063 (O_4063,N_47133,N_43055);
xor UO_4064 (O_4064,N_44398,N_40569);
nand UO_4065 (O_4065,N_44300,N_45843);
or UO_4066 (O_4066,N_41445,N_45123);
nand UO_4067 (O_4067,N_43978,N_42998);
nor UO_4068 (O_4068,N_41932,N_47727);
nand UO_4069 (O_4069,N_45803,N_45187);
or UO_4070 (O_4070,N_47417,N_43905);
and UO_4071 (O_4071,N_45913,N_45059);
and UO_4072 (O_4072,N_48719,N_41213);
xnor UO_4073 (O_4073,N_49156,N_48077);
nor UO_4074 (O_4074,N_48374,N_43422);
nor UO_4075 (O_4075,N_47256,N_49785);
nand UO_4076 (O_4076,N_44594,N_47602);
nor UO_4077 (O_4077,N_40871,N_49199);
and UO_4078 (O_4078,N_47303,N_48309);
or UO_4079 (O_4079,N_48018,N_47752);
and UO_4080 (O_4080,N_43721,N_40227);
xnor UO_4081 (O_4081,N_42862,N_46903);
and UO_4082 (O_4082,N_49442,N_47491);
or UO_4083 (O_4083,N_47548,N_42631);
and UO_4084 (O_4084,N_41850,N_42248);
nand UO_4085 (O_4085,N_42928,N_44580);
and UO_4086 (O_4086,N_42343,N_43729);
xnor UO_4087 (O_4087,N_45973,N_47164);
nand UO_4088 (O_4088,N_46526,N_45740);
nor UO_4089 (O_4089,N_46103,N_42612);
xnor UO_4090 (O_4090,N_41058,N_46388);
xor UO_4091 (O_4091,N_40626,N_48470);
or UO_4092 (O_4092,N_47485,N_47763);
and UO_4093 (O_4093,N_49400,N_49239);
and UO_4094 (O_4094,N_47907,N_48174);
nor UO_4095 (O_4095,N_42739,N_44292);
nand UO_4096 (O_4096,N_44809,N_46973);
xnor UO_4097 (O_4097,N_47317,N_44271);
nor UO_4098 (O_4098,N_42243,N_47543);
nand UO_4099 (O_4099,N_41670,N_44465);
nor UO_4100 (O_4100,N_46430,N_44885);
nand UO_4101 (O_4101,N_42676,N_42042);
and UO_4102 (O_4102,N_43647,N_47983);
or UO_4103 (O_4103,N_40596,N_40260);
nor UO_4104 (O_4104,N_41094,N_41138);
or UO_4105 (O_4105,N_49626,N_49397);
xnor UO_4106 (O_4106,N_47496,N_45217);
and UO_4107 (O_4107,N_41180,N_46058);
xor UO_4108 (O_4108,N_48332,N_48854);
nor UO_4109 (O_4109,N_46012,N_43390);
nor UO_4110 (O_4110,N_44007,N_42159);
nor UO_4111 (O_4111,N_49051,N_47482);
nand UO_4112 (O_4112,N_42455,N_49149);
xnor UO_4113 (O_4113,N_49742,N_46059);
nand UO_4114 (O_4114,N_46993,N_46931);
nor UO_4115 (O_4115,N_44334,N_41020);
or UO_4116 (O_4116,N_46604,N_43018);
and UO_4117 (O_4117,N_45253,N_41038);
nand UO_4118 (O_4118,N_48675,N_44457);
xor UO_4119 (O_4119,N_47254,N_43706);
nand UO_4120 (O_4120,N_47457,N_49472);
and UO_4121 (O_4121,N_49343,N_42507);
and UO_4122 (O_4122,N_44734,N_43604);
xor UO_4123 (O_4123,N_45763,N_41054);
xor UO_4124 (O_4124,N_40866,N_42424);
or UO_4125 (O_4125,N_46943,N_41390);
nor UO_4126 (O_4126,N_49717,N_41857);
nor UO_4127 (O_4127,N_43392,N_40966);
or UO_4128 (O_4128,N_46774,N_46900);
and UO_4129 (O_4129,N_44301,N_48541);
or UO_4130 (O_4130,N_48290,N_42530);
nand UO_4131 (O_4131,N_44203,N_44083);
and UO_4132 (O_4132,N_47735,N_47076);
or UO_4133 (O_4133,N_40195,N_48870);
or UO_4134 (O_4134,N_48482,N_44677);
and UO_4135 (O_4135,N_49658,N_48130);
nor UO_4136 (O_4136,N_49538,N_42287);
and UO_4137 (O_4137,N_43000,N_42749);
nor UO_4138 (O_4138,N_46651,N_42736);
xnor UO_4139 (O_4139,N_43240,N_41306);
and UO_4140 (O_4140,N_45783,N_47542);
nand UO_4141 (O_4141,N_48663,N_48224);
nand UO_4142 (O_4142,N_48000,N_46006);
nor UO_4143 (O_4143,N_48915,N_44684);
nand UO_4144 (O_4144,N_45911,N_44257);
or UO_4145 (O_4145,N_49992,N_41924);
nor UO_4146 (O_4146,N_42936,N_44035);
or UO_4147 (O_4147,N_40080,N_47384);
xnor UO_4148 (O_4148,N_47947,N_45245);
or UO_4149 (O_4149,N_41756,N_49925);
nand UO_4150 (O_4150,N_46092,N_41168);
xor UO_4151 (O_4151,N_42250,N_46881);
nor UO_4152 (O_4152,N_42668,N_47261);
nand UO_4153 (O_4153,N_49625,N_43506);
nor UO_4154 (O_4154,N_43395,N_45881);
or UO_4155 (O_4155,N_48022,N_40633);
nor UO_4156 (O_4156,N_46586,N_42479);
nand UO_4157 (O_4157,N_41729,N_49774);
xnor UO_4158 (O_4158,N_43085,N_42392);
or UO_4159 (O_4159,N_43804,N_43680);
xnor UO_4160 (O_4160,N_40086,N_49771);
or UO_4161 (O_4161,N_44419,N_43702);
nand UO_4162 (O_4162,N_43540,N_40879);
or UO_4163 (O_4163,N_46531,N_40576);
and UO_4164 (O_4164,N_41579,N_49985);
nor UO_4165 (O_4165,N_43714,N_47694);
nor UO_4166 (O_4166,N_41736,N_46628);
nand UO_4167 (O_4167,N_42223,N_48692);
and UO_4168 (O_4168,N_42013,N_46566);
or UO_4169 (O_4169,N_44191,N_49013);
or UO_4170 (O_4170,N_42306,N_40446);
or UO_4171 (O_4171,N_43554,N_41545);
nor UO_4172 (O_4172,N_47975,N_44689);
or UO_4173 (O_4173,N_49446,N_49912);
nand UO_4174 (O_4174,N_40876,N_46278);
or UO_4175 (O_4175,N_43857,N_44888);
nand UO_4176 (O_4176,N_46893,N_49762);
nor UO_4177 (O_4177,N_45656,N_45048);
and UO_4178 (O_4178,N_48072,N_47755);
or UO_4179 (O_4179,N_40230,N_41139);
or UO_4180 (O_4180,N_42270,N_41315);
and UO_4181 (O_4181,N_40173,N_45782);
nand UO_4182 (O_4182,N_49797,N_40937);
nand UO_4183 (O_4183,N_48516,N_44699);
nand UO_4184 (O_4184,N_41633,N_48626);
and UO_4185 (O_4185,N_45231,N_42999);
nand UO_4186 (O_4186,N_44544,N_43656);
nand UO_4187 (O_4187,N_44467,N_45599);
or UO_4188 (O_4188,N_42743,N_40062);
nand UO_4189 (O_4189,N_43227,N_40210);
or UO_4190 (O_4190,N_47204,N_40730);
xor UO_4191 (O_4191,N_43620,N_43176);
or UO_4192 (O_4192,N_41908,N_40884);
nand UO_4193 (O_4193,N_49362,N_48099);
xor UO_4194 (O_4194,N_46254,N_46743);
nand UO_4195 (O_4195,N_40539,N_47313);
or UO_4196 (O_4196,N_42842,N_46328);
nand UO_4197 (O_4197,N_44872,N_43126);
and UO_4198 (O_4198,N_42191,N_42600);
or UO_4199 (O_4199,N_46838,N_45503);
and UO_4200 (O_4200,N_49979,N_48888);
or UO_4201 (O_4201,N_42022,N_44928);
and UO_4202 (O_4202,N_41148,N_40531);
or UO_4203 (O_4203,N_41906,N_48116);
nor UO_4204 (O_4204,N_46276,N_44704);
nor UO_4205 (O_4205,N_45683,N_47577);
nand UO_4206 (O_4206,N_40203,N_45251);
nor UO_4207 (O_4207,N_44749,N_44918);
or UO_4208 (O_4208,N_42912,N_43683);
nor UO_4209 (O_4209,N_44034,N_46294);
nor UO_4210 (O_4210,N_45849,N_45546);
nand UO_4211 (O_4211,N_47040,N_45582);
and UO_4212 (O_4212,N_44503,N_42174);
and UO_4213 (O_4213,N_43095,N_44415);
or UO_4214 (O_4214,N_43910,N_41393);
and UO_4215 (O_4215,N_40788,N_41127);
or UO_4216 (O_4216,N_42127,N_42101);
and UO_4217 (O_4217,N_42814,N_48223);
or UO_4218 (O_4218,N_49827,N_43877);
nor UO_4219 (O_4219,N_40619,N_43241);
or UO_4220 (O_4220,N_44972,N_48829);
and UO_4221 (O_4221,N_48612,N_42367);
nor UO_4222 (O_4222,N_47340,N_40168);
or UO_4223 (O_4223,N_40889,N_45743);
and UO_4224 (O_4224,N_42423,N_43602);
and UO_4225 (O_4225,N_42003,N_44165);
nand UO_4226 (O_4226,N_46205,N_41740);
nand UO_4227 (O_4227,N_42897,N_43670);
and UO_4228 (O_4228,N_43575,N_43896);
nor UO_4229 (O_4229,N_42791,N_40614);
nand UO_4230 (O_4230,N_47711,N_49132);
nand UO_4231 (O_4231,N_47306,N_45955);
and UO_4232 (O_4232,N_47210,N_40254);
nand UO_4233 (O_4233,N_45833,N_40257);
and UO_4234 (O_4234,N_44800,N_44466);
xnor UO_4235 (O_4235,N_43556,N_44727);
nand UO_4236 (O_4236,N_40598,N_43288);
and UO_4237 (O_4237,N_44946,N_44940);
or UO_4238 (O_4238,N_43955,N_48940);
nand UO_4239 (O_4239,N_44970,N_44361);
nor UO_4240 (O_4240,N_43257,N_49629);
nand UO_4241 (O_4241,N_44474,N_45484);
xnor UO_4242 (O_4242,N_43951,N_40893);
or UO_4243 (O_4243,N_46664,N_46003);
and UO_4244 (O_4244,N_40146,N_41839);
and UO_4245 (O_4245,N_41510,N_41781);
or UO_4246 (O_4246,N_45252,N_41008);
nand UO_4247 (O_4247,N_45291,N_45998);
nor UO_4248 (O_4248,N_43614,N_48233);
nor UO_4249 (O_4249,N_49398,N_43162);
and UO_4250 (O_4250,N_49953,N_48868);
or UO_4251 (O_4251,N_41650,N_44542);
or UO_4252 (O_4252,N_46480,N_47793);
nor UO_4253 (O_4253,N_42856,N_45345);
nand UO_4254 (O_4254,N_47379,N_47900);
and UO_4255 (O_4255,N_42576,N_45781);
nand UO_4256 (O_4256,N_48590,N_42259);
nor UO_4257 (O_4257,N_45080,N_45635);
and UO_4258 (O_4258,N_41934,N_45949);
and UO_4259 (O_4259,N_42984,N_41027);
nor UO_4260 (O_4260,N_43668,N_40685);
nand UO_4261 (O_4261,N_49859,N_40844);
nand UO_4262 (O_4262,N_49118,N_49408);
nand UO_4263 (O_4263,N_47257,N_42663);
or UO_4264 (O_4264,N_42019,N_42675);
nand UO_4265 (O_4265,N_46064,N_41637);
nand UO_4266 (O_4266,N_47364,N_42863);
nor UO_4267 (O_4267,N_48878,N_49467);
nor UO_4268 (O_4268,N_47038,N_43201);
nand UO_4269 (O_4269,N_42871,N_43230);
nand UO_4270 (O_4270,N_43370,N_43784);
nand UO_4271 (O_4271,N_42916,N_44863);
nand UO_4272 (O_4272,N_43639,N_42381);
nor UO_4273 (O_4273,N_48379,N_46063);
nor UO_4274 (O_4274,N_43547,N_43281);
and UO_4275 (O_4275,N_41272,N_40351);
nand UO_4276 (O_4276,N_44604,N_45125);
nand UO_4277 (O_4277,N_41425,N_47478);
nor UO_4278 (O_4278,N_41170,N_43307);
or UO_4279 (O_4279,N_42027,N_42433);
and UO_4280 (O_4280,N_44904,N_46171);
nor UO_4281 (O_4281,N_49661,N_42567);
or UO_4282 (O_4282,N_44859,N_47495);
nor UO_4283 (O_4283,N_48872,N_44624);
nand UO_4284 (O_4284,N_44576,N_44383);
or UO_4285 (O_4285,N_49496,N_43576);
nand UO_4286 (O_4286,N_47186,N_40247);
nand UO_4287 (O_4287,N_40299,N_44753);
nand UO_4288 (O_4288,N_44603,N_40785);
nand UO_4289 (O_4289,N_45994,N_44084);
or UO_4290 (O_4290,N_45052,N_44773);
nand UO_4291 (O_4291,N_47994,N_47224);
or UO_4292 (O_4292,N_44185,N_47439);
xnor UO_4293 (O_4293,N_41572,N_48021);
nand UO_4294 (O_4294,N_40632,N_44736);
xor UO_4295 (O_4295,N_45586,N_42852);
nand UO_4296 (O_4296,N_40607,N_43876);
xnor UO_4297 (O_4297,N_48258,N_43204);
and UO_4298 (O_4298,N_45553,N_47963);
nor UO_4299 (O_4299,N_41403,N_48842);
nor UO_4300 (O_4300,N_46239,N_41489);
nor UO_4301 (O_4301,N_48615,N_49414);
nand UO_4302 (O_4302,N_46023,N_43834);
nor UO_4303 (O_4303,N_43878,N_41304);
and UO_4304 (O_4304,N_40741,N_45406);
or UO_4305 (O_4305,N_42305,N_49335);
or UO_4306 (O_4306,N_49539,N_45004);
or UO_4307 (O_4307,N_49251,N_40426);
nor UO_4308 (O_4308,N_41962,N_41235);
nor UO_4309 (O_4309,N_48631,N_43926);
nor UO_4310 (O_4310,N_47031,N_43094);
nor UO_4311 (O_4311,N_45901,N_47289);
nand UO_4312 (O_4312,N_40149,N_48006);
xor UO_4313 (O_4313,N_46535,N_44321);
nor UO_4314 (O_4314,N_42919,N_47232);
nor UO_4315 (O_4315,N_42500,N_42751);
and UO_4316 (O_4316,N_47147,N_43006);
nand UO_4317 (O_4317,N_48237,N_43021);
nor UO_4318 (O_4318,N_40863,N_45719);
nand UO_4319 (O_4319,N_42589,N_44307);
nand UO_4320 (O_4320,N_40620,N_41721);
nor UO_4321 (O_4321,N_43898,N_49684);
or UO_4322 (O_4322,N_49523,N_49443);
nand UO_4323 (O_4323,N_48618,N_45468);
nor UO_4324 (O_4324,N_45896,N_44698);
nand UO_4325 (O_4325,N_42949,N_44177);
nand UO_4326 (O_4326,N_43746,N_49996);
nand UO_4327 (O_4327,N_47648,N_43601);
nand UO_4328 (O_4328,N_46343,N_40853);
or UO_4329 (O_4329,N_49377,N_41254);
and UO_4330 (O_4330,N_45210,N_45812);
nor UO_4331 (O_4331,N_49192,N_46770);
nor UO_4332 (O_4332,N_49864,N_49001);
nor UO_4333 (O_4333,N_49853,N_40472);
and UO_4334 (O_4334,N_45662,N_40130);
nand UO_4335 (O_4335,N_43198,N_41262);
xor UO_4336 (O_4336,N_47512,N_48566);
or UO_4337 (O_4337,N_42226,N_43479);
and UO_4338 (O_4338,N_48557,N_47925);
xnor UO_4339 (O_4339,N_43949,N_49518);
xnor UO_4340 (O_4340,N_44999,N_42673);
xnor UO_4341 (O_4341,N_48240,N_40114);
nand UO_4342 (O_4342,N_48794,N_44654);
nand UO_4343 (O_4343,N_49254,N_42921);
nand UO_4344 (O_4344,N_42493,N_49144);
or UO_4345 (O_4345,N_48193,N_40116);
nor UO_4346 (O_4346,N_42227,N_44656);
or UO_4347 (O_4347,N_48311,N_44135);
and UO_4348 (O_4348,N_49115,N_44517);
and UO_4349 (O_4349,N_47139,N_45947);
or UO_4350 (O_4350,N_46539,N_47065);
nor UO_4351 (O_4351,N_47578,N_48410);
or UO_4352 (O_4352,N_40052,N_45072);
nor UO_4353 (O_4353,N_42623,N_49815);
or UO_4354 (O_4354,N_40425,N_41705);
nor UO_4355 (O_4355,N_46114,N_44772);
and UO_4356 (O_4356,N_44413,N_47635);
nand UO_4357 (O_4357,N_40352,N_45083);
nor UO_4358 (O_4358,N_42029,N_47001);
and UO_4359 (O_4359,N_42508,N_49285);
nand UO_4360 (O_4360,N_43768,N_41975);
nand UO_4361 (O_4361,N_45005,N_40608);
nand UO_4362 (O_4362,N_47358,N_48998);
nand UO_4363 (O_4363,N_43871,N_41980);
and UO_4364 (O_4364,N_43233,N_42694);
or UO_4365 (O_4365,N_43159,N_40573);
nor UO_4366 (O_4366,N_48894,N_42588);
or UO_4367 (O_4367,N_48214,N_48681);
nand UO_4368 (O_4368,N_43851,N_40381);
nand UO_4369 (O_4369,N_47129,N_46141);
nand UO_4370 (O_4370,N_42282,N_41706);
and UO_4371 (O_4371,N_43342,N_47629);
nor UO_4372 (O_4372,N_40698,N_49883);
xor UO_4373 (O_4373,N_45311,N_41149);
nand UO_4374 (O_4374,N_44272,N_48373);
nor UO_4375 (O_4375,N_42097,N_47556);
and UO_4376 (O_4376,N_42804,N_48790);
and UO_4377 (O_4377,N_48360,N_49709);
nor UO_4378 (O_4378,N_40000,N_47302);
nor UO_4379 (O_4379,N_44526,N_40095);
nand UO_4380 (O_4380,N_49601,N_45248);
or UO_4381 (O_4381,N_46049,N_41446);
or UO_4382 (O_4382,N_41771,N_49511);
nand UO_4383 (O_4383,N_48091,N_40860);
and UO_4384 (O_4384,N_43504,N_47846);
nand UO_4385 (O_4385,N_46405,N_43163);
or UO_4386 (O_4386,N_47611,N_41519);
or UO_4387 (O_4387,N_46042,N_43210);
nor UO_4388 (O_4388,N_45897,N_41249);
and UO_4389 (O_4389,N_45521,N_42648);
and UO_4390 (O_4390,N_48029,N_48226);
nand UO_4391 (O_4391,N_45701,N_41398);
nor UO_4392 (O_4392,N_43755,N_41500);
or UO_4393 (O_4393,N_47219,N_47192);
nor UO_4394 (O_4394,N_49028,N_49775);
nand UO_4395 (O_4395,N_41297,N_49759);
and UO_4396 (O_4396,N_42590,N_48039);
nand UO_4397 (O_4397,N_44046,N_46843);
and UO_4398 (O_4398,N_42758,N_48069);
xor UO_4399 (O_4399,N_41101,N_42902);
nand UO_4400 (O_4400,N_48519,N_41401);
or UO_4401 (O_4401,N_46142,N_45145);
nand UO_4402 (O_4402,N_45749,N_46291);
and UO_4403 (O_4403,N_48450,N_45909);
and UO_4404 (O_4404,N_41295,N_43446);
or UO_4405 (O_4405,N_44806,N_45475);
nor UO_4406 (O_4406,N_43039,N_41122);
and UO_4407 (O_4407,N_42888,N_44097);
and UO_4408 (O_4408,N_41220,N_40182);
and UO_4409 (O_4409,N_47967,N_48680);
nor UO_4410 (O_4410,N_47480,N_41570);
and UO_4411 (O_4411,N_41710,N_49852);
xnor UO_4412 (O_4412,N_44511,N_42618);
nor UO_4413 (O_4413,N_41773,N_47448);
and UO_4414 (O_4414,N_48317,N_46721);
xor UO_4415 (O_4415,N_43562,N_40017);
nor UO_4416 (O_4416,N_40506,N_45882);
nor UO_4417 (O_4417,N_48575,N_47746);
and UO_4418 (O_4418,N_43070,N_47919);
and UO_4419 (O_4419,N_44195,N_48306);
and UO_4420 (O_4420,N_42490,N_44080);
nor UO_4421 (O_4421,N_43536,N_41216);
or UO_4422 (O_4422,N_44114,N_48905);
nor UO_4423 (O_4423,N_47558,N_45774);
nor UO_4424 (O_4424,N_41345,N_42651);
nand UO_4425 (O_4425,N_44495,N_41448);
nor UO_4426 (O_4426,N_40546,N_44320);
nor UO_4427 (O_4427,N_43362,N_48735);
nor UO_4428 (O_4428,N_44662,N_42153);
nor UO_4429 (O_4429,N_49643,N_42043);
and UO_4430 (O_4430,N_41720,N_47890);
nor UO_4431 (O_4431,N_41965,N_46610);
xor UO_4432 (O_4432,N_48823,N_47898);
nand UO_4433 (O_4433,N_45154,N_44081);
nor UO_4434 (O_4434,N_42063,N_43117);
nor UO_4435 (O_4435,N_45835,N_46397);
and UO_4436 (O_4436,N_43561,N_42391);
or UO_4437 (O_4437,N_40864,N_41918);
nand UO_4438 (O_4438,N_47716,N_46227);
nand UO_4439 (O_4439,N_40836,N_47760);
and UO_4440 (O_4440,N_41136,N_40839);
or UO_4441 (O_4441,N_47853,N_40486);
nor UO_4442 (O_4442,N_46756,N_47443);
nand UO_4443 (O_4443,N_45240,N_42834);
nor UO_4444 (O_4444,N_41486,N_43336);
nor UO_4445 (O_4445,N_47465,N_41995);
nor UO_4446 (O_4446,N_45013,N_43024);
nor UO_4447 (O_4447,N_41668,N_41909);
nor UO_4448 (O_4448,N_48220,N_44204);
nand UO_4449 (O_4449,N_47190,N_43106);
and UO_4450 (O_4450,N_42772,N_44746);
or UO_4451 (O_4451,N_40601,N_41253);
nand UO_4452 (O_4452,N_44173,N_48717);
and UO_4453 (O_4453,N_46281,N_49739);
and UO_4454 (O_4454,N_43931,N_49994);
and UO_4455 (O_4455,N_41391,N_45158);
and UO_4456 (O_4456,N_45100,N_44756);
or UO_4457 (O_4457,N_48330,N_49901);
and UO_4458 (O_4458,N_45900,N_43616);
and UO_4459 (O_4459,N_44373,N_49230);
or UO_4460 (O_4460,N_48395,N_41159);
and UO_4461 (O_4461,N_49733,N_44793);
xnor UO_4462 (O_4462,N_48508,N_46877);
nand UO_4463 (O_4463,N_46591,N_42012);
or UO_4464 (O_4464,N_43597,N_44142);
and UO_4465 (O_4465,N_48887,N_47725);
xor UO_4466 (O_4466,N_43794,N_48441);
xnor UO_4467 (O_4467,N_48070,N_44348);
xor UO_4468 (O_4468,N_49152,N_45866);
nor UO_4469 (O_4469,N_45670,N_41954);
nand UO_4470 (O_4470,N_47288,N_48312);
nand UO_4471 (O_4471,N_46926,N_44294);
nand UO_4472 (O_4472,N_41483,N_43173);
or UO_4473 (O_4473,N_47819,N_48921);
nand UO_4474 (O_4474,N_46752,N_44217);
and UO_4475 (O_4475,N_41587,N_47134);
xor UO_4476 (O_4476,N_43762,N_49935);
or UO_4477 (O_4477,N_45512,N_47700);
nand UO_4478 (O_4478,N_40867,N_45459);
nand UO_4479 (O_4479,N_41433,N_42018);
or UO_4480 (O_4480,N_41963,N_41632);
nand UO_4481 (O_4481,N_42793,N_40285);
nand UO_4482 (O_4482,N_48924,N_46094);
and UO_4483 (O_4483,N_48281,N_49222);
nor UO_4484 (O_4484,N_42810,N_41392);
or UO_4485 (O_4485,N_48078,N_44739);
nand UO_4486 (O_4486,N_43615,N_46209);
nor UO_4487 (O_4487,N_45970,N_48139);
nor UO_4488 (O_4488,N_41463,N_43571);
xnor UO_4489 (O_4489,N_40107,N_44420);
xor UO_4490 (O_4490,N_43492,N_47467);
nand UO_4491 (O_4491,N_44519,N_44775);
and UO_4492 (O_4492,N_48113,N_43573);
nor UO_4493 (O_4493,N_42628,N_44066);
or UO_4494 (O_4494,N_41388,N_45076);
nor UO_4495 (O_4495,N_48028,N_47554);
and UO_4496 (O_4496,N_43705,N_44824);
and UO_4497 (O_4497,N_47613,N_40374);
nor UO_4498 (O_4498,N_46863,N_42908);
nand UO_4499 (O_4499,N_46192,N_48911);
or UO_4500 (O_4500,N_43698,N_43751);
nor UO_4501 (O_4501,N_40371,N_42471);
or UO_4502 (O_4502,N_49018,N_43580);
nand UO_4503 (O_4503,N_45702,N_42769);
or UO_4504 (O_4504,N_48187,N_46980);
xnor UO_4505 (O_4505,N_44984,N_48504);
nand UO_4506 (O_4506,N_44078,N_43622);
nor UO_4507 (O_4507,N_40029,N_45364);
nor UO_4508 (O_4508,N_41207,N_45426);
and UO_4509 (O_4509,N_41423,N_45711);
nor UO_4510 (O_4510,N_40777,N_42669);
and UO_4511 (O_4511,N_46833,N_42214);
and UO_4512 (O_4512,N_47785,N_49065);
xnor UO_4513 (O_4513,N_48067,N_46622);
or UO_4514 (O_4514,N_48755,N_42370);
nor UO_4515 (O_4515,N_46386,N_42472);
nor UO_4516 (O_4516,N_46195,N_48799);
nand UO_4517 (O_4517,N_48185,N_48153);
nor UO_4518 (O_4518,N_48751,N_41997);
and UO_4519 (O_4519,N_49908,N_43496);
nor UO_4520 (O_4520,N_41046,N_41903);
and UO_4521 (O_4521,N_43246,N_45432);
and UO_4522 (O_4522,N_48457,N_41222);
xor UO_4523 (O_4523,N_45614,N_47258);
nor UO_4524 (O_4524,N_41040,N_46101);
nor UO_4525 (O_4525,N_49627,N_43648);
nor UO_4526 (O_4526,N_42523,N_40125);
or UO_4527 (O_4527,N_47110,N_44549);
or UO_4528 (O_4528,N_41606,N_47910);
nor UO_4529 (O_4529,N_44386,N_47479);
or UO_4530 (O_4530,N_47913,N_46233);
nor UO_4531 (O_4531,N_45348,N_46285);
xnor UO_4532 (O_4532,N_42801,N_42698);
xnor UO_4533 (O_4533,N_47671,N_45098);
and UO_4534 (O_4534,N_43929,N_43769);
nor UO_4535 (O_4535,N_44444,N_40384);
nor UO_4536 (O_4536,N_47585,N_46849);
nor UO_4537 (O_4537,N_40651,N_46210);
nand UO_4538 (O_4538,N_42964,N_44996);
or UO_4539 (O_4539,N_43924,N_42313);
nor UO_4540 (O_4540,N_46600,N_40832);
nor UO_4541 (O_4541,N_48211,N_45969);
nand UO_4542 (O_4542,N_45313,N_41760);
nand UO_4543 (O_4543,N_49615,N_42026);
nand UO_4544 (O_4544,N_45550,N_46411);
and UO_4545 (O_4545,N_44428,N_49971);
nor UO_4546 (O_4546,N_49754,N_40156);
nand UO_4547 (O_4547,N_49309,N_47751);
nor UO_4548 (O_4548,N_48700,N_40528);
nor UO_4549 (O_4549,N_44119,N_46123);
nor UO_4550 (O_4550,N_46920,N_40786);
or UO_4551 (O_4551,N_41115,N_48722);
nor UO_4552 (O_4552,N_40705,N_48283);
nor UO_4553 (O_4553,N_48966,N_40512);
nand UO_4554 (O_4554,N_40379,N_40470);
or UO_4555 (O_4555,N_48629,N_42481);
nand UO_4556 (O_4556,N_41967,N_42545);
and UO_4557 (O_4557,N_44127,N_44400);
nand UO_4558 (O_4558,N_48007,N_47764);
nand UO_4559 (O_4559,N_48596,N_44438);
nand UO_4560 (O_4560,N_48916,N_46961);
nor UO_4561 (O_4561,N_49877,N_41628);
xor UO_4562 (O_4562,N_46352,N_48102);
nor UO_4563 (O_4563,N_41905,N_40093);
and UO_4564 (O_4564,N_41327,N_42204);
nor UO_4565 (O_4565,N_49727,N_47278);
and UO_4566 (O_4566,N_49662,N_49059);
nand UO_4567 (O_4567,N_48529,N_48404);
and UO_4568 (O_4568,N_49752,N_49665);
xnor UO_4569 (O_4569,N_48115,N_48446);
xnor UO_4570 (O_4570,N_47463,N_46342);
nor UO_4571 (O_4571,N_42398,N_40883);
nor UO_4572 (O_4572,N_42036,N_49184);
or UO_4573 (O_4573,N_47704,N_49509);
and UO_4574 (O_4574,N_42413,N_41418);
nor UO_4575 (O_4575,N_41817,N_45164);
and UO_4576 (O_4576,N_49934,N_45513);
nor UO_4577 (O_4577,N_45332,N_40219);
and UO_4578 (O_4578,N_48537,N_47879);
and UO_4579 (O_4579,N_47990,N_43139);
nor UO_4580 (O_4580,N_45730,N_47993);
nand UO_4581 (O_4581,N_40393,N_45259);
nor UO_4582 (O_4582,N_46772,N_44472);
xor UO_4583 (O_4583,N_44202,N_42869);
and UO_4584 (O_4584,N_45647,N_42234);
or UO_4585 (O_4585,N_46614,N_47788);
nor UO_4586 (O_4586,N_44868,N_44404);
nor UO_4587 (O_4587,N_46154,N_45936);
and UO_4588 (O_4588,N_45862,N_42569);
nor UO_4589 (O_4589,N_41191,N_46793);
nand UO_4590 (O_4590,N_41996,N_48906);
or UO_4591 (O_4591,N_40686,N_47800);
nand UO_4592 (O_4592,N_41684,N_41950);
nand UO_4593 (O_4593,N_46924,N_41051);
nand UO_4594 (O_4594,N_40723,N_43795);
or UO_4595 (O_4595,N_46056,N_46862);
nor UO_4596 (O_4596,N_40205,N_41064);
nand UO_4597 (O_4597,N_41948,N_41037);
or UO_4598 (O_4598,N_49454,N_41171);
or UO_4599 (O_4599,N_43481,N_48785);
nor UO_4600 (O_4600,N_48147,N_45858);
nor UO_4601 (O_4601,N_41041,N_49640);
xor UO_4602 (O_4602,N_48127,N_48601);
nand UO_4603 (O_4603,N_44461,N_46819);
or UO_4604 (O_4604,N_43903,N_42575);
nand UO_4605 (O_4605,N_49685,N_46969);
nand UO_4606 (O_4606,N_48811,N_45378);
and UO_4607 (O_4607,N_40238,N_46540);
nor UO_4608 (O_4608,N_47770,N_47709);
or UO_4609 (O_4609,N_49682,N_44290);
nor UO_4610 (O_4610,N_49960,N_48926);
nor UO_4611 (O_4611,N_44575,N_48577);
or UO_4612 (O_4612,N_48881,N_47987);
nand UO_4613 (O_4613,N_48807,N_42685);
nor UO_4614 (O_4614,N_48278,N_43130);
nand UO_4615 (O_4615,N_45093,N_43361);
xor UO_4616 (O_4616,N_42807,N_42906);
and UO_4617 (O_4617,N_40553,N_47736);
and UO_4618 (O_4618,N_49620,N_46174);
and UO_4619 (O_4619,N_48573,N_44285);
and UO_4620 (O_4620,N_48146,N_41878);
nand UO_4621 (O_4621,N_47710,N_44719);
nor UO_4622 (O_4622,N_45149,N_46251);
or UO_4623 (O_4623,N_43344,N_49923);
nor UO_4624 (O_4624,N_42334,N_41504);
xor UO_4625 (O_4625,N_45530,N_41317);
nand UO_4626 (O_4626,N_45899,N_43260);
nor UO_4627 (O_4627,N_40190,N_41205);
and UO_4628 (O_4628,N_44490,N_40455);
nor UO_4629 (O_4629,N_46175,N_42186);
and UO_4630 (O_4630,N_45377,N_41440);
and UO_4631 (O_4631,N_45078,N_48101);
xor UO_4632 (O_4632,N_42613,N_46312);
or UO_4633 (O_4633,N_49404,N_48399);
nor UO_4634 (O_4634,N_40789,N_48633);
and UO_4635 (O_4635,N_44880,N_44158);
and UO_4636 (O_4636,N_49416,N_42124);
nand UO_4637 (O_4637,N_44479,N_49331);
nand UO_4638 (O_4638,N_47855,N_41242);
and UO_4639 (O_4639,N_44543,N_44625);
and UO_4640 (O_4640,N_46603,N_42028);
or UO_4641 (O_4641,N_47809,N_41334);
nor UO_4642 (O_4642,N_42337,N_42564);
and UO_4643 (O_4643,N_44275,N_46915);
nand UO_4644 (O_4644,N_48266,N_42816);
nand UO_4645 (O_4645,N_49127,N_48743);
and UO_4646 (O_4646,N_43691,N_46631);
and UO_4647 (O_4647,N_47041,N_40852);
xor UO_4648 (O_4648,N_41513,N_48723);
and UO_4649 (O_4649,N_46314,N_43396);
nand UO_4650 (O_4650,N_49474,N_48979);
nor UO_4651 (O_4651,N_44132,N_41121);
xor UO_4652 (O_4652,N_45828,N_44961);
nor UO_4653 (O_4653,N_42965,N_40011);
and UO_4654 (O_4654,N_41852,N_48289);
xor UO_4655 (O_4655,N_43657,N_48438);
nand UO_4656 (O_4656,N_49534,N_45661);
nor UO_4657 (O_4657,N_45105,N_45360);
or UO_4658 (O_4658,N_41951,N_47836);
nand UO_4659 (O_4659,N_47864,N_49540);
nand UO_4660 (O_4660,N_42262,N_42065);
or UO_4661 (O_4661,N_46391,N_44579);
nand UO_4662 (O_4662,N_43432,N_44192);
or UO_4663 (O_4663,N_43129,N_48424);
and UO_4664 (O_4664,N_49029,N_42178);
nor UO_4665 (O_4665,N_48405,N_40261);
or UO_4666 (O_4666,N_43730,N_45212);
and UO_4667 (O_4667,N_44694,N_48376);
nand UO_4668 (O_4668,N_40318,N_48064);
and UO_4669 (O_4669,N_44427,N_44055);
xnor UO_4670 (O_4670,N_46950,N_43141);
xor UO_4671 (O_4671,N_42076,N_40010);
xnor UO_4672 (O_4672,N_43788,N_45902);
nand UO_4673 (O_4673,N_47327,N_46632);
or UO_4674 (O_4674,N_40724,N_43076);
or UO_4675 (O_4675,N_41944,N_41241);
nand UO_4676 (O_4676,N_40221,N_43433);
nand UO_4677 (O_4677,N_49057,N_49498);
and UO_4678 (O_4678,N_42163,N_44138);
nand UO_4679 (O_4679,N_44821,N_44917);
and UO_4680 (O_4680,N_40432,N_41711);
nand UO_4681 (O_4681,N_47681,N_45201);
nand UO_4682 (O_4682,N_41356,N_41412);
or UO_4683 (O_4683,N_48440,N_44830);
or UO_4684 (O_4684,N_45215,N_40537);
nor UO_4685 (O_4685,N_42541,N_46824);
and UO_4686 (O_4686,N_42581,N_45779);
xnor UO_4687 (O_4687,N_47370,N_44891);
or UO_4688 (O_4688,N_46713,N_45706);
or UO_4689 (O_4689,N_45420,N_40265);
nor UO_4690 (O_4690,N_42597,N_40479);
and UO_4691 (O_4691,N_41984,N_46832);
or UO_4692 (O_4692,N_44215,N_42599);
nor UO_4693 (O_4693,N_41983,N_48121);
or UO_4694 (O_4694,N_46668,N_44778);
and UO_4695 (O_4695,N_45593,N_40180);
nand UO_4696 (O_4696,N_40289,N_49814);
nor UO_4697 (O_4697,N_47502,N_40949);
nand UO_4698 (O_4698,N_49750,N_43791);
or UO_4699 (O_4699,N_49214,N_40081);
nand UO_4700 (O_4700,N_49564,N_44421);
nand UO_4701 (O_4701,N_49470,N_48898);
nor UO_4702 (O_4702,N_40347,N_43516);
and UO_4703 (O_4703,N_42200,N_43986);
or UO_4704 (O_4704,N_44218,N_46996);
or UO_4705 (O_4705,N_42645,N_40373);
and UO_4706 (O_4706,N_41719,N_44462);
or UO_4707 (O_4707,N_42418,N_48804);
nand UO_4708 (O_4708,N_41512,N_40641);
nor UO_4709 (O_4709,N_44003,N_44344);
xor UO_4710 (O_4710,N_45414,N_45448);
xor UO_4711 (O_4711,N_43676,N_46518);
or UO_4712 (O_4712,N_44981,N_44234);
nor UO_4713 (O_4713,N_44633,N_48472);
or UO_4714 (O_4714,N_47052,N_43609);
or UO_4715 (O_4715,N_42506,N_45450);
nor UO_4716 (O_4716,N_49777,N_48105);
and UO_4717 (O_4717,N_48918,N_48300);
nand UO_4718 (O_4718,N_47165,N_40978);
nor UO_4719 (O_4719,N_44896,N_47969);
xor UO_4720 (O_4720,N_48235,N_46295);
and UO_4721 (O_4721,N_47783,N_42453);
and UO_4722 (O_4722,N_47405,N_48613);
or UO_4723 (O_4723,N_40637,N_40166);
and UO_4724 (O_4724,N_48221,N_48086);
or UO_4725 (O_4725,N_48795,N_40496);
or UO_4726 (O_4726,N_43560,N_43292);
nor UO_4727 (O_4727,N_46317,N_42372);
or UO_4728 (O_4728,N_47382,N_48184);
or UO_4729 (O_4729,N_45588,N_43617);
nand UO_4730 (O_4730,N_49379,N_43065);
and UO_4731 (O_4731,N_43069,N_42686);
and UO_4732 (O_4732,N_47533,N_46412);
or UO_4733 (O_4733,N_45569,N_44452);
nand UO_4734 (O_4734,N_43864,N_40215);
nand UO_4735 (O_4735,N_40829,N_49151);
nor UO_4736 (O_4736,N_40900,N_41582);
nor UO_4737 (O_4737,N_44013,N_47017);
nand UO_4738 (O_4738,N_46986,N_43827);
xor UO_4739 (O_4739,N_40603,N_44130);
nor UO_4740 (O_4740,N_46009,N_40940);
or UO_4741 (O_4741,N_41044,N_47677);
or UO_4742 (O_4742,N_45436,N_43923);
nor UO_4743 (O_4743,N_48995,N_40420);
or UO_4744 (O_4744,N_46346,N_48920);
xnor UO_4745 (O_4745,N_49208,N_48344);
or UO_4746 (O_4746,N_44683,N_45267);
nor UO_4747 (O_4747,N_42940,N_48382);
and UO_4748 (O_4748,N_48485,N_48431);
nand UO_4749 (O_4749,N_41067,N_43652);
nand UO_4750 (O_4750,N_47453,N_42379);
nor UO_4751 (O_4751,N_48453,N_47739);
nand UO_4752 (O_4752,N_41256,N_41066);
xor UO_4753 (O_4753,N_41977,N_49899);
nor UO_4754 (O_4754,N_40566,N_48270);
nand UO_4755 (O_4755,N_47082,N_47726);
or UO_4756 (O_4756,N_41488,N_41089);
nor UO_4757 (O_4757,N_46368,N_47862);
and UO_4758 (O_4758,N_41444,N_45699);
and UO_4759 (O_4759,N_42414,N_40865);
nand UO_4760 (O_4760,N_40548,N_47209);
or UO_4761 (O_4761,N_44430,N_44567);
nand UO_4762 (O_4762,N_46948,N_48433);
and UO_4763 (O_4763,N_44367,N_48316);
or UO_4764 (O_4764,N_49165,N_41436);
and UO_4765 (O_4765,N_46451,N_44554);
nor UO_4766 (O_4766,N_45634,N_48594);
or UO_4767 (O_4767,N_43645,N_49856);
and UO_4768 (O_4768,N_43066,N_40720);
nand UO_4769 (O_4769,N_46623,N_46884);
nor UO_4770 (O_4770,N_43720,N_40309);
nand UO_4771 (O_4771,N_49936,N_42741);
nor UO_4772 (O_4772,N_44520,N_49212);
nor UO_4773 (O_4773,N_42454,N_45999);
and UO_4774 (O_4774,N_48654,N_45237);
and UO_4775 (O_4775,N_46682,N_43740);
and UO_4776 (O_4776,N_48189,N_41573);
nor UO_4777 (O_4777,N_48004,N_40074);
xnor UO_4778 (O_4778,N_46644,N_43799);
or UO_4779 (O_4779,N_42811,N_42274);
nand UO_4780 (O_4780,N_47046,N_43552);
nor UO_4781 (O_4781,N_42484,N_49188);
and UO_4782 (O_4782,N_43399,N_43214);
nor UO_4783 (O_4783,N_48925,N_45619);
nand UO_4784 (O_4784,N_46021,N_42323);
and UO_4785 (O_4785,N_49806,N_47588);
and UO_4786 (O_4786,N_44038,N_45817);
and UO_4787 (O_4787,N_45465,N_48988);
nor UO_4788 (O_4788,N_47080,N_45523);
or UO_4789 (O_4789,N_46923,N_41698);
or UO_4790 (O_4790,N_45735,N_46825);
nor UO_4791 (O_4791,N_41568,N_45140);
nand UO_4792 (O_4792,N_43789,N_45710);
and UO_4793 (O_4793,N_44593,N_42134);
or UO_4794 (O_4794,N_41335,N_44445);
nor UO_4795 (O_4795,N_46124,N_49000);
nor UO_4796 (O_4796,N_49154,N_44784);
nand UO_4797 (O_4797,N_43277,N_40102);
or UO_4798 (O_4798,N_43046,N_42692);
nor UO_4799 (O_4799,N_46991,N_40198);
and UO_4800 (O_4800,N_49623,N_48897);
nor UO_4801 (O_4801,N_44120,N_49288);
nand UO_4802 (O_4802,N_48093,N_44710);
xor UO_4803 (O_4803,N_44788,N_48444);
nor UO_4804 (O_4804,N_40063,N_43368);
and UO_4805 (O_4805,N_44513,N_42328);
and UO_4806 (O_4806,N_40225,N_43511);
or UO_4807 (O_4807,N_45686,N_41746);
or UO_4808 (O_4808,N_42705,N_47575);
or UO_4809 (O_4809,N_45498,N_42329);
nor UO_4810 (O_4810,N_49671,N_45451);
nand UO_4811 (O_4811,N_46670,N_47452);
or UO_4812 (O_4812,N_49479,N_45075);
nor UO_4813 (O_4813,N_49635,N_49067);
or UO_4814 (O_4814,N_45234,N_40695);
nand UO_4815 (O_4815,N_46886,N_48207);
nor UO_4816 (O_4816,N_43856,N_45777);
nand UO_4817 (O_4817,N_41558,N_48591);
nand UO_4818 (O_4818,N_42544,N_48798);
nor UO_4819 (O_4819,N_41597,N_48839);
and UO_4820 (O_4820,N_46004,N_45655);
or UO_4821 (O_4821,N_43958,N_47396);
nor UO_4822 (O_4822,N_46149,N_42755);
nor UO_4823 (O_4823,N_47193,N_47010);
nand UO_4824 (O_4824,N_48181,N_40440);
xor UO_4825 (O_4825,N_41599,N_45143);
nor UO_4826 (O_4826,N_49887,N_49845);
and UO_4827 (O_4827,N_46906,N_45336);
or UO_4828 (O_4828,N_46321,N_44111);
and UO_4829 (O_4829,N_42285,N_44448);
and UO_4830 (O_4830,N_42556,N_40606);
and UO_4831 (O_4831,N_40992,N_40281);
and UO_4832 (O_4832,N_47410,N_42199);
or UO_4833 (O_4833,N_45547,N_41913);
nand UO_4834 (O_4834,N_41480,N_46469);
or UO_4835 (O_4835,N_45760,N_47904);
nor UO_4836 (O_4836,N_44693,N_49502);
and UO_4837 (O_4837,N_42872,N_43308);
nor UO_4838 (O_4838,N_40941,N_49263);
nand UO_4839 (O_4839,N_48866,N_42267);
or UO_4840 (O_4840,N_40311,N_45594);
and UO_4841 (O_4841,N_43415,N_46939);
or UO_4842 (O_4842,N_49895,N_42515);
or UO_4843 (O_4843,N_48096,N_48230);
or UO_4844 (O_4844,N_44596,N_49320);
or UO_4845 (O_4845,N_48414,N_44846);
or UO_4846 (O_4846,N_47367,N_49818);
nor UO_4847 (O_4847,N_41466,N_43550);
nor UO_4848 (O_4848,N_42797,N_43772);
nor UO_4849 (O_4849,N_42657,N_47674);
and UO_4850 (O_4850,N_47273,N_49882);
nand UO_4851 (O_4851,N_46871,N_47651);
or UO_4852 (O_4852,N_45768,N_47697);
and UO_4853 (O_4853,N_45314,N_40996);
nand UO_4854 (O_4854,N_47424,N_43682);
nor UO_4855 (O_4855,N_41487,N_40919);
or UO_4856 (O_4856,N_42535,N_41447);
nor UO_4857 (O_4857,N_46537,N_45329);
nor UO_4858 (O_4858,N_49773,N_47092);
nor UO_4859 (O_4859,N_41117,N_49312);
nor UO_4860 (O_4860,N_40729,N_49751);
nand UO_4861 (O_4861,N_41693,N_44297);
xor UO_4862 (O_4862,N_49862,N_41449);
nor UO_4863 (O_4863,N_47162,N_40164);
and UO_4864 (O_4864,N_41098,N_40077);
nand UO_4865 (O_4865,N_41202,N_49097);
xnor UO_4866 (O_4866,N_44237,N_43155);
xor UO_4867 (O_4867,N_44649,N_45385);
nand UO_4868 (O_4868,N_48838,N_47125);
xnor UO_4869 (O_4869,N_40154,N_40119);
or UO_4870 (O_4870,N_46226,N_46813);
and UO_4871 (O_4871,N_45959,N_42375);
nor UO_4872 (O_4872,N_40742,N_46665);
nand UO_4873 (O_4873,N_40033,N_44634);
and UO_4874 (O_4874,N_46549,N_44086);
or UO_4875 (O_4875,N_44664,N_41898);
and UO_4876 (O_4876,N_49209,N_49600);
xor UO_4877 (O_4877,N_49050,N_47707);
nand UO_4878 (O_4878,N_45548,N_44475);
xnor UO_4879 (O_4879,N_41976,N_43023);
nor UO_4880 (O_4880,N_40861,N_41269);
nor UO_4881 (O_4881,N_40414,N_44655);
or UO_4882 (O_4882,N_48025,N_40101);
nand UO_4883 (O_4883,N_45698,N_46255);
or UO_4884 (O_4884,N_47587,N_43836);
or UO_4885 (O_4885,N_44978,N_44803);
nor UO_4886 (O_4886,N_49432,N_45506);
or UO_4887 (O_4887,N_44555,N_48041);
nand UO_4888 (O_4888,N_47294,N_40412);
and UO_4889 (O_4889,N_41753,N_46120);
or UO_4890 (O_4890,N_42242,N_46723);
nand UO_4891 (O_4891,N_41318,N_49837);
and UO_4892 (O_4892,N_43968,N_48766);
or UO_4893 (O_4893,N_44759,N_42105);
nand UO_4894 (O_4894,N_43373,N_47519);
nor UO_4895 (O_4895,N_44763,N_42622);
and UO_4896 (O_4896,N_49425,N_44358);
xor UO_4897 (O_4897,N_44540,N_49618);
nand UO_4898 (O_4898,N_40345,N_41292);
and UO_4899 (O_4899,N_48016,N_47402);
or UO_4900 (O_4900,N_42296,N_45062);
xor UO_4901 (O_4901,N_41333,N_40571);
nand UO_4902 (O_4902,N_44266,N_48917);
or UO_4903 (O_4903,N_48292,N_49652);
nor UO_4904 (O_4904,N_47318,N_41421);
xnor UO_4905 (O_4905,N_43235,N_44525);
nor UO_4906 (O_4906,N_45705,N_45373);
or UO_4907 (O_4907,N_43660,N_46559);
nor UO_4908 (O_4908,N_47325,N_41731);
nand UO_4909 (O_4909,N_42620,N_45966);
or UO_4910 (O_4910,N_42503,N_40298);
nand UO_4911 (O_4911,N_45094,N_48471);
or UO_4912 (O_4912,N_42573,N_42703);
nor UO_4913 (O_4913,N_44547,N_43883);
nand UO_4914 (O_4914,N_49940,N_45489);
nand UO_4915 (O_4915,N_45572,N_47178);
nand UO_4916 (O_4916,N_43297,N_44020);
nand UO_4917 (O_4917,N_46260,N_46967);
nand UO_4918 (O_4918,N_43642,N_47149);
nand UO_4919 (O_4919,N_40591,N_44048);
nand UO_4920 (O_4920,N_44282,N_40679);
xor UO_4921 (O_4921,N_41419,N_43973);
xnor UO_4922 (O_4922,N_49122,N_40252);
nor UO_4923 (O_4923,N_40036,N_46360);
or UO_4924 (O_4924,N_46888,N_46470);
xor UO_4925 (O_4925,N_48364,N_47095);
and UO_4926 (O_4926,N_41226,N_49812);
or UO_4927 (O_4927,N_47970,N_49535);
xor UO_4928 (O_4928,N_43727,N_40947);
or UO_4929 (O_4929,N_49036,N_45002);
and UO_4930 (O_4930,N_48272,N_48980);
nor UO_4931 (O_4931,N_49046,N_49366);
or UO_4932 (O_4932,N_48608,N_43850);
nand UO_4933 (O_4933,N_45405,N_40460);
nor UO_4934 (O_4934,N_42796,N_49964);
nor UO_4935 (O_4935,N_45207,N_41376);
nor UO_4936 (O_4936,N_42354,N_46577);
or UO_4937 (O_4937,N_48148,N_43860);
xnor UO_4938 (O_4938,N_48669,N_40818);
nor UO_4939 (O_4939,N_46215,N_44725);
nand UO_4940 (O_4940,N_46037,N_43914);
or UO_4941 (O_4941,N_49634,N_49701);
or UO_4942 (O_4942,N_47239,N_43732);
nor UO_4943 (O_4943,N_44835,N_41355);
and UO_4944 (O_4944,N_42371,N_48648);
nor UO_4945 (O_4945,N_42000,N_44469);
xor UO_4946 (O_4946,N_42232,N_49927);
nand UO_4947 (O_4947,N_49452,N_49997);
and UO_4948 (O_4948,N_44069,N_42727);
and UO_4949 (O_4949,N_47075,N_49549);
or UO_4950 (O_4950,N_42528,N_44509);
nand UO_4951 (O_4951,N_46196,N_49159);
and UO_4952 (O_4952,N_49264,N_46130);
nor UO_4953 (O_4953,N_41451,N_46704);
nor UO_4954 (O_4954,N_43254,N_47843);
nor UO_4955 (O_4955,N_45570,N_41417);
nor UO_4956 (O_4956,N_48302,N_44497);
nor UO_4957 (O_4957,N_49102,N_46737);
nor UO_4958 (O_4958,N_45316,N_49892);
nor UO_4959 (O_4959,N_47870,N_45208);
or UO_4960 (O_4960,N_45794,N_48242);
nand UO_4961 (O_4961,N_49676,N_46110);
and UO_4962 (O_4962,N_46608,N_49012);
or UO_4963 (O_4963,N_48641,N_42374);
or UO_4964 (O_4964,N_45722,N_47518);
and UO_4965 (O_4965,N_47369,N_40441);
and UO_4966 (O_4966,N_47552,N_45046);
and UO_4967 (O_4967,N_48848,N_46760);
or UO_4968 (O_4968,N_47571,N_49321);
or UO_4969 (O_4969,N_46247,N_48155);
nor UO_4970 (O_4970,N_45340,N_42822);
and UO_4971 (O_4971,N_46872,N_44058);
and UO_4972 (O_4972,N_42893,N_47893);
or UO_4973 (O_4973,N_41522,N_48701);
nor UO_4974 (O_4974,N_45980,N_47932);
or UO_4975 (O_4975,N_40032,N_42899);
and UO_4976 (O_4976,N_49418,N_49481);
nand UO_4977 (O_4977,N_46800,N_43270);
xor UO_4978 (O_4978,N_48892,N_45334);
nor UO_4979 (O_4979,N_49191,N_46859);
or UO_4980 (O_4980,N_49712,N_42877);
nor UO_4981 (O_4981,N_47023,N_40848);
or UO_4982 (O_4982,N_42111,N_45931);
nand UO_4983 (O_4983,N_41077,N_40756);
or UO_4984 (O_4984,N_49124,N_48257);
nand UO_4985 (O_4985,N_44295,N_49596);
nor UO_4986 (O_4986,N_47513,N_48262);
and UO_4987 (O_4987,N_49995,N_46207);
or UO_4988 (O_4988,N_45692,N_40461);
or UO_4989 (O_4989,N_45088,N_42671);
nor UO_4990 (O_4990,N_40613,N_46402);
nand UO_4991 (O_4991,N_40188,N_44949);
or UO_4992 (O_4992,N_47416,N_43880);
nor UO_4993 (O_4993,N_44958,N_40954);
or UO_4994 (O_4994,N_48845,N_46652);
and UO_4995 (O_4995,N_45063,N_49407);
or UO_4996 (O_4996,N_42948,N_46885);
nor UO_4997 (O_4997,N_43452,N_49921);
nand UO_4998 (O_4998,N_46941,N_49609);
or UO_4999 (O_4999,N_47332,N_47657);
endmodule