module basic_1000_10000_1500_10_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_163,In_899);
nor U1 (N_1,In_945,In_278);
or U2 (N_2,In_702,In_492);
or U3 (N_3,In_108,In_437);
xor U4 (N_4,In_963,In_58);
nand U5 (N_5,In_410,In_799);
and U6 (N_6,In_472,In_753);
and U7 (N_7,In_33,In_478);
nand U8 (N_8,In_442,In_955);
xor U9 (N_9,In_719,In_351);
and U10 (N_10,In_981,In_110);
and U11 (N_11,In_463,In_75);
or U12 (N_12,In_560,In_857);
nand U13 (N_13,In_996,In_666);
xnor U14 (N_14,In_407,In_859);
and U15 (N_15,In_867,In_23);
or U16 (N_16,In_215,In_700);
xnor U17 (N_17,In_992,In_723);
nand U18 (N_18,In_482,In_658);
nand U19 (N_19,In_161,In_412);
or U20 (N_20,In_481,In_291);
nor U21 (N_21,In_571,In_748);
xnor U22 (N_22,In_872,In_132);
nand U23 (N_23,In_912,In_611);
and U24 (N_24,In_404,In_352);
nand U25 (N_25,In_375,In_852);
xor U26 (N_26,In_251,In_489);
nand U27 (N_27,In_928,In_145);
or U28 (N_28,In_320,In_592);
nor U29 (N_29,In_676,In_526);
or U30 (N_30,In_988,In_897);
and U31 (N_31,In_121,In_72);
nand U32 (N_32,In_956,In_757);
nor U33 (N_33,In_847,In_711);
or U34 (N_34,In_669,In_494);
xnor U35 (N_35,In_67,In_538);
xor U36 (N_36,In_16,In_573);
or U37 (N_37,In_281,In_331);
and U38 (N_38,In_306,In_721);
and U39 (N_39,In_200,In_791);
nor U40 (N_40,In_754,In_623);
or U41 (N_41,In_158,In_539);
nand U42 (N_42,In_429,In_732);
and U43 (N_43,In_810,In_172);
nand U44 (N_44,In_54,In_191);
nand U45 (N_45,In_22,In_706);
nor U46 (N_46,In_850,In_443);
nor U47 (N_47,In_973,In_903);
nor U48 (N_48,In_220,In_357);
and U49 (N_49,In_905,In_186);
nand U50 (N_50,In_814,In_484);
nand U51 (N_51,In_940,In_391);
or U52 (N_52,In_42,In_683);
xor U53 (N_53,In_679,In_486);
nor U54 (N_54,In_885,In_752);
or U55 (N_55,In_376,In_873);
or U56 (N_56,In_646,In_902);
and U57 (N_57,In_11,In_977);
xnor U58 (N_58,In_267,In_212);
or U59 (N_59,In_262,In_659);
and U60 (N_60,In_136,In_383);
or U61 (N_61,In_672,In_587);
nor U62 (N_62,In_246,In_173);
nand U63 (N_63,In_74,In_235);
nor U64 (N_64,In_257,In_910);
or U65 (N_65,In_835,In_73);
and U66 (N_66,In_284,In_275);
and U67 (N_67,In_598,In_112);
and U68 (N_68,In_451,In_690);
xor U69 (N_69,In_50,In_896);
nand U70 (N_70,In_809,In_709);
nor U71 (N_71,In_315,In_848);
and U72 (N_72,In_400,In_89);
and U73 (N_73,In_332,In_990);
nand U74 (N_74,In_579,In_796);
nor U75 (N_75,In_764,In_185);
and U76 (N_76,In_188,In_553);
or U77 (N_77,In_156,In_368);
nand U78 (N_78,In_530,In_864);
nor U79 (N_79,In_552,In_529);
xor U80 (N_80,In_44,In_199);
xnor U81 (N_81,In_877,In_787);
xor U82 (N_82,In_182,In_290);
and U83 (N_83,In_607,In_783);
or U84 (N_84,In_584,In_310);
nor U85 (N_85,In_625,In_164);
nor U86 (N_86,In_248,In_935);
nand U87 (N_87,In_642,In_414);
nor U88 (N_88,In_534,In_915);
or U89 (N_89,In_171,In_862);
nor U90 (N_90,In_344,In_562);
nor U91 (N_91,In_69,In_405);
xor U92 (N_92,In_399,In_986);
or U93 (N_93,In_435,In_942);
or U94 (N_94,In_464,In_581);
xnor U95 (N_95,In_675,In_204);
and U96 (N_96,In_631,In_293);
or U97 (N_97,In_323,In_4);
and U98 (N_98,In_545,In_947);
xor U99 (N_99,In_403,In_37);
nand U100 (N_100,In_227,In_677);
or U101 (N_101,In_636,In_575);
and U102 (N_102,In_6,In_203);
nand U103 (N_103,In_969,In_496);
nand U104 (N_104,In_205,In_28);
or U105 (N_105,In_697,In_760);
xnor U106 (N_106,In_510,In_167);
nand U107 (N_107,In_301,In_934);
and U108 (N_108,In_370,In_548);
and U109 (N_109,In_56,In_430);
nand U110 (N_110,In_390,In_479);
nor U111 (N_111,In_184,In_718);
or U112 (N_112,In_866,In_427);
and U113 (N_113,In_296,In_682);
nor U114 (N_114,In_604,In_244);
or U115 (N_115,In_381,In_766);
and U116 (N_116,In_725,In_855);
xor U117 (N_117,In_114,In_468);
and U118 (N_118,In_314,In_355);
and U119 (N_119,In_453,In_819);
or U120 (N_120,In_507,In_389);
and U121 (N_121,In_216,In_989);
or U122 (N_122,In_837,In_392);
nor U123 (N_123,In_289,In_789);
nor U124 (N_124,In_459,In_868);
nor U125 (N_125,In_603,In_888);
and U126 (N_126,In_727,In_749);
or U127 (N_127,In_117,In_738);
or U128 (N_128,In_999,In_506);
nor U129 (N_129,In_187,In_544);
nor U130 (N_130,In_909,In_843);
nor U131 (N_131,In_350,In_214);
nor U132 (N_132,In_580,In_151);
nor U133 (N_133,In_273,In_739);
nor U134 (N_134,In_124,In_378);
nor U135 (N_135,In_66,In_129);
or U136 (N_136,In_113,In_209);
nand U137 (N_137,In_870,In_433);
nor U138 (N_138,In_193,In_586);
and U139 (N_139,In_798,In_266);
and U140 (N_140,In_360,In_882);
nor U141 (N_141,In_432,In_970);
or U142 (N_142,In_475,In_190);
nand U143 (N_143,In_851,In_569);
nor U144 (N_144,In_624,In_19);
or U145 (N_145,In_7,In_0);
nand U146 (N_146,In_629,In_364);
xor U147 (N_147,In_250,In_338);
nor U148 (N_148,In_68,In_865);
nor U149 (N_149,In_728,In_619);
and U150 (N_150,In_635,In_150);
nor U151 (N_151,In_588,In_313);
nor U152 (N_152,In_962,In_703);
or U153 (N_153,In_861,In_409);
and U154 (N_154,In_192,In_232);
nor U155 (N_155,In_336,In_197);
and U156 (N_156,In_794,In_35);
nor U157 (N_157,In_265,In_20);
or U158 (N_158,In_576,In_680);
and U159 (N_159,In_373,In_450);
and U160 (N_160,In_369,In_933);
and U161 (N_161,In_564,In_651);
nand U162 (N_162,In_133,In_308);
nand U163 (N_163,In_974,In_39);
or U164 (N_164,In_931,In_456);
and U165 (N_165,In_547,In_751);
nand U166 (N_166,In_226,In_599);
and U167 (N_167,In_64,In_480);
xor U168 (N_168,In_518,In_239);
and U169 (N_169,In_511,In_218);
and U170 (N_170,In_347,In_29);
nand U171 (N_171,In_162,In_477);
and U172 (N_172,In_609,In_12);
or U173 (N_173,In_627,In_950);
and U174 (N_174,In_128,In_965);
nand U175 (N_175,In_516,In_330);
or U176 (N_176,In_665,In_833);
and U177 (N_177,In_813,In_528);
xnor U178 (N_178,In_997,In_233);
nor U179 (N_179,In_946,In_640);
and U180 (N_180,In_123,In_966);
nor U181 (N_181,In_803,In_844);
and U182 (N_182,In_998,In_527);
or U183 (N_183,In_297,In_109);
nor U184 (N_184,In_107,In_729);
xor U185 (N_185,In_127,In_43);
or U186 (N_186,In_470,In_842);
nand U187 (N_187,In_555,In_52);
nor U188 (N_188,In_660,In_979);
xor U189 (N_189,In_202,In_380);
xnor U190 (N_190,In_856,In_53);
nor U191 (N_191,In_303,In_637);
nor U192 (N_192,In_175,In_15);
and U193 (N_193,In_149,In_206);
and U194 (N_194,In_148,In_82);
nor U195 (N_195,In_140,In_438);
xor U196 (N_196,In_964,In_696);
nand U197 (N_197,In_322,In_225);
and U198 (N_198,In_119,In_142);
and U199 (N_199,In_169,In_889);
and U200 (N_200,In_230,In_643);
nand U201 (N_201,In_921,In_525);
xor U202 (N_202,In_532,In_595);
and U203 (N_203,In_439,In_522);
nand U204 (N_204,In_854,In_906);
or U205 (N_205,In_601,In_255);
nor U206 (N_206,In_740,In_812);
or U207 (N_207,In_670,In_499);
xnor U208 (N_208,In_210,In_566);
nor U209 (N_209,In_231,In_756);
and U210 (N_210,In_632,In_420);
nand U211 (N_211,In_245,In_334);
nand U212 (N_212,In_79,In_504);
nand U213 (N_213,In_773,In_978);
or U214 (N_214,In_356,In_514);
nor U215 (N_215,In_36,In_201);
or U216 (N_216,In_495,In_448);
and U217 (N_217,In_734,In_243);
nor U218 (N_218,In_177,In_820);
and U219 (N_219,In_473,In_772);
nor U220 (N_220,In_421,In_176);
nand U221 (N_221,In_874,In_881);
and U222 (N_222,In_104,In_40);
nor U223 (N_223,In_893,In_980);
or U224 (N_224,In_372,In_605);
and U225 (N_225,In_827,In_274);
and U226 (N_226,In_616,In_384);
or U227 (N_227,In_917,In_490);
nor U228 (N_228,In_497,In_45);
or U229 (N_229,In_491,In_523);
and U230 (N_230,In_223,In_304);
xor U231 (N_231,In_594,In_704);
xor U232 (N_232,In_25,In_673);
xnor U233 (N_233,In_508,In_860);
or U234 (N_234,In_247,In_471);
and U235 (N_235,In_120,In_606);
or U236 (N_236,In_259,In_620);
nor U237 (N_237,In_792,In_345);
nand U238 (N_238,In_103,In_319);
and U239 (N_239,In_335,In_716);
nor U240 (N_240,In_249,In_654);
or U241 (N_241,In_118,In_900);
nand U242 (N_242,In_180,In_805);
and U243 (N_243,In_241,In_894);
nand U244 (N_244,In_519,In_326);
nand U245 (N_245,In_645,In_396);
and U246 (N_246,In_687,In_712);
xnor U247 (N_247,In_24,In_691);
nand U248 (N_248,In_277,In_260);
nand U249 (N_249,In_467,In_808);
xnor U250 (N_250,In_48,In_457);
and U251 (N_251,In_288,In_353);
and U252 (N_252,In_558,In_1);
and U253 (N_253,In_134,In_823);
or U254 (N_254,In_811,In_630);
nand U255 (N_255,In_318,In_512);
or U256 (N_256,In_328,In_87);
nor U257 (N_257,In_655,In_836);
and U258 (N_258,In_939,In_890);
xnor U259 (N_259,In_570,In_689);
xnor U260 (N_260,In_994,In_612);
nor U261 (N_261,In_454,In_165);
or U262 (N_262,In_685,In_641);
nor U263 (N_263,In_661,In_726);
nand U264 (N_264,In_287,In_818);
nor U265 (N_265,In_130,In_366);
nor U266 (N_266,In_500,In_261);
and U267 (N_267,In_47,In_198);
xnor U268 (N_268,In_937,In_572);
or U269 (N_269,In_325,In_436);
nor U270 (N_270,In_160,In_31);
nor U271 (N_271,In_838,In_398);
nor U272 (N_272,In_583,In_228);
nor U273 (N_273,In_664,In_578);
and U274 (N_274,In_388,In_717);
or U275 (N_275,In_417,In_395);
nand U276 (N_276,In_840,In_549);
nor U277 (N_277,In_406,In_194);
nor U278 (N_278,In_735,In_268);
xnor U279 (N_279,In_83,In_920);
nor U280 (N_280,In_466,In_849);
xnor U281 (N_281,In_705,In_286);
and U282 (N_282,In_731,In_600);
or U283 (N_283,In_770,In_876);
and U284 (N_284,In_122,In_822);
and U285 (N_285,In_487,In_256);
or U286 (N_286,In_299,In_125);
and U287 (N_287,In_144,In_116);
nand U288 (N_288,In_458,In_307);
or U289 (N_289,In_621,In_189);
or U290 (N_290,In_46,In_714);
nor U291 (N_291,In_785,In_141);
or U292 (N_292,In_270,In_63);
or U293 (N_293,In_556,In_542);
nor U294 (N_294,In_741,In_730);
nand U295 (N_295,In_744,In_300);
nor U296 (N_296,In_264,In_991);
and U297 (N_297,In_419,In_745);
nand U298 (N_298,In_90,In_829);
xnor U299 (N_299,In_385,In_317);
nand U300 (N_300,In_359,In_14);
and U301 (N_301,In_348,In_217);
nand U302 (N_302,In_667,In_904);
nor U303 (N_303,In_340,In_62);
xnor U304 (N_304,In_927,In_807);
nand U305 (N_305,In_648,In_423);
nand U306 (N_306,In_957,In_901);
xnor U307 (N_307,In_449,In_111);
or U308 (N_308,In_343,In_61);
or U309 (N_309,In_138,In_804);
or U310 (N_310,In_153,In_887);
nand U311 (N_311,In_85,In_561);
nand U312 (N_312,In_688,In_768);
and U313 (N_313,In_613,In_137);
or U314 (N_314,In_115,In_183);
nor U315 (N_315,In_276,In_181);
xor U316 (N_316,In_543,In_361);
or U317 (N_317,In_80,In_771);
nand U318 (N_318,In_483,In_26);
or U319 (N_319,In_413,In_958);
nor U320 (N_320,In_147,In_354);
or U321 (N_321,In_5,In_455);
nor U322 (N_322,In_746,In_38);
and U323 (N_323,In_460,In_678);
or U324 (N_324,In_238,In_639);
nor U325 (N_325,In_221,In_663);
and U326 (N_326,In_778,In_476);
or U327 (N_327,In_96,In_242);
nor U328 (N_328,In_784,In_941);
nand U329 (N_329,In_10,In_444);
and U330 (N_330,In_918,In_57);
nand U331 (N_331,In_608,In_657);
nand U332 (N_332,In_258,In_960);
or U333 (N_333,In_196,In_84);
xnor U334 (N_334,In_763,In_788);
nor U335 (N_335,In_793,In_541);
and U336 (N_336,In_311,In_485);
nand U337 (N_337,In_563,In_49);
or U338 (N_338,In_891,In_701);
xnor U339 (N_339,In_537,In_652);
nor U340 (N_340,In_411,In_101);
xor U341 (N_341,In_628,In_815);
nor U342 (N_342,In_674,In_422);
xor U343 (N_343,In_146,In_397);
nor U344 (N_344,In_386,In_948);
nand U345 (N_345,In_961,In_327);
xnor U346 (N_346,In_428,In_825);
and U347 (N_347,In_309,In_285);
nor U348 (N_348,In_213,In_211);
nand U349 (N_349,In_377,In_758);
nand U350 (N_350,In_924,In_736);
and U351 (N_351,In_425,In_321);
nand U352 (N_352,In_790,In_70);
or U353 (N_353,In_416,In_166);
nand U354 (N_354,In_174,In_229);
nor U355 (N_355,In_30,In_95);
nand U356 (N_356,In_312,In_907);
and U357 (N_357,In_155,In_565);
or U358 (N_358,In_589,In_597);
and U359 (N_359,In_761,In_106);
nand U360 (N_360,In_94,In_86);
nand U361 (N_361,In_925,In_681);
and U362 (N_362,In_60,In_590);
xor U363 (N_363,In_767,In_853);
and U364 (N_364,In_295,In_699);
and U365 (N_365,In_708,In_898);
xnor U366 (N_366,In_349,In_932);
nor U367 (N_367,In_878,In_17);
nand U368 (N_368,In_720,In_875);
nor U369 (N_369,In_447,In_618);
or U370 (N_370,In_32,In_984);
or U371 (N_371,In_402,In_333);
or U372 (N_372,In_953,In_445);
and U373 (N_373,In_971,In_554);
nand U374 (N_374,In_170,In_294);
xor U375 (N_375,In_208,In_615);
nor U376 (N_376,In_929,In_776);
or U377 (N_377,In_236,In_952);
or U378 (N_378,In_41,In_59);
nand U379 (N_379,In_341,In_883);
and U380 (N_380,In_21,In_98);
xor U381 (N_381,In_207,In_55);
nand U382 (N_382,In_533,In_342);
and U383 (N_383,In_520,In_282);
nand U384 (N_384,In_707,In_858);
nand U385 (N_385,In_936,In_493);
and U386 (N_386,In_252,In_653);
nor U387 (N_387,In_817,In_895);
and U388 (N_388,In_78,In_759);
nand U389 (N_389,In_824,In_668);
and U390 (N_390,In_938,In_710);
nand U391 (N_391,In_18,In_684);
nand U392 (N_392,In_644,In_71);
or U393 (N_393,In_846,In_135);
or U394 (N_394,In_362,In_926);
nand U395 (N_395,In_92,In_13);
nor U396 (N_396,In_656,In_195);
or U397 (N_397,In_271,In_298);
and U398 (N_398,In_551,In_540);
nor U399 (N_399,In_509,In_949);
nor U400 (N_400,In_880,In_408);
and U401 (N_401,In_126,In_845);
and U402 (N_402,In_346,In_152);
nand U403 (N_403,In_394,In_367);
or U404 (N_404,In_585,In_724);
nor U405 (N_405,In_77,In_801);
and U406 (N_406,In_168,In_452);
nor U407 (N_407,In_610,In_503);
nand U408 (N_408,In_800,In_462);
nand U409 (N_409,In_263,In_777);
and U410 (N_410,In_821,In_374);
xnor U411 (N_411,In_944,In_99);
or U412 (N_412,In_647,In_302);
and U413 (N_413,In_831,In_976);
or U414 (N_414,In_329,In_987);
or U415 (N_415,In_983,In_401);
xor U416 (N_416,In_339,In_916);
nor U417 (N_417,In_828,In_972);
nor U418 (N_418,In_418,In_531);
xor U419 (N_419,In_982,In_634);
nand U420 (N_420,In_662,In_967);
nand U421 (N_421,In_81,In_283);
nor U422 (N_422,In_713,In_426);
nor U423 (N_423,In_686,In_816);
and U424 (N_424,In_786,In_517);
or U425 (N_425,In_365,In_97);
nor U426 (N_426,In_100,In_715);
nand U427 (N_427,In_424,In_305);
nor U428 (N_428,In_596,In_280);
nor U429 (N_429,In_649,In_105);
nor U430 (N_430,In_324,In_51);
or U431 (N_431,In_559,In_622);
and U432 (N_432,In_650,In_919);
nor U433 (N_433,In_782,In_968);
xor U434 (N_434,In_694,In_886);
or U435 (N_435,In_775,In_536);
or U436 (N_436,In_502,In_550);
and U437 (N_437,In_363,In_951);
or U438 (N_438,In_591,In_567);
or U439 (N_439,In_469,In_693);
and U440 (N_440,In_993,In_358);
nor U441 (N_441,In_671,In_3);
and U442 (N_442,In_501,In_779);
or U443 (N_443,In_157,In_780);
or U444 (N_444,In_546,In_737);
nor U445 (N_445,In_577,In_626);
xnor U446 (N_446,In_498,In_863);
nand U447 (N_447,In_441,In_513);
nor U448 (N_448,In_269,In_943);
xnor U449 (N_449,In_337,In_750);
nor U450 (N_450,In_922,In_154);
nor U451 (N_451,In_774,In_892);
nor U452 (N_452,In_521,In_869);
and U453 (N_453,In_179,In_9);
nand U454 (N_454,In_879,In_434);
xor U455 (N_455,In_830,In_292);
and U456 (N_456,In_695,In_839);
or U457 (N_457,In_393,In_914);
xnor U458 (N_458,In_568,In_841);
and U459 (N_459,In_614,In_832);
nand U460 (N_460,In_781,In_461);
nand U461 (N_461,In_692,In_985);
nand U462 (N_462,In_582,In_995);
and U463 (N_463,In_382,In_747);
or U464 (N_464,In_638,In_959);
xor U465 (N_465,In_698,In_440);
or U466 (N_466,In_743,In_765);
nand U467 (N_467,In_224,In_272);
nor U468 (N_468,In_802,In_139);
nand U469 (N_469,In_911,In_143);
nand U470 (N_470,In_387,In_234);
nand U471 (N_471,In_755,In_431);
nand U472 (N_472,In_913,In_253);
or U473 (N_473,In_733,In_593);
nand U474 (N_474,In_826,In_76);
and U475 (N_475,In_371,In_633);
or U476 (N_476,In_2,In_806);
and U477 (N_477,In_574,In_316);
nor U478 (N_478,In_159,In_954);
xor U479 (N_479,In_446,In_722);
nand U480 (N_480,In_91,In_535);
nand U481 (N_481,In_415,In_488);
or U482 (N_482,In_34,In_884);
nand U483 (N_483,In_834,In_8);
and U484 (N_484,In_465,In_908);
nor U485 (N_485,In_515,In_219);
nand U486 (N_486,In_279,In_871);
nor U487 (N_487,In_762,In_254);
nor U488 (N_488,In_524,In_93);
nand U489 (N_489,In_88,In_240);
nand U490 (N_490,In_557,In_742);
nand U491 (N_491,In_505,In_102);
nand U492 (N_492,In_795,In_65);
and U493 (N_493,In_617,In_602);
or U494 (N_494,In_975,In_379);
nand U495 (N_495,In_923,In_237);
nand U496 (N_496,In_769,In_474);
nor U497 (N_497,In_131,In_930);
and U498 (N_498,In_797,In_27);
xnor U499 (N_499,In_178,In_222);
or U500 (N_500,In_70,In_615);
and U501 (N_501,In_469,In_993);
xnor U502 (N_502,In_426,In_237);
nor U503 (N_503,In_911,In_37);
nand U504 (N_504,In_348,In_231);
nor U505 (N_505,In_88,In_131);
nand U506 (N_506,In_600,In_575);
nor U507 (N_507,In_327,In_257);
or U508 (N_508,In_930,In_901);
and U509 (N_509,In_563,In_470);
nor U510 (N_510,In_3,In_520);
and U511 (N_511,In_407,In_276);
nor U512 (N_512,In_503,In_981);
or U513 (N_513,In_874,In_801);
nand U514 (N_514,In_666,In_894);
or U515 (N_515,In_795,In_918);
and U516 (N_516,In_529,In_218);
nor U517 (N_517,In_358,In_165);
xor U518 (N_518,In_306,In_887);
or U519 (N_519,In_967,In_796);
or U520 (N_520,In_813,In_702);
nor U521 (N_521,In_416,In_207);
and U522 (N_522,In_764,In_65);
and U523 (N_523,In_460,In_201);
nor U524 (N_524,In_866,In_523);
nand U525 (N_525,In_648,In_821);
and U526 (N_526,In_690,In_797);
nand U527 (N_527,In_303,In_137);
or U528 (N_528,In_287,In_942);
nand U529 (N_529,In_365,In_330);
xnor U530 (N_530,In_41,In_609);
nor U531 (N_531,In_427,In_953);
and U532 (N_532,In_561,In_422);
and U533 (N_533,In_731,In_63);
nand U534 (N_534,In_853,In_216);
or U535 (N_535,In_679,In_439);
xnor U536 (N_536,In_527,In_98);
nand U537 (N_537,In_218,In_231);
nor U538 (N_538,In_741,In_866);
or U539 (N_539,In_685,In_337);
and U540 (N_540,In_162,In_970);
nand U541 (N_541,In_874,In_157);
and U542 (N_542,In_209,In_923);
nand U543 (N_543,In_960,In_511);
nand U544 (N_544,In_747,In_120);
xor U545 (N_545,In_74,In_641);
xor U546 (N_546,In_136,In_508);
and U547 (N_547,In_387,In_749);
xor U548 (N_548,In_913,In_327);
nand U549 (N_549,In_860,In_795);
and U550 (N_550,In_300,In_938);
and U551 (N_551,In_117,In_621);
or U552 (N_552,In_779,In_532);
or U553 (N_553,In_379,In_610);
nor U554 (N_554,In_875,In_985);
nor U555 (N_555,In_591,In_53);
nor U556 (N_556,In_103,In_961);
and U557 (N_557,In_87,In_908);
and U558 (N_558,In_833,In_691);
or U559 (N_559,In_421,In_441);
or U560 (N_560,In_106,In_813);
and U561 (N_561,In_32,In_301);
xnor U562 (N_562,In_791,In_977);
or U563 (N_563,In_146,In_101);
nand U564 (N_564,In_239,In_660);
nand U565 (N_565,In_231,In_746);
nor U566 (N_566,In_358,In_879);
and U567 (N_567,In_843,In_382);
or U568 (N_568,In_476,In_89);
and U569 (N_569,In_394,In_513);
and U570 (N_570,In_729,In_465);
nand U571 (N_571,In_239,In_991);
or U572 (N_572,In_353,In_466);
nor U573 (N_573,In_869,In_674);
or U574 (N_574,In_381,In_10);
or U575 (N_575,In_730,In_51);
or U576 (N_576,In_330,In_501);
nand U577 (N_577,In_50,In_521);
nor U578 (N_578,In_695,In_625);
nor U579 (N_579,In_986,In_506);
or U580 (N_580,In_908,In_291);
and U581 (N_581,In_628,In_936);
and U582 (N_582,In_364,In_514);
and U583 (N_583,In_849,In_278);
nand U584 (N_584,In_933,In_700);
nand U585 (N_585,In_365,In_316);
nor U586 (N_586,In_252,In_827);
nor U587 (N_587,In_202,In_96);
xor U588 (N_588,In_36,In_987);
nand U589 (N_589,In_219,In_753);
or U590 (N_590,In_794,In_448);
or U591 (N_591,In_638,In_283);
or U592 (N_592,In_843,In_652);
or U593 (N_593,In_545,In_809);
nor U594 (N_594,In_328,In_50);
xnor U595 (N_595,In_535,In_322);
or U596 (N_596,In_391,In_448);
or U597 (N_597,In_615,In_934);
nand U598 (N_598,In_883,In_808);
nand U599 (N_599,In_416,In_119);
and U600 (N_600,In_476,In_364);
and U601 (N_601,In_638,In_609);
xor U602 (N_602,In_360,In_665);
nor U603 (N_603,In_65,In_135);
xnor U604 (N_604,In_479,In_43);
and U605 (N_605,In_853,In_421);
or U606 (N_606,In_876,In_409);
xnor U607 (N_607,In_318,In_54);
or U608 (N_608,In_918,In_425);
and U609 (N_609,In_720,In_528);
or U610 (N_610,In_241,In_511);
nor U611 (N_611,In_914,In_366);
or U612 (N_612,In_854,In_142);
nor U613 (N_613,In_818,In_340);
and U614 (N_614,In_564,In_559);
nor U615 (N_615,In_426,In_503);
nand U616 (N_616,In_771,In_809);
xnor U617 (N_617,In_183,In_895);
or U618 (N_618,In_669,In_483);
xor U619 (N_619,In_658,In_531);
xor U620 (N_620,In_92,In_166);
nand U621 (N_621,In_650,In_65);
or U622 (N_622,In_290,In_507);
and U623 (N_623,In_327,In_5);
or U624 (N_624,In_503,In_187);
and U625 (N_625,In_230,In_642);
and U626 (N_626,In_176,In_110);
or U627 (N_627,In_297,In_239);
xnor U628 (N_628,In_46,In_944);
or U629 (N_629,In_71,In_196);
and U630 (N_630,In_385,In_930);
nor U631 (N_631,In_951,In_604);
xnor U632 (N_632,In_713,In_766);
nand U633 (N_633,In_643,In_5);
or U634 (N_634,In_184,In_939);
or U635 (N_635,In_259,In_661);
xnor U636 (N_636,In_787,In_823);
xnor U637 (N_637,In_695,In_171);
nor U638 (N_638,In_167,In_221);
nor U639 (N_639,In_951,In_313);
nor U640 (N_640,In_642,In_606);
xnor U641 (N_641,In_571,In_775);
and U642 (N_642,In_271,In_723);
nand U643 (N_643,In_456,In_684);
or U644 (N_644,In_300,In_155);
and U645 (N_645,In_667,In_446);
nand U646 (N_646,In_889,In_27);
nor U647 (N_647,In_734,In_410);
or U648 (N_648,In_699,In_32);
xnor U649 (N_649,In_707,In_727);
and U650 (N_650,In_496,In_797);
and U651 (N_651,In_816,In_521);
nor U652 (N_652,In_872,In_500);
or U653 (N_653,In_582,In_242);
or U654 (N_654,In_878,In_535);
or U655 (N_655,In_537,In_717);
or U656 (N_656,In_798,In_199);
or U657 (N_657,In_266,In_134);
and U658 (N_658,In_376,In_897);
nor U659 (N_659,In_244,In_739);
nor U660 (N_660,In_855,In_448);
nor U661 (N_661,In_832,In_984);
xor U662 (N_662,In_164,In_825);
or U663 (N_663,In_472,In_181);
or U664 (N_664,In_99,In_810);
or U665 (N_665,In_717,In_309);
or U666 (N_666,In_0,In_842);
nand U667 (N_667,In_193,In_534);
nor U668 (N_668,In_235,In_88);
nand U669 (N_669,In_949,In_81);
and U670 (N_670,In_217,In_561);
or U671 (N_671,In_721,In_293);
xor U672 (N_672,In_531,In_91);
or U673 (N_673,In_418,In_454);
or U674 (N_674,In_180,In_914);
xor U675 (N_675,In_978,In_785);
nor U676 (N_676,In_716,In_290);
and U677 (N_677,In_292,In_770);
nor U678 (N_678,In_578,In_642);
or U679 (N_679,In_731,In_583);
xor U680 (N_680,In_774,In_831);
or U681 (N_681,In_750,In_920);
or U682 (N_682,In_113,In_603);
or U683 (N_683,In_692,In_100);
or U684 (N_684,In_929,In_991);
and U685 (N_685,In_210,In_209);
nor U686 (N_686,In_584,In_433);
nor U687 (N_687,In_939,In_775);
or U688 (N_688,In_326,In_841);
nor U689 (N_689,In_684,In_692);
nand U690 (N_690,In_411,In_292);
xnor U691 (N_691,In_178,In_604);
and U692 (N_692,In_701,In_121);
nor U693 (N_693,In_59,In_909);
nand U694 (N_694,In_394,In_730);
and U695 (N_695,In_648,In_511);
nor U696 (N_696,In_692,In_44);
nor U697 (N_697,In_474,In_411);
nor U698 (N_698,In_631,In_940);
nor U699 (N_699,In_170,In_204);
nor U700 (N_700,In_890,In_363);
and U701 (N_701,In_900,In_973);
nor U702 (N_702,In_957,In_792);
nand U703 (N_703,In_79,In_873);
xor U704 (N_704,In_242,In_965);
or U705 (N_705,In_249,In_360);
and U706 (N_706,In_281,In_55);
or U707 (N_707,In_584,In_739);
or U708 (N_708,In_572,In_727);
nand U709 (N_709,In_382,In_673);
nor U710 (N_710,In_397,In_362);
nor U711 (N_711,In_112,In_439);
xor U712 (N_712,In_834,In_113);
nor U713 (N_713,In_24,In_670);
xor U714 (N_714,In_600,In_208);
nor U715 (N_715,In_177,In_724);
nor U716 (N_716,In_217,In_925);
nor U717 (N_717,In_558,In_432);
xor U718 (N_718,In_791,In_236);
nand U719 (N_719,In_9,In_724);
xnor U720 (N_720,In_537,In_217);
or U721 (N_721,In_965,In_756);
xnor U722 (N_722,In_779,In_484);
or U723 (N_723,In_469,In_51);
nand U724 (N_724,In_830,In_89);
xor U725 (N_725,In_767,In_314);
nor U726 (N_726,In_843,In_994);
nand U727 (N_727,In_813,In_174);
xnor U728 (N_728,In_258,In_792);
nand U729 (N_729,In_515,In_127);
nor U730 (N_730,In_22,In_747);
nand U731 (N_731,In_631,In_587);
nand U732 (N_732,In_241,In_925);
nor U733 (N_733,In_225,In_156);
or U734 (N_734,In_140,In_252);
and U735 (N_735,In_243,In_521);
or U736 (N_736,In_331,In_13);
nor U737 (N_737,In_555,In_747);
and U738 (N_738,In_662,In_356);
xnor U739 (N_739,In_864,In_184);
xnor U740 (N_740,In_624,In_262);
xnor U741 (N_741,In_68,In_332);
nor U742 (N_742,In_303,In_6);
nand U743 (N_743,In_51,In_338);
nor U744 (N_744,In_469,In_210);
and U745 (N_745,In_414,In_15);
nor U746 (N_746,In_406,In_58);
xnor U747 (N_747,In_73,In_588);
or U748 (N_748,In_424,In_942);
and U749 (N_749,In_757,In_947);
or U750 (N_750,In_121,In_101);
and U751 (N_751,In_711,In_448);
or U752 (N_752,In_798,In_365);
nand U753 (N_753,In_43,In_153);
nor U754 (N_754,In_794,In_313);
nand U755 (N_755,In_299,In_407);
nor U756 (N_756,In_632,In_255);
nand U757 (N_757,In_59,In_604);
nor U758 (N_758,In_987,In_880);
and U759 (N_759,In_807,In_770);
and U760 (N_760,In_491,In_544);
and U761 (N_761,In_259,In_281);
nand U762 (N_762,In_158,In_82);
xnor U763 (N_763,In_882,In_654);
or U764 (N_764,In_322,In_103);
and U765 (N_765,In_850,In_396);
or U766 (N_766,In_655,In_174);
nand U767 (N_767,In_66,In_636);
or U768 (N_768,In_902,In_457);
or U769 (N_769,In_580,In_5);
or U770 (N_770,In_787,In_691);
and U771 (N_771,In_208,In_227);
and U772 (N_772,In_139,In_95);
nand U773 (N_773,In_177,In_738);
nor U774 (N_774,In_150,In_894);
xnor U775 (N_775,In_267,In_766);
nor U776 (N_776,In_104,In_47);
nand U777 (N_777,In_210,In_963);
or U778 (N_778,In_176,In_86);
and U779 (N_779,In_946,In_618);
and U780 (N_780,In_632,In_975);
and U781 (N_781,In_195,In_951);
and U782 (N_782,In_365,In_210);
nor U783 (N_783,In_316,In_222);
nand U784 (N_784,In_938,In_859);
nand U785 (N_785,In_720,In_908);
nand U786 (N_786,In_417,In_939);
nor U787 (N_787,In_203,In_641);
nor U788 (N_788,In_429,In_122);
nor U789 (N_789,In_633,In_830);
and U790 (N_790,In_844,In_456);
and U791 (N_791,In_398,In_250);
or U792 (N_792,In_973,In_889);
or U793 (N_793,In_592,In_767);
nor U794 (N_794,In_513,In_515);
or U795 (N_795,In_888,In_365);
nand U796 (N_796,In_982,In_220);
xnor U797 (N_797,In_938,In_26);
nand U798 (N_798,In_418,In_321);
nand U799 (N_799,In_489,In_811);
or U800 (N_800,In_248,In_108);
xor U801 (N_801,In_772,In_721);
and U802 (N_802,In_936,In_522);
and U803 (N_803,In_107,In_222);
nor U804 (N_804,In_454,In_441);
nor U805 (N_805,In_106,In_315);
or U806 (N_806,In_869,In_695);
or U807 (N_807,In_348,In_208);
or U808 (N_808,In_671,In_983);
nand U809 (N_809,In_526,In_182);
and U810 (N_810,In_342,In_31);
nand U811 (N_811,In_3,In_685);
nand U812 (N_812,In_702,In_999);
nor U813 (N_813,In_521,In_650);
nand U814 (N_814,In_989,In_835);
or U815 (N_815,In_288,In_200);
and U816 (N_816,In_591,In_342);
nand U817 (N_817,In_757,In_419);
nor U818 (N_818,In_291,In_723);
or U819 (N_819,In_327,In_791);
and U820 (N_820,In_459,In_244);
nor U821 (N_821,In_589,In_352);
nand U822 (N_822,In_624,In_755);
or U823 (N_823,In_239,In_885);
nand U824 (N_824,In_207,In_541);
or U825 (N_825,In_762,In_751);
and U826 (N_826,In_199,In_252);
nor U827 (N_827,In_324,In_18);
and U828 (N_828,In_851,In_37);
or U829 (N_829,In_303,In_195);
and U830 (N_830,In_455,In_193);
xor U831 (N_831,In_904,In_150);
xor U832 (N_832,In_983,In_397);
nor U833 (N_833,In_861,In_459);
and U834 (N_834,In_586,In_257);
and U835 (N_835,In_93,In_75);
or U836 (N_836,In_203,In_968);
and U837 (N_837,In_125,In_16);
and U838 (N_838,In_833,In_607);
and U839 (N_839,In_98,In_314);
nor U840 (N_840,In_715,In_916);
nand U841 (N_841,In_802,In_263);
nor U842 (N_842,In_996,In_852);
or U843 (N_843,In_387,In_373);
nor U844 (N_844,In_476,In_973);
and U845 (N_845,In_156,In_934);
and U846 (N_846,In_900,In_51);
nor U847 (N_847,In_136,In_374);
xnor U848 (N_848,In_231,In_623);
nor U849 (N_849,In_947,In_446);
nor U850 (N_850,In_880,In_54);
or U851 (N_851,In_279,In_351);
nand U852 (N_852,In_330,In_31);
xnor U853 (N_853,In_769,In_402);
nor U854 (N_854,In_135,In_574);
and U855 (N_855,In_914,In_775);
nand U856 (N_856,In_703,In_56);
nor U857 (N_857,In_482,In_560);
and U858 (N_858,In_159,In_851);
and U859 (N_859,In_954,In_998);
nand U860 (N_860,In_849,In_597);
xnor U861 (N_861,In_668,In_701);
nand U862 (N_862,In_894,In_40);
and U863 (N_863,In_431,In_530);
or U864 (N_864,In_768,In_568);
nand U865 (N_865,In_954,In_167);
or U866 (N_866,In_115,In_338);
nand U867 (N_867,In_913,In_627);
and U868 (N_868,In_632,In_497);
nand U869 (N_869,In_129,In_730);
nand U870 (N_870,In_205,In_814);
nand U871 (N_871,In_204,In_196);
or U872 (N_872,In_369,In_522);
and U873 (N_873,In_81,In_516);
or U874 (N_874,In_796,In_368);
and U875 (N_875,In_230,In_1);
nor U876 (N_876,In_564,In_237);
and U877 (N_877,In_730,In_582);
nand U878 (N_878,In_753,In_397);
xnor U879 (N_879,In_634,In_599);
nand U880 (N_880,In_192,In_48);
or U881 (N_881,In_691,In_151);
nor U882 (N_882,In_869,In_575);
xor U883 (N_883,In_325,In_45);
nand U884 (N_884,In_471,In_229);
and U885 (N_885,In_315,In_127);
and U886 (N_886,In_981,In_784);
or U887 (N_887,In_704,In_223);
nor U888 (N_888,In_64,In_714);
or U889 (N_889,In_969,In_101);
nand U890 (N_890,In_939,In_176);
and U891 (N_891,In_985,In_974);
or U892 (N_892,In_81,In_464);
nor U893 (N_893,In_95,In_613);
and U894 (N_894,In_129,In_127);
or U895 (N_895,In_161,In_990);
and U896 (N_896,In_185,In_431);
nor U897 (N_897,In_431,In_322);
xnor U898 (N_898,In_596,In_405);
nand U899 (N_899,In_486,In_234);
nor U900 (N_900,In_473,In_146);
nand U901 (N_901,In_41,In_10);
nand U902 (N_902,In_576,In_741);
nor U903 (N_903,In_216,In_846);
nand U904 (N_904,In_710,In_430);
and U905 (N_905,In_380,In_458);
or U906 (N_906,In_608,In_394);
or U907 (N_907,In_899,In_908);
or U908 (N_908,In_869,In_707);
and U909 (N_909,In_206,In_167);
and U910 (N_910,In_565,In_700);
nor U911 (N_911,In_346,In_272);
and U912 (N_912,In_344,In_149);
nand U913 (N_913,In_929,In_327);
nor U914 (N_914,In_162,In_325);
and U915 (N_915,In_896,In_806);
or U916 (N_916,In_92,In_658);
nor U917 (N_917,In_164,In_808);
nand U918 (N_918,In_964,In_642);
nand U919 (N_919,In_531,In_773);
nand U920 (N_920,In_15,In_848);
nand U921 (N_921,In_505,In_332);
and U922 (N_922,In_449,In_31);
xnor U923 (N_923,In_166,In_927);
or U924 (N_924,In_255,In_678);
and U925 (N_925,In_664,In_840);
and U926 (N_926,In_555,In_74);
and U927 (N_927,In_27,In_573);
nor U928 (N_928,In_763,In_547);
nor U929 (N_929,In_524,In_614);
nor U930 (N_930,In_731,In_103);
and U931 (N_931,In_606,In_841);
nor U932 (N_932,In_760,In_951);
nand U933 (N_933,In_615,In_817);
xnor U934 (N_934,In_130,In_196);
xor U935 (N_935,In_133,In_362);
or U936 (N_936,In_246,In_826);
or U937 (N_937,In_490,In_677);
and U938 (N_938,In_112,In_714);
nand U939 (N_939,In_122,In_82);
or U940 (N_940,In_225,In_104);
nand U941 (N_941,In_776,In_817);
and U942 (N_942,In_609,In_713);
and U943 (N_943,In_889,In_284);
nor U944 (N_944,In_236,In_811);
or U945 (N_945,In_868,In_179);
and U946 (N_946,In_303,In_840);
and U947 (N_947,In_851,In_545);
nor U948 (N_948,In_822,In_29);
or U949 (N_949,In_865,In_277);
or U950 (N_950,In_808,In_17);
or U951 (N_951,In_593,In_332);
and U952 (N_952,In_315,In_323);
nor U953 (N_953,In_748,In_143);
nand U954 (N_954,In_35,In_271);
xnor U955 (N_955,In_828,In_337);
nor U956 (N_956,In_847,In_301);
nor U957 (N_957,In_894,In_235);
nor U958 (N_958,In_836,In_215);
nor U959 (N_959,In_13,In_810);
and U960 (N_960,In_415,In_726);
nor U961 (N_961,In_782,In_361);
nand U962 (N_962,In_564,In_265);
and U963 (N_963,In_615,In_110);
nand U964 (N_964,In_149,In_873);
nand U965 (N_965,In_636,In_301);
and U966 (N_966,In_651,In_877);
or U967 (N_967,In_202,In_801);
or U968 (N_968,In_717,In_225);
nand U969 (N_969,In_387,In_49);
or U970 (N_970,In_148,In_585);
and U971 (N_971,In_373,In_19);
and U972 (N_972,In_784,In_897);
and U973 (N_973,In_213,In_106);
nand U974 (N_974,In_192,In_768);
and U975 (N_975,In_940,In_406);
nor U976 (N_976,In_877,In_236);
nor U977 (N_977,In_485,In_513);
or U978 (N_978,In_12,In_606);
nor U979 (N_979,In_966,In_572);
xnor U980 (N_980,In_660,In_751);
nor U981 (N_981,In_419,In_714);
or U982 (N_982,In_537,In_374);
and U983 (N_983,In_685,In_918);
nor U984 (N_984,In_722,In_885);
or U985 (N_985,In_656,In_885);
nand U986 (N_986,In_608,In_23);
xor U987 (N_987,In_216,In_968);
and U988 (N_988,In_927,In_66);
nor U989 (N_989,In_725,In_907);
and U990 (N_990,In_787,In_125);
nand U991 (N_991,In_4,In_888);
xnor U992 (N_992,In_496,In_273);
and U993 (N_993,In_628,In_849);
and U994 (N_994,In_938,In_274);
nor U995 (N_995,In_672,In_451);
or U996 (N_996,In_774,In_512);
or U997 (N_997,In_357,In_572);
and U998 (N_998,In_796,In_224);
nor U999 (N_999,In_655,In_696);
nor U1000 (N_1000,N_299,N_503);
and U1001 (N_1001,N_649,N_209);
nor U1002 (N_1002,N_787,N_386);
and U1003 (N_1003,N_981,N_32);
nor U1004 (N_1004,N_656,N_492);
nor U1005 (N_1005,N_817,N_126);
or U1006 (N_1006,N_17,N_947);
nand U1007 (N_1007,N_292,N_364);
and U1008 (N_1008,N_185,N_362);
or U1009 (N_1009,N_844,N_142);
xnor U1010 (N_1010,N_574,N_406);
nand U1011 (N_1011,N_339,N_360);
nor U1012 (N_1012,N_198,N_448);
nand U1013 (N_1013,N_805,N_419);
nand U1014 (N_1014,N_978,N_83);
and U1015 (N_1015,N_992,N_745);
or U1016 (N_1016,N_834,N_720);
or U1017 (N_1017,N_679,N_626);
nand U1018 (N_1018,N_59,N_527);
nand U1019 (N_1019,N_277,N_550);
or U1020 (N_1020,N_107,N_622);
nor U1021 (N_1021,N_862,N_639);
nand U1022 (N_1022,N_483,N_251);
or U1023 (N_1023,N_352,N_506);
nand U1024 (N_1024,N_623,N_691);
xnor U1025 (N_1025,N_463,N_554);
and U1026 (N_1026,N_263,N_405);
and U1027 (N_1027,N_994,N_797);
nor U1028 (N_1028,N_301,N_984);
nor U1029 (N_1029,N_243,N_157);
or U1030 (N_1030,N_792,N_865);
nand U1031 (N_1031,N_616,N_786);
and U1032 (N_1032,N_849,N_693);
xor U1033 (N_1033,N_82,N_872);
or U1034 (N_1034,N_516,N_235);
nand U1035 (N_1035,N_831,N_612);
and U1036 (N_1036,N_400,N_72);
nor U1037 (N_1037,N_784,N_373);
or U1038 (N_1038,N_174,N_827);
xnor U1039 (N_1039,N_881,N_426);
or U1040 (N_1040,N_972,N_968);
or U1041 (N_1041,N_13,N_206);
or U1042 (N_1042,N_23,N_504);
or U1043 (N_1043,N_782,N_214);
and U1044 (N_1044,N_930,N_764);
xnor U1045 (N_1045,N_919,N_906);
nand U1046 (N_1046,N_618,N_788);
or U1047 (N_1047,N_848,N_159);
nand U1048 (N_1048,N_27,N_594);
nor U1049 (N_1049,N_886,N_954);
xnor U1050 (N_1050,N_98,N_599);
xnor U1051 (N_1051,N_517,N_60);
nand U1052 (N_1052,N_401,N_888);
nand U1053 (N_1053,N_293,N_4);
nand U1054 (N_1054,N_986,N_800);
nand U1055 (N_1055,N_20,N_697);
nor U1056 (N_1056,N_948,N_634);
nor U1057 (N_1057,N_790,N_999);
nand U1058 (N_1058,N_897,N_49);
xnor U1059 (N_1059,N_450,N_26);
and U1060 (N_1060,N_348,N_140);
nor U1061 (N_1061,N_253,N_873);
or U1062 (N_1062,N_603,N_260);
or U1063 (N_1063,N_573,N_188);
nand U1064 (N_1064,N_974,N_507);
or U1065 (N_1065,N_257,N_808);
or U1066 (N_1066,N_590,N_536);
nand U1067 (N_1067,N_624,N_628);
nor U1068 (N_1068,N_902,N_957);
or U1069 (N_1069,N_338,N_486);
or U1070 (N_1070,N_543,N_208);
or U1071 (N_1071,N_581,N_767);
xor U1072 (N_1072,N_71,N_215);
or U1073 (N_1073,N_712,N_130);
or U1074 (N_1074,N_168,N_997);
nor U1075 (N_1075,N_588,N_990);
and U1076 (N_1076,N_964,N_548);
or U1077 (N_1077,N_751,N_278);
xnor U1078 (N_1078,N_180,N_891);
and U1079 (N_1079,N_920,N_171);
nand U1080 (N_1080,N_773,N_217);
nor U1081 (N_1081,N_681,N_452);
xor U1082 (N_1082,N_914,N_696);
or U1083 (N_1083,N_949,N_525);
or U1084 (N_1084,N_498,N_789);
and U1085 (N_1085,N_714,N_116);
xor U1086 (N_1086,N_2,N_899);
nand U1087 (N_1087,N_99,N_495);
nor U1088 (N_1088,N_207,N_88);
and U1089 (N_1089,N_763,N_982);
xnor U1090 (N_1090,N_381,N_416);
nor U1091 (N_1091,N_65,N_979);
or U1092 (N_1092,N_371,N_935);
and U1093 (N_1093,N_708,N_93);
and U1094 (N_1094,N_520,N_380);
or U1095 (N_1095,N_79,N_295);
or U1096 (N_1096,N_660,N_843);
nand U1097 (N_1097,N_212,N_0);
nor U1098 (N_1098,N_155,N_201);
or U1099 (N_1099,N_250,N_723);
nor U1100 (N_1100,N_48,N_756);
and U1101 (N_1101,N_801,N_666);
nand U1102 (N_1102,N_804,N_650);
or U1103 (N_1103,N_923,N_10);
nor U1104 (N_1104,N_749,N_956);
nor U1105 (N_1105,N_665,N_465);
and U1106 (N_1106,N_728,N_560);
or U1107 (N_1107,N_78,N_327);
nand U1108 (N_1108,N_910,N_74);
nor U1109 (N_1109,N_427,N_247);
nand U1110 (N_1110,N_42,N_170);
and U1111 (N_1111,N_993,N_272);
nor U1112 (N_1112,N_908,N_839);
and U1113 (N_1113,N_490,N_601);
or U1114 (N_1114,N_633,N_669);
xnor U1115 (N_1115,N_153,N_298);
xor U1116 (N_1116,N_90,N_425);
and U1117 (N_1117,N_877,N_423);
nand U1118 (N_1118,N_567,N_703);
nor U1119 (N_1119,N_346,N_397);
and U1120 (N_1120,N_562,N_264);
nand U1121 (N_1121,N_551,N_772);
nand U1122 (N_1122,N_694,N_619);
and U1123 (N_1123,N_532,N_641);
nor U1124 (N_1124,N_630,N_621);
and U1125 (N_1125,N_175,N_112);
or U1126 (N_1126,N_62,N_706);
nand U1127 (N_1127,N_682,N_803);
and U1128 (N_1128,N_100,N_457);
nor U1129 (N_1129,N_584,N_882);
or U1130 (N_1130,N_722,N_456);
or U1131 (N_1131,N_819,N_91);
nor U1132 (N_1132,N_462,N_991);
and U1133 (N_1133,N_814,N_85);
or U1134 (N_1134,N_145,N_953);
nor U1135 (N_1135,N_137,N_775);
nor U1136 (N_1136,N_342,N_746);
and U1137 (N_1137,N_221,N_307);
xor U1138 (N_1138,N_202,N_771);
and U1139 (N_1139,N_45,N_296);
nand U1140 (N_1140,N_119,N_859);
nand U1141 (N_1141,N_927,N_273);
and U1142 (N_1142,N_36,N_675);
or U1143 (N_1143,N_904,N_702);
nor U1144 (N_1144,N_256,N_709);
nand U1145 (N_1145,N_768,N_545);
xnor U1146 (N_1146,N_283,N_579);
and U1147 (N_1147,N_876,N_439);
and U1148 (N_1148,N_152,N_480);
nand U1149 (N_1149,N_35,N_387);
nor U1150 (N_1150,N_729,N_353);
or U1151 (N_1151,N_396,N_356);
and U1152 (N_1152,N_370,N_289);
or U1153 (N_1153,N_388,N_55);
nor U1154 (N_1154,N_530,N_950);
nor U1155 (N_1155,N_580,N_181);
and U1156 (N_1156,N_661,N_690);
nor U1157 (N_1157,N_333,N_258);
nor U1158 (N_1158,N_916,N_674);
nand U1159 (N_1159,N_928,N_821);
and U1160 (N_1160,N_280,N_328);
or U1161 (N_1161,N_512,N_985);
and U1162 (N_1162,N_673,N_571);
or U1163 (N_1163,N_197,N_191);
and U1164 (N_1164,N_730,N_522);
or U1165 (N_1165,N_826,N_758);
xor U1166 (N_1166,N_879,N_149);
and U1167 (N_1167,N_76,N_643);
or U1168 (N_1168,N_487,N_615);
nand U1169 (N_1169,N_592,N_645);
nand U1170 (N_1170,N_636,N_854);
xnor U1171 (N_1171,N_12,N_811);
nor U1172 (N_1172,N_239,N_858);
or U1173 (N_1173,N_200,N_719);
nor U1174 (N_1174,N_828,N_837);
nand U1175 (N_1175,N_499,N_655);
and U1176 (N_1176,N_309,N_585);
nand U1177 (N_1177,N_686,N_315);
nand U1178 (N_1178,N_306,N_971);
nand U1179 (N_1179,N_566,N_223);
nand U1180 (N_1180,N_704,N_736);
nand U1181 (N_1181,N_196,N_22);
xor U1182 (N_1182,N_795,N_14);
nand U1183 (N_1183,N_248,N_81);
and U1184 (N_1184,N_493,N_582);
or U1185 (N_1185,N_446,N_358);
xnor U1186 (N_1186,N_163,N_102);
nand U1187 (N_1187,N_374,N_1);
and U1188 (N_1188,N_430,N_458);
nand U1189 (N_1189,N_864,N_798);
or U1190 (N_1190,N_451,N_903);
xor U1191 (N_1191,N_220,N_791);
nand U1192 (N_1192,N_147,N_262);
nand U1193 (N_1193,N_510,N_528);
nor U1194 (N_1194,N_127,N_938);
nand U1195 (N_1195,N_101,N_933);
nand U1196 (N_1196,N_351,N_939);
and U1197 (N_1197,N_187,N_179);
nand U1198 (N_1198,N_382,N_820);
xor U1199 (N_1199,N_866,N_818);
nand U1200 (N_1200,N_835,N_907);
nor U1201 (N_1201,N_945,N_754);
nor U1202 (N_1202,N_762,N_39);
nand U1203 (N_1203,N_631,N_932);
and U1204 (N_1204,N_408,N_402);
nand U1205 (N_1205,N_173,N_322);
and U1206 (N_1206,N_57,N_336);
or U1207 (N_1207,N_51,N_638);
and U1208 (N_1208,N_249,N_29);
nand U1209 (N_1209,N_195,N_150);
and U1210 (N_1210,N_549,N_604);
nor U1211 (N_1211,N_853,N_193);
or U1212 (N_1212,N_414,N_610);
nor U1213 (N_1213,N_213,N_438);
xnor U1214 (N_1214,N_437,N_880);
nor U1215 (N_1215,N_25,N_529);
nor U1216 (N_1216,N_648,N_505);
and U1217 (N_1217,N_218,N_963);
nor U1218 (N_1218,N_940,N_114);
nor U1219 (N_1219,N_44,N_806);
nand U1220 (N_1220,N_350,N_917);
or U1221 (N_1221,N_915,N_887);
and U1222 (N_1222,N_472,N_657);
or U1223 (N_1223,N_318,N_189);
nor U1224 (N_1224,N_761,N_61);
xnor U1225 (N_1225,N_468,N_169);
nand U1226 (N_1226,N_6,N_434);
nor U1227 (N_1227,N_976,N_54);
or U1228 (N_1228,N_108,N_593);
nand U1229 (N_1229,N_347,N_357);
xnor U1230 (N_1230,N_52,N_670);
nor U1231 (N_1231,N_28,N_46);
or U1232 (N_1232,N_575,N_883);
xor U1233 (N_1233,N_67,N_205);
or U1234 (N_1234,N_534,N_418);
and U1235 (N_1235,N_41,N_11);
or U1236 (N_1236,N_676,N_470);
and U1237 (N_1237,N_341,N_874);
xnor U1238 (N_1238,N_732,N_747);
nor U1239 (N_1239,N_894,N_905);
nand U1240 (N_1240,N_422,N_365);
and U1241 (N_1241,N_139,N_228);
or U1242 (N_1242,N_598,N_809);
or U1243 (N_1243,N_931,N_606);
nand U1244 (N_1244,N_447,N_276);
xor U1245 (N_1245,N_118,N_832);
or U1246 (N_1246,N_469,N_429);
or U1247 (N_1247,N_122,N_836);
nor U1248 (N_1248,N_494,N_227);
or U1249 (N_1249,N_748,N_436);
or U1250 (N_1250,N_392,N_411);
nor U1251 (N_1251,N_496,N_449);
nand U1252 (N_1252,N_737,N_319);
and U1253 (N_1253,N_268,N_368);
or U1254 (N_1254,N_440,N_334);
nor U1255 (N_1255,N_491,N_160);
nand U1256 (N_1256,N_165,N_410);
and U1257 (N_1257,N_216,N_552);
nand U1258 (N_1258,N_15,N_186);
and U1259 (N_1259,N_497,N_428);
xnor U1260 (N_1260,N_889,N_110);
and U1261 (N_1261,N_294,N_952);
nand U1262 (N_1262,N_308,N_199);
or U1263 (N_1263,N_533,N_312);
nor U1264 (N_1264,N_501,N_518);
xor U1265 (N_1265,N_725,N_106);
and U1266 (N_1266,N_852,N_21);
or U1267 (N_1267,N_476,N_521);
xnor U1268 (N_1268,N_325,N_683);
nand U1269 (N_1269,N_30,N_445);
nand U1270 (N_1270,N_861,N_829);
or U1271 (N_1271,N_526,N_688);
and U1272 (N_1272,N_245,N_369);
nand U1273 (N_1273,N_18,N_750);
nand U1274 (N_1274,N_53,N_846);
nand U1275 (N_1275,N_123,N_799);
or U1276 (N_1276,N_868,N_658);
or U1277 (N_1277,N_611,N_323);
nand U1278 (N_1278,N_409,N_359);
nor U1279 (N_1279,N_838,N_75);
nand U1280 (N_1280,N_524,N_664);
nor U1281 (N_1281,N_995,N_134);
or U1282 (N_1282,N_166,N_176);
xor U1283 (N_1283,N_484,N_812);
or U1284 (N_1284,N_103,N_744);
nand U1285 (N_1285,N_538,N_64);
nand U1286 (N_1286,N_934,N_461);
nand U1287 (N_1287,N_869,N_488);
nor U1288 (N_1288,N_105,N_133);
nand U1289 (N_1289,N_698,N_475);
nand U1290 (N_1290,N_766,N_361);
nor U1291 (N_1291,N_509,N_344);
nor U1292 (N_1292,N_711,N_959);
xor U1293 (N_1293,N_871,N_672);
nor U1294 (N_1294,N_557,N_659);
nand U1295 (N_1295,N_313,N_69);
nand U1296 (N_1296,N_845,N_231);
or U1297 (N_1297,N_282,N_407);
or U1298 (N_1298,N_464,N_547);
nor U1299 (N_1299,N_893,N_254);
nand U1300 (N_1300,N_810,N_678);
or U1301 (N_1301,N_577,N_183);
nand U1302 (N_1302,N_779,N_471);
nand U1303 (N_1303,N_31,N_514);
xnor U1304 (N_1304,N_331,N_332);
nand U1305 (N_1305,N_987,N_366);
nor U1306 (N_1306,N_420,N_742);
or U1307 (N_1307,N_87,N_337);
nor U1308 (N_1308,N_544,N_667);
or U1309 (N_1309,N_415,N_569);
xnor U1310 (N_1310,N_937,N_211);
and U1311 (N_1311,N_303,N_695);
nand U1312 (N_1312,N_572,N_700);
nand U1313 (N_1313,N_378,N_261);
and U1314 (N_1314,N_115,N_909);
and U1315 (N_1315,N_851,N_317);
or U1316 (N_1316,N_395,N_304);
xor U1317 (N_1317,N_620,N_885);
nand U1318 (N_1318,N_625,N_241);
nor U1319 (N_1319,N_857,N_390);
or U1320 (N_1320,N_715,N_489);
xnor U1321 (N_1321,N_975,N_285);
nor U1322 (N_1322,N_738,N_80);
and U1323 (N_1323,N_33,N_617);
or U1324 (N_1324,N_825,N_399);
nor U1325 (N_1325,N_727,N_240);
and U1326 (N_1326,N_274,N_965);
and U1327 (N_1327,N_109,N_340);
nand U1328 (N_1328,N_19,N_117);
nand U1329 (N_1329,N_988,N_559);
or U1330 (N_1330,N_757,N_345);
nand U1331 (N_1331,N_314,N_895);
or U1332 (N_1332,N_925,N_977);
nand U1333 (N_1333,N_929,N_961);
xnor U1334 (N_1334,N_343,N_454);
and U1335 (N_1335,N_589,N_607);
nor U1336 (N_1336,N_774,N_73);
xnor U1337 (N_1337,N_958,N_8);
and U1338 (N_1338,N_967,N_329);
xnor U1339 (N_1339,N_890,N_546);
nand U1340 (N_1340,N_43,N_7);
nor U1341 (N_1341,N_413,N_113);
or U1342 (N_1342,N_781,N_271);
nand U1343 (N_1343,N_431,N_467);
nor U1344 (N_1344,N_111,N_637);
nand U1345 (N_1345,N_63,N_167);
nand U1346 (N_1346,N_741,N_383);
nor U1347 (N_1347,N_878,N_473);
and U1348 (N_1348,N_275,N_398);
xnor U1349 (N_1349,N_238,N_586);
nor U1350 (N_1350,N_717,N_924);
xor U1351 (N_1351,N_391,N_219);
nand U1352 (N_1352,N_482,N_367);
nor U1353 (N_1353,N_677,N_287);
nand U1354 (N_1354,N_203,N_684);
nor U1355 (N_1355,N_234,N_726);
nand U1356 (N_1356,N_230,N_125);
or U1357 (N_1357,N_148,N_297);
nand U1358 (N_1358,N_860,N_376);
or U1359 (N_1359,N_237,N_266);
xnor U1360 (N_1360,N_896,N_403);
and U1361 (N_1361,N_640,N_870);
or U1362 (N_1362,N_783,N_962);
xnor U1363 (N_1363,N_780,N_823);
nand U1364 (N_1364,N_680,N_596);
nand U1365 (N_1365,N_855,N_647);
nand U1366 (N_1366,N_47,N_535);
nand U1367 (N_1367,N_740,N_379);
nor U1368 (N_1368,N_989,N_833);
and U1369 (N_1369,N_943,N_983);
and U1370 (N_1370,N_841,N_94);
nand U1371 (N_1371,N_970,N_537);
and U1372 (N_1372,N_229,N_605);
and U1373 (N_1373,N_807,N_842);
xor U1374 (N_1374,N_120,N_9);
nor U1375 (N_1375,N_394,N_755);
or U1376 (N_1376,N_37,N_960);
xor U1377 (N_1377,N_595,N_66);
or U1378 (N_1378,N_608,N_417);
xnor U1379 (N_1379,N_389,N_587);
or U1380 (N_1380,N_246,N_922);
xnor U1381 (N_1381,N_459,N_162);
nand U1382 (N_1382,N_478,N_190);
nand U1383 (N_1383,N_92,N_671);
nor U1384 (N_1384,N_901,N_561);
or U1385 (N_1385,N_918,N_583);
or U1386 (N_1386,N_921,N_286);
nor U1387 (N_1387,N_178,N_713);
nor U1388 (N_1388,N_270,N_5);
nor U1389 (N_1389,N_531,N_455);
nor U1390 (N_1390,N_564,N_996);
nor U1391 (N_1391,N_466,N_511);
nor U1392 (N_1392,N_710,N_384);
nand U1393 (N_1393,N_156,N_863);
nand U1394 (N_1394,N_777,N_184);
or U1395 (N_1395,N_128,N_716);
nor U1396 (N_1396,N_84,N_479);
and U1397 (N_1397,N_316,N_305);
nand U1398 (N_1398,N_335,N_542);
nor U1399 (N_1399,N_760,N_330);
or U1400 (N_1400,N_508,N_627);
xor U1401 (N_1401,N_259,N_355);
nor U1402 (N_1402,N_265,N_281);
or U1403 (N_1403,N_393,N_38);
and U1404 (N_1404,N_144,N_513);
xor U1405 (N_1405,N_776,N_210);
nand U1406 (N_1406,N_541,N_444);
nor U1407 (N_1407,N_941,N_724);
and U1408 (N_1408,N_652,N_375);
nand U1409 (N_1409,N_802,N_913);
xor U1410 (N_1410,N_632,N_143);
nor U1411 (N_1411,N_785,N_138);
or U1412 (N_1412,N_752,N_68);
or U1413 (N_1413,N_926,N_500);
and U1414 (N_1414,N_847,N_70);
nor U1415 (N_1415,N_856,N_385);
or U1416 (N_1416,N_687,N_136);
xor U1417 (N_1417,N_553,N_558);
and U1418 (N_1418,N_441,N_16);
nand U1419 (N_1419,N_867,N_481);
and U1420 (N_1420,N_460,N_89);
nand U1421 (N_1421,N_154,N_609);
nand U1422 (N_1422,N_321,N_326);
nor U1423 (N_1423,N_721,N_796);
nand U1424 (N_1424,N_96,N_646);
and U1425 (N_1425,N_291,N_668);
or U1426 (N_1426,N_824,N_735);
nand U1427 (N_1427,N_226,N_600);
nor U1428 (N_1428,N_944,N_815);
and U1429 (N_1429,N_222,N_377);
nor U1430 (N_1430,N_320,N_912);
nand U1431 (N_1431,N_689,N_502);
or U1432 (N_1432,N_523,N_290);
nand U1433 (N_1433,N_421,N_565);
nor U1434 (N_1434,N_95,N_734);
or U1435 (N_1435,N_232,N_435);
or U1436 (N_1436,N_840,N_432);
nand U1437 (N_1437,N_759,N_955);
nor U1438 (N_1438,N_651,N_363);
or U1439 (N_1439,N_311,N_310);
or U1440 (N_1440,N_50,N_34);
xnor U1441 (N_1441,N_765,N_477);
nand U1442 (N_1442,N_568,N_58);
nand U1443 (N_1443,N_443,N_242);
or U1444 (N_1444,N_830,N_300);
and U1445 (N_1445,N_642,N_892);
and U1446 (N_1446,N_131,N_692);
nand U1447 (N_1447,N_233,N_86);
nand U1448 (N_1448,N_354,N_753);
and U1449 (N_1449,N_284,N_822);
nand U1450 (N_1450,N_97,N_424);
nand U1451 (N_1451,N_158,N_77);
or U1452 (N_1452,N_404,N_591);
nor U1453 (N_1453,N_412,N_662);
nor U1454 (N_1454,N_172,N_124);
nor U1455 (N_1455,N_349,N_244);
and U1456 (N_1456,N_279,N_911);
nor U1457 (N_1457,N_204,N_578);
xor U1458 (N_1458,N_850,N_519);
or U1459 (N_1459,N_302,N_685);
or U1460 (N_1460,N_998,N_653);
nand U1461 (N_1461,N_898,N_485);
nand U1462 (N_1462,N_56,N_324);
nand U1463 (N_1463,N_900,N_739);
and U1464 (N_1464,N_515,N_973);
xor U1465 (N_1465,N_161,N_556);
and U1466 (N_1466,N_570,N_252);
or U1467 (N_1467,N_733,N_224);
and U1468 (N_1468,N_769,N_936);
nand U1469 (N_1469,N_236,N_705);
nand U1470 (N_1470,N_951,N_743);
nor U1471 (N_1471,N_875,N_225);
nor U1472 (N_1472,N_576,N_555);
and U1473 (N_1473,N_182,N_194);
nor U1474 (N_1474,N_613,N_718);
nand U1475 (N_1475,N_731,N_597);
nor U1476 (N_1476,N_644,N_474);
and U1477 (N_1477,N_602,N_942);
nor U1478 (N_1478,N_980,N_40);
or U1479 (N_1479,N_24,N_3);
and U1480 (N_1480,N_453,N_129);
and U1481 (N_1481,N_969,N_563);
and U1482 (N_1482,N_813,N_794);
or U1483 (N_1483,N_540,N_433);
and U1484 (N_1484,N_793,N_146);
and U1485 (N_1485,N_816,N_654);
xnor U1486 (N_1486,N_629,N_701);
nand U1487 (N_1487,N_121,N_132);
and U1488 (N_1488,N_966,N_770);
and U1489 (N_1489,N_177,N_267);
or U1490 (N_1490,N_135,N_104);
or U1491 (N_1491,N_663,N_699);
or U1492 (N_1492,N_707,N_442);
nand U1493 (N_1493,N_372,N_141);
and U1494 (N_1494,N_635,N_269);
and U1495 (N_1495,N_884,N_539);
and U1496 (N_1496,N_614,N_192);
nor U1497 (N_1497,N_255,N_946);
nand U1498 (N_1498,N_778,N_151);
nand U1499 (N_1499,N_164,N_288);
and U1500 (N_1500,N_741,N_339);
xnor U1501 (N_1501,N_998,N_257);
nor U1502 (N_1502,N_64,N_875);
or U1503 (N_1503,N_70,N_86);
xor U1504 (N_1504,N_266,N_770);
xor U1505 (N_1505,N_464,N_775);
xnor U1506 (N_1506,N_646,N_682);
or U1507 (N_1507,N_407,N_333);
and U1508 (N_1508,N_305,N_675);
nor U1509 (N_1509,N_372,N_712);
or U1510 (N_1510,N_467,N_963);
nor U1511 (N_1511,N_992,N_437);
and U1512 (N_1512,N_903,N_428);
nand U1513 (N_1513,N_197,N_742);
xor U1514 (N_1514,N_871,N_178);
or U1515 (N_1515,N_571,N_865);
or U1516 (N_1516,N_75,N_22);
nand U1517 (N_1517,N_733,N_923);
and U1518 (N_1518,N_11,N_316);
nor U1519 (N_1519,N_713,N_110);
nand U1520 (N_1520,N_497,N_855);
nor U1521 (N_1521,N_62,N_304);
and U1522 (N_1522,N_86,N_756);
or U1523 (N_1523,N_959,N_541);
or U1524 (N_1524,N_876,N_3);
or U1525 (N_1525,N_776,N_259);
or U1526 (N_1526,N_443,N_138);
and U1527 (N_1527,N_309,N_254);
xor U1528 (N_1528,N_496,N_31);
or U1529 (N_1529,N_673,N_96);
and U1530 (N_1530,N_297,N_448);
nor U1531 (N_1531,N_284,N_825);
and U1532 (N_1532,N_681,N_328);
xnor U1533 (N_1533,N_667,N_964);
nor U1534 (N_1534,N_508,N_419);
or U1535 (N_1535,N_389,N_433);
and U1536 (N_1536,N_289,N_648);
nand U1537 (N_1537,N_356,N_335);
xor U1538 (N_1538,N_277,N_513);
or U1539 (N_1539,N_953,N_839);
nor U1540 (N_1540,N_594,N_854);
nand U1541 (N_1541,N_419,N_946);
nand U1542 (N_1542,N_104,N_373);
nor U1543 (N_1543,N_922,N_773);
nand U1544 (N_1544,N_868,N_810);
nand U1545 (N_1545,N_925,N_481);
xnor U1546 (N_1546,N_51,N_156);
nor U1547 (N_1547,N_140,N_28);
nand U1548 (N_1548,N_78,N_107);
nor U1549 (N_1549,N_433,N_19);
nand U1550 (N_1550,N_511,N_650);
or U1551 (N_1551,N_527,N_512);
nand U1552 (N_1552,N_323,N_215);
or U1553 (N_1553,N_648,N_600);
nand U1554 (N_1554,N_763,N_242);
nor U1555 (N_1555,N_851,N_533);
xor U1556 (N_1556,N_471,N_272);
or U1557 (N_1557,N_408,N_941);
nand U1558 (N_1558,N_622,N_91);
and U1559 (N_1559,N_579,N_442);
nor U1560 (N_1560,N_983,N_959);
nor U1561 (N_1561,N_795,N_708);
nand U1562 (N_1562,N_802,N_869);
nor U1563 (N_1563,N_347,N_577);
nor U1564 (N_1564,N_618,N_115);
nand U1565 (N_1565,N_655,N_397);
nand U1566 (N_1566,N_911,N_267);
nor U1567 (N_1567,N_872,N_87);
nor U1568 (N_1568,N_580,N_487);
and U1569 (N_1569,N_380,N_579);
nand U1570 (N_1570,N_203,N_476);
or U1571 (N_1571,N_990,N_500);
or U1572 (N_1572,N_121,N_209);
nand U1573 (N_1573,N_731,N_294);
and U1574 (N_1574,N_125,N_774);
or U1575 (N_1575,N_252,N_673);
xnor U1576 (N_1576,N_548,N_660);
or U1577 (N_1577,N_688,N_735);
xnor U1578 (N_1578,N_103,N_73);
or U1579 (N_1579,N_533,N_679);
and U1580 (N_1580,N_818,N_814);
nor U1581 (N_1581,N_115,N_711);
nor U1582 (N_1582,N_16,N_324);
nand U1583 (N_1583,N_679,N_61);
nand U1584 (N_1584,N_592,N_492);
nand U1585 (N_1585,N_902,N_461);
nor U1586 (N_1586,N_52,N_65);
nor U1587 (N_1587,N_748,N_605);
xor U1588 (N_1588,N_641,N_427);
and U1589 (N_1589,N_328,N_690);
and U1590 (N_1590,N_396,N_251);
nand U1591 (N_1591,N_561,N_673);
nor U1592 (N_1592,N_471,N_846);
nand U1593 (N_1593,N_669,N_515);
or U1594 (N_1594,N_282,N_924);
and U1595 (N_1595,N_177,N_474);
nand U1596 (N_1596,N_991,N_951);
nor U1597 (N_1597,N_973,N_882);
nand U1598 (N_1598,N_284,N_926);
nand U1599 (N_1599,N_921,N_689);
and U1600 (N_1600,N_941,N_182);
or U1601 (N_1601,N_230,N_873);
xor U1602 (N_1602,N_635,N_713);
and U1603 (N_1603,N_754,N_306);
nand U1604 (N_1604,N_655,N_488);
nor U1605 (N_1605,N_670,N_752);
nand U1606 (N_1606,N_281,N_483);
or U1607 (N_1607,N_650,N_369);
nand U1608 (N_1608,N_818,N_939);
nand U1609 (N_1609,N_216,N_395);
nand U1610 (N_1610,N_194,N_59);
xnor U1611 (N_1611,N_548,N_565);
nand U1612 (N_1612,N_737,N_200);
and U1613 (N_1613,N_556,N_356);
nor U1614 (N_1614,N_797,N_101);
nor U1615 (N_1615,N_665,N_323);
and U1616 (N_1616,N_895,N_936);
nand U1617 (N_1617,N_463,N_473);
nor U1618 (N_1618,N_252,N_626);
or U1619 (N_1619,N_344,N_963);
and U1620 (N_1620,N_804,N_908);
nand U1621 (N_1621,N_351,N_147);
nand U1622 (N_1622,N_338,N_305);
or U1623 (N_1623,N_208,N_599);
nor U1624 (N_1624,N_860,N_560);
or U1625 (N_1625,N_560,N_294);
nor U1626 (N_1626,N_563,N_818);
nand U1627 (N_1627,N_205,N_964);
xor U1628 (N_1628,N_625,N_614);
xnor U1629 (N_1629,N_746,N_293);
nor U1630 (N_1630,N_949,N_370);
or U1631 (N_1631,N_815,N_541);
nor U1632 (N_1632,N_562,N_45);
and U1633 (N_1633,N_899,N_146);
or U1634 (N_1634,N_798,N_151);
nor U1635 (N_1635,N_353,N_968);
or U1636 (N_1636,N_601,N_13);
and U1637 (N_1637,N_560,N_819);
or U1638 (N_1638,N_709,N_446);
nand U1639 (N_1639,N_242,N_453);
nor U1640 (N_1640,N_87,N_452);
nor U1641 (N_1641,N_300,N_27);
or U1642 (N_1642,N_444,N_815);
and U1643 (N_1643,N_664,N_915);
nor U1644 (N_1644,N_225,N_366);
and U1645 (N_1645,N_678,N_92);
and U1646 (N_1646,N_555,N_440);
nand U1647 (N_1647,N_709,N_871);
nand U1648 (N_1648,N_888,N_160);
and U1649 (N_1649,N_291,N_138);
xor U1650 (N_1650,N_477,N_421);
nand U1651 (N_1651,N_629,N_601);
nor U1652 (N_1652,N_34,N_934);
xnor U1653 (N_1653,N_462,N_183);
nor U1654 (N_1654,N_618,N_375);
nor U1655 (N_1655,N_602,N_279);
nor U1656 (N_1656,N_532,N_251);
nand U1657 (N_1657,N_422,N_9);
nand U1658 (N_1658,N_738,N_438);
or U1659 (N_1659,N_220,N_51);
or U1660 (N_1660,N_924,N_73);
nand U1661 (N_1661,N_724,N_631);
nor U1662 (N_1662,N_900,N_902);
or U1663 (N_1663,N_10,N_449);
nor U1664 (N_1664,N_367,N_973);
and U1665 (N_1665,N_326,N_40);
nor U1666 (N_1666,N_721,N_829);
nor U1667 (N_1667,N_580,N_625);
and U1668 (N_1668,N_114,N_35);
nor U1669 (N_1669,N_700,N_876);
and U1670 (N_1670,N_596,N_638);
or U1671 (N_1671,N_442,N_753);
nand U1672 (N_1672,N_96,N_405);
xnor U1673 (N_1673,N_418,N_21);
and U1674 (N_1674,N_629,N_784);
nand U1675 (N_1675,N_4,N_822);
nand U1676 (N_1676,N_566,N_570);
nor U1677 (N_1677,N_55,N_806);
nand U1678 (N_1678,N_719,N_885);
and U1679 (N_1679,N_688,N_125);
nand U1680 (N_1680,N_555,N_57);
and U1681 (N_1681,N_650,N_868);
xor U1682 (N_1682,N_664,N_272);
or U1683 (N_1683,N_140,N_534);
nand U1684 (N_1684,N_814,N_446);
and U1685 (N_1685,N_596,N_908);
or U1686 (N_1686,N_77,N_312);
nand U1687 (N_1687,N_218,N_431);
nor U1688 (N_1688,N_369,N_255);
xor U1689 (N_1689,N_958,N_111);
nand U1690 (N_1690,N_214,N_290);
xnor U1691 (N_1691,N_693,N_667);
or U1692 (N_1692,N_785,N_399);
xnor U1693 (N_1693,N_334,N_365);
and U1694 (N_1694,N_414,N_960);
nand U1695 (N_1695,N_649,N_782);
nor U1696 (N_1696,N_103,N_222);
or U1697 (N_1697,N_452,N_432);
nor U1698 (N_1698,N_154,N_459);
nand U1699 (N_1699,N_4,N_448);
or U1700 (N_1700,N_863,N_393);
nand U1701 (N_1701,N_321,N_242);
nand U1702 (N_1702,N_713,N_283);
or U1703 (N_1703,N_437,N_740);
nor U1704 (N_1704,N_270,N_751);
nor U1705 (N_1705,N_142,N_75);
nand U1706 (N_1706,N_460,N_782);
nand U1707 (N_1707,N_867,N_488);
and U1708 (N_1708,N_120,N_113);
nand U1709 (N_1709,N_59,N_389);
or U1710 (N_1710,N_31,N_1);
nand U1711 (N_1711,N_691,N_525);
or U1712 (N_1712,N_108,N_51);
nand U1713 (N_1713,N_847,N_456);
or U1714 (N_1714,N_985,N_618);
nor U1715 (N_1715,N_745,N_837);
nand U1716 (N_1716,N_313,N_299);
xnor U1717 (N_1717,N_175,N_890);
or U1718 (N_1718,N_799,N_143);
or U1719 (N_1719,N_257,N_272);
xor U1720 (N_1720,N_534,N_30);
nand U1721 (N_1721,N_810,N_299);
or U1722 (N_1722,N_281,N_585);
and U1723 (N_1723,N_829,N_493);
nand U1724 (N_1724,N_455,N_607);
nand U1725 (N_1725,N_192,N_743);
xor U1726 (N_1726,N_488,N_532);
and U1727 (N_1727,N_839,N_937);
nand U1728 (N_1728,N_8,N_674);
nor U1729 (N_1729,N_671,N_100);
or U1730 (N_1730,N_133,N_365);
nor U1731 (N_1731,N_402,N_896);
xor U1732 (N_1732,N_143,N_804);
and U1733 (N_1733,N_75,N_706);
and U1734 (N_1734,N_773,N_13);
xor U1735 (N_1735,N_870,N_167);
nor U1736 (N_1736,N_58,N_179);
xor U1737 (N_1737,N_10,N_661);
xor U1738 (N_1738,N_524,N_509);
or U1739 (N_1739,N_29,N_287);
nand U1740 (N_1740,N_939,N_529);
and U1741 (N_1741,N_309,N_723);
or U1742 (N_1742,N_980,N_956);
nand U1743 (N_1743,N_958,N_470);
nor U1744 (N_1744,N_11,N_434);
and U1745 (N_1745,N_731,N_319);
nor U1746 (N_1746,N_798,N_910);
nor U1747 (N_1747,N_859,N_84);
nor U1748 (N_1748,N_360,N_908);
and U1749 (N_1749,N_391,N_395);
nor U1750 (N_1750,N_454,N_67);
nand U1751 (N_1751,N_40,N_226);
nor U1752 (N_1752,N_736,N_678);
nor U1753 (N_1753,N_660,N_11);
and U1754 (N_1754,N_189,N_919);
xnor U1755 (N_1755,N_307,N_931);
nand U1756 (N_1756,N_749,N_738);
and U1757 (N_1757,N_267,N_671);
nor U1758 (N_1758,N_991,N_578);
or U1759 (N_1759,N_512,N_98);
nand U1760 (N_1760,N_531,N_452);
nor U1761 (N_1761,N_777,N_891);
xor U1762 (N_1762,N_689,N_245);
nor U1763 (N_1763,N_921,N_120);
nor U1764 (N_1764,N_415,N_681);
nor U1765 (N_1765,N_426,N_519);
nor U1766 (N_1766,N_735,N_513);
or U1767 (N_1767,N_37,N_801);
and U1768 (N_1768,N_342,N_437);
nor U1769 (N_1769,N_562,N_853);
or U1770 (N_1770,N_235,N_767);
or U1771 (N_1771,N_592,N_714);
or U1772 (N_1772,N_271,N_440);
xnor U1773 (N_1773,N_395,N_708);
nor U1774 (N_1774,N_814,N_750);
nor U1775 (N_1775,N_249,N_722);
or U1776 (N_1776,N_730,N_292);
nor U1777 (N_1777,N_627,N_482);
xnor U1778 (N_1778,N_492,N_850);
and U1779 (N_1779,N_233,N_606);
nand U1780 (N_1780,N_21,N_751);
nor U1781 (N_1781,N_383,N_7);
nand U1782 (N_1782,N_252,N_959);
or U1783 (N_1783,N_342,N_553);
and U1784 (N_1784,N_779,N_293);
or U1785 (N_1785,N_120,N_493);
or U1786 (N_1786,N_652,N_970);
nand U1787 (N_1787,N_493,N_674);
nand U1788 (N_1788,N_550,N_945);
nand U1789 (N_1789,N_156,N_98);
or U1790 (N_1790,N_145,N_987);
and U1791 (N_1791,N_946,N_124);
xnor U1792 (N_1792,N_370,N_673);
and U1793 (N_1793,N_710,N_677);
or U1794 (N_1794,N_335,N_515);
xor U1795 (N_1795,N_379,N_731);
or U1796 (N_1796,N_766,N_250);
xnor U1797 (N_1797,N_314,N_738);
or U1798 (N_1798,N_972,N_861);
nor U1799 (N_1799,N_988,N_51);
and U1800 (N_1800,N_619,N_601);
xnor U1801 (N_1801,N_93,N_893);
and U1802 (N_1802,N_417,N_225);
or U1803 (N_1803,N_730,N_215);
or U1804 (N_1804,N_38,N_80);
xnor U1805 (N_1805,N_481,N_434);
nand U1806 (N_1806,N_755,N_933);
and U1807 (N_1807,N_270,N_108);
and U1808 (N_1808,N_715,N_166);
and U1809 (N_1809,N_812,N_583);
or U1810 (N_1810,N_206,N_396);
nand U1811 (N_1811,N_928,N_861);
nand U1812 (N_1812,N_240,N_951);
nand U1813 (N_1813,N_932,N_309);
and U1814 (N_1814,N_277,N_143);
xnor U1815 (N_1815,N_27,N_522);
and U1816 (N_1816,N_702,N_290);
and U1817 (N_1817,N_920,N_262);
or U1818 (N_1818,N_664,N_80);
nand U1819 (N_1819,N_420,N_873);
and U1820 (N_1820,N_249,N_951);
nand U1821 (N_1821,N_224,N_33);
and U1822 (N_1822,N_711,N_241);
or U1823 (N_1823,N_835,N_35);
nand U1824 (N_1824,N_175,N_302);
nand U1825 (N_1825,N_238,N_691);
or U1826 (N_1826,N_724,N_401);
nor U1827 (N_1827,N_431,N_479);
nor U1828 (N_1828,N_661,N_944);
nand U1829 (N_1829,N_497,N_890);
nand U1830 (N_1830,N_60,N_962);
nand U1831 (N_1831,N_294,N_386);
or U1832 (N_1832,N_670,N_213);
or U1833 (N_1833,N_607,N_630);
nand U1834 (N_1834,N_980,N_823);
nor U1835 (N_1835,N_825,N_978);
and U1836 (N_1836,N_604,N_816);
or U1837 (N_1837,N_91,N_544);
nand U1838 (N_1838,N_397,N_614);
or U1839 (N_1839,N_653,N_151);
nor U1840 (N_1840,N_847,N_628);
nand U1841 (N_1841,N_389,N_653);
and U1842 (N_1842,N_892,N_819);
nand U1843 (N_1843,N_536,N_290);
nor U1844 (N_1844,N_64,N_573);
or U1845 (N_1845,N_80,N_780);
nor U1846 (N_1846,N_681,N_701);
or U1847 (N_1847,N_336,N_288);
or U1848 (N_1848,N_192,N_381);
or U1849 (N_1849,N_208,N_233);
or U1850 (N_1850,N_76,N_884);
nand U1851 (N_1851,N_613,N_968);
and U1852 (N_1852,N_420,N_107);
nand U1853 (N_1853,N_858,N_922);
or U1854 (N_1854,N_558,N_236);
or U1855 (N_1855,N_645,N_447);
and U1856 (N_1856,N_959,N_52);
or U1857 (N_1857,N_222,N_290);
nor U1858 (N_1858,N_317,N_541);
xnor U1859 (N_1859,N_27,N_541);
xnor U1860 (N_1860,N_567,N_929);
nand U1861 (N_1861,N_516,N_834);
nand U1862 (N_1862,N_492,N_269);
nand U1863 (N_1863,N_198,N_502);
and U1864 (N_1864,N_306,N_463);
nor U1865 (N_1865,N_463,N_693);
nor U1866 (N_1866,N_664,N_687);
nand U1867 (N_1867,N_545,N_401);
or U1868 (N_1868,N_13,N_429);
nand U1869 (N_1869,N_85,N_697);
nor U1870 (N_1870,N_571,N_941);
or U1871 (N_1871,N_277,N_543);
or U1872 (N_1872,N_763,N_476);
nor U1873 (N_1873,N_487,N_59);
and U1874 (N_1874,N_643,N_911);
or U1875 (N_1875,N_622,N_505);
nand U1876 (N_1876,N_799,N_896);
or U1877 (N_1877,N_137,N_540);
or U1878 (N_1878,N_823,N_393);
nand U1879 (N_1879,N_538,N_847);
nor U1880 (N_1880,N_790,N_507);
or U1881 (N_1881,N_728,N_586);
and U1882 (N_1882,N_478,N_932);
or U1883 (N_1883,N_250,N_413);
or U1884 (N_1884,N_276,N_615);
and U1885 (N_1885,N_935,N_290);
or U1886 (N_1886,N_172,N_897);
and U1887 (N_1887,N_600,N_507);
nor U1888 (N_1888,N_836,N_245);
or U1889 (N_1889,N_188,N_263);
and U1890 (N_1890,N_108,N_581);
or U1891 (N_1891,N_633,N_76);
nor U1892 (N_1892,N_783,N_184);
and U1893 (N_1893,N_737,N_678);
nor U1894 (N_1894,N_402,N_200);
or U1895 (N_1895,N_569,N_335);
nor U1896 (N_1896,N_565,N_499);
or U1897 (N_1897,N_899,N_510);
nand U1898 (N_1898,N_483,N_951);
nand U1899 (N_1899,N_844,N_611);
or U1900 (N_1900,N_998,N_865);
xor U1901 (N_1901,N_487,N_911);
and U1902 (N_1902,N_986,N_509);
nand U1903 (N_1903,N_75,N_466);
or U1904 (N_1904,N_643,N_10);
and U1905 (N_1905,N_90,N_139);
and U1906 (N_1906,N_451,N_418);
and U1907 (N_1907,N_279,N_516);
or U1908 (N_1908,N_878,N_417);
nand U1909 (N_1909,N_442,N_278);
or U1910 (N_1910,N_890,N_552);
nor U1911 (N_1911,N_506,N_492);
and U1912 (N_1912,N_299,N_51);
or U1913 (N_1913,N_758,N_998);
nand U1914 (N_1914,N_155,N_240);
nand U1915 (N_1915,N_344,N_463);
nand U1916 (N_1916,N_888,N_68);
or U1917 (N_1917,N_348,N_709);
and U1918 (N_1918,N_325,N_40);
nand U1919 (N_1919,N_501,N_836);
or U1920 (N_1920,N_263,N_453);
and U1921 (N_1921,N_50,N_867);
nand U1922 (N_1922,N_931,N_619);
or U1923 (N_1923,N_810,N_110);
or U1924 (N_1924,N_221,N_389);
nand U1925 (N_1925,N_80,N_541);
nor U1926 (N_1926,N_620,N_817);
nand U1927 (N_1927,N_154,N_855);
or U1928 (N_1928,N_374,N_285);
nand U1929 (N_1929,N_649,N_358);
or U1930 (N_1930,N_377,N_103);
nand U1931 (N_1931,N_530,N_40);
and U1932 (N_1932,N_726,N_588);
and U1933 (N_1933,N_936,N_484);
and U1934 (N_1934,N_984,N_112);
xor U1935 (N_1935,N_289,N_3);
and U1936 (N_1936,N_579,N_903);
and U1937 (N_1937,N_67,N_338);
and U1938 (N_1938,N_572,N_597);
xnor U1939 (N_1939,N_399,N_438);
or U1940 (N_1940,N_501,N_885);
xor U1941 (N_1941,N_244,N_202);
and U1942 (N_1942,N_738,N_257);
nor U1943 (N_1943,N_256,N_125);
xnor U1944 (N_1944,N_599,N_608);
or U1945 (N_1945,N_540,N_124);
nand U1946 (N_1946,N_817,N_982);
nand U1947 (N_1947,N_631,N_968);
or U1948 (N_1948,N_551,N_439);
and U1949 (N_1949,N_933,N_314);
or U1950 (N_1950,N_89,N_927);
or U1951 (N_1951,N_883,N_125);
nor U1952 (N_1952,N_440,N_124);
nor U1953 (N_1953,N_516,N_445);
and U1954 (N_1954,N_765,N_717);
nor U1955 (N_1955,N_948,N_422);
and U1956 (N_1956,N_615,N_368);
or U1957 (N_1957,N_316,N_541);
nand U1958 (N_1958,N_762,N_248);
nand U1959 (N_1959,N_64,N_278);
and U1960 (N_1960,N_415,N_103);
nor U1961 (N_1961,N_162,N_694);
or U1962 (N_1962,N_957,N_358);
xor U1963 (N_1963,N_517,N_399);
nand U1964 (N_1964,N_964,N_495);
nand U1965 (N_1965,N_261,N_438);
nor U1966 (N_1966,N_318,N_187);
nor U1967 (N_1967,N_870,N_95);
and U1968 (N_1968,N_719,N_224);
or U1969 (N_1969,N_528,N_997);
or U1970 (N_1970,N_751,N_146);
and U1971 (N_1971,N_224,N_810);
and U1972 (N_1972,N_414,N_310);
or U1973 (N_1973,N_728,N_865);
nor U1974 (N_1974,N_924,N_499);
xnor U1975 (N_1975,N_208,N_849);
and U1976 (N_1976,N_484,N_124);
nand U1977 (N_1977,N_869,N_378);
nand U1978 (N_1978,N_169,N_148);
xor U1979 (N_1979,N_158,N_754);
nor U1980 (N_1980,N_890,N_353);
nand U1981 (N_1981,N_427,N_567);
nand U1982 (N_1982,N_725,N_703);
or U1983 (N_1983,N_769,N_217);
or U1984 (N_1984,N_543,N_155);
and U1985 (N_1985,N_474,N_989);
or U1986 (N_1986,N_42,N_432);
and U1987 (N_1987,N_149,N_858);
xnor U1988 (N_1988,N_371,N_396);
and U1989 (N_1989,N_730,N_639);
or U1990 (N_1990,N_614,N_842);
xor U1991 (N_1991,N_558,N_754);
nand U1992 (N_1992,N_685,N_203);
nand U1993 (N_1993,N_69,N_488);
nand U1994 (N_1994,N_822,N_416);
nand U1995 (N_1995,N_849,N_361);
and U1996 (N_1996,N_899,N_280);
and U1997 (N_1997,N_654,N_275);
or U1998 (N_1998,N_311,N_775);
and U1999 (N_1999,N_968,N_246);
and U2000 (N_2000,N_1579,N_1289);
and U2001 (N_2001,N_1799,N_1550);
and U2002 (N_2002,N_1998,N_1153);
nor U2003 (N_2003,N_1232,N_1065);
or U2004 (N_2004,N_1192,N_1657);
nor U2005 (N_2005,N_1880,N_1202);
or U2006 (N_2006,N_1188,N_1593);
xor U2007 (N_2007,N_1312,N_1043);
nand U2008 (N_2008,N_1166,N_1104);
nand U2009 (N_2009,N_1221,N_1546);
nor U2010 (N_2010,N_1840,N_1870);
nand U2011 (N_2011,N_1989,N_1055);
nand U2012 (N_2012,N_1162,N_1747);
and U2013 (N_2013,N_1673,N_1950);
or U2014 (N_2014,N_1234,N_1525);
and U2015 (N_2015,N_1246,N_1150);
nand U2016 (N_2016,N_1122,N_1767);
nor U2017 (N_2017,N_1855,N_1013);
nand U2018 (N_2018,N_1488,N_1031);
nand U2019 (N_2019,N_1968,N_1597);
or U2020 (N_2020,N_1443,N_1270);
nor U2021 (N_2021,N_1596,N_1844);
nand U2022 (N_2022,N_1372,N_1274);
xnor U2023 (N_2023,N_1460,N_1308);
and U2024 (N_2024,N_1155,N_1782);
and U2025 (N_2025,N_1002,N_1029);
xor U2026 (N_2026,N_1563,N_1207);
or U2027 (N_2027,N_1867,N_1336);
nor U2028 (N_2028,N_1101,N_1120);
and U2029 (N_2029,N_1824,N_1461);
or U2030 (N_2030,N_1536,N_1981);
or U2031 (N_2031,N_1740,N_1046);
nor U2032 (N_2032,N_1904,N_1821);
and U2033 (N_2033,N_1204,N_1247);
nand U2034 (N_2034,N_1718,N_1353);
nor U2035 (N_2035,N_1023,N_1455);
and U2036 (N_2036,N_1032,N_1492);
and U2037 (N_2037,N_1709,N_1705);
or U2038 (N_2038,N_1068,N_1377);
xnor U2039 (N_2039,N_1351,N_1267);
or U2040 (N_2040,N_1158,N_1343);
nor U2041 (N_2041,N_1766,N_1292);
and U2042 (N_2042,N_1729,N_1807);
nand U2043 (N_2043,N_1639,N_1746);
nor U2044 (N_2044,N_1518,N_1070);
nor U2045 (N_2045,N_1708,N_1058);
or U2046 (N_2046,N_1344,N_1466);
nor U2047 (N_2047,N_1285,N_1277);
and U2048 (N_2048,N_1215,N_1745);
nand U2049 (N_2049,N_1589,N_1795);
nor U2050 (N_2050,N_1739,N_1364);
and U2051 (N_2051,N_1811,N_1973);
or U2052 (N_2052,N_1763,N_1691);
nor U2053 (N_2053,N_1303,N_1540);
or U2054 (N_2054,N_1385,N_1863);
nor U2055 (N_2055,N_1912,N_1113);
nor U2056 (N_2056,N_1637,N_1809);
and U2057 (N_2057,N_1846,N_1642);
and U2058 (N_2058,N_1400,N_1357);
xor U2059 (N_2059,N_1626,N_1131);
and U2060 (N_2060,N_1045,N_1059);
nor U2061 (N_2061,N_1648,N_1940);
nand U2062 (N_2062,N_1585,N_1420);
nand U2063 (N_2063,N_1792,N_1905);
and U2064 (N_2064,N_1275,N_1810);
nand U2065 (N_2065,N_1520,N_1230);
or U2066 (N_2066,N_1114,N_1895);
nor U2067 (N_2067,N_1581,N_1759);
xor U2068 (N_2068,N_1765,N_1095);
and U2069 (N_2069,N_1697,N_1146);
or U2070 (N_2070,N_1110,N_1618);
or U2071 (N_2071,N_1926,N_1298);
and U2072 (N_2072,N_1318,N_1812);
and U2073 (N_2073,N_1768,N_1568);
and U2074 (N_2074,N_1373,N_1435);
and U2075 (N_2075,N_1238,N_1136);
nor U2076 (N_2076,N_1554,N_1872);
nand U2077 (N_2077,N_1814,N_1719);
or U2078 (N_2078,N_1877,N_1080);
xor U2079 (N_2079,N_1201,N_1873);
nor U2080 (N_2080,N_1272,N_1409);
nor U2081 (N_2081,N_1199,N_1701);
and U2082 (N_2082,N_1044,N_1832);
xnor U2083 (N_2083,N_1355,N_1086);
nor U2084 (N_2084,N_1493,N_1082);
nand U2085 (N_2085,N_1995,N_1137);
and U2086 (N_2086,N_1220,N_1035);
nor U2087 (N_2087,N_1416,N_1943);
nor U2088 (N_2088,N_1026,N_1311);
xnor U2089 (N_2089,N_1963,N_1453);
nand U2090 (N_2090,N_1576,N_1197);
nand U2091 (N_2091,N_1392,N_1572);
or U2092 (N_2092,N_1301,N_1389);
or U2093 (N_2093,N_1452,N_1957);
or U2094 (N_2094,N_1669,N_1454);
nand U2095 (N_2095,N_1564,N_1128);
nand U2096 (N_2096,N_1027,N_1854);
nor U2097 (N_2097,N_1674,N_1501);
nor U2098 (N_2098,N_1240,N_1291);
and U2099 (N_2099,N_1864,N_1819);
nor U2100 (N_2100,N_1874,N_1297);
nand U2101 (N_2101,N_1347,N_1015);
and U2102 (N_2102,N_1481,N_1789);
and U2103 (N_2103,N_1670,N_1426);
nand U2104 (N_2104,N_1735,N_1195);
or U2105 (N_2105,N_1219,N_1555);
xnor U2106 (N_2106,N_1052,N_1316);
or U2107 (N_2107,N_1173,N_1030);
nand U2108 (N_2108,N_1259,N_1667);
nand U2109 (N_2109,N_1714,N_1099);
nand U2110 (N_2110,N_1093,N_1020);
nor U2111 (N_2111,N_1974,N_1494);
and U2112 (N_2112,N_1817,N_1092);
or U2113 (N_2113,N_1793,N_1543);
nand U2114 (N_2114,N_1914,N_1006);
or U2115 (N_2115,N_1764,N_1894);
nand U2116 (N_2116,N_1279,N_1898);
nand U2117 (N_2117,N_1041,N_1539);
and U2118 (N_2118,N_1360,N_1982);
and U2119 (N_2119,N_1504,N_1791);
or U2120 (N_2120,N_1323,N_1081);
nor U2121 (N_2121,N_1375,N_1008);
nand U2122 (N_2122,N_1242,N_1861);
nor U2123 (N_2123,N_1731,N_1076);
nor U2124 (N_2124,N_1510,N_1482);
nand U2125 (N_2125,N_1439,N_1251);
nand U2126 (N_2126,N_1775,N_1448);
nor U2127 (N_2127,N_1848,N_1176);
nand U2128 (N_2128,N_1147,N_1630);
nor U2129 (N_2129,N_1613,N_1690);
nand U2130 (N_2130,N_1953,N_1395);
and U2131 (N_2131,N_1037,N_1227);
nor U2132 (N_2132,N_1515,N_1533);
or U2133 (N_2133,N_1498,N_1975);
and U2134 (N_2134,N_1988,N_1784);
or U2135 (N_2135,N_1712,N_1605);
nand U2136 (N_2136,N_1748,N_1915);
or U2137 (N_2137,N_1551,N_1217);
or U2138 (N_2138,N_1643,N_1154);
xnor U2139 (N_2139,N_1228,N_1529);
or U2140 (N_2140,N_1567,N_1857);
nand U2141 (N_2141,N_1858,N_1899);
or U2142 (N_2142,N_1485,N_1004);
nand U2143 (N_2143,N_1646,N_1370);
nand U2144 (N_2144,N_1206,N_1315);
nor U2145 (N_2145,N_1437,N_1334);
and U2146 (N_2146,N_1946,N_1557);
nand U2147 (N_2147,N_1066,N_1189);
xnor U2148 (N_2148,N_1332,N_1139);
and U2149 (N_2149,N_1363,N_1813);
nor U2150 (N_2150,N_1619,N_1060);
nor U2151 (N_2151,N_1777,N_1036);
or U2152 (N_2152,N_1650,N_1786);
nand U2153 (N_2153,N_1394,N_1773);
and U2154 (N_2154,N_1964,N_1440);
and U2155 (N_2155,N_1842,N_1129);
or U2156 (N_2156,N_1598,N_1752);
nand U2157 (N_2157,N_1205,N_1888);
nand U2158 (N_2158,N_1398,N_1329);
or U2159 (N_2159,N_1921,N_1404);
or U2160 (N_2160,N_1505,N_1829);
or U2161 (N_2161,N_1871,N_1760);
or U2162 (N_2162,N_1959,N_1361);
nand U2163 (N_2163,N_1951,N_1330);
nor U2164 (N_2164,N_1127,N_1732);
nor U2165 (N_2165,N_1530,N_1063);
and U2166 (N_2166,N_1552,N_1226);
nand U2167 (N_2167,N_1157,N_1427);
nor U2168 (N_2168,N_1256,N_1999);
and U2169 (N_2169,N_1417,N_1487);
and U2170 (N_2170,N_1790,N_1491);
and U2171 (N_2171,N_1341,N_1756);
or U2172 (N_2172,N_1457,N_1947);
and U2173 (N_2173,N_1741,N_1933);
xnor U2174 (N_2174,N_1293,N_1273);
and U2175 (N_2175,N_1475,N_1314);
nor U2176 (N_2176,N_1098,N_1660);
nand U2177 (N_2177,N_1352,N_1879);
or U2178 (N_2178,N_1604,N_1423);
or U2179 (N_2179,N_1366,N_1796);
nor U2180 (N_2180,N_1997,N_1362);
nand U2181 (N_2181,N_1901,N_1700);
nor U2182 (N_2182,N_1930,N_1755);
or U2183 (N_2183,N_1507,N_1378);
and U2184 (N_2184,N_1024,N_1499);
and U2185 (N_2185,N_1566,N_1354);
and U2186 (N_2186,N_1213,N_1662);
and U2187 (N_2187,N_1727,N_1265);
xor U2188 (N_2188,N_1818,N_1069);
nor U2189 (N_2189,N_1209,N_1614);
nor U2190 (N_2190,N_1680,N_1382);
or U2191 (N_2191,N_1805,N_1252);
and U2192 (N_2192,N_1218,N_1838);
and U2193 (N_2193,N_1853,N_1028);
xnor U2194 (N_2194,N_1428,N_1433);
nor U2195 (N_2195,N_1236,N_1991);
xor U2196 (N_2196,N_1283,N_1050);
nor U2197 (N_2197,N_1235,N_1806);
nor U2198 (N_2198,N_1606,N_1387);
or U2199 (N_2199,N_1284,N_1627);
nand U2200 (N_2200,N_1526,N_1359);
or U2201 (N_2201,N_1112,N_1425);
and U2202 (N_2202,N_1422,N_1469);
nor U2203 (N_2203,N_1725,N_1911);
nor U2204 (N_2204,N_1135,N_1983);
xor U2205 (N_2205,N_1307,N_1609);
and U2206 (N_2206,N_1115,N_1304);
nor U2207 (N_2207,N_1671,N_1945);
nor U2208 (N_2208,N_1480,N_1445);
nand U2209 (N_2209,N_1118,N_1734);
or U2210 (N_2210,N_1502,N_1056);
nand U2211 (N_2211,N_1278,N_1094);
and U2212 (N_2212,N_1358,N_1726);
nand U2213 (N_2213,N_1021,N_1703);
or U2214 (N_2214,N_1684,N_1184);
xnor U2215 (N_2215,N_1165,N_1241);
xnor U2216 (N_2216,N_1477,N_1584);
or U2217 (N_2217,N_1776,N_1621);
nor U2218 (N_2218,N_1418,N_1411);
nor U2219 (N_2219,N_1152,N_1509);
nand U2220 (N_2220,N_1191,N_1414);
xor U2221 (N_2221,N_1084,N_1682);
or U2222 (N_2222,N_1441,N_1778);
nand U2223 (N_2223,N_1010,N_1716);
xor U2224 (N_2224,N_1990,N_1723);
or U2225 (N_2225,N_1062,N_1996);
or U2226 (N_2226,N_1048,N_1808);
and U2227 (N_2227,N_1771,N_1512);
nor U2228 (N_2228,N_1071,N_1223);
nor U2229 (N_2229,N_1229,N_1722);
or U2230 (N_2230,N_1476,N_1847);
nor U2231 (N_2231,N_1449,N_1560);
nand U2232 (N_2232,N_1276,N_1845);
nor U2233 (N_2233,N_1587,N_1841);
or U2234 (N_2234,N_1761,N_1144);
and U2235 (N_2235,N_1908,N_1051);
xnor U2236 (N_2236,N_1750,N_1622);
and U2237 (N_2237,N_1875,N_1710);
and U2238 (N_2238,N_1194,N_1590);
nand U2239 (N_2239,N_1169,N_1280);
nand U2240 (N_2240,N_1713,N_1887);
nor U2241 (N_2241,N_1936,N_1390);
and U2242 (N_2242,N_1295,N_1683);
nand U2243 (N_2243,N_1299,N_1478);
and U2244 (N_2244,N_1583,N_1625);
nor U2245 (N_2245,N_1876,N_1090);
xnor U2246 (N_2246,N_1751,N_1016);
or U2247 (N_2247,N_1233,N_1769);
nand U2248 (N_2248,N_1571,N_1346);
or U2249 (N_2249,N_1126,N_1672);
nand U2250 (N_2250,N_1985,N_1405);
or U2251 (N_2251,N_1506,N_1349);
and U2252 (N_2252,N_1788,N_1151);
nor U2253 (N_2253,N_1954,N_1290);
and U2254 (N_2254,N_1500,N_1214);
or U2255 (N_2255,N_1117,N_1248);
or U2256 (N_2256,N_1816,N_1025);
xor U2257 (N_2257,N_1827,N_1629);
and U2258 (N_2258,N_1203,N_1286);
nand U2259 (N_2259,N_1388,N_1730);
or U2260 (N_2260,N_1497,N_1900);
and U2261 (N_2261,N_1631,N_1532);
xor U2262 (N_2262,N_1687,N_1800);
nand U2263 (N_2263,N_1326,N_1869);
nor U2264 (N_2264,N_1456,N_1595);
or U2265 (N_2265,N_1486,N_1091);
and U2266 (N_2266,N_1224,N_1211);
nor U2267 (N_2267,N_1379,N_1038);
nand U2268 (N_2268,N_1922,N_1801);
xor U2269 (N_2269,N_1431,N_1143);
and U2270 (N_2270,N_1849,N_1075);
nand U2271 (N_2271,N_1941,N_1715);
or U2272 (N_2272,N_1823,N_1770);
nand U2273 (N_2273,N_1462,N_1891);
nand U2274 (N_2274,N_1432,N_1496);
and U2275 (N_2275,N_1340,N_1434);
xnor U2276 (N_2276,N_1017,N_1685);
nor U2277 (N_2277,N_1369,N_1815);
and U2278 (N_2278,N_1067,N_1545);
or U2279 (N_2279,N_1257,N_1464);
and U2280 (N_2280,N_1072,N_1706);
nand U2281 (N_2281,N_1516,N_1742);
nand U2282 (N_2282,N_1935,N_1885);
nand U2283 (N_2283,N_1222,N_1012);
or U2284 (N_2284,N_1523,N_1266);
xor U2285 (N_2285,N_1960,N_1696);
and U2286 (N_2286,N_1707,N_1702);
xor U2287 (N_2287,N_1612,N_1061);
and U2288 (N_2288,N_1651,N_1883);
nand U2289 (N_2289,N_1663,N_1649);
or U2290 (N_2290,N_1079,N_1603);
xor U2291 (N_2291,N_1961,N_1172);
and U2292 (N_2292,N_1243,N_1635);
and U2293 (N_2293,N_1163,N_1264);
nor U2294 (N_2294,N_1294,N_1822);
and U2295 (N_2295,N_1843,N_1837);
nand U2296 (N_2296,N_1890,N_1100);
and U2297 (N_2297,N_1738,N_1728);
and U2298 (N_2298,N_1049,N_1802);
and U2299 (N_2299,N_1820,N_1513);
nand U2300 (N_2300,N_1878,N_1231);
or U2301 (N_2301,N_1190,N_1178);
xor U2302 (N_2302,N_1884,N_1397);
nand U2303 (N_2303,N_1288,N_1889);
and U2304 (N_2304,N_1446,N_1720);
and U2305 (N_2305,N_1000,N_1447);
and U2306 (N_2306,N_1830,N_1956);
and U2307 (N_2307,N_1949,N_1893);
nand U2308 (N_2308,N_1666,N_1468);
nand U2309 (N_2309,N_1521,N_1296);
nand U2310 (N_2310,N_1653,N_1383);
and U2311 (N_2311,N_1556,N_1969);
nor U2312 (N_2312,N_1535,N_1503);
or U2313 (N_2313,N_1133,N_1850);
or U2314 (N_2314,N_1438,N_1164);
or U2315 (N_2315,N_1979,N_1717);
and U2316 (N_2316,N_1785,N_1967);
or U2317 (N_2317,N_1421,N_1313);
nor U2318 (N_2318,N_1125,N_1356);
and U2319 (N_2319,N_1575,N_1675);
nand U2320 (N_2320,N_1966,N_1106);
and U2321 (N_2321,N_1976,N_1862);
and U2322 (N_2322,N_1401,N_1328);
nor U2323 (N_2323,N_1287,N_1001);
or U2324 (N_2324,N_1470,N_1138);
nor U2325 (N_2325,N_1721,N_1955);
or U2326 (N_2326,N_1616,N_1774);
and U2327 (N_2327,N_1465,N_1054);
nand U2328 (N_2328,N_1569,N_1319);
nand U2329 (N_2329,N_1402,N_1711);
nor U2330 (N_2330,N_1342,N_1263);
nand U2331 (N_2331,N_1828,N_1928);
nor U2332 (N_2332,N_1519,N_1327);
nor U2333 (N_2333,N_1524,N_1306);
nand U2334 (N_2334,N_1656,N_1170);
nand U2335 (N_2335,N_1317,N_1534);
nor U2336 (N_2336,N_1537,N_1833);
and U2337 (N_2337,N_1255,N_1085);
nor U2338 (N_2338,N_1910,N_1570);
xor U2339 (N_2339,N_1305,N_1261);
nand U2340 (N_2340,N_1177,N_1182);
nand U2341 (N_2341,N_1856,N_1365);
nand U2342 (N_2342,N_1577,N_1559);
nand U2343 (N_2343,N_1473,N_1187);
and U2344 (N_2344,N_1632,N_1958);
nor U2345 (N_2345,N_1130,N_1664);
xnor U2346 (N_2346,N_1033,N_1436);
and U2347 (N_2347,N_1262,N_1097);
and U2348 (N_2348,N_1757,N_1514);
or U2349 (N_2349,N_1628,N_1088);
nor U2350 (N_2350,N_1479,N_1271);
and U2351 (N_2351,N_1798,N_1624);
and U2352 (N_2352,N_1978,N_1574);
nor U2353 (N_2353,N_1733,N_1918);
nand U2354 (N_2354,N_1923,N_1210);
nor U2355 (N_2355,N_1167,N_1665);
and U2356 (N_2356,N_1804,N_1580);
nand U2357 (N_2357,N_1623,N_1548);
nor U2358 (N_2358,N_1860,N_1474);
or U2359 (N_2359,N_1407,N_1645);
nand U2360 (N_2360,N_1859,N_1986);
nor U2361 (N_2361,N_1924,N_1932);
nor U2362 (N_2362,N_1089,N_1348);
nand U2363 (N_2363,N_1934,N_1371);
xnor U2364 (N_2364,N_1018,N_1592);
and U2365 (N_2365,N_1927,N_1198);
xor U2366 (N_2366,N_1588,N_1429);
or U2367 (N_2367,N_1600,N_1825);
or U2368 (N_2368,N_1471,N_1483);
nor U2369 (N_2369,N_1057,N_1331);
nand U2370 (N_2370,N_1109,N_1517);
nand U2371 (N_2371,N_1522,N_1148);
nand U2372 (N_2372,N_1410,N_1542);
xnor U2373 (N_2373,N_1450,N_1931);
or U2374 (N_2374,N_1852,N_1042);
nand U2375 (N_2375,N_1064,N_1909);
nand U2376 (N_2376,N_1458,N_1607);
nand U2377 (N_2377,N_1938,N_1463);
nor U2378 (N_2378,N_1972,N_1495);
xnor U2379 (N_2379,N_1123,N_1345);
nor U2380 (N_2380,N_1538,N_1881);
or U2381 (N_2381,N_1424,N_1391);
nand U2382 (N_2382,N_1942,N_1302);
nand U2383 (N_2383,N_1678,N_1337);
and U2384 (N_2384,N_1868,N_1142);
nand U2385 (N_2385,N_1467,N_1965);
and U2386 (N_2386,N_1937,N_1237);
or U2387 (N_2387,N_1459,N_1962);
nor U2388 (N_2388,N_1269,N_1834);
or U2389 (N_2389,N_1300,N_1386);
or U2390 (N_2390,N_1594,N_1260);
xor U2391 (N_2391,N_1661,N_1381);
or U2392 (N_2392,N_1333,N_1339);
nor U2393 (N_2393,N_1781,N_1971);
xnor U2394 (N_2394,N_1655,N_1633);
nand U2395 (N_2395,N_1641,N_1107);
nand U2396 (N_2396,N_1039,N_1758);
nand U2397 (N_2397,N_1249,N_1212);
nand U2398 (N_2398,N_1014,N_1586);
or U2399 (N_2399,N_1254,N_1040);
and U2400 (N_2400,N_1698,N_1886);
and U2401 (N_2401,N_1121,N_1620);
nor U2402 (N_2402,N_1797,N_1073);
and U2403 (N_2403,N_1906,N_1749);
and U2404 (N_2404,N_1321,N_1693);
nor U2405 (N_2405,N_1022,N_1737);
or U2406 (N_2406,N_1980,N_1490);
and U2407 (N_2407,N_1694,N_1528);
or U2408 (N_2408,N_1772,N_1527);
nor U2409 (N_2409,N_1511,N_1689);
or U2410 (N_2410,N_1408,N_1245);
nor U2411 (N_2411,N_1994,N_1156);
nor U2412 (N_2412,N_1601,N_1181);
nor U2413 (N_2413,N_1826,N_1179);
or U2414 (N_2414,N_1688,N_1145);
xnor U2415 (N_2415,N_1987,N_1952);
xnor U2416 (N_2416,N_1335,N_1610);
and U2417 (N_2417,N_1406,N_1917);
nor U2418 (N_2418,N_1896,N_1562);
nor U2419 (N_2419,N_1677,N_1944);
nand U2420 (N_2420,N_1116,N_1380);
nand U2421 (N_2421,N_1268,N_1892);
nor U2422 (N_2422,N_1047,N_1686);
nand U2423 (N_2423,N_1149,N_1216);
nor U2424 (N_2424,N_1108,N_1704);
and U2425 (N_2425,N_1168,N_1103);
or U2426 (N_2426,N_1558,N_1376);
and U2427 (N_2427,N_1134,N_1430);
nor U2428 (N_2428,N_1668,N_1310);
nor U2429 (N_2429,N_1743,N_1374);
nor U2430 (N_2430,N_1615,N_1882);
and U2431 (N_2431,N_1367,N_1929);
nor U2432 (N_2432,N_1925,N_1442);
and U2433 (N_2433,N_1865,N_1762);
nand U2434 (N_2434,N_1992,N_1561);
nand U2435 (N_2435,N_1659,N_1654);
nand U2436 (N_2436,N_1083,N_1508);
nor U2437 (N_2437,N_1403,N_1907);
nor U2438 (N_2438,N_1591,N_1602);
and U2439 (N_2439,N_1578,N_1611);
or U2440 (N_2440,N_1866,N_1320);
and U2441 (N_2441,N_1250,N_1444);
and U2442 (N_2442,N_1258,N_1325);
and U2443 (N_2443,N_1180,N_1282);
and U2444 (N_2444,N_1019,N_1489);
and U2445 (N_2445,N_1077,N_1984);
xor U2446 (N_2446,N_1413,N_1836);
nor U2447 (N_2447,N_1553,N_1903);
nor U2448 (N_2448,N_1699,N_1787);
or U2449 (N_2449,N_1599,N_1281);
nand U2450 (N_2450,N_1053,N_1253);
and U2451 (N_2451,N_1183,N_1636);
nand U2452 (N_2452,N_1412,N_1652);
nor U2453 (N_2453,N_1225,N_1839);
and U2454 (N_2454,N_1644,N_1547);
nor U2455 (N_2455,N_1851,N_1124);
nor U2456 (N_2456,N_1384,N_1679);
or U2457 (N_2457,N_1753,N_1913);
and U2458 (N_2458,N_1658,N_1119);
or U2459 (N_2459,N_1074,N_1140);
and U2460 (N_2460,N_1803,N_1920);
nand U2461 (N_2461,N_1640,N_1565);
nor U2462 (N_2462,N_1780,N_1175);
xnor U2463 (N_2463,N_1835,N_1159);
nor U2464 (N_2464,N_1368,N_1695);
and U2465 (N_2465,N_1132,N_1977);
nand U2466 (N_2466,N_1034,N_1322);
xor U2467 (N_2467,N_1309,N_1902);
and U2468 (N_2468,N_1003,N_1007);
nor U2469 (N_2469,N_1174,N_1239);
nand U2470 (N_2470,N_1111,N_1171);
nand U2471 (N_2471,N_1638,N_1744);
xnor U2472 (N_2472,N_1608,N_1993);
xnor U2473 (N_2473,N_1919,N_1338);
xnor U2474 (N_2474,N_1970,N_1185);
nand U2475 (N_2475,N_1009,N_1415);
and U2476 (N_2476,N_1005,N_1939);
nand U2477 (N_2477,N_1484,N_1102);
nor U2478 (N_2478,N_1573,N_1779);
nor U2479 (N_2479,N_1647,N_1324);
nand U2480 (N_2480,N_1676,N_1549);
or U2481 (N_2481,N_1350,N_1897);
nand U2482 (N_2482,N_1916,N_1200);
and U2483 (N_2483,N_1161,N_1736);
nand U2484 (N_2484,N_1419,N_1196);
nand U2485 (N_2485,N_1105,N_1244);
or U2486 (N_2486,N_1160,N_1754);
xnor U2487 (N_2487,N_1096,N_1724);
or U2488 (N_2488,N_1541,N_1472);
nand U2489 (N_2489,N_1399,N_1393);
and U2490 (N_2490,N_1831,N_1078);
or U2491 (N_2491,N_1208,N_1617);
or U2492 (N_2492,N_1634,N_1011);
nand U2493 (N_2493,N_1794,N_1186);
xor U2494 (N_2494,N_1692,N_1681);
xor U2495 (N_2495,N_1141,N_1396);
or U2496 (N_2496,N_1783,N_1193);
and U2497 (N_2497,N_1582,N_1544);
or U2498 (N_2498,N_1948,N_1087);
and U2499 (N_2499,N_1451,N_1531);
or U2500 (N_2500,N_1242,N_1839);
and U2501 (N_2501,N_1073,N_1796);
nand U2502 (N_2502,N_1627,N_1756);
nor U2503 (N_2503,N_1161,N_1073);
and U2504 (N_2504,N_1484,N_1788);
nand U2505 (N_2505,N_1112,N_1293);
or U2506 (N_2506,N_1229,N_1483);
nor U2507 (N_2507,N_1780,N_1711);
and U2508 (N_2508,N_1800,N_1216);
and U2509 (N_2509,N_1424,N_1943);
and U2510 (N_2510,N_1396,N_1945);
and U2511 (N_2511,N_1531,N_1694);
or U2512 (N_2512,N_1626,N_1429);
nand U2513 (N_2513,N_1044,N_1084);
xnor U2514 (N_2514,N_1859,N_1528);
or U2515 (N_2515,N_1758,N_1121);
and U2516 (N_2516,N_1801,N_1513);
or U2517 (N_2517,N_1943,N_1811);
or U2518 (N_2518,N_1205,N_1925);
nor U2519 (N_2519,N_1078,N_1412);
xor U2520 (N_2520,N_1535,N_1540);
and U2521 (N_2521,N_1426,N_1269);
or U2522 (N_2522,N_1133,N_1294);
or U2523 (N_2523,N_1596,N_1258);
nand U2524 (N_2524,N_1163,N_1448);
nor U2525 (N_2525,N_1142,N_1726);
nand U2526 (N_2526,N_1676,N_1689);
xnor U2527 (N_2527,N_1533,N_1403);
nand U2528 (N_2528,N_1629,N_1775);
and U2529 (N_2529,N_1596,N_1392);
nand U2530 (N_2530,N_1580,N_1172);
nand U2531 (N_2531,N_1470,N_1480);
and U2532 (N_2532,N_1259,N_1000);
nor U2533 (N_2533,N_1747,N_1095);
nand U2534 (N_2534,N_1384,N_1587);
and U2535 (N_2535,N_1264,N_1241);
or U2536 (N_2536,N_1712,N_1576);
nor U2537 (N_2537,N_1133,N_1374);
or U2538 (N_2538,N_1771,N_1280);
nand U2539 (N_2539,N_1192,N_1151);
nor U2540 (N_2540,N_1044,N_1778);
nand U2541 (N_2541,N_1243,N_1432);
nand U2542 (N_2542,N_1466,N_1529);
xor U2543 (N_2543,N_1368,N_1737);
or U2544 (N_2544,N_1458,N_1112);
or U2545 (N_2545,N_1784,N_1610);
nand U2546 (N_2546,N_1702,N_1274);
nor U2547 (N_2547,N_1011,N_1418);
nand U2548 (N_2548,N_1536,N_1613);
nor U2549 (N_2549,N_1297,N_1726);
and U2550 (N_2550,N_1662,N_1730);
and U2551 (N_2551,N_1582,N_1100);
nand U2552 (N_2552,N_1176,N_1610);
nor U2553 (N_2553,N_1227,N_1767);
or U2554 (N_2554,N_1261,N_1369);
and U2555 (N_2555,N_1491,N_1455);
nand U2556 (N_2556,N_1742,N_1869);
and U2557 (N_2557,N_1704,N_1828);
nor U2558 (N_2558,N_1815,N_1069);
or U2559 (N_2559,N_1073,N_1401);
nor U2560 (N_2560,N_1730,N_1887);
nor U2561 (N_2561,N_1228,N_1288);
or U2562 (N_2562,N_1454,N_1599);
nand U2563 (N_2563,N_1100,N_1748);
nand U2564 (N_2564,N_1046,N_1192);
and U2565 (N_2565,N_1908,N_1829);
or U2566 (N_2566,N_1066,N_1999);
and U2567 (N_2567,N_1069,N_1678);
nand U2568 (N_2568,N_1547,N_1134);
and U2569 (N_2569,N_1519,N_1366);
nor U2570 (N_2570,N_1970,N_1361);
and U2571 (N_2571,N_1404,N_1432);
xnor U2572 (N_2572,N_1059,N_1103);
and U2573 (N_2573,N_1584,N_1924);
and U2574 (N_2574,N_1185,N_1475);
or U2575 (N_2575,N_1510,N_1642);
nor U2576 (N_2576,N_1358,N_1326);
nor U2577 (N_2577,N_1219,N_1753);
nor U2578 (N_2578,N_1371,N_1202);
nand U2579 (N_2579,N_1509,N_1903);
nor U2580 (N_2580,N_1805,N_1380);
and U2581 (N_2581,N_1089,N_1510);
xnor U2582 (N_2582,N_1596,N_1414);
nand U2583 (N_2583,N_1454,N_1135);
nor U2584 (N_2584,N_1767,N_1163);
nor U2585 (N_2585,N_1641,N_1395);
and U2586 (N_2586,N_1458,N_1117);
nor U2587 (N_2587,N_1623,N_1533);
and U2588 (N_2588,N_1750,N_1379);
and U2589 (N_2589,N_1737,N_1665);
nand U2590 (N_2590,N_1456,N_1550);
nor U2591 (N_2591,N_1559,N_1015);
or U2592 (N_2592,N_1014,N_1146);
or U2593 (N_2593,N_1616,N_1910);
nor U2594 (N_2594,N_1403,N_1008);
nand U2595 (N_2595,N_1398,N_1033);
and U2596 (N_2596,N_1054,N_1955);
nand U2597 (N_2597,N_1870,N_1543);
or U2598 (N_2598,N_1104,N_1940);
and U2599 (N_2599,N_1647,N_1445);
xor U2600 (N_2600,N_1749,N_1293);
nand U2601 (N_2601,N_1926,N_1820);
or U2602 (N_2602,N_1556,N_1884);
nor U2603 (N_2603,N_1813,N_1859);
nand U2604 (N_2604,N_1539,N_1521);
or U2605 (N_2605,N_1575,N_1775);
and U2606 (N_2606,N_1938,N_1850);
nor U2607 (N_2607,N_1031,N_1041);
nor U2608 (N_2608,N_1979,N_1850);
or U2609 (N_2609,N_1308,N_1905);
nor U2610 (N_2610,N_1352,N_1966);
nor U2611 (N_2611,N_1388,N_1161);
or U2612 (N_2612,N_1104,N_1993);
xor U2613 (N_2613,N_1119,N_1028);
and U2614 (N_2614,N_1544,N_1352);
or U2615 (N_2615,N_1221,N_1857);
nor U2616 (N_2616,N_1737,N_1775);
or U2617 (N_2617,N_1646,N_1788);
nand U2618 (N_2618,N_1012,N_1958);
and U2619 (N_2619,N_1470,N_1656);
xnor U2620 (N_2620,N_1229,N_1936);
xnor U2621 (N_2621,N_1970,N_1229);
or U2622 (N_2622,N_1217,N_1017);
nand U2623 (N_2623,N_1899,N_1896);
or U2624 (N_2624,N_1207,N_1847);
nor U2625 (N_2625,N_1863,N_1315);
nor U2626 (N_2626,N_1797,N_1220);
nand U2627 (N_2627,N_1744,N_1441);
and U2628 (N_2628,N_1255,N_1399);
nand U2629 (N_2629,N_1443,N_1419);
nand U2630 (N_2630,N_1803,N_1092);
nand U2631 (N_2631,N_1268,N_1023);
and U2632 (N_2632,N_1508,N_1756);
nor U2633 (N_2633,N_1017,N_1912);
nor U2634 (N_2634,N_1755,N_1164);
nand U2635 (N_2635,N_1836,N_1332);
xor U2636 (N_2636,N_1697,N_1257);
nand U2637 (N_2637,N_1029,N_1193);
nor U2638 (N_2638,N_1749,N_1190);
or U2639 (N_2639,N_1629,N_1065);
nor U2640 (N_2640,N_1492,N_1625);
or U2641 (N_2641,N_1237,N_1117);
nand U2642 (N_2642,N_1260,N_1772);
xnor U2643 (N_2643,N_1871,N_1856);
and U2644 (N_2644,N_1585,N_1677);
nor U2645 (N_2645,N_1258,N_1132);
nand U2646 (N_2646,N_1093,N_1391);
nand U2647 (N_2647,N_1104,N_1382);
nor U2648 (N_2648,N_1884,N_1246);
and U2649 (N_2649,N_1153,N_1116);
and U2650 (N_2650,N_1241,N_1288);
and U2651 (N_2651,N_1311,N_1748);
xnor U2652 (N_2652,N_1938,N_1667);
nor U2653 (N_2653,N_1735,N_1592);
nor U2654 (N_2654,N_1768,N_1559);
or U2655 (N_2655,N_1853,N_1929);
nand U2656 (N_2656,N_1295,N_1589);
and U2657 (N_2657,N_1294,N_1337);
or U2658 (N_2658,N_1882,N_1819);
nor U2659 (N_2659,N_1314,N_1076);
nand U2660 (N_2660,N_1011,N_1329);
or U2661 (N_2661,N_1395,N_1557);
nand U2662 (N_2662,N_1068,N_1924);
or U2663 (N_2663,N_1589,N_1103);
and U2664 (N_2664,N_1494,N_1539);
nor U2665 (N_2665,N_1906,N_1828);
nand U2666 (N_2666,N_1238,N_1756);
or U2667 (N_2667,N_1563,N_1992);
xnor U2668 (N_2668,N_1542,N_1298);
xnor U2669 (N_2669,N_1073,N_1354);
xor U2670 (N_2670,N_1307,N_1469);
nand U2671 (N_2671,N_1215,N_1603);
xor U2672 (N_2672,N_1186,N_1586);
xnor U2673 (N_2673,N_1678,N_1781);
nor U2674 (N_2674,N_1408,N_1072);
or U2675 (N_2675,N_1674,N_1460);
nand U2676 (N_2676,N_1903,N_1951);
nor U2677 (N_2677,N_1539,N_1317);
or U2678 (N_2678,N_1386,N_1076);
nand U2679 (N_2679,N_1930,N_1671);
nor U2680 (N_2680,N_1689,N_1173);
and U2681 (N_2681,N_1708,N_1773);
and U2682 (N_2682,N_1981,N_1574);
nor U2683 (N_2683,N_1619,N_1794);
nor U2684 (N_2684,N_1613,N_1519);
and U2685 (N_2685,N_1856,N_1082);
and U2686 (N_2686,N_1409,N_1408);
nand U2687 (N_2687,N_1786,N_1192);
nand U2688 (N_2688,N_1715,N_1741);
nand U2689 (N_2689,N_1035,N_1123);
nand U2690 (N_2690,N_1019,N_1112);
nor U2691 (N_2691,N_1659,N_1502);
and U2692 (N_2692,N_1295,N_1108);
or U2693 (N_2693,N_1823,N_1349);
and U2694 (N_2694,N_1314,N_1960);
xor U2695 (N_2695,N_1634,N_1480);
and U2696 (N_2696,N_1699,N_1453);
nand U2697 (N_2697,N_1442,N_1333);
or U2698 (N_2698,N_1702,N_1415);
and U2699 (N_2699,N_1568,N_1360);
nor U2700 (N_2700,N_1500,N_1212);
and U2701 (N_2701,N_1513,N_1972);
and U2702 (N_2702,N_1845,N_1762);
or U2703 (N_2703,N_1735,N_1835);
xnor U2704 (N_2704,N_1358,N_1788);
or U2705 (N_2705,N_1931,N_1299);
and U2706 (N_2706,N_1689,N_1574);
and U2707 (N_2707,N_1236,N_1093);
nand U2708 (N_2708,N_1593,N_1189);
and U2709 (N_2709,N_1367,N_1645);
nor U2710 (N_2710,N_1517,N_1824);
or U2711 (N_2711,N_1115,N_1138);
nand U2712 (N_2712,N_1763,N_1702);
nor U2713 (N_2713,N_1101,N_1316);
nor U2714 (N_2714,N_1916,N_1804);
or U2715 (N_2715,N_1951,N_1843);
and U2716 (N_2716,N_1425,N_1952);
nand U2717 (N_2717,N_1328,N_1165);
or U2718 (N_2718,N_1437,N_1419);
nor U2719 (N_2719,N_1842,N_1550);
or U2720 (N_2720,N_1022,N_1612);
nor U2721 (N_2721,N_1624,N_1044);
nor U2722 (N_2722,N_1499,N_1250);
and U2723 (N_2723,N_1304,N_1152);
nand U2724 (N_2724,N_1451,N_1964);
xnor U2725 (N_2725,N_1125,N_1174);
nand U2726 (N_2726,N_1821,N_1388);
nand U2727 (N_2727,N_1021,N_1839);
xnor U2728 (N_2728,N_1930,N_1017);
and U2729 (N_2729,N_1245,N_1508);
or U2730 (N_2730,N_1513,N_1561);
and U2731 (N_2731,N_1603,N_1266);
and U2732 (N_2732,N_1054,N_1096);
and U2733 (N_2733,N_1023,N_1232);
and U2734 (N_2734,N_1590,N_1236);
or U2735 (N_2735,N_1566,N_1275);
nor U2736 (N_2736,N_1968,N_1583);
nor U2737 (N_2737,N_1600,N_1516);
nor U2738 (N_2738,N_1517,N_1942);
nor U2739 (N_2739,N_1792,N_1475);
nand U2740 (N_2740,N_1799,N_1710);
nand U2741 (N_2741,N_1562,N_1489);
nor U2742 (N_2742,N_1044,N_1506);
nand U2743 (N_2743,N_1390,N_1653);
nand U2744 (N_2744,N_1086,N_1476);
or U2745 (N_2745,N_1899,N_1155);
or U2746 (N_2746,N_1571,N_1653);
nor U2747 (N_2747,N_1817,N_1210);
and U2748 (N_2748,N_1119,N_1039);
or U2749 (N_2749,N_1749,N_1902);
and U2750 (N_2750,N_1441,N_1748);
and U2751 (N_2751,N_1549,N_1568);
nor U2752 (N_2752,N_1003,N_1013);
or U2753 (N_2753,N_1287,N_1191);
and U2754 (N_2754,N_1033,N_1508);
and U2755 (N_2755,N_1651,N_1565);
nand U2756 (N_2756,N_1304,N_1326);
or U2757 (N_2757,N_1888,N_1312);
nor U2758 (N_2758,N_1249,N_1094);
and U2759 (N_2759,N_1700,N_1846);
nand U2760 (N_2760,N_1053,N_1210);
or U2761 (N_2761,N_1785,N_1375);
or U2762 (N_2762,N_1918,N_1764);
and U2763 (N_2763,N_1580,N_1176);
nand U2764 (N_2764,N_1718,N_1520);
or U2765 (N_2765,N_1873,N_1609);
or U2766 (N_2766,N_1259,N_1002);
and U2767 (N_2767,N_1579,N_1524);
xor U2768 (N_2768,N_1347,N_1411);
or U2769 (N_2769,N_1126,N_1035);
or U2770 (N_2770,N_1677,N_1404);
nand U2771 (N_2771,N_1162,N_1440);
nand U2772 (N_2772,N_1246,N_1569);
or U2773 (N_2773,N_1380,N_1875);
nor U2774 (N_2774,N_1865,N_1980);
nand U2775 (N_2775,N_1303,N_1291);
nand U2776 (N_2776,N_1021,N_1057);
nor U2777 (N_2777,N_1637,N_1560);
and U2778 (N_2778,N_1598,N_1946);
and U2779 (N_2779,N_1050,N_1907);
nand U2780 (N_2780,N_1471,N_1836);
nor U2781 (N_2781,N_1815,N_1206);
nor U2782 (N_2782,N_1054,N_1829);
nor U2783 (N_2783,N_1637,N_1675);
nor U2784 (N_2784,N_1770,N_1243);
and U2785 (N_2785,N_1343,N_1943);
nor U2786 (N_2786,N_1054,N_1995);
xnor U2787 (N_2787,N_1674,N_1819);
xor U2788 (N_2788,N_1905,N_1110);
xnor U2789 (N_2789,N_1887,N_1798);
and U2790 (N_2790,N_1076,N_1588);
and U2791 (N_2791,N_1790,N_1613);
xor U2792 (N_2792,N_1905,N_1401);
or U2793 (N_2793,N_1453,N_1278);
xnor U2794 (N_2794,N_1976,N_1992);
and U2795 (N_2795,N_1307,N_1872);
xnor U2796 (N_2796,N_1364,N_1686);
nand U2797 (N_2797,N_1576,N_1707);
nor U2798 (N_2798,N_1098,N_1831);
or U2799 (N_2799,N_1190,N_1074);
and U2800 (N_2800,N_1853,N_1310);
xnor U2801 (N_2801,N_1965,N_1789);
and U2802 (N_2802,N_1534,N_1590);
and U2803 (N_2803,N_1617,N_1616);
or U2804 (N_2804,N_1003,N_1201);
or U2805 (N_2805,N_1440,N_1306);
nor U2806 (N_2806,N_1267,N_1260);
nand U2807 (N_2807,N_1047,N_1098);
nor U2808 (N_2808,N_1304,N_1896);
xor U2809 (N_2809,N_1854,N_1363);
xnor U2810 (N_2810,N_1899,N_1656);
and U2811 (N_2811,N_1488,N_1612);
or U2812 (N_2812,N_1663,N_1893);
and U2813 (N_2813,N_1350,N_1782);
nand U2814 (N_2814,N_1691,N_1232);
nor U2815 (N_2815,N_1725,N_1337);
xnor U2816 (N_2816,N_1083,N_1271);
nor U2817 (N_2817,N_1963,N_1022);
and U2818 (N_2818,N_1683,N_1921);
nand U2819 (N_2819,N_1050,N_1823);
and U2820 (N_2820,N_1690,N_1472);
nor U2821 (N_2821,N_1527,N_1133);
nand U2822 (N_2822,N_1789,N_1307);
nand U2823 (N_2823,N_1925,N_1116);
and U2824 (N_2824,N_1875,N_1817);
or U2825 (N_2825,N_1488,N_1813);
nand U2826 (N_2826,N_1338,N_1987);
or U2827 (N_2827,N_1541,N_1387);
nor U2828 (N_2828,N_1686,N_1822);
nand U2829 (N_2829,N_1132,N_1868);
or U2830 (N_2830,N_1061,N_1418);
xnor U2831 (N_2831,N_1551,N_1819);
or U2832 (N_2832,N_1603,N_1535);
nor U2833 (N_2833,N_1249,N_1082);
nand U2834 (N_2834,N_1761,N_1585);
nor U2835 (N_2835,N_1671,N_1455);
and U2836 (N_2836,N_1821,N_1070);
nor U2837 (N_2837,N_1543,N_1177);
and U2838 (N_2838,N_1402,N_1796);
and U2839 (N_2839,N_1791,N_1891);
nand U2840 (N_2840,N_1462,N_1853);
or U2841 (N_2841,N_1530,N_1618);
or U2842 (N_2842,N_1484,N_1357);
nand U2843 (N_2843,N_1448,N_1441);
and U2844 (N_2844,N_1592,N_1523);
nand U2845 (N_2845,N_1096,N_1851);
or U2846 (N_2846,N_1217,N_1452);
and U2847 (N_2847,N_1110,N_1775);
nor U2848 (N_2848,N_1584,N_1035);
and U2849 (N_2849,N_1593,N_1507);
or U2850 (N_2850,N_1148,N_1334);
nand U2851 (N_2851,N_1544,N_1131);
and U2852 (N_2852,N_1946,N_1171);
nand U2853 (N_2853,N_1637,N_1879);
nor U2854 (N_2854,N_1953,N_1031);
nand U2855 (N_2855,N_1390,N_1672);
nand U2856 (N_2856,N_1465,N_1739);
nand U2857 (N_2857,N_1963,N_1473);
nor U2858 (N_2858,N_1744,N_1468);
nand U2859 (N_2859,N_1493,N_1305);
xor U2860 (N_2860,N_1649,N_1260);
nor U2861 (N_2861,N_1503,N_1884);
nor U2862 (N_2862,N_1756,N_1114);
nand U2863 (N_2863,N_1468,N_1980);
or U2864 (N_2864,N_1599,N_1416);
nand U2865 (N_2865,N_1061,N_1833);
nor U2866 (N_2866,N_1483,N_1141);
nor U2867 (N_2867,N_1379,N_1551);
or U2868 (N_2868,N_1854,N_1468);
and U2869 (N_2869,N_1763,N_1657);
xor U2870 (N_2870,N_1842,N_1665);
and U2871 (N_2871,N_1985,N_1373);
nor U2872 (N_2872,N_1698,N_1787);
nand U2873 (N_2873,N_1315,N_1170);
nand U2874 (N_2874,N_1277,N_1213);
nand U2875 (N_2875,N_1905,N_1099);
and U2876 (N_2876,N_1287,N_1782);
and U2877 (N_2877,N_1433,N_1088);
nand U2878 (N_2878,N_1148,N_1674);
nand U2879 (N_2879,N_1842,N_1513);
nor U2880 (N_2880,N_1382,N_1423);
xnor U2881 (N_2881,N_1596,N_1371);
xnor U2882 (N_2882,N_1418,N_1113);
nor U2883 (N_2883,N_1415,N_1978);
nand U2884 (N_2884,N_1258,N_1309);
nand U2885 (N_2885,N_1421,N_1424);
nand U2886 (N_2886,N_1289,N_1848);
nand U2887 (N_2887,N_1275,N_1907);
nand U2888 (N_2888,N_1206,N_1954);
and U2889 (N_2889,N_1919,N_1334);
and U2890 (N_2890,N_1259,N_1144);
or U2891 (N_2891,N_1524,N_1971);
nor U2892 (N_2892,N_1850,N_1124);
or U2893 (N_2893,N_1808,N_1854);
nand U2894 (N_2894,N_1397,N_1759);
xor U2895 (N_2895,N_1993,N_1594);
and U2896 (N_2896,N_1782,N_1617);
and U2897 (N_2897,N_1841,N_1385);
xnor U2898 (N_2898,N_1053,N_1193);
and U2899 (N_2899,N_1494,N_1717);
and U2900 (N_2900,N_1044,N_1123);
nand U2901 (N_2901,N_1893,N_1362);
nand U2902 (N_2902,N_1732,N_1811);
and U2903 (N_2903,N_1374,N_1872);
and U2904 (N_2904,N_1128,N_1957);
or U2905 (N_2905,N_1896,N_1310);
or U2906 (N_2906,N_1339,N_1213);
nor U2907 (N_2907,N_1223,N_1096);
nor U2908 (N_2908,N_1275,N_1616);
nand U2909 (N_2909,N_1583,N_1373);
xnor U2910 (N_2910,N_1446,N_1637);
or U2911 (N_2911,N_1730,N_1563);
nor U2912 (N_2912,N_1874,N_1162);
nor U2913 (N_2913,N_1265,N_1090);
nand U2914 (N_2914,N_1849,N_1575);
nand U2915 (N_2915,N_1725,N_1822);
and U2916 (N_2916,N_1893,N_1662);
nor U2917 (N_2917,N_1190,N_1843);
nand U2918 (N_2918,N_1715,N_1991);
and U2919 (N_2919,N_1933,N_1092);
nor U2920 (N_2920,N_1867,N_1938);
nand U2921 (N_2921,N_1598,N_1703);
or U2922 (N_2922,N_1879,N_1943);
and U2923 (N_2923,N_1651,N_1939);
nand U2924 (N_2924,N_1058,N_1122);
nor U2925 (N_2925,N_1413,N_1533);
nor U2926 (N_2926,N_1884,N_1308);
nor U2927 (N_2927,N_1769,N_1808);
nand U2928 (N_2928,N_1045,N_1501);
nor U2929 (N_2929,N_1934,N_1804);
or U2930 (N_2930,N_1533,N_1270);
and U2931 (N_2931,N_1124,N_1790);
or U2932 (N_2932,N_1197,N_1261);
nor U2933 (N_2933,N_1665,N_1457);
and U2934 (N_2934,N_1718,N_1121);
nor U2935 (N_2935,N_1375,N_1266);
xor U2936 (N_2936,N_1119,N_1394);
or U2937 (N_2937,N_1818,N_1755);
or U2938 (N_2938,N_1651,N_1722);
nor U2939 (N_2939,N_1723,N_1985);
nand U2940 (N_2940,N_1296,N_1886);
and U2941 (N_2941,N_1133,N_1843);
nor U2942 (N_2942,N_1880,N_1697);
nand U2943 (N_2943,N_1234,N_1631);
or U2944 (N_2944,N_1221,N_1707);
or U2945 (N_2945,N_1714,N_1855);
nor U2946 (N_2946,N_1783,N_1887);
xnor U2947 (N_2947,N_1141,N_1170);
or U2948 (N_2948,N_1577,N_1368);
and U2949 (N_2949,N_1804,N_1203);
nand U2950 (N_2950,N_1813,N_1124);
or U2951 (N_2951,N_1802,N_1115);
and U2952 (N_2952,N_1695,N_1883);
nor U2953 (N_2953,N_1190,N_1290);
or U2954 (N_2954,N_1125,N_1185);
and U2955 (N_2955,N_1501,N_1250);
xnor U2956 (N_2956,N_1550,N_1603);
and U2957 (N_2957,N_1080,N_1221);
or U2958 (N_2958,N_1252,N_1533);
or U2959 (N_2959,N_1111,N_1107);
or U2960 (N_2960,N_1925,N_1724);
or U2961 (N_2961,N_1896,N_1805);
nor U2962 (N_2962,N_1202,N_1612);
or U2963 (N_2963,N_1695,N_1514);
or U2964 (N_2964,N_1618,N_1317);
or U2965 (N_2965,N_1462,N_1281);
and U2966 (N_2966,N_1393,N_1321);
xnor U2967 (N_2967,N_1239,N_1120);
or U2968 (N_2968,N_1604,N_1591);
or U2969 (N_2969,N_1038,N_1808);
xor U2970 (N_2970,N_1809,N_1901);
nor U2971 (N_2971,N_1530,N_1313);
nand U2972 (N_2972,N_1938,N_1310);
or U2973 (N_2973,N_1530,N_1582);
or U2974 (N_2974,N_1695,N_1858);
nor U2975 (N_2975,N_1157,N_1303);
and U2976 (N_2976,N_1167,N_1894);
or U2977 (N_2977,N_1019,N_1825);
nand U2978 (N_2978,N_1457,N_1659);
and U2979 (N_2979,N_1585,N_1610);
nor U2980 (N_2980,N_1145,N_1052);
xor U2981 (N_2981,N_1787,N_1732);
nand U2982 (N_2982,N_1770,N_1857);
or U2983 (N_2983,N_1636,N_1467);
or U2984 (N_2984,N_1802,N_1605);
nor U2985 (N_2985,N_1585,N_1944);
and U2986 (N_2986,N_1315,N_1810);
nand U2987 (N_2987,N_1018,N_1312);
and U2988 (N_2988,N_1387,N_1895);
or U2989 (N_2989,N_1494,N_1936);
and U2990 (N_2990,N_1543,N_1676);
and U2991 (N_2991,N_1586,N_1490);
xor U2992 (N_2992,N_1495,N_1935);
and U2993 (N_2993,N_1854,N_1963);
and U2994 (N_2994,N_1768,N_1277);
xnor U2995 (N_2995,N_1952,N_1518);
nand U2996 (N_2996,N_1828,N_1212);
and U2997 (N_2997,N_1003,N_1353);
nand U2998 (N_2998,N_1764,N_1547);
nor U2999 (N_2999,N_1173,N_1256);
and U3000 (N_3000,N_2893,N_2876);
xnor U3001 (N_3001,N_2092,N_2496);
and U3002 (N_3002,N_2756,N_2918);
and U3003 (N_3003,N_2619,N_2524);
nand U3004 (N_3004,N_2487,N_2314);
xnor U3005 (N_3005,N_2713,N_2825);
xor U3006 (N_3006,N_2646,N_2689);
and U3007 (N_3007,N_2174,N_2266);
and U3008 (N_3008,N_2955,N_2145);
xor U3009 (N_3009,N_2963,N_2760);
nor U3010 (N_3010,N_2187,N_2981);
nor U3011 (N_3011,N_2320,N_2896);
and U3012 (N_3012,N_2767,N_2178);
nand U3013 (N_3013,N_2434,N_2199);
or U3014 (N_3014,N_2383,N_2543);
nor U3015 (N_3015,N_2623,N_2054);
or U3016 (N_3016,N_2761,N_2891);
nor U3017 (N_3017,N_2557,N_2155);
nor U3018 (N_3018,N_2657,N_2639);
nor U3019 (N_3019,N_2341,N_2871);
nor U3020 (N_3020,N_2438,N_2656);
and U3021 (N_3021,N_2203,N_2824);
or U3022 (N_3022,N_2947,N_2762);
xor U3023 (N_3023,N_2584,N_2753);
and U3024 (N_3024,N_2363,N_2396);
xor U3025 (N_3025,N_2351,N_2879);
nand U3026 (N_3026,N_2594,N_2969);
nor U3027 (N_3027,N_2764,N_2915);
nand U3028 (N_3028,N_2538,N_2348);
or U3029 (N_3029,N_2360,N_2294);
nand U3030 (N_3030,N_2186,N_2384);
nor U3031 (N_3031,N_2143,N_2062);
nand U3032 (N_3032,N_2215,N_2666);
and U3033 (N_3033,N_2710,N_2603);
or U3034 (N_3034,N_2122,N_2688);
nor U3035 (N_3035,N_2711,N_2447);
and U3036 (N_3036,N_2738,N_2707);
nor U3037 (N_3037,N_2651,N_2058);
nand U3038 (N_3038,N_2050,N_2458);
nand U3039 (N_3039,N_2392,N_2884);
nor U3040 (N_3040,N_2339,N_2826);
or U3041 (N_3041,N_2387,N_2974);
nor U3042 (N_3042,N_2614,N_2908);
nand U3043 (N_3043,N_2902,N_2250);
nor U3044 (N_3044,N_2324,N_2751);
nand U3045 (N_3045,N_2198,N_2532);
or U3046 (N_3046,N_2925,N_2616);
nor U3047 (N_3047,N_2223,N_2179);
and U3048 (N_3048,N_2425,N_2717);
nand U3049 (N_3049,N_2232,N_2003);
and U3050 (N_3050,N_2916,N_2863);
and U3051 (N_3051,N_2926,N_2681);
nand U3052 (N_3052,N_2725,N_2935);
nand U3053 (N_3053,N_2456,N_2497);
nand U3054 (N_3054,N_2726,N_2217);
and U3055 (N_3055,N_2796,N_2797);
xnor U3056 (N_3056,N_2774,N_2870);
nor U3057 (N_3057,N_2197,N_2428);
or U3058 (N_3058,N_2548,N_2106);
and U3059 (N_3059,N_2486,N_2427);
nor U3060 (N_3060,N_2752,N_2812);
and U3061 (N_3061,N_2983,N_2192);
nor U3062 (N_3062,N_2480,N_2373);
nand U3063 (N_3063,N_2057,N_2086);
nand U3064 (N_3064,N_2793,N_2953);
and U3065 (N_3065,N_2783,N_2512);
nor U3066 (N_3066,N_2431,N_2099);
nor U3067 (N_3067,N_2887,N_2677);
nand U3068 (N_3068,N_2801,N_2951);
nor U3069 (N_3069,N_2274,N_2968);
and U3070 (N_3070,N_2407,N_2813);
or U3071 (N_3071,N_2516,N_2967);
xnor U3072 (N_3072,N_2653,N_2188);
or U3073 (N_3073,N_2328,N_2088);
xor U3074 (N_3074,N_2031,N_2006);
nor U3075 (N_3075,N_2780,N_2271);
nand U3076 (N_3076,N_2593,N_2270);
nor U3077 (N_3077,N_2345,N_2355);
nand U3078 (N_3078,N_2704,N_2528);
or U3079 (N_3079,N_2181,N_2941);
nor U3080 (N_3080,N_2148,N_2892);
or U3081 (N_3081,N_2123,N_2462);
and U3082 (N_3082,N_2504,N_2119);
or U3083 (N_3083,N_2372,N_2165);
and U3084 (N_3084,N_2381,N_2109);
nor U3085 (N_3085,N_2452,N_2036);
xnor U3086 (N_3086,N_2575,N_2869);
nor U3087 (N_3087,N_2976,N_2218);
or U3088 (N_3088,N_2133,N_2544);
xor U3089 (N_3089,N_2263,N_2698);
or U3090 (N_3090,N_2262,N_2558);
or U3091 (N_3091,N_2402,N_2077);
or U3092 (N_3092,N_2567,N_2990);
and U3093 (N_3093,N_2747,N_2632);
xnor U3094 (N_3094,N_2134,N_2325);
or U3095 (N_3095,N_2105,N_2770);
nand U3096 (N_3096,N_2131,N_2081);
nand U3097 (N_3097,N_2549,N_2530);
nor U3098 (N_3098,N_2859,N_2301);
nand U3099 (N_3099,N_2588,N_2421);
and U3100 (N_3100,N_2288,N_2598);
or U3101 (N_3101,N_2872,N_2874);
xnor U3102 (N_3102,N_2553,N_2861);
nor U3103 (N_3103,N_2676,N_2000);
or U3104 (N_3104,N_2286,N_2479);
or U3105 (N_3105,N_2540,N_2478);
or U3106 (N_3106,N_2715,N_2811);
nor U3107 (N_3107,N_2107,N_2032);
or U3108 (N_3108,N_2267,N_2459);
nand U3109 (N_3109,N_2757,N_2749);
nand U3110 (N_3110,N_2848,N_2937);
nand U3111 (N_3111,N_2911,N_2536);
nand U3112 (N_3112,N_2844,N_2508);
xnor U3113 (N_3113,N_2437,N_2009);
nor U3114 (N_3114,N_2035,N_2611);
nand U3115 (N_3115,N_2405,N_2505);
xnor U3116 (N_3116,N_2889,N_2578);
nand U3117 (N_3117,N_2815,N_2858);
nand U3118 (N_3118,N_2950,N_2239);
nand U3119 (N_3119,N_2592,N_2307);
nor U3120 (N_3120,N_2230,N_2514);
and U3121 (N_3121,N_2568,N_2996);
nand U3122 (N_3122,N_2207,N_2555);
nor U3123 (N_3123,N_2928,N_2771);
and U3124 (N_3124,N_2117,N_2924);
nor U3125 (N_3125,N_2506,N_2112);
nand U3126 (N_3126,N_2150,N_2474);
nor U3127 (N_3127,N_2680,N_2455);
and U3128 (N_3128,N_2873,N_2944);
xnor U3129 (N_3129,N_2597,N_2070);
or U3130 (N_3130,N_2068,N_2913);
and U3131 (N_3131,N_2346,N_2991);
or U3132 (N_3132,N_2766,N_2529);
nand U3133 (N_3133,N_2875,N_2097);
nand U3134 (N_3134,N_2708,N_2862);
or U3135 (N_3135,N_2473,N_2962);
nor U3136 (N_3136,N_2393,N_2570);
nand U3137 (N_3137,N_2227,N_2450);
nand U3138 (N_3138,N_2451,N_2406);
nor U3139 (N_3139,N_2792,N_2278);
nor U3140 (N_3140,N_2183,N_2214);
nor U3141 (N_3141,N_2807,N_2040);
nor U3142 (N_3142,N_2556,N_2659);
nor U3143 (N_3143,N_2140,N_2443);
or U3144 (N_3144,N_2213,N_2901);
and U3145 (N_3145,N_2489,N_2814);
nand U3146 (N_3146,N_2055,N_2017);
xnor U3147 (N_3147,N_2258,N_2520);
nand U3148 (N_3148,N_2854,N_2587);
and U3149 (N_3149,N_2599,N_2609);
xnor U3150 (N_3150,N_2519,N_2180);
xor U3151 (N_3151,N_2775,N_2746);
and U3152 (N_3152,N_2354,N_2045);
and U3153 (N_3153,N_2216,N_2413);
and U3154 (N_3154,N_2485,N_2137);
or U3155 (N_3155,N_2021,N_2564);
nor U3156 (N_3156,N_2033,N_2238);
or U3157 (N_3157,N_2690,N_2159);
or U3158 (N_3158,N_2272,N_2731);
xor U3159 (N_3159,N_2836,N_2240);
and U3160 (N_3160,N_2997,N_2574);
and U3161 (N_3161,N_2222,N_2161);
and U3162 (N_3162,N_2102,N_2552);
xor U3163 (N_3163,N_2259,N_2034);
nand U3164 (N_3164,N_2053,N_2633);
and U3165 (N_3165,N_2369,N_2791);
and U3166 (N_3166,N_2498,N_2295);
nand U3167 (N_3167,N_2298,N_2171);
nor U3168 (N_3168,N_2679,N_2987);
or U3169 (N_3169,N_2481,N_2810);
nand U3170 (N_3170,N_2444,N_2454);
nand U3171 (N_3171,N_2601,N_2299);
xnor U3172 (N_3172,N_2291,N_2560);
nand U3173 (N_3173,N_2353,N_2125);
and U3174 (N_3174,N_2210,N_2025);
xor U3175 (N_3175,N_2781,N_2965);
or U3176 (N_3176,N_2841,N_2643);
and U3177 (N_3177,N_2201,N_2970);
nor U3178 (N_3178,N_2477,N_2082);
or U3179 (N_3179,N_2417,N_2763);
xor U3180 (N_3180,N_2265,N_2920);
nand U3181 (N_3181,N_2284,N_2663);
or U3182 (N_3182,N_2631,N_2020);
or U3183 (N_3183,N_2471,N_2583);
or U3184 (N_3184,N_2847,N_2596);
nor U3185 (N_3185,N_2304,N_2337);
nor U3186 (N_3186,N_2957,N_2042);
xor U3187 (N_3187,N_2590,N_2061);
or U3188 (N_3188,N_2248,N_2418);
nor U3189 (N_3189,N_2789,N_2577);
xnor U3190 (N_3190,N_2157,N_2765);
nand U3191 (N_3191,N_2185,N_2897);
nor U3192 (N_3192,N_2476,N_2388);
nand U3193 (N_3193,N_2500,N_2261);
nand U3194 (N_3194,N_2175,N_2467);
nand U3195 (N_3195,N_2051,N_2395);
or U3196 (N_3196,N_2310,N_2401);
nor U3197 (N_3197,N_2482,N_2358);
or U3198 (N_3198,N_2151,N_2678);
xnor U3199 (N_3199,N_2224,N_2943);
and U3200 (N_3200,N_2211,N_2805);
or U3201 (N_3201,N_2542,N_2121);
nand U3202 (N_3202,N_2727,N_2977);
and U3203 (N_3203,N_2315,N_2705);
and U3204 (N_3204,N_2090,N_2758);
nor U3205 (N_3205,N_2827,N_2436);
nor U3206 (N_3206,N_2404,N_2886);
or U3207 (N_3207,N_2022,N_2745);
or U3208 (N_3208,N_2285,N_2243);
xnor U3209 (N_3209,N_2703,N_2275);
xor U3210 (N_3210,N_2682,N_2980);
and U3211 (N_3211,N_2629,N_2300);
nand U3212 (N_3212,N_2586,N_2683);
nor U3213 (N_3213,N_2819,N_2670);
nor U3214 (N_3214,N_2978,N_2961);
nor U3215 (N_3215,N_2909,N_2029);
nand U3216 (N_3216,N_2279,N_2956);
nand U3217 (N_3217,N_2039,N_2209);
nor U3218 (N_3218,N_2537,N_2648);
and U3219 (N_3219,N_2076,N_2959);
or U3220 (N_3220,N_2290,N_2101);
nor U3221 (N_3221,N_2469,N_2533);
and U3222 (N_3222,N_2817,N_2219);
or U3223 (N_3223,N_2857,N_2675);
and U3224 (N_3224,N_2719,N_2010);
or U3225 (N_3225,N_2853,N_2297);
nor U3226 (N_3226,N_2332,N_2024);
or U3227 (N_3227,N_2546,N_2184);
or U3228 (N_3228,N_2610,N_2895);
and U3229 (N_3229,N_2226,N_2917);
or U3230 (N_3230,N_2787,N_2687);
or U3231 (N_3231,N_2289,N_2347);
nor U3232 (N_3232,N_2655,N_2241);
nand U3233 (N_3233,N_2015,N_2843);
nand U3234 (N_3234,N_2168,N_2940);
or U3235 (N_3235,N_2931,N_2132);
xnor U3236 (N_3236,N_2306,N_2379);
nor U3237 (N_3237,N_2495,N_2435);
nand U3238 (N_3238,N_2439,N_2625);
nor U3239 (N_3239,N_2466,N_2626);
nor U3240 (N_3240,N_2449,N_2382);
nor U3241 (N_3241,N_2292,N_2788);
and U3242 (N_3242,N_2880,N_2249);
or U3243 (N_3243,N_2453,N_2499);
and U3244 (N_3244,N_2463,N_2782);
nand U3245 (N_3245,N_2182,N_2044);
nand U3246 (N_3246,N_2850,N_2565);
or U3247 (N_3247,N_2733,N_2773);
nor U3248 (N_3248,N_2697,N_2135);
and U3249 (N_3249,N_2147,N_2692);
or U3250 (N_3250,N_2194,N_2995);
nand U3251 (N_3251,N_2089,N_2163);
nand U3252 (N_3252,N_2400,N_2942);
nor U3253 (N_3253,N_2576,N_2430);
xor U3254 (N_3254,N_2080,N_2741);
nor U3255 (N_3255,N_2833,N_2864);
xnor U3256 (N_3256,N_2110,N_2330);
and U3257 (N_3257,N_2866,N_2635);
nand U3258 (N_3258,N_2634,N_2362);
nand U3259 (N_3259,N_2309,N_2612);
nor U3260 (N_3260,N_2027,N_2883);
nand U3261 (N_3261,N_2998,N_2321);
or U3262 (N_3262,N_2167,N_2359);
nand U3263 (N_3263,N_2885,N_2714);
and U3264 (N_3264,N_2842,N_2100);
and U3265 (N_3265,N_2515,N_2964);
nor U3266 (N_3266,N_2313,N_2377);
or U3267 (N_3267,N_2988,N_2484);
nor U3268 (N_3268,N_2699,N_2242);
or U3269 (N_3269,N_2510,N_2342);
nand U3270 (N_3270,N_2475,N_2046);
and U3271 (N_3271,N_2293,N_2637);
xor U3272 (N_3272,N_2803,N_2316);
or U3273 (N_3273,N_2344,N_2281);
or U3274 (N_3274,N_2525,N_2144);
nand U3275 (N_3275,N_2971,N_2349);
and U3276 (N_3276,N_2071,N_2820);
nand U3277 (N_3277,N_2038,N_2790);
and U3278 (N_3278,N_2067,N_2531);
nand U3279 (N_3279,N_2412,N_2221);
nor U3280 (N_3280,N_2335,N_2702);
xor U3281 (N_3281,N_2849,N_2865);
and U3282 (N_3282,N_2855,N_2028);
nand U3283 (N_3283,N_2389,N_2317);
or U3284 (N_3284,N_2527,N_2252);
and U3285 (N_3285,N_2492,N_2411);
xnor U3286 (N_3286,N_2312,N_2694);
xor U3287 (N_3287,N_2257,N_2882);
or U3288 (N_3288,N_2986,N_2580);
nor U3289 (N_3289,N_2160,N_2483);
nor U3290 (N_3290,N_2472,N_2319);
nand U3291 (N_3291,N_2828,N_2253);
and U3292 (N_3292,N_2907,N_2126);
nor U3293 (N_3293,N_2246,N_2534);
nand U3294 (N_3294,N_2936,N_2660);
nand U3295 (N_3295,N_2838,N_2742);
nand U3296 (N_3296,N_2602,N_2740);
nand U3297 (N_3297,N_2685,N_2419);
nor U3298 (N_3298,N_2975,N_2972);
nor U3299 (N_3299,N_2014,N_2644);
nor U3300 (N_3300,N_2366,N_2691);
nor U3301 (N_3301,N_2989,N_2769);
xnor U3302 (N_3302,N_2390,N_2056);
nor U3303 (N_3303,N_2894,N_2674);
or U3304 (N_3304,N_2254,N_2701);
or U3305 (N_3305,N_2662,N_2060);
nand U3306 (N_3306,N_2939,N_2878);
nor U3307 (N_3307,N_2938,N_2063);
or U3308 (N_3308,N_2851,N_2146);
nand U3309 (N_3309,N_2108,N_2468);
nand U3310 (N_3310,N_2343,N_2370);
nor U3311 (N_3311,N_2999,N_2730);
nor U3312 (N_3312,N_2172,N_2799);
nor U3313 (N_3313,N_2138,N_2904);
and U3314 (N_3314,N_2754,N_2607);
or U3315 (N_3315,N_2994,N_2164);
or U3316 (N_3316,N_2948,N_2043);
and U3317 (N_3317,N_2296,N_2728);
nand U3318 (N_3318,N_2268,N_2423);
and U3319 (N_3319,N_2759,N_2890);
nand U3320 (N_3320,N_2804,N_2664);
xnor U3321 (N_3321,N_2591,N_2352);
or U3322 (N_3322,N_2367,N_2103);
nand U3323 (N_3323,N_2903,N_2059);
and U3324 (N_3324,N_2120,N_2712);
and U3325 (N_3325,N_2834,N_2166);
and U3326 (N_3326,N_2195,N_2011);
nor U3327 (N_3327,N_2618,N_2276);
and U3328 (N_3328,N_2706,N_2013);
nand U3329 (N_3329,N_2949,N_2735);
or U3330 (N_3330,N_2244,N_2114);
or U3331 (N_3331,N_2709,N_2193);
nor U3332 (N_3332,N_2128,N_2426);
and U3333 (N_3333,N_2008,N_2613);
nand U3334 (N_3334,N_2642,N_2432);
xor U3335 (N_3335,N_2667,N_2093);
nand U3336 (N_3336,N_2269,N_2399);
xor U3337 (N_3337,N_2303,N_2808);
or U3338 (N_3338,N_2661,N_2397);
and U3339 (N_3339,N_2104,N_2569);
or U3340 (N_3340,N_2260,N_2311);
xnor U3341 (N_3341,N_2624,N_2518);
and U3342 (N_3342,N_2772,N_2212);
and U3343 (N_3343,N_2566,N_2173);
nand U3344 (N_3344,N_2069,N_2608);
nor U3345 (N_3345,N_2460,N_2235);
xor U3346 (N_3346,N_2647,N_2502);
nand U3347 (N_3347,N_2340,N_2073);
and U3348 (N_3348,N_2922,N_2493);
xnor U3349 (N_3349,N_2433,N_2605);
and U3350 (N_3350,N_2323,N_2445);
and U3351 (N_3351,N_2784,N_2231);
nor U3352 (N_3352,N_2734,N_2934);
and U3353 (N_3353,N_2318,N_2153);
or U3354 (N_3354,N_2620,N_2336);
nand U3355 (N_3355,N_2049,N_2795);
and U3356 (N_3356,N_2572,N_2600);
xnor U3357 (N_3357,N_2139,N_2357);
nand U3358 (N_3358,N_2012,N_2441);
nor U3359 (N_3359,N_2127,N_2507);
nand U3360 (N_3360,N_2744,N_2442);
and U3361 (N_3361,N_2521,N_2946);
and U3362 (N_3362,N_2394,N_2408);
and U3363 (N_3363,N_2729,N_2554);
or U3364 (N_3364,N_2041,N_2118);
xnor U3365 (N_3365,N_2004,N_2914);
or U3366 (N_3366,N_2736,N_2162);
and U3367 (N_3367,N_2881,N_2721);
nor U3368 (N_3368,N_2465,N_2490);
nor U3369 (N_3369,N_2416,N_2535);
or U3370 (N_3370,N_2491,N_2562);
and U3371 (N_3371,N_2169,N_2415);
nand U3372 (N_3372,N_2818,N_2005);
xor U3373 (N_3373,N_2375,N_2654);
nand U3374 (N_3374,N_2154,N_2900);
and U3375 (N_3375,N_2779,N_2800);
or U3376 (N_3376,N_2066,N_2037);
or U3377 (N_3377,N_2846,N_2350);
xnor U3378 (N_3378,N_2563,N_2722);
and U3379 (N_3379,N_2589,N_2755);
nor U3380 (N_3380,N_2440,N_2693);
nor U3381 (N_3381,N_2200,N_2420);
and U3382 (N_3382,N_2116,N_2237);
nor U3383 (N_3383,N_2585,N_2982);
and U3384 (N_3384,N_2595,N_2856);
nand U3385 (N_3385,N_2047,N_2503);
nor U3386 (N_3386,N_2398,N_2177);
nor U3387 (N_3387,N_2509,N_2158);
or U3388 (N_3388,N_2684,N_2615);
nor U3389 (N_3389,N_2391,N_2671);
nor U3390 (N_3390,N_2115,N_2929);
nor U3391 (N_3391,N_2196,N_2026);
xnor U3392 (N_3392,N_2973,N_2628);
or U3393 (N_3393,N_2446,N_2225);
nor U3394 (N_3394,N_2550,N_2287);
or U3395 (N_3395,N_2737,N_2966);
or U3396 (N_3396,N_2280,N_2526);
and U3397 (N_3397,N_2424,N_2945);
nand U3398 (N_3398,N_2927,N_2686);
nor U3399 (N_3399,N_2724,N_2149);
nor U3400 (N_3400,N_2905,N_2837);
and U3401 (N_3401,N_2582,N_2672);
nand U3402 (N_3402,N_2448,N_2501);
nor U3403 (N_3403,N_2621,N_2233);
nor U3404 (N_3404,N_2302,N_2777);
nor U3405 (N_3405,N_2830,N_2356);
and U3406 (N_3406,N_2256,N_2839);
nand U3407 (N_3407,N_2282,N_2739);
or U3408 (N_3408,N_2522,N_2523);
nor U3409 (N_3409,N_2930,N_2305);
or U3410 (N_3410,N_2627,N_2136);
and U3411 (N_3411,N_2668,N_2130);
and U3412 (N_3412,N_2932,N_2673);
or U3413 (N_3413,N_2912,N_2494);
nand U3414 (N_3414,N_2064,N_2539);
and U3415 (N_3415,N_2561,N_2852);
or U3416 (N_3416,N_2993,N_2001);
nand U3417 (N_3417,N_2919,N_2716);
or U3418 (N_3418,N_2923,N_2979);
nand U3419 (N_3419,N_2630,N_2802);
or U3420 (N_3420,N_2072,N_2338);
nor U3421 (N_3421,N_2720,N_2984);
nor U3422 (N_3422,N_2208,N_2579);
and U3423 (N_3423,N_2868,N_2331);
xnor U3424 (N_3424,N_2308,N_2541);
nand U3425 (N_3425,N_2176,N_2786);
nand U3426 (N_3426,N_2084,N_2617);
and U3427 (N_3427,N_2124,N_2245);
nand U3428 (N_3428,N_2236,N_2111);
or U3429 (N_3429,N_2141,N_2910);
nand U3430 (N_3430,N_2002,N_2085);
nor U3431 (N_3431,N_2189,N_2083);
or U3432 (N_3432,N_2571,N_2547);
nor U3433 (N_3433,N_2096,N_2018);
nand U3434 (N_3434,N_2142,N_2652);
or U3435 (N_3435,N_2954,N_2094);
nor U3436 (N_3436,N_2906,N_2277);
xnor U3437 (N_3437,N_2374,N_2079);
nor U3438 (N_3438,N_2640,N_2016);
nor U3439 (N_3439,N_2750,N_2732);
xnor U3440 (N_3440,N_2414,N_2649);
and U3441 (N_3441,N_2958,N_2898);
nor U3442 (N_3442,N_2933,N_2075);
and U3443 (N_3443,N_2422,N_2511);
nor U3444 (N_3444,N_2205,N_2778);
nand U3445 (N_3445,N_2985,N_2821);
nand U3446 (N_3446,N_2385,N_2087);
or U3447 (N_3447,N_2835,N_2513);
nor U3448 (N_3448,N_2251,N_2470);
nand U3449 (N_3449,N_2326,N_2461);
nand U3450 (N_3450,N_2464,N_2113);
nand U3451 (N_3451,N_2921,N_2641);
nand U3452 (N_3452,N_2604,N_2723);
nand U3453 (N_3453,N_2074,N_2368);
xor U3454 (N_3454,N_2380,N_2403);
nand U3455 (N_3455,N_2091,N_2156);
and U3456 (N_3456,N_2007,N_2329);
xor U3457 (N_3457,N_2860,N_2545);
and U3458 (N_3458,N_2098,N_2264);
xor U3459 (N_3459,N_2371,N_2899);
nand U3460 (N_3460,N_2992,N_2322);
or U3461 (N_3461,N_2206,N_2283);
or U3462 (N_3462,N_2831,N_2361);
or U3463 (N_3463,N_2832,N_2798);
nand U3464 (N_3464,N_2204,N_2748);
or U3465 (N_3465,N_2768,N_2816);
nand U3466 (N_3466,N_2867,N_2845);
nor U3467 (N_3467,N_2327,N_2573);
or U3468 (N_3468,N_2228,N_2065);
or U3469 (N_3469,N_2365,N_2095);
nand U3470 (N_3470,N_2220,N_2273);
xor U3471 (N_3471,N_2364,N_2078);
nor U3472 (N_3472,N_2809,N_2247);
xor U3473 (N_3473,N_2960,N_2658);
or U3474 (N_3474,N_2019,N_2052);
or U3475 (N_3475,N_2888,N_2234);
nor U3476 (N_3476,N_2170,N_2255);
or U3477 (N_3477,N_2696,N_2794);
and U3478 (N_3478,N_2202,N_2829);
and U3479 (N_3479,N_2129,N_2776);
nor U3480 (N_3480,N_2023,N_2650);
or U3481 (N_3481,N_2743,N_2606);
nor U3482 (N_3482,N_2378,N_2669);
or U3483 (N_3483,N_2665,N_2559);
nand U3484 (N_3484,N_2806,N_2822);
nor U3485 (N_3485,N_2376,N_2638);
nand U3486 (N_3486,N_2840,N_2622);
and U3487 (N_3487,N_2229,N_2409);
xnor U3488 (N_3488,N_2190,N_2386);
or U3489 (N_3489,N_2952,N_2700);
and U3490 (N_3490,N_2030,N_2191);
or U3491 (N_3491,N_2410,N_2048);
or U3492 (N_3492,N_2785,N_2152);
nand U3493 (N_3493,N_2695,N_2581);
xnor U3494 (N_3494,N_2517,N_2333);
nand U3495 (N_3495,N_2718,N_2488);
xnor U3496 (N_3496,N_2636,N_2877);
nor U3497 (N_3497,N_2551,N_2645);
and U3498 (N_3498,N_2334,N_2823);
nand U3499 (N_3499,N_2429,N_2457);
nor U3500 (N_3500,N_2231,N_2147);
or U3501 (N_3501,N_2810,N_2602);
nand U3502 (N_3502,N_2550,N_2763);
and U3503 (N_3503,N_2577,N_2747);
nor U3504 (N_3504,N_2260,N_2098);
nor U3505 (N_3505,N_2215,N_2732);
xnor U3506 (N_3506,N_2382,N_2627);
or U3507 (N_3507,N_2207,N_2570);
or U3508 (N_3508,N_2067,N_2583);
nor U3509 (N_3509,N_2789,N_2594);
and U3510 (N_3510,N_2569,N_2417);
nor U3511 (N_3511,N_2499,N_2360);
or U3512 (N_3512,N_2214,N_2934);
and U3513 (N_3513,N_2549,N_2019);
nor U3514 (N_3514,N_2748,N_2797);
xor U3515 (N_3515,N_2195,N_2149);
nor U3516 (N_3516,N_2683,N_2579);
nand U3517 (N_3517,N_2573,N_2800);
xor U3518 (N_3518,N_2993,N_2236);
nand U3519 (N_3519,N_2478,N_2502);
nand U3520 (N_3520,N_2907,N_2675);
nor U3521 (N_3521,N_2401,N_2004);
or U3522 (N_3522,N_2007,N_2365);
nand U3523 (N_3523,N_2965,N_2338);
nor U3524 (N_3524,N_2503,N_2110);
or U3525 (N_3525,N_2152,N_2631);
and U3526 (N_3526,N_2490,N_2230);
xor U3527 (N_3527,N_2185,N_2872);
nor U3528 (N_3528,N_2864,N_2869);
or U3529 (N_3529,N_2432,N_2295);
nand U3530 (N_3530,N_2716,N_2773);
nand U3531 (N_3531,N_2137,N_2478);
nand U3532 (N_3532,N_2300,N_2526);
or U3533 (N_3533,N_2947,N_2204);
or U3534 (N_3534,N_2944,N_2597);
and U3535 (N_3535,N_2064,N_2108);
nand U3536 (N_3536,N_2015,N_2610);
and U3537 (N_3537,N_2733,N_2836);
nand U3538 (N_3538,N_2276,N_2190);
and U3539 (N_3539,N_2540,N_2616);
or U3540 (N_3540,N_2252,N_2635);
and U3541 (N_3541,N_2007,N_2033);
nor U3542 (N_3542,N_2233,N_2527);
and U3543 (N_3543,N_2823,N_2012);
nand U3544 (N_3544,N_2039,N_2506);
nand U3545 (N_3545,N_2956,N_2392);
and U3546 (N_3546,N_2984,N_2070);
and U3547 (N_3547,N_2491,N_2533);
and U3548 (N_3548,N_2630,N_2840);
nor U3549 (N_3549,N_2925,N_2664);
and U3550 (N_3550,N_2217,N_2096);
nor U3551 (N_3551,N_2665,N_2607);
and U3552 (N_3552,N_2588,N_2674);
xnor U3553 (N_3553,N_2735,N_2198);
or U3554 (N_3554,N_2022,N_2477);
xnor U3555 (N_3555,N_2644,N_2717);
nor U3556 (N_3556,N_2701,N_2804);
and U3557 (N_3557,N_2158,N_2290);
nand U3558 (N_3558,N_2056,N_2399);
or U3559 (N_3559,N_2923,N_2536);
or U3560 (N_3560,N_2220,N_2320);
or U3561 (N_3561,N_2431,N_2623);
nand U3562 (N_3562,N_2897,N_2100);
and U3563 (N_3563,N_2428,N_2062);
or U3564 (N_3564,N_2895,N_2813);
and U3565 (N_3565,N_2790,N_2129);
and U3566 (N_3566,N_2944,N_2386);
nor U3567 (N_3567,N_2915,N_2226);
nor U3568 (N_3568,N_2548,N_2131);
nor U3569 (N_3569,N_2429,N_2001);
nor U3570 (N_3570,N_2410,N_2324);
nand U3571 (N_3571,N_2840,N_2417);
or U3572 (N_3572,N_2250,N_2813);
or U3573 (N_3573,N_2683,N_2551);
and U3574 (N_3574,N_2823,N_2155);
nand U3575 (N_3575,N_2973,N_2654);
nand U3576 (N_3576,N_2991,N_2747);
nand U3577 (N_3577,N_2650,N_2052);
nand U3578 (N_3578,N_2124,N_2332);
or U3579 (N_3579,N_2141,N_2953);
or U3580 (N_3580,N_2161,N_2300);
or U3581 (N_3581,N_2331,N_2393);
nor U3582 (N_3582,N_2422,N_2342);
xor U3583 (N_3583,N_2298,N_2473);
nand U3584 (N_3584,N_2529,N_2515);
xnor U3585 (N_3585,N_2158,N_2931);
and U3586 (N_3586,N_2730,N_2179);
and U3587 (N_3587,N_2982,N_2833);
nor U3588 (N_3588,N_2072,N_2048);
nor U3589 (N_3589,N_2568,N_2796);
nand U3590 (N_3590,N_2123,N_2730);
and U3591 (N_3591,N_2889,N_2697);
or U3592 (N_3592,N_2719,N_2173);
nand U3593 (N_3593,N_2902,N_2211);
nor U3594 (N_3594,N_2300,N_2041);
and U3595 (N_3595,N_2293,N_2920);
and U3596 (N_3596,N_2109,N_2997);
or U3597 (N_3597,N_2880,N_2082);
or U3598 (N_3598,N_2489,N_2497);
or U3599 (N_3599,N_2450,N_2084);
nor U3600 (N_3600,N_2619,N_2012);
nor U3601 (N_3601,N_2399,N_2268);
or U3602 (N_3602,N_2409,N_2254);
nand U3603 (N_3603,N_2696,N_2706);
nand U3604 (N_3604,N_2556,N_2105);
or U3605 (N_3605,N_2215,N_2975);
and U3606 (N_3606,N_2471,N_2065);
xor U3607 (N_3607,N_2437,N_2146);
and U3608 (N_3608,N_2063,N_2163);
xor U3609 (N_3609,N_2812,N_2447);
xnor U3610 (N_3610,N_2886,N_2200);
and U3611 (N_3611,N_2442,N_2992);
xor U3612 (N_3612,N_2459,N_2707);
nor U3613 (N_3613,N_2819,N_2886);
or U3614 (N_3614,N_2747,N_2006);
or U3615 (N_3615,N_2741,N_2915);
xor U3616 (N_3616,N_2898,N_2625);
nand U3617 (N_3617,N_2283,N_2785);
nor U3618 (N_3618,N_2111,N_2158);
or U3619 (N_3619,N_2112,N_2076);
and U3620 (N_3620,N_2424,N_2506);
nand U3621 (N_3621,N_2674,N_2089);
xor U3622 (N_3622,N_2451,N_2957);
or U3623 (N_3623,N_2835,N_2270);
and U3624 (N_3624,N_2192,N_2576);
and U3625 (N_3625,N_2000,N_2747);
nor U3626 (N_3626,N_2137,N_2301);
nor U3627 (N_3627,N_2369,N_2776);
xnor U3628 (N_3628,N_2909,N_2441);
nand U3629 (N_3629,N_2346,N_2814);
or U3630 (N_3630,N_2014,N_2318);
or U3631 (N_3631,N_2829,N_2957);
nor U3632 (N_3632,N_2502,N_2716);
nand U3633 (N_3633,N_2084,N_2236);
and U3634 (N_3634,N_2332,N_2185);
nor U3635 (N_3635,N_2925,N_2899);
and U3636 (N_3636,N_2995,N_2387);
nor U3637 (N_3637,N_2291,N_2266);
nand U3638 (N_3638,N_2085,N_2683);
or U3639 (N_3639,N_2308,N_2901);
and U3640 (N_3640,N_2440,N_2194);
and U3641 (N_3641,N_2058,N_2562);
or U3642 (N_3642,N_2072,N_2357);
or U3643 (N_3643,N_2236,N_2166);
or U3644 (N_3644,N_2543,N_2617);
or U3645 (N_3645,N_2262,N_2361);
or U3646 (N_3646,N_2966,N_2491);
xor U3647 (N_3647,N_2247,N_2109);
or U3648 (N_3648,N_2049,N_2842);
nor U3649 (N_3649,N_2148,N_2172);
nand U3650 (N_3650,N_2388,N_2482);
and U3651 (N_3651,N_2070,N_2863);
or U3652 (N_3652,N_2783,N_2464);
nor U3653 (N_3653,N_2117,N_2554);
or U3654 (N_3654,N_2456,N_2044);
nand U3655 (N_3655,N_2857,N_2517);
or U3656 (N_3656,N_2508,N_2623);
and U3657 (N_3657,N_2416,N_2538);
nor U3658 (N_3658,N_2084,N_2090);
xor U3659 (N_3659,N_2962,N_2823);
nand U3660 (N_3660,N_2342,N_2905);
and U3661 (N_3661,N_2536,N_2327);
nor U3662 (N_3662,N_2955,N_2611);
or U3663 (N_3663,N_2796,N_2113);
nor U3664 (N_3664,N_2524,N_2232);
nand U3665 (N_3665,N_2525,N_2310);
nand U3666 (N_3666,N_2256,N_2858);
nor U3667 (N_3667,N_2646,N_2459);
and U3668 (N_3668,N_2262,N_2826);
xor U3669 (N_3669,N_2721,N_2764);
xnor U3670 (N_3670,N_2813,N_2831);
nand U3671 (N_3671,N_2023,N_2713);
nand U3672 (N_3672,N_2233,N_2224);
nand U3673 (N_3673,N_2627,N_2018);
or U3674 (N_3674,N_2068,N_2923);
nand U3675 (N_3675,N_2950,N_2746);
or U3676 (N_3676,N_2030,N_2882);
nand U3677 (N_3677,N_2258,N_2941);
nor U3678 (N_3678,N_2832,N_2825);
nand U3679 (N_3679,N_2149,N_2891);
and U3680 (N_3680,N_2852,N_2058);
and U3681 (N_3681,N_2292,N_2669);
and U3682 (N_3682,N_2777,N_2141);
nor U3683 (N_3683,N_2523,N_2208);
or U3684 (N_3684,N_2586,N_2860);
nor U3685 (N_3685,N_2932,N_2356);
or U3686 (N_3686,N_2019,N_2425);
xnor U3687 (N_3687,N_2203,N_2910);
and U3688 (N_3688,N_2863,N_2384);
nor U3689 (N_3689,N_2810,N_2761);
or U3690 (N_3690,N_2952,N_2683);
and U3691 (N_3691,N_2074,N_2347);
and U3692 (N_3692,N_2860,N_2613);
and U3693 (N_3693,N_2355,N_2449);
nor U3694 (N_3694,N_2822,N_2015);
nand U3695 (N_3695,N_2934,N_2059);
and U3696 (N_3696,N_2191,N_2971);
nor U3697 (N_3697,N_2968,N_2145);
and U3698 (N_3698,N_2758,N_2962);
or U3699 (N_3699,N_2373,N_2924);
nor U3700 (N_3700,N_2165,N_2604);
or U3701 (N_3701,N_2910,N_2500);
nor U3702 (N_3702,N_2780,N_2051);
and U3703 (N_3703,N_2597,N_2891);
xnor U3704 (N_3704,N_2501,N_2427);
nor U3705 (N_3705,N_2212,N_2416);
nor U3706 (N_3706,N_2382,N_2216);
or U3707 (N_3707,N_2253,N_2374);
xnor U3708 (N_3708,N_2185,N_2967);
nor U3709 (N_3709,N_2131,N_2055);
nor U3710 (N_3710,N_2245,N_2688);
nand U3711 (N_3711,N_2312,N_2911);
nand U3712 (N_3712,N_2032,N_2061);
and U3713 (N_3713,N_2481,N_2409);
nand U3714 (N_3714,N_2257,N_2744);
nor U3715 (N_3715,N_2713,N_2831);
and U3716 (N_3716,N_2632,N_2991);
and U3717 (N_3717,N_2337,N_2778);
xor U3718 (N_3718,N_2482,N_2429);
and U3719 (N_3719,N_2600,N_2303);
and U3720 (N_3720,N_2549,N_2646);
or U3721 (N_3721,N_2605,N_2552);
nand U3722 (N_3722,N_2936,N_2323);
and U3723 (N_3723,N_2402,N_2631);
and U3724 (N_3724,N_2922,N_2616);
nor U3725 (N_3725,N_2649,N_2360);
xnor U3726 (N_3726,N_2597,N_2978);
xnor U3727 (N_3727,N_2840,N_2629);
nand U3728 (N_3728,N_2444,N_2213);
and U3729 (N_3729,N_2885,N_2926);
or U3730 (N_3730,N_2423,N_2338);
xnor U3731 (N_3731,N_2094,N_2320);
or U3732 (N_3732,N_2130,N_2444);
or U3733 (N_3733,N_2176,N_2833);
xnor U3734 (N_3734,N_2878,N_2637);
nor U3735 (N_3735,N_2456,N_2394);
nor U3736 (N_3736,N_2527,N_2588);
and U3737 (N_3737,N_2440,N_2423);
and U3738 (N_3738,N_2345,N_2438);
xor U3739 (N_3739,N_2057,N_2779);
and U3740 (N_3740,N_2026,N_2915);
or U3741 (N_3741,N_2560,N_2667);
xnor U3742 (N_3742,N_2252,N_2295);
nor U3743 (N_3743,N_2081,N_2124);
and U3744 (N_3744,N_2609,N_2834);
nor U3745 (N_3745,N_2632,N_2474);
nand U3746 (N_3746,N_2971,N_2150);
nand U3747 (N_3747,N_2867,N_2085);
and U3748 (N_3748,N_2260,N_2949);
nand U3749 (N_3749,N_2401,N_2125);
xor U3750 (N_3750,N_2777,N_2649);
nor U3751 (N_3751,N_2101,N_2569);
nand U3752 (N_3752,N_2708,N_2507);
or U3753 (N_3753,N_2652,N_2153);
and U3754 (N_3754,N_2388,N_2519);
xor U3755 (N_3755,N_2386,N_2932);
nand U3756 (N_3756,N_2183,N_2494);
or U3757 (N_3757,N_2919,N_2781);
or U3758 (N_3758,N_2814,N_2633);
or U3759 (N_3759,N_2892,N_2164);
or U3760 (N_3760,N_2807,N_2734);
or U3761 (N_3761,N_2041,N_2441);
nor U3762 (N_3762,N_2494,N_2240);
nand U3763 (N_3763,N_2456,N_2918);
and U3764 (N_3764,N_2377,N_2020);
and U3765 (N_3765,N_2659,N_2361);
and U3766 (N_3766,N_2248,N_2939);
and U3767 (N_3767,N_2596,N_2783);
nand U3768 (N_3768,N_2769,N_2863);
and U3769 (N_3769,N_2248,N_2405);
and U3770 (N_3770,N_2816,N_2480);
nor U3771 (N_3771,N_2164,N_2611);
or U3772 (N_3772,N_2114,N_2349);
and U3773 (N_3773,N_2098,N_2618);
xnor U3774 (N_3774,N_2343,N_2628);
nand U3775 (N_3775,N_2488,N_2043);
and U3776 (N_3776,N_2336,N_2146);
or U3777 (N_3777,N_2382,N_2859);
xor U3778 (N_3778,N_2100,N_2419);
xor U3779 (N_3779,N_2911,N_2224);
nor U3780 (N_3780,N_2327,N_2931);
and U3781 (N_3781,N_2828,N_2784);
or U3782 (N_3782,N_2532,N_2589);
and U3783 (N_3783,N_2708,N_2063);
xnor U3784 (N_3784,N_2873,N_2835);
nand U3785 (N_3785,N_2702,N_2171);
and U3786 (N_3786,N_2894,N_2124);
xor U3787 (N_3787,N_2477,N_2089);
or U3788 (N_3788,N_2018,N_2338);
or U3789 (N_3789,N_2632,N_2597);
or U3790 (N_3790,N_2179,N_2960);
nor U3791 (N_3791,N_2277,N_2909);
and U3792 (N_3792,N_2556,N_2891);
nand U3793 (N_3793,N_2143,N_2040);
and U3794 (N_3794,N_2528,N_2910);
and U3795 (N_3795,N_2139,N_2606);
nand U3796 (N_3796,N_2466,N_2806);
or U3797 (N_3797,N_2914,N_2885);
nand U3798 (N_3798,N_2558,N_2211);
xnor U3799 (N_3799,N_2831,N_2635);
xnor U3800 (N_3800,N_2031,N_2765);
nand U3801 (N_3801,N_2236,N_2891);
or U3802 (N_3802,N_2976,N_2842);
or U3803 (N_3803,N_2335,N_2928);
or U3804 (N_3804,N_2334,N_2816);
or U3805 (N_3805,N_2202,N_2780);
or U3806 (N_3806,N_2844,N_2527);
and U3807 (N_3807,N_2031,N_2753);
and U3808 (N_3808,N_2004,N_2471);
and U3809 (N_3809,N_2968,N_2598);
or U3810 (N_3810,N_2364,N_2604);
and U3811 (N_3811,N_2769,N_2319);
nor U3812 (N_3812,N_2194,N_2864);
and U3813 (N_3813,N_2410,N_2718);
nand U3814 (N_3814,N_2779,N_2084);
nand U3815 (N_3815,N_2767,N_2255);
nand U3816 (N_3816,N_2405,N_2109);
nand U3817 (N_3817,N_2624,N_2774);
nor U3818 (N_3818,N_2426,N_2110);
and U3819 (N_3819,N_2248,N_2222);
nor U3820 (N_3820,N_2991,N_2191);
nor U3821 (N_3821,N_2196,N_2646);
nand U3822 (N_3822,N_2958,N_2071);
or U3823 (N_3823,N_2816,N_2739);
xnor U3824 (N_3824,N_2959,N_2389);
or U3825 (N_3825,N_2982,N_2244);
nor U3826 (N_3826,N_2345,N_2523);
and U3827 (N_3827,N_2184,N_2582);
nand U3828 (N_3828,N_2138,N_2243);
or U3829 (N_3829,N_2987,N_2087);
and U3830 (N_3830,N_2271,N_2728);
or U3831 (N_3831,N_2925,N_2393);
and U3832 (N_3832,N_2772,N_2672);
and U3833 (N_3833,N_2431,N_2476);
and U3834 (N_3834,N_2293,N_2500);
xor U3835 (N_3835,N_2714,N_2744);
or U3836 (N_3836,N_2760,N_2878);
and U3837 (N_3837,N_2154,N_2881);
nor U3838 (N_3838,N_2626,N_2362);
nand U3839 (N_3839,N_2888,N_2233);
nor U3840 (N_3840,N_2247,N_2231);
and U3841 (N_3841,N_2355,N_2144);
and U3842 (N_3842,N_2702,N_2734);
nor U3843 (N_3843,N_2237,N_2085);
xor U3844 (N_3844,N_2391,N_2935);
xnor U3845 (N_3845,N_2313,N_2721);
nand U3846 (N_3846,N_2989,N_2345);
and U3847 (N_3847,N_2079,N_2647);
or U3848 (N_3848,N_2262,N_2503);
nor U3849 (N_3849,N_2892,N_2063);
nand U3850 (N_3850,N_2310,N_2209);
nand U3851 (N_3851,N_2566,N_2073);
nand U3852 (N_3852,N_2570,N_2488);
or U3853 (N_3853,N_2114,N_2799);
and U3854 (N_3854,N_2992,N_2955);
xnor U3855 (N_3855,N_2200,N_2500);
or U3856 (N_3856,N_2279,N_2805);
nand U3857 (N_3857,N_2609,N_2349);
and U3858 (N_3858,N_2303,N_2968);
nor U3859 (N_3859,N_2295,N_2731);
nor U3860 (N_3860,N_2765,N_2441);
or U3861 (N_3861,N_2365,N_2280);
nor U3862 (N_3862,N_2211,N_2330);
xor U3863 (N_3863,N_2821,N_2049);
nor U3864 (N_3864,N_2191,N_2862);
xor U3865 (N_3865,N_2523,N_2809);
nor U3866 (N_3866,N_2437,N_2796);
nor U3867 (N_3867,N_2847,N_2900);
and U3868 (N_3868,N_2977,N_2159);
nand U3869 (N_3869,N_2495,N_2276);
nand U3870 (N_3870,N_2975,N_2754);
xnor U3871 (N_3871,N_2950,N_2805);
and U3872 (N_3872,N_2964,N_2043);
nor U3873 (N_3873,N_2591,N_2635);
nand U3874 (N_3874,N_2955,N_2404);
nand U3875 (N_3875,N_2444,N_2164);
or U3876 (N_3876,N_2615,N_2705);
nor U3877 (N_3877,N_2837,N_2228);
and U3878 (N_3878,N_2870,N_2137);
xnor U3879 (N_3879,N_2477,N_2256);
and U3880 (N_3880,N_2136,N_2976);
or U3881 (N_3881,N_2795,N_2201);
xnor U3882 (N_3882,N_2868,N_2905);
nor U3883 (N_3883,N_2054,N_2415);
and U3884 (N_3884,N_2358,N_2823);
nor U3885 (N_3885,N_2742,N_2848);
nor U3886 (N_3886,N_2414,N_2788);
and U3887 (N_3887,N_2476,N_2957);
nor U3888 (N_3888,N_2264,N_2550);
nand U3889 (N_3889,N_2844,N_2662);
nor U3890 (N_3890,N_2375,N_2708);
and U3891 (N_3891,N_2836,N_2424);
nor U3892 (N_3892,N_2569,N_2020);
nor U3893 (N_3893,N_2497,N_2206);
nand U3894 (N_3894,N_2584,N_2519);
or U3895 (N_3895,N_2189,N_2197);
nor U3896 (N_3896,N_2081,N_2364);
and U3897 (N_3897,N_2326,N_2328);
nor U3898 (N_3898,N_2630,N_2666);
nor U3899 (N_3899,N_2744,N_2538);
and U3900 (N_3900,N_2428,N_2120);
nor U3901 (N_3901,N_2070,N_2996);
nor U3902 (N_3902,N_2325,N_2700);
or U3903 (N_3903,N_2359,N_2256);
and U3904 (N_3904,N_2128,N_2642);
and U3905 (N_3905,N_2838,N_2505);
nand U3906 (N_3906,N_2837,N_2929);
xor U3907 (N_3907,N_2999,N_2023);
xnor U3908 (N_3908,N_2893,N_2709);
nand U3909 (N_3909,N_2115,N_2986);
and U3910 (N_3910,N_2052,N_2318);
and U3911 (N_3911,N_2714,N_2756);
or U3912 (N_3912,N_2579,N_2877);
and U3913 (N_3913,N_2988,N_2349);
and U3914 (N_3914,N_2812,N_2033);
nand U3915 (N_3915,N_2514,N_2595);
nand U3916 (N_3916,N_2331,N_2655);
or U3917 (N_3917,N_2226,N_2233);
xor U3918 (N_3918,N_2196,N_2220);
and U3919 (N_3919,N_2591,N_2878);
or U3920 (N_3920,N_2562,N_2564);
and U3921 (N_3921,N_2571,N_2568);
nand U3922 (N_3922,N_2442,N_2589);
or U3923 (N_3923,N_2888,N_2513);
nand U3924 (N_3924,N_2568,N_2547);
xor U3925 (N_3925,N_2070,N_2724);
nor U3926 (N_3926,N_2790,N_2824);
nor U3927 (N_3927,N_2137,N_2842);
nand U3928 (N_3928,N_2674,N_2505);
or U3929 (N_3929,N_2139,N_2027);
nand U3930 (N_3930,N_2814,N_2399);
nand U3931 (N_3931,N_2420,N_2683);
nor U3932 (N_3932,N_2315,N_2334);
and U3933 (N_3933,N_2718,N_2782);
or U3934 (N_3934,N_2606,N_2873);
xnor U3935 (N_3935,N_2709,N_2473);
or U3936 (N_3936,N_2180,N_2020);
or U3937 (N_3937,N_2610,N_2219);
or U3938 (N_3938,N_2789,N_2549);
or U3939 (N_3939,N_2932,N_2505);
nand U3940 (N_3940,N_2822,N_2784);
and U3941 (N_3941,N_2392,N_2005);
or U3942 (N_3942,N_2883,N_2016);
nor U3943 (N_3943,N_2932,N_2472);
xnor U3944 (N_3944,N_2508,N_2465);
and U3945 (N_3945,N_2873,N_2044);
and U3946 (N_3946,N_2232,N_2983);
nand U3947 (N_3947,N_2799,N_2146);
and U3948 (N_3948,N_2373,N_2681);
nand U3949 (N_3949,N_2463,N_2875);
nor U3950 (N_3950,N_2645,N_2982);
nor U3951 (N_3951,N_2262,N_2387);
nor U3952 (N_3952,N_2261,N_2203);
xnor U3953 (N_3953,N_2401,N_2708);
or U3954 (N_3954,N_2428,N_2763);
or U3955 (N_3955,N_2000,N_2567);
xnor U3956 (N_3956,N_2956,N_2659);
or U3957 (N_3957,N_2044,N_2941);
and U3958 (N_3958,N_2709,N_2326);
xor U3959 (N_3959,N_2531,N_2370);
nor U3960 (N_3960,N_2433,N_2666);
nand U3961 (N_3961,N_2460,N_2157);
or U3962 (N_3962,N_2028,N_2558);
or U3963 (N_3963,N_2890,N_2390);
nand U3964 (N_3964,N_2757,N_2326);
nor U3965 (N_3965,N_2618,N_2539);
and U3966 (N_3966,N_2598,N_2251);
and U3967 (N_3967,N_2508,N_2961);
or U3968 (N_3968,N_2311,N_2304);
nor U3969 (N_3969,N_2389,N_2560);
nor U3970 (N_3970,N_2151,N_2829);
or U3971 (N_3971,N_2633,N_2272);
and U3972 (N_3972,N_2358,N_2803);
nand U3973 (N_3973,N_2752,N_2046);
and U3974 (N_3974,N_2248,N_2140);
and U3975 (N_3975,N_2880,N_2473);
xor U3976 (N_3976,N_2261,N_2812);
and U3977 (N_3977,N_2804,N_2670);
or U3978 (N_3978,N_2057,N_2273);
and U3979 (N_3979,N_2973,N_2724);
and U3980 (N_3980,N_2969,N_2261);
or U3981 (N_3981,N_2007,N_2696);
nand U3982 (N_3982,N_2495,N_2738);
and U3983 (N_3983,N_2939,N_2094);
nand U3984 (N_3984,N_2003,N_2507);
or U3985 (N_3985,N_2069,N_2126);
xnor U3986 (N_3986,N_2932,N_2251);
and U3987 (N_3987,N_2279,N_2266);
or U3988 (N_3988,N_2171,N_2187);
and U3989 (N_3989,N_2039,N_2933);
nand U3990 (N_3990,N_2538,N_2688);
xnor U3991 (N_3991,N_2979,N_2016);
xor U3992 (N_3992,N_2776,N_2120);
and U3993 (N_3993,N_2055,N_2458);
nor U3994 (N_3994,N_2227,N_2797);
nand U3995 (N_3995,N_2283,N_2453);
or U3996 (N_3996,N_2605,N_2920);
and U3997 (N_3997,N_2390,N_2071);
nand U3998 (N_3998,N_2730,N_2636);
or U3999 (N_3999,N_2353,N_2838);
or U4000 (N_4000,N_3771,N_3321);
nor U4001 (N_4001,N_3862,N_3107);
nor U4002 (N_4002,N_3911,N_3625);
or U4003 (N_4003,N_3880,N_3653);
or U4004 (N_4004,N_3474,N_3543);
nand U4005 (N_4005,N_3071,N_3858);
or U4006 (N_4006,N_3808,N_3641);
or U4007 (N_4007,N_3832,N_3831);
and U4008 (N_4008,N_3667,N_3461);
nand U4009 (N_4009,N_3523,N_3914);
nor U4010 (N_4010,N_3773,N_3782);
nand U4011 (N_4011,N_3665,N_3293);
nand U4012 (N_4012,N_3567,N_3555);
nor U4013 (N_4013,N_3256,N_3556);
nor U4014 (N_4014,N_3302,N_3372);
and U4015 (N_4015,N_3851,N_3693);
and U4016 (N_4016,N_3162,N_3766);
xnor U4017 (N_4017,N_3136,N_3134);
nor U4018 (N_4018,N_3888,N_3675);
and U4019 (N_4019,N_3287,N_3092);
nand U4020 (N_4020,N_3096,N_3337);
and U4021 (N_4021,N_3339,N_3307);
nand U4022 (N_4022,N_3102,N_3030);
nor U4023 (N_4023,N_3519,N_3809);
xnor U4024 (N_4024,N_3342,N_3769);
xnor U4025 (N_4025,N_3963,N_3095);
nor U4026 (N_4026,N_3229,N_3081);
or U4027 (N_4027,N_3724,N_3278);
nor U4028 (N_4028,N_3195,N_3261);
and U4029 (N_4029,N_3300,N_3944);
nor U4030 (N_4030,N_3252,N_3750);
or U4031 (N_4031,N_3871,N_3759);
nand U4032 (N_4032,N_3251,N_3082);
nand U4033 (N_4033,N_3013,N_3715);
or U4034 (N_4034,N_3466,N_3617);
xor U4035 (N_4035,N_3920,N_3786);
xnor U4036 (N_4036,N_3838,N_3646);
nand U4037 (N_4037,N_3533,N_3717);
nand U4038 (N_4038,N_3046,N_3634);
nor U4039 (N_4039,N_3507,N_3189);
or U4040 (N_4040,N_3159,N_3311);
and U4041 (N_4041,N_3805,N_3345);
nand U4042 (N_4042,N_3070,N_3012);
or U4043 (N_4043,N_3131,N_3062);
or U4044 (N_4044,N_3089,N_3347);
or U4045 (N_4045,N_3719,N_3577);
nor U4046 (N_4046,N_3129,N_3812);
or U4047 (N_4047,N_3488,N_3177);
nand U4048 (N_4048,N_3609,N_3649);
or U4049 (N_4049,N_3643,N_3192);
and U4050 (N_4050,N_3975,N_3432);
nand U4051 (N_4051,N_3363,N_3670);
or U4052 (N_4052,N_3477,N_3040);
nor U4053 (N_4053,N_3591,N_3420);
nand U4054 (N_4054,N_3542,N_3493);
xor U4055 (N_4055,N_3984,N_3268);
nand U4056 (N_4056,N_3530,N_3451);
or U4057 (N_4057,N_3502,N_3018);
or U4058 (N_4058,N_3428,N_3978);
nor U4059 (N_4059,N_3020,N_3566);
nand U4060 (N_4060,N_3601,N_3448);
and U4061 (N_4061,N_3032,N_3811);
or U4062 (N_4062,N_3043,N_3604);
or U4063 (N_4063,N_3970,N_3789);
and U4064 (N_4064,N_3411,N_3352);
and U4065 (N_4065,N_3000,N_3234);
and U4066 (N_4066,N_3708,N_3343);
nor U4067 (N_4067,N_3045,N_3479);
nand U4068 (N_4068,N_3657,N_3151);
nor U4069 (N_4069,N_3833,N_3796);
nor U4070 (N_4070,N_3740,N_3517);
and U4071 (N_4071,N_3156,N_3438);
and U4072 (N_4072,N_3351,N_3205);
or U4073 (N_4073,N_3338,N_3763);
xor U4074 (N_4074,N_3024,N_3679);
nand U4075 (N_4075,N_3879,N_3385);
xor U4076 (N_4076,N_3623,N_3377);
nor U4077 (N_4077,N_3235,N_3168);
and U4078 (N_4078,N_3494,N_3931);
or U4079 (N_4079,N_3607,N_3481);
or U4080 (N_4080,N_3050,N_3768);
and U4081 (N_4081,N_3854,N_3619);
xnor U4082 (N_4082,N_3285,N_3837);
nor U4083 (N_4083,N_3696,N_3439);
nor U4084 (N_4084,N_3305,N_3605);
or U4085 (N_4085,N_3584,N_3611);
and U4086 (N_4086,N_3572,N_3153);
and U4087 (N_4087,N_3335,N_3928);
xnor U4088 (N_4088,N_3721,N_3125);
nor U4089 (N_4089,N_3262,N_3797);
and U4090 (N_4090,N_3067,N_3196);
or U4091 (N_4091,N_3425,N_3840);
and U4092 (N_4092,N_3830,N_3937);
and U4093 (N_4093,N_3441,N_3956);
and U4094 (N_4094,N_3506,N_3224);
xnor U4095 (N_4095,N_3402,N_3829);
nand U4096 (N_4096,N_3462,N_3201);
and U4097 (N_4097,N_3473,N_3558);
xor U4098 (N_4098,N_3689,N_3650);
nand U4099 (N_4099,N_3539,N_3254);
nor U4100 (N_4100,N_3424,N_3645);
nand U4101 (N_4101,N_3207,N_3265);
and U4102 (N_4102,N_3968,N_3714);
or U4103 (N_4103,N_3144,N_3846);
nand U4104 (N_4104,N_3504,N_3765);
nand U4105 (N_4105,N_3427,N_3048);
nor U4106 (N_4106,N_3999,N_3915);
nor U4107 (N_4107,N_3280,N_3110);
xnor U4108 (N_4108,N_3528,N_3757);
or U4109 (N_4109,N_3158,N_3482);
xor U4110 (N_4110,N_3529,N_3998);
nor U4111 (N_4111,N_3817,N_3487);
nand U4112 (N_4112,N_3957,N_3686);
nor U4113 (N_4113,N_3974,N_3097);
or U4114 (N_4114,N_3222,N_3713);
nand U4115 (N_4115,N_3329,N_3250);
nor U4116 (N_4116,N_3258,N_3510);
and U4117 (N_4117,N_3374,N_3866);
and U4118 (N_4118,N_3935,N_3722);
nor U4119 (N_4119,N_3575,N_3867);
nand U4120 (N_4120,N_3630,N_3171);
xnor U4121 (N_4121,N_3106,N_3274);
nor U4122 (N_4122,N_3035,N_3170);
nor U4123 (N_4123,N_3631,N_3692);
or U4124 (N_4124,N_3146,N_3899);
and U4125 (N_4125,N_3112,N_3085);
or U4126 (N_4126,N_3232,N_3264);
nor U4127 (N_4127,N_3340,N_3108);
nand U4128 (N_4128,N_3676,N_3615);
nand U4129 (N_4129,N_3036,N_3279);
nand U4130 (N_4130,N_3289,N_3621);
xnor U4131 (N_4131,N_3620,N_3955);
nor U4132 (N_4132,N_3313,N_3799);
and U4133 (N_4133,N_3728,N_3739);
nand U4134 (N_4134,N_3359,N_3415);
and U4135 (N_4135,N_3301,N_3516);
or U4136 (N_4136,N_3038,N_3044);
nor U4137 (N_4137,N_3027,N_3456);
nand U4138 (N_4138,N_3560,N_3749);
and U4139 (N_4139,N_3225,N_3009);
nand U4140 (N_4140,N_3291,N_3212);
nand U4141 (N_4141,N_3354,N_3988);
and U4142 (N_4142,N_3981,N_3864);
nor U4143 (N_4143,N_3730,N_3476);
and U4144 (N_4144,N_3094,N_3458);
nand U4145 (N_4145,N_3319,N_3820);
and U4146 (N_4146,N_3122,N_3348);
and U4147 (N_4147,N_3698,N_3105);
xor U4148 (N_4148,N_3016,N_3685);
and U4149 (N_4149,N_3671,N_3887);
xnor U4150 (N_4150,N_3148,N_3467);
nor U4151 (N_4151,N_3794,N_3894);
nand U4152 (N_4152,N_3142,N_3564);
and U4153 (N_4153,N_3227,N_3622);
and U4154 (N_4154,N_3169,N_3160);
nand U4155 (N_4155,N_3384,N_3953);
and U4156 (N_4156,N_3248,N_3612);
nor U4157 (N_4157,N_3497,N_3901);
xnor U4158 (N_4158,N_3541,N_3525);
nor U4159 (N_4159,N_3892,N_3545);
nand U4160 (N_4160,N_3104,N_3677);
xor U4161 (N_4161,N_3720,N_3025);
and U4162 (N_4162,N_3538,N_3752);
nor U4163 (N_4163,N_3632,N_3777);
nor U4164 (N_4164,N_3513,N_3190);
nor U4165 (N_4165,N_3404,N_3128);
nor U4166 (N_4166,N_3309,N_3526);
or U4167 (N_4167,N_3961,N_3276);
nand U4168 (N_4168,N_3578,N_3852);
nand U4169 (N_4169,N_3221,N_3783);
nand U4170 (N_4170,N_3996,N_3850);
or U4171 (N_4171,N_3270,N_3853);
and U4172 (N_4172,N_3760,N_3198);
and U4173 (N_4173,N_3945,N_3163);
and U4174 (N_4174,N_3772,N_3660);
or U4175 (N_4175,N_3336,N_3491);
nand U4176 (N_4176,N_3596,N_3369);
xnor U4177 (N_4177,N_3006,N_3551);
nor U4178 (N_4178,N_3445,N_3465);
xor U4179 (N_4179,N_3399,N_3091);
nor U4180 (N_4180,N_3303,N_3930);
and U4181 (N_4181,N_3073,N_3554);
nand U4182 (N_4182,N_3470,N_3845);
nor U4183 (N_4183,N_3534,N_3992);
or U4184 (N_4184,N_3063,N_3787);
nand U4185 (N_4185,N_3921,N_3580);
xnor U4186 (N_4186,N_3848,N_3594);
or U4187 (N_4187,N_3100,N_3536);
or U4188 (N_4188,N_3219,N_3994);
nand U4189 (N_4189,N_3614,N_3124);
or U4190 (N_4190,N_3468,N_3946);
nand U4191 (N_4191,N_3241,N_3599);
nor U4192 (N_4192,N_3193,N_3231);
nor U4193 (N_4193,N_3127,N_3903);
or U4194 (N_4194,N_3544,N_3881);
nor U4195 (N_4195,N_3446,N_3877);
xnor U4196 (N_4196,N_3678,N_3098);
xnor U4197 (N_4197,N_3332,N_3496);
nor U4198 (N_4198,N_3857,N_3403);
and U4199 (N_4199,N_3985,N_3767);
xor U4200 (N_4200,N_3725,N_3712);
nand U4201 (N_4201,N_3120,N_3793);
nand U4202 (N_4202,N_3362,N_3115);
and U4203 (N_4203,N_3865,N_3933);
nand U4204 (N_4204,N_3346,N_3426);
and U4205 (N_4205,N_3795,N_3015);
or U4206 (N_4206,N_3531,N_3639);
xor U4207 (N_4207,N_3898,N_3041);
or U4208 (N_4208,N_3977,N_3989);
xnor U4209 (N_4209,N_3061,N_3075);
xor U4210 (N_4210,N_3029,N_3316);
nor U4211 (N_4211,N_3272,N_3701);
nor U4212 (N_4212,N_3825,N_3243);
nor U4213 (N_4213,N_3906,N_3770);
or U4214 (N_4214,N_3469,N_3669);
nor U4215 (N_4215,N_3870,N_3742);
or U4216 (N_4216,N_3618,N_3435);
nor U4217 (N_4217,N_3357,N_3139);
nor U4218 (N_4218,N_3406,N_3246);
or U4219 (N_4219,N_3079,N_3822);
and U4220 (N_4220,N_3801,N_3341);
xnor U4221 (N_4221,N_3932,N_3896);
xor U4222 (N_4222,N_3202,N_3548);
and U4223 (N_4223,N_3306,N_3269);
nand U4224 (N_4224,N_3034,N_3317);
nand U4225 (N_4225,N_3214,N_3668);
and U4226 (N_4226,N_3296,N_3042);
and U4227 (N_4227,N_3421,N_3187);
xor U4228 (N_4228,N_3386,N_3813);
nand U4229 (N_4229,N_3123,N_3064);
nand U4230 (N_4230,N_3113,N_3059);
nand U4231 (N_4231,N_3355,N_3429);
nor U4232 (N_4232,N_3464,N_3520);
nand U4233 (N_4233,N_3155,N_3382);
and U4234 (N_4234,N_3400,N_3026);
or U4235 (N_4235,N_3966,N_3133);
and U4236 (N_4236,N_3731,N_3109);
or U4237 (N_4237,N_3051,N_3226);
and U4238 (N_4238,N_3925,N_3590);
xor U4239 (N_4239,N_3310,N_3360);
xor U4240 (N_4240,N_3373,N_3138);
or U4241 (N_4241,N_3288,N_3707);
and U4242 (N_4242,N_3705,N_3052);
nand U4243 (N_4243,N_3947,N_3764);
or U4244 (N_4244,N_3856,N_3500);
or U4245 (N_4245,N_3281,N_3674);
and U4246 (N_4246,N_3616,N_3242);
or U4247 (N_4247,N_3283,N_3489);
or U4248 (N_4248,N_3353,N_3188);
xnor U4249 (N_4249,N_3819,N_3778);
nand U4250 (N_4250,N_3077,N_3726);
nand U4251 (N_4251,N_3861,N_3565);
or U4252 (N_4252,N_3943,N_3613);
nand U4253 (N_4253,N_3217,N_3074);
xnor U4254 (N_4254,N_3333,N_3185);
nand U4255 (N_4255,N_3495,N_3640);
and U4256 (N_4256,N_3552,N_3878);
nand U4257 (N_4257,N_3602,N_3397);
nor U4258 (N_4258,N_3121,N_3501);
or U4259 (N_4259,N_3161,N_3508);
or U4260 (N_4260,N_3271,N_3883);
or U4261 (N_4261,N_3798,N_3290);
xnor U4262 (N_4262,N_3150,N_3732);
or U4263 (N_4263,N_3413,N_3304);
nor U4264 (N_4264,N_3628,N_3587);
or U4265 (N_4265,N_3320,N_3068);
or U4266 (N_4266,N_3266,N_3367);
or U4267 (N_4267,N_3755,N_3563);
nor U4268 (N_4268,N_3758,N_3747);
and U4269 (N_4269,N_3648,N_3093);
and U4270 (N_4270,N_3003,N_3284);
and U4271 (N_4271,N_3659,N_3550);
nor U4272 (N_4272,N_3983,N_3330);
nor U4273 (N_4273,N_3736,N_3573);
xnor U4274 (N_4274,N_3661,N_3691);
nor U4275 (N_4275,N_3005,N_3130);
nor U4276 (N_4276,N_3637,N_3200);
and U4277 (N_4277,N_3282,N_3344);
and U4278 (N_4278,N_3593,N_3084);
nand U4279 (N_4279,N_3512,N_3350);
nand U4280 (N_4280,N_3547,N_3743);
nor U4281 (N_4281,N_3318,N_3328);
xnor U4282 (N_4282,N_3610,N_3595);
and U4283 (N_4283,N_3314,N_3422);
nand U4284 (N_4284,N_3117,N_3509);
nand U4285 (N_4285,N_3066,N_3334);
nand U4286 (N_4286,N_3823,N_3847);
xnor U4287 (N_4287,N_3499,N_3004);
nand U4288 (N_4288,N_3626,N_3804);
and U4289 (N_4289,N_3561,N_3600);
nand U4290 (N_4290,N_3119,N_3603);
nand U4291 (N_4291,N_3080,N_3514);
xnor U4292 (N_4292,N_3588,N_3390);
or U4293 (N_4293,N_3295,N_3941);
nor U4294 (N_4294,N_3598,N_3088);
xnor U4295 (N_4295,N_3680,N_3203);
nor U4296 (N_4296,N_3371,N_3821);
and U4297 (N_4297,N_3748,N_3729);
nand U4298 (N_4298,N_3902,N_3886);
nand U4299 (N_4299,N_3849,N_3683);
or U4300 (N_4300,N_3802,N_3298);
nor U4301 (N_4301,N_3292,N_3518);
and U4302 (N_4302,N_3065,N_3228);
nand U4303 (N_4303,N_3002,N_3909);
nand U4304 (N_4304,N_3206,N_3568);
nor U4305 (N_4305,N_3391,N_3450);
nor U4306 (N_4306,N_3718,N_3672);
xor U4307 (N_4307,N_3021,N_3788);
xnor U4308 (N_4308,N_3299,N_3037);
and U4309 (N_4309,N_3987,N_3746);
and U4310 (N_4310,N_3559,N_3960);
and U4311 (N_4311,N_3204,N_3405);
and U4312 (N_4312,N_3826,N_3140);
xor U4313 (N_4313,N_3267,N_3055);
nand U4314 (N_4314,N_3836,N_3485);
nand U4315 (N_4315,N_3913,N_3498);
nor U4316 (N_4316,N_3194,N_3664);
nor U4317 (N_4317,N_3452,N_3257);
nor U4318 (N_4318,N_3690,N_3841);
and U4319 (N_4319,N_3597,N_3331);
or U4320 (N_4320,N_3997,N_3761);
nand U4321 (N_4321,N_3608,N_3019);
nor U4322 (N_4322,N_3143,N_3582);
or U4323 (N_4323,N_3638,N_3173);
or U4324 (N_4324,N_3900,N_3135);
and U4325 (N_4325,N_3023,N_3855);
and U4326 (N_4326,N_3358,N_3844);
and U4327 (N_4327,N_3907,N_3443);
or U4328 (N_4328,N_3924,N_3751);
or U4329 (N_4329,N_3401,N_3815);
nand U4330 (N_4330,N_3741,N_3629);
or U4331 (N_4331,N_3964,N_3753);
or U4332 (N_4332,N_3408,N_3286);
nand U4333 (N_4333,N_3581,N_3571);
nor U4334 (N_4334,N_3001,N_3430);
and U4335 (N_4335,N_3735,N_3380);
and U4336 (N_4336,N_3209,N_3392);
nor U4337 (N_4337,N_3532,N_3505);
nor U4338 (N_4338,N_3673,N_3586);
and U4339 (N_4339,N_3215,N_3118);
and U4340 (N_4340,N_3835,N_3436);
xor U4341 (N_4341,N_3375,N_3263);
or U4342 (N_4342,N_3967,N_3585);
nor U4343 (N_4343,N_3434,N_3076);
nor U4344 (N_4344,N_3583,N_3549);
xnor U4345 (N_4345,N_3694,N_3323);
and U4346 (N_4346,N_3570,N_3368);
or U4347 (N_4347,N_3260,N_3174);
nor U4348 (N_4348,N_3412,N_3398);
and U4349 (N_4349,N_3651,N_3954);
and U4350 (N_4350,N_3240,N_3882);
or U4351 (N_4351,N_3463,N_3167);
xnor U4352 (N_4352,N_3184,N_3972);
nor U4353 (N_4353,N_3475,N_3927);
nor U4354 (N_4354,N_3860,N_3383);
nor U4355 (N_4355,N_3060,N_3951);
or U4356 (N_4356,N_3654,N_3589);
nand U4357 (N_4357,N_3624,N_3255);
xor U4358 (N_4358,N_3010,N_3917);
and U4359 (N_4359,N_3410,N_3175);
nand U4360 (N_4360,N_3447,N_3387);
or U4361 (N_4361,N_3535,N_3419);
or U4362 (N_4362,N_3103,N_3982);
or U4363 (N_4363,N_3950,N_3165);
and U4364 (N_4364,N_3524,N_3949);
nand U4365 (N_4365,N_3039,N_3433);
xnor U4366 (N_4366,N_3157,N_3111);
xnor U4367 (N_4367,N_3592,N_3546);
nor U4368 (N_4368,N_3365,N_3014);
nand U4369 (N_4369,N_3409,N_3483);
nand U4370 (N_4370,N_3275,N_3440);
or U4371 (N_4371,N_3008,N_3503);
nand U4372 (N_4372,N_3868,N_3775);
or U4373 (N_4373,N_3457,N_3810);
nor U4374 (N_4374,N_3416,N_3356);
and U4375 (N_4375,N_3414,N_3239);
nand U4376 (N_4376,N_3576,N_3484);
or U4377 (N_4377,N_3049,N_3366);
xnor U4378 (N_4378,N_3893,N_3197);
and U4379 (N_4379,N_3557,N_3993);
and U4380 (N_4380,N_3181,N_3942);
nor U4381 (N_4381,N_3897,N_3486);
nor U4382 (N_4382,N_3824,N_3172);
nand U4383 (N_4383,N_3253,N_3948);
nand U4384 (N_4384,N_3431,N_3273);
nor U4385 (N_4385,N_3969,N_3114);
nor U4386 (N_4386,N_3918,N_3297);
nor U4387 (N_4387,N_3976,N_3863);
nor U4388 (N_4388,N_3929,N_3449);
and U4389 (N_4389,N_3223,N_3381);
nand U4390 (N_4390,N_3213,N_3521);
nand U4391 (N_4391,N_3723,N_3734);
nor U4392 (N_4392,N_3635,N_3540);
xnor U4393 (N_4393,N_3818,N_3791);
or U4394 (N_4394,N_3827,N_3727);
or U4395 (N_4395,N_3912,N_3069);
and U4396 (N_4396,N_3908,N_3326);
nand U4397 (N_4397,N_3574,N_3806);
or U4398 (N_4398,N_3843,N_3378);
nand U4399 (N_4399,N_3834,N_3986);
and U4400 (N_4400,N_3078,N_3182);
and U4401 (N_4401,N_3472,N_3176);
nand U4402 (N_4402,N_3703,N_3249);
or U4403 (N_4403,N_3396,N_3057);
xor U4404 (N_4404,N_3774,N_3816);
nor U4405 (N_4405,N_3839,N_3460);
nand U4406 (N_4406,N_3706,N_3453);
nor U4407 (N_4407,N_3859,N_3756);
and U4408 (N_4408,N_3754,N_3154);
nand U4409 (N_4409,N_3022,N_3058);
and U4410 (N_4410,N_3238,N_3145);
xnor U4411 (N_4411,N_3166,N_3697);
or U4412 (N_4412,N_3803,N_3511);
and U4413 (N_4413,N_3733,N_3418);
or U4414 (N_4414,N_3562,N_3247);
and U4415 (N_4415,N_3776,N_3872);
and U4416 (N_4416,N_3031,N_3388);
and U4417 (N_4417,N_3186,N_3642);
xnor U4418 (N_4418,N_3349,N_3308);
nand U4419 (N_4419,N_3370,N_3407);
nand U4420 (N_4420,N_3393,N_3889);
nor U4421 (N_4421,N_3979,N_3716);
nand U4422 (N_4422,N_3442,N_3710);
or U4423 (N_4423,N_3666,N_3905);
nand U4424 (N_4424,N_3086,N_3245);
nor U4425 (N_4425,N_3444,N_3910);
and U4426 (N_4426,N_3828,N_3965);
or U4427 (N_4427,N_3737,N_3785);
and U4428 (N_4428,N_3047,N_3938);
and U4429 (N_4429,N_3934,N_3962);
xnor U4430 (N_4430,N_3904,N_3379);
nor U4431 (N_4431,N_3191,N_3952);
nand U4432 (N_4432,N_3980,N_3790);
and U4433 (N_4433,N_3515,N_3395);
nand U4434 (N_4434,N_3149,N_3033);
and U4435 (N_4435,N_3738,N_3922);
nor U4436 (N_4436,N_3394,N_3842);
and U4437 (N_4437,N_3216,N_3807);
or U4438 (N_4438,N_3180,N_3211);
nor U4439 (N_4439,N_3210,N_3876);
nand U4440 (N_4440,N_3312,N_3417);
nor U4441 (N_4441,N_3579,N_3711);
or U4442 (N_4442,N_3147,N_3325);
nand U4443 (N_4443,N_3480,N_3990);
and U4444 (N_4444,N_3891,N_3814);
or U4445 (N_4445,N_3152,N_3662);
xor U4446 (N_4446,N_3315,N_3101);
xnor U4447 (N_4447,N_3361,N_3681);
and U4448 (N_4448,N_3244,N_3087);
nor U4449 (N_4449,N_3800,N_3655);
nor U4450 (N_4450,N_3874,N_3537);
and U4451 (N_4451,N_3569,N_3090);
nor U4452 (N_4452,N_3490,N_3183);
and U4453 (N_4453,N_3164,N_3884);
nand U4454 (N_4454,N_3873,N_3700);
or U4455 (N_4455,N_3017,N_3199);
and U4456 (N_4456,N_3885,N_3423);
or U4457 (N_4457,N_3895,N_3784);
and U4458 (N_4458,N_3652,N_3437);
and U4459 (N_4459,N_3455,N_3959);
or U4460 (N_4460,N_3277,N_3656);
nand U4461 (N_4461,N_3940,N_3792);
or U4462 (N_4462,N_3324,N_3072);
nor U4463 (N_4463,N_3553,N_3083);
or U4464 (N_4464,N_3178,N_3237);
and U4465 (N_4465,N_3126,N_3471);
or U4466 (N_4466,N_3606,N_3364);
nand U4467 (N_4467,N_3699,N_3702);
nand U4468 (N_4468,N_3663,N_3230);
nand U4469 (N_4469,N_3054,N_3633);
nor U4470 (N_4470,N_3522,N_3688);
and U4471 (N_4471,N_3053,N_3208);
or U4472 (N_4472,N_3971,N_3919);
or U4473 (N_4473,N_3762,N_3695);
or U4474 (N_4474,N_3939,N_3916);
nor U4475 (N_4475,N_3220,N_3007);
nand U4476 (N_4476,N_3644,N_3647);
nor U4477 (N_4477,N_3991,N_3099);
nand U4478 (N_4478,N_3236,N_3869);
or U4479 (N_4479,N_3322,N_3958);
and U4480 (N_4480,N_3875,N_3137);
nand U4481 (N_4481,N_3627,N_3923);
nor U4482 (N_4482,N_3492,N_3926);
nand U4483 (N_4483,N_3056,N_3779);
nand U4484 (N_4484,N_3995,N_3781);
and U4485 (N_4485,N_3218,N_3780);
nor U4486 (N_4486,N_3454,N_3259);
or U4487 (N_4487,N_3745,N_3116);
or U4488 (N_4488,N_3704,N_3011);
xnor U4489 (N_4489,N_3294,N_3684);
or U4490 (N_4490,N_3744,N_3233);
xor U4491 (N_4491,N_3028,N_3682);
and U4492 (N_4492,N_3687,N_3527);
or U4493 (N_4493,N_3179,N_3459);
and U4494 (N_4494,N_3709,N_3132);
nor U4495 (N_4495,N_3327,N_3890);
nor U4496 (N_4496,N_3636,N_3658);
or U4497 (N_4497,N_3478,N_3389);
nor U4498 (N_4498,N_3936,N_3141);
and U4499 (N_4499,N_3973,N_3376);
and U4500 (N_4500,N_3737,N_3579);
nor U4501 (N_4501,N_3168,N_3248);
or U4502 (N_4502,N_3571,N_3376);
xnor U4503 (N_4503,N_3380,N_3818);
or U4504 (N_4504,N_3801,N_3128);
and U4505 (N_4505,N_3076,N_3296);
xor U4506 (N_4506,N_3344,N_3899);
nor U4507 (N_4507,N_3969,N_3098);
nand U4508 (N_4508,N_3658,N_3626);
and U4509 (N_4509,N_3932,N_3015);
nor U4510 (N_4510,N_3369,N_3290);
nor U4511 (N_4511,N_3540,N_3527);
and U4512 (N_4512,N_3112,N_3104);
nand U4513 (N_4513,N_3660,N_3742);
xnor U4514 (N_4514,N_3900,N_3409);
nor U4515 (N_4515,N_3550,N_3288);
or U4516 (N_4516,N_3300,N_3738);
or U4517 (N_4517,N_3281,N_3663);
xnor U4518 (N_4518,N_3883,N_3471);
nand U4519 (N_4519,N_3674,N_3105);
xnor U4520 (N_4520,N_3410,N_3606);
nand U4521 (N_4521,N_3854,N_3591);
xor U4522 (N_4522,N_3786,N_3110);
or U4523 (N_4523,N_3145,N_3764);
xor U4524 (N_4524,N_3408,N_3748);
nand U4525 (N_4525,N_3807,N_3626);
nor U4526 (N_4526,N_3192,N_3005);
or U4527 (N_4527,N_3075,N_3661);
nor U4528 (N_4528,N_3201,N_3544);
nor U4529 (N_4529,N_3012,N_3175);
nor U4530 (N_4530,N_3787,N_3189);
or U4531 (N_4531,N_3688,N_3254);
and U4532 (N_4532,N_3947,N_3255);
and U4533 (N_4533,N_3409,N_3237);
or U4534 (N_4534,N_3572,N_3264);
nor U4535 (N_4535,N_3402,N_3305);
nor U4536 (N_4536,N_3360,N_3408);
or U4537 (N_4537,N_3045,N_3756);
and U4538 (N_4538,N_3004,N_3799);
xor U4539 (N_4539,N_3460,N_3736);
nor U4540 (N_4540,N_3047,N_3086);
and U4541 (N_4541,N_3172,N_3860);
nand U4542 (N_4542,N_3446,N_3264);
xor U4543 (N_4543,N_3200,N_3290);
and U4544 (N_4544,N_3174,N_3044);
xor U4545 (N_4545,N_3653,N_3800);
xnor U4546 (N_4546,N_3684,N_3016);
or U4547 (N_4547,N_3941,N_3483);
and U4548 (N_4548,N_3460,N_3141);
nor U4549 (N_4549,N_3739,N_3035);
or U4550 (N_4550,N_3456,N_3532);
nand U4551 (N_4551,N_3548,N_3752);
and U4552 (N_4552,N_3624,N_3362);
nor U4553 (N_4553,N_3274,N_3356);
nand U4554 (N_4554,N_3511,N_3213);
nand U4555 (N_4555,N_3228,N_3691);
nand U4556 (N_4556,N_3648,N_3646);
or U4557 (N_4557,N_3775,N_3733);
and U4558 (N_4558,N_3901,N_3599);
or U4559 (N_4559,N_3889,N_3218);
xor U4560 (N_4560,N_3087,N_3335);
or U4561 (N_4561,N_3238,N_3509);
nand U4562 (N_4562,N_3930,N_3323);
or U4563 (N_4563,N_3579,N_3971);
or U4564 (N_4564,N_3183,N_3904);
nor U4565 (N_4565,N_3596,N_3106);
and U4566 (N_4566,N_3069,N_3643);
or U4567 (N_4567,N_3253,N_3188);
nand U4568 (N_4568,N_3464,N_3188);
nor U4569 (N_4569,N_3459,N_3881);
and U4570 (N_4570,N_3869,N_3924);
nor U4571 (N_4571,N_3410,N_3032);
and U4572 (N_4572,N_3475,N_3365);
nor U4573 (N_4573,N_3055,N_3804);
nor U4574 (N_4574,N_3921,N_3851);
nor U4575 (N_4575,N_3897,N_3410);
xnor U4576 (N_4576,N_3917,N_3088);
nor U4577 (N_4577,N_3417,N_3949);
nor U4578 (N_4578,N_3142,N_3330);
xnor U4579 (N_4579,N_3157,N_3014);
xnor U4580 (N_4580,N_3451,N_3676);
or U4581 (N_4581,N_3608,N_3924);
nand U4582 (N_4582,N_3911,N_3028);
nor U4583 (N_4583,N_3061,N_3806);
or U4584 (N_4584,N_3960,N_3682);
nand U4585 (N_4585,N_3142,N_3240);
nor U4586 (N_4586,N_3085,N_3957);
xor U4587 (N_4587,N_3776,N_3787);
or U4588 (N_4588,N_3218,N_3857);
and U4589 (N_4589,N_3729,N_3862);
nor U4590 (N_4590,N_3954,N_3349);
nand U4591 (N_4591,N_3352,N_3486);
nand U4592 (N_4592,N_3599,N_3922);
and U4593 (N_4593,N_3903,N_3063);
nand U4594 (N_4594,N_3746,N_3605);
and U4595 (N_4595,N_3844,N_3326);
nand U4596 (N_4596,N_3114,N_3957);
or U4597 (N_4597,N_3395,N_3652);
and U4598 (N_4598,N_3601,N_3282);
and U4599 (N_4599,N_3550,N_3794);
and U4600 (N_4600,N_3868,N_3178);
nand U4601 (N_4601,N_3743,N_3227);
nor U4602 (N_4602,N_3553,N_3404);
or U4603 (N_4603,N_3054,N_3444);
nand U4604 (N_4604,N_3235,N_3843);
and U4605 (N_4605,N_3961,N_3095);
or U4606 (N_4606,N_3531,N_3856);
xnor U4607 (N_4607,N_3328,N_3741);
nand U4608 (N_4608,N_3940,N_3320);
nor U4609 (N_4609,N_3373,N_3890);
or U4610 (N_4610,N_3321,N_3251);
and U4611 (N_4611,N_3763,N_3660);
nand U4612 (N_4612,N_3332,N_3012);
and U4613 (N_4613,N_3413,N_3230);
nand U4614 (N_4614,N_3091,N_3705);
nand U4615 (N_4615,N_3171,N_3983);
nand U4616 (N_4616,N_3284,N_3768);
xor U4617 (N_4617,N_3869,N_3651);
and U4618 (N_4618,N_3209,N_3707);
nand U4619 (N_4619,N_3215,N_3796);
or U4620 (N_4620,N_3126,N_3006);
xor U4621 (N_4621,N_3309,N_3478);
nor U4622 (N_4622,N_3866,N_3048);
nor U4623 (N_4623,N_3472,N_3185);
nor U4624 (N_4624,N_3279,N_3524);
nor U4625 (N_4625,N_3066,N_3866);
and U4626 (N_4626,N_3829,N_3488);
xnor U4627 (N_4627,N_3632,N_3173);
nor U4628 (N_4628,N_3692,N_3406);
nand U4629 (N_4629,N_3966,N_3501);
or U4630 (N_4630,N_3453,N_3963);
xnor U4631 (N_4631,N_3926,N_3660);
xor U4632 (N_4632,N_3445,N_3588);
or U4633 (N_4633,N_3770,N_3351);
nand U4634 (N_4634,N_3720,N_3365);
and U4635 (N_4635,N_3463,N_3740);
or U4636 (N_4636,N_3533,N_3850);
nor U4637 (N_4637,N_3256,N_3216);
or U4638 (N_4638,N_3677,N_3374);
nand U4639 (N_4639,N_3895,N_3468);
and U4640 (N_4640,N_3599,N_3970);
nor U4641 (N_4641,N_3050,N_3258);
xor U4642 (N_4642,N_3873,N_3444);
nor U4643 (N_4643,N_3155,N_3214);
nand U4644 (N_4644,N_3849,N_3730);
or U4645 (N_4645,N_3172,N_3193);
and U4646 (N_4646,N_3546,N_3018);
or U4647 (N_4647,N_3338,N_3825);
xor U4648 (N_4648,N_3703,N_3841);
and U4649 (N_4649,N_3091,N_3387);
xnor U4650 (N_4650,N_3747,N_3589);
nor U4651 (N_4651,N_3765,N_3923);
nor U4652 (N_4652,N_3870,N_3097);
nor U4653 (N_4653,N_3547,N_3307);
nand U4654 (N_4654,N_3858,N_3544);
or U4655 (N_4655,N_3951,N_3654);
and U4656 (N_4656,N_3486,N_3025);
nor U4657 (N_4657,N_3576,N_3176);
or U4658 (N_4658,N_3853,N_3133);
nand U4659 (N_4659,N_3551,N_3425);
nor U4660 (N_4660,N_3808,N_3930);
nand U4661 (N_4661,N_3223,N_3213);
and U4662 (N_4662,N_3141,N_3125);
nand U4663 (N_4663,N_3038,N_3215);
nand U4664 (N_4664,N_3146,N_3571);
and U4665 (N_4665,N_3459,N_3096);
and U4666 (N_4666,N_3811,N_3431);
nor U4667 (N_4667,N_3970,N_3779);
or U4668 (N_4668,N_3888,N_3834);
nand U4669 (N_4669,N_3241,N_3632);
and U4670 (N_4670,N_3590,N_3568);
nor U4671 (N_4671,N_3975,N_3244);
nor U4672 (N_4672,N_3709,N_3189);
xnor U4673 (N_4673,N_3148,N_3656);
or U4674 (N_4674,N_3343,N_3882);
nor U4675 (N_4675,N_3240,N_3420);
nor U4676 (N_4676,N_3050,N_3437);
nand U4677 (N_4677,N_3237,N_3873);
or U4678 (N_4678,N_3492,N_3191);
and U4679 (N_4679,N_3879,N_3289);
xor U4680 (N_4680,N_3863,N_3176);
and U4681 (N_4681,N_3843,N_3326);
nor U4682 (N_4682,N_3520,N_3582);
or U4683 (N_4683,N_3929,N_3349);
and U4684 (N_4684,N_3926,N_3467);
xor U4685 (N_4685,N_3388,N_3046);
nand U4686 (N_4686,N_3309,N_3776);
nand U4687 (N_4687,N_3160,N_3320);
nand U4688 (N_4688,N_3131,N_3821);
or U4689 (N_4689,N_3068,N_3533);
and U4690 (N_4690,N_3348,N_3976);
or U4691 (N_4691,N_3916,N_3690);
nand U4692 (N_4692,N_3028,N_3355);
nor U4693 (N_4693,N_3680,N_3623);
and U4694 (N_4694,N_3325,N_3698);
and U4695 (N_4695,N_3143,N_3573);
nand U4696 (N_4696,N_3062,N_3000);
or U4697 (N_4697,N_3974,N_3502);
or U4698 (N_4698,N_3830,N_3693);
or U4699 (N_4699,N_3028,N_3300);
and U4700 (N_4700,N_3746,N_3367);
or U4701 (N_4701,N_3672,N_3964);
and U4702 (N_4702,N_3319,N_3133);
nand U4703 (N_4703,N_3638,N_3100);
nand U4704 (N_4704,N_3666,N_3096);
and U4705 (N_4705,N_3238,N_3068);
and U4706 (N_4706,N_3945,N_3739);
nand U4707 (N_4707,N_3404,N_3935);
nor U4708 (N_4708,N_3168,N_3707);
nand U4709 (N_4709,N_3250,N_3650);
and U4710 (N_4710,N_3335,N_3504);
nor U4711 (N_4711,N_3261,N_3659);
nand U4712 (N_4712,N_3254,N_3513);
xnor U4713 (N_4713,N_3858,N_3862);
nand U4714 (N_4714,N_3166,N_3142);
nand U4715 (N_4715,N_3069,N_3001);
nor U4716 (N_4716,N_3152,N_3785);
and U4717 (N_4717,N_3259,N_3530);
nor U4718 (N_4718,N_3807,N_3549);
or U4719 (N_4719,N_3513,N_3976);
or U4720 (N_4720,N_3458,N_3422);
nor U4721 (N_4721,N_3425,N_3993);
nand U4722 (N_4722,N_3801,N_3103);
and U4723 (N_4723,N_3268,N_3817);
and U4724 (N_4724,N_3065,N_3344);
nand U4725 (N_4725,N_3071,N_3309);
or U4726 (N_4726,N_3604,N_3827);
and U4727 (N_4727,N_3143,N_3429);
and U4728 (N_4728,N_3249,N_3182);
nand U4729 (N_4729,N_3861,N_3249);
and U4730 (N_4730,N_3577,N_3438);
and U4731 (N_4731,N_3461,N_3005);
nand U4732 (N_4732,N_3592,N_3141);
or U4733 (N_4733,N_3971,N_3486);
nor U4734 (N_4734,N_3664,N_3511);
or U4735 (N_4735,N_3413,N_3864);
and U4736 (N_4736,N_3403,N_3914);
nor U4737 (N_4737,N_3900,N_3269);
nor U4738 (N_4738,N_3747,N_3783);
and U4739 (N_4739,N_3106,N_3703);
and U4740 (N_4740,N_3679,N_3216);
nand U4741 (N_4741,N_3468,N_3058);
nand U4742 (N_4742,N_3323,N_3295);
or U4743 (N_4743,N_3508,N_3475);
and U4744 (N_4744,N_3522,N_3929);
and U4745 (N_4745,N_3668,N_3554);
and U4746 (N_4746,N_3965,N_3873);
nor U4747 (N_4747,N_3304,N_3429);
and U4748 (N_4748,N_3539,N_3625);
and U4749 (N_4749,N_3889,N_3940);
nor U4750 (N_4750,N_3223,N_3856);
and U4751 (N_4751,N_3268,N_3605);
nor U4752 (N_4752,N_3571,N_3901);
or U4753 (N_4753,N_3641,N_3760);
and U4754 (N_4754,N_3955,N_3504);
xor U4755 (N_4755,N_3564,N_3973);
or U4756 (N_4756,N_3245,N_3851);
or U4757 (N_4757,N_3085,N_3966);
and U4758 (N_4758,N_3439,N_3068);
or U4759 (N_4759,N_3581,N_3346);
and U4760 (N_4760,N_3799,N_3215);
nand U4761 (N_4761,N_3169,N_3526);
xnor U4762 (N_4762,N_3693,N_3954);
and U4763 (N_4763,N_3269,N_3168);
and U4764 (N_4764,N_3227,N_3056);
or U4765 (N_4765,N_3448,N_3283);
xor U4766 (N_4766,N_3376,N_3455);
and U4767 (N_4767,N_3667,N_3899);
nand U4768 (N_4768,N_3191,N_3430);
or U4769 (N_4769,N_3670,N_3604);
and U4770 (N_4770,N_3777,N_3443);
nor U4771 (N_4771,N_3627,N_3753);
and U4772 (N_4772,N_3221,N_3908);
and U4773 (N_4773,N_3234,N_3194);
nor U4774 (N_4774,N_3266,N_3080);
nor U4775 (N_4775,N_3948,N_3327);
nor U4776 (N_4776,N_3796,N_3770);
and U4777 (N_4777,N_3785,N_3881);
or U4778 (N_4778,N_3292,N_3266);
and U4779 (N_4779,N_3232,N_3817);
nor U4780 (N_4780,N_3039,N_3782);
and U4781 (N_4781,N_3565,N_3763);
and U4782 (N_4782,N_3872,N_3117);
nor U4783 (N_4783,N_3176,N_3416);
nor U4784 (N_4784,N_3352,N_3359);
or U4785 (N_4785,N_3242,N_3247);
nor U4786 (N_4786,N_3173,N_3864);
nor U4787 (N_4787,N_3415,N_3578);
nand U4788 (N_4788,N_3696,N_3301);
nor U4789 (N_4789,N_3709,N_3615);
or U4790 (N_4790,N_3286,N_3815);
nand U4791 (N_4791,N_3605,N_3299);
and U4792 (N_4792,N_3677,N_3902);
nand U4793 (N_4793,N_3970,N_3051);
nand U4794 (N_4794,N_3386,N_3501);
or U4795 (N_4795,N_3937,N_3076);
or U4796 (N_4796,N_3480,N_3627);
nor U4797 (N_4797,N_3485,N_3120);
nand U4798 (N_4798,N_3568,N_3198);
nand U4799 (N_4799,N_3047,N_3489);
nor U4800 (N_4800,N_3250,N_3442);
nand U4801 (N_4801,N_3135,N_3976);
nor U4802 (N_4802,N_3431,N_3543);
or U4803 (N_4803,N_3498,N_3593);
and U4804 (N_4804,N_3146,N_3396);
and U4805 (N_4805,N_3592,N_3624);
and U4806 (N_4806,N_3844,N_3765);
and U4807 (N_4807,N_3882,N_3708);
or U4808 (N_4808,N_3255,N_3416);
nor U4809 (N_4809,N_3290,N_3757);
or U4810 (N_4810,N_3972,N_3489);
nor U4811 (N_4811,N_3173,N_3521);
nand U4812 (N_4812,N_3316,N_3255);
nor U4813 (N_4813,N_3153,N_3320);
nand U4814 (N_4814,N_3954,N_3893);
or U4815 (N_4815,N_3431,N_3747);
or U4816 (N_4816,N_3855,N_3832);
nand U4817 (N_4817,N_3067,N_3408);
nor U4818 (N_4818,N_3036,N_3309);
or U4819 (N_4819,N_3747,N_3122);
nand U4820 (N_4820,N_3787,N_3002);
nand U4821 (N_4821,N_3472,N_3587);
nand U4822 (N_4822,N_3346,N_3377);
nor U4823 (N_4823,N_3756,N_3326);
nand U4824 (N_4824,N_3544,N_3760);
or U4825 (N_4825,N_3936,N_3892);
nand U4826 (N_4826,N_3670,N_3771);
nand U4827 (N_4827,N_3212,N_3783);
nand U4828 (N_4828,N_3189,N_3543);
nand U4829 (N_4829,N_3583,N_3785);
nor U4830 (N_4830,N_3410,N_3294);
nand U4831 (N_4831,N_3289,N_3766);
or U4832 (N_4832,N_3733,N_3249);
or U4833 (N_4833,N_3722,N_3952);
nand U4834 (N_4834,N_3275,N_3917);
nand U4835 (N_4835,N_3023,N_3789);
xnor U4836 (N_4836,N_3922,N_3981);
and U4837 (N_4837,N_3141,N_3269);
nor U4838 (N_4838,N_3312,N_3805);
nand U4839 (N_4839,N_3117,N_3940);
nand U4840 (N_4840,N_3930,N_3425);
nor U4841 (N_4841,N_3351,N_3212);
nor U4842 (N_4842,N_3463,N_3609);
nor U4843 (N_4843,N_3274,N_3096);
nor U4844 (N_4844,N_3136,N_3234);
xnor U4845 (N_4845,N_3837,N_3711);
nor U4846 (N_4846,N_3832,N_3759);
nor U4847 (N_4847,N_3859,N_3337);
nand U4848 (N_4848,N_3338,N_3608);
or U4849 (N_4849,N_3028,N_3510);
nor U4850 (N_4850,N_3313,N_3124);
nor U4851 (N_4851,N_3391,N_3952);
and U4852 (N_4852,N_3419,N_3809);
xor U4853 (N_4853,N_3119,N_3416);
nand U4854 (N_4854,N_3150,N_3669);
and U4855 (N_4855,N_3049,N_3189);
and U4856 (N_4856,N_3557,N_3130);
nor U4857 (N_4857,N_3304,N_3602);
nor U4858 (N_4858,N_3168,N_3619);
or U4859 (N_4859,N_3149,N_3565);
nor U4860 (N_4860,N_3948,N_3031);
nor U4861 (N_4861,N_3755,N_3712);
xor U4862 (N_4862,N_3932,N_3923);
or U4863 (N_4863,N_3414,N_3997);
nand U4864 (N_4864,N_3497,N_3714);
nand U4865 (N_4865,N_3927,N_3469);
nand U4866 (N_4866,N_3568,N_3028);
nor U4867 (N_4867,N_3228,N_3620);
xnor U4868 (N_4868,N_3938,N_3848);
nand U4869 (N_4869,N_3579,N_3536);
and U4870 (N_4870,N_3628,N_3980);
xnor U4871 (N_4871,N_3518,N_3983);
nand U4872 (N_4872,N_3066,N_3705);
xor U4873 (N_4873,N_3643,N_3868);
nand U4874 (N_4874,N_3566,N_3679);
or U4875 (N_4875,N_3630,N_3871);
or U4876 (N_4876,N_3693,N_3174);
or U4877 (N_4877,N_3941,N_3849);
and U4878 (N_4878,N_3343,N_3912);
nor U4879 (N_4879,N_3071,N_3099);
or U4880 (N_4880,N_3292,N_3763);
nor U4881 (N_4881,N_3261,N_3958);
nand U4882 (N_4882,N_3851,N_3377);
nand U4883 (N_4883,N_3476,N_3598);
nor U4884 (N_4884,N_3456,N_3145);
and U4885 (N_4885,N_3772,N_3512);
nand U4886 (N_4886,N_3347,N_3882);
or U4887 (N_4887,N_3005,N_3972);
and U4888 (N_4888,N_3608,N_3896);
nor U4889 (N_4889,N_3980,N_3487);
nor U4890 (N_4890,N_3890,N_3130);
nor U4891 (N_4891,N_3799,N_3728);
nor U4892 (N_4892,N_3110,N_3370);
nor U4893 (N_4893,N_3528,N_3600);
nor U4894 (N_4894,N_3978,N_3172);
nand U4895 (N_4895,N_3232,N_3555);
nor U4896 (N_4896,N_3525,N_3914);
nand U4897 (N_4897,N_3613,N_3038);
xnor U4898 (N_4898,N_3502,N_3722);
xor U4899 (N_4899,N_3306,N_3394);
nor U4900 (N_4900,N_3381,N_3888);
nand U4901 (N_4901,N_3565,N_3457);
nor U4902 (N_4902,N_3072,N_3053);
nor U4903 (N_4903,N_3717,N_3438);
and U4904 (N_4904,N_3732,N_3591);
nor U4905 (N_4905,N_3520,N_3588);
or U4906 (N_4906,N_3968,N_3865);
nand U4907 (N_4907,N_3012,N_3577);
and U4908 (N_4908,N_3983,N_3821);
nor U4909 (N_4909,N_3779,N_3277);
xor U4910 (N_4910,N_3561,N_3441);
and U4911 (N_4911,N_3027,N_3510);
nand U4912 (N_4912,N_3211,N_3430);
and U4913 (N_4913,N_3287,N_3900);
nand U4914 (N_4914,N_3937,N_3945);
and U4915 (N_4915,N_3307,N_3030);
or U4916 (N_4916,N_3197,N_3497);
nor U4917 (N_4917,N_3234,N_3072);
xnor U4918 (N_4918,N_3917,N_3204);
and U4919 (N_4919,N_3439,N_3709);
nor U4920 (N_4920,N_3074,N_3774);
nor U4921 (N_4921,N_3516,N_3387);
nor U4922 (N_4922,N_3083,N_3994);
nor U4923 (N_4923,N_3658,N_3572);
and U4924 (N_4924,N_3948,N_3632);
nor U4925 (N_4925,N_3985,N_3325);
or U4926 (N_4926,N_3620,N_3898);
xor U4927 (N_4927,N_3724,N_3782);
and U4928 (N_4928,N_3103,N_3579);
nand U4929 (N_4929,N_3624,N_3906);
nor U4930 (N_4930,N_3716,N_3747);
xnor U4931 (N_4931,N_3302,N_3066);
nor U4932 (N_4932,N_3275,N_3479);
nor U4933 (N_4933,N_3047,N_3295);
and U4934 (N_4934,N_3310,N_3507);
xor U4935 (N_4935,N_3861,N_3856);
nor U4936 (N_4936,N_3576,N_3465);
nand U4937 (N_4937,N_3469,N_3668);
nor U4938 (N_4938,N_3802,N_3631);
and U4939 (N_4939,N_3121,N_3186);
or U4940 (N_4940,N_3343,N_3416);
nand U4941 (N_4941,N_3022,N_3804);
or U4942 (N_4942,N_3942,N_3854);
or U4943 (N_4943,N_3606,N_3680);
nand U4944 (N_4944,N_3358,N_3964);
and U4945 (N_4945,N_3155,N_3340);
nor U4946 (N_4946,N_3598,N_3585);
nor U4947 (N_4947,N_3463,N_3275);
nand U4948 (N_4948,N_3741,N_3106);
xor U4949 (N_4949,N_3491,N_3360);
nor U4950 (N_4950,N_3653,N_3537);
nand U4951 (N_4951,N_3006,N_3998);
nand U4952 (N_4952,N_3820,N_3541);
or U4953 (N_4953,N_3820,N_3219);
and U4954 (N_4954,N_3829,N_3778);
and U4955 (N_4955,N_3306,N_3760);
nand U4956 (N_4956,N_3404,N_3874);
and U4957 (N_4957,N_3890,N_3817);
and U4958 (N_4958,N_3385,N_3387);
nand U4959 (N_4959,N_3025,N_3302);
nor U4960 (N_4960,N_3815,N_3549);
or U4961 (N_4961,N_3240,N_3840);
nor U4962 (N_4962,N_3127,N_3228);
or U4963 (N_4963,N_3582,N_3137);
or U4964 (N_4964,N_3258,N_3759);
nand U4965 (N_4965,N_3828,N_3744);
nor U4966 (N_4966,N_3313,N_3350);
nor U4967 (N_4967,N_3303,N_3921);
or U4968 (N_4968,N_3882,N_3425);
nor U4969 (N_4969,N_3395,N_3513);
and U4970 (N_4970,N_3142,N_3719);
nor U4971 (N_4971,N_3872,N_3119);
or U4972 (N_4972,N_3205,N_3294);
or U4973 (N_4973,N_3738,N_3174);
nand U4974 (N_4974,N_3712,N_3866);
nand U4975 (N_4975,N_3926,N_3218);
nand U4976 (N_4976,N_3401,N_3726);
or U4977 (N_4977,N_3474,N_3546);
nand U4978 (N_4978,N_3523,N_3805);
or U4979 (N_4979,N_3677,N_3237);
nand U4980 (N_4980,N_3147,N_3941);
nand U4981 (N_4981,N_3332,N_3114);
or U4982 (N_4982,N_3770,N_3206);
and U4983 (N_4983,N_3381,N_3727);
nand U4984 (N_4984,N_3264,N_3820);
nor U4985 (N_4985,N_3984,N_3509);
nor U4986 (N_4986,N_3336,N_3892);
nand U4987 (N_4987,N_3591,N_3879);
and U4988 (N_4988,N_3873,N_3323);
nor U4989 (N_4989,N_3146,N_3448);
or U4990 (N_4990,N_3205,N_3968);
nand U4991 (N_4991,N_3577,N_3848);
xnor U4992 (N_4992,N_3488,N_3274);
nor U4993 (N_4993,N_3645,N_3731);
or U4994 (N_4994,N_3403,N_3439);
nand U4995 (N_4995,N_3034,N_3745);
and U4996 (N_4996,N_3363,N_3889);
or U4997 (N_4997,N_3531,N_3241);
nand U4998 (N_4998,N_3799,N_3741);
nand U4999 (N_4999,N_3405,N_3089);
nor U5000 (N_5000,N_4568,N_4247);
or U5001 (N_5001,N_4779,N_4735);
xnor U5002 (N_5002,N_4418,N_4271);
and U5003 (N_5003,N_4887,N_4209);
and U5004 (N_5004,N_4205,N_4954);
and U5005 (N_5005,N_4280,N_4763);
and U5006 (N_5006,N_4404,N_4594);
xnor U5007 (N_5007,N_4210,N_4429);
and U5008 (N_5008,N_4761,N_4500);
nor U5009 (N_5009,N_4879,N_4553);
nor U5010 (N_5010,N_4614,N_4387);
xnor U5011 (N_5011,N_4913,N_4499);
or U5012 (N_5012,N_4972,N_4762);
and U5013 (N_5013,N_4377,N_4077);
nand U5014 (N_5014,N_4883,N_4385);
nand U5015 (N_5015,N_4218,N_4263);
nand U5016 (N_5016,N_4923,N_4215);
nor U5017 (N_5017,N_4356,N_4912);
xnor U5018 (N_5018,N_4015,N_4004);
nand U5019 (N_5019,N_4078,N_4283);
and U5020 (N_5020,N_4425,N_4135);
and U5021 (N_5021,N_4213,N_4606);
xor U5022 (N_5022,N_4663,N_4770);
nor U5023 (N_5023,N_4371,N_4650);
nor U5024 (N_5024,N_4460,N_4658);
and U5025 (N_5025,N_4128,N_4997);
and U5026 (N_5026,N_4511,N_4060);
nor U5027 (N_5027,N_4296,N_4054);
nor U5028 (N_5028,N_4829,N_4701);
and U5029 (N_5029,N_4709,N_4345);
or U5030 (N_5030,N_4707,N_4148);
nor U5031 (N_5031,N_4277,N_4091);
or U5032 (N_5032,N_4417,N_4420);
nor U5033 (N_5033,N_4047,N_4502);
nand U5034 (N_5034,N_4375,N_4051);
nor U5035 (N_5035,N_4539,N_4522);
nor U5036 (N_5036,N_4605,N_4619);
nand U5037 (N_5037,N_4145,N_4293);
xor U5038 (N_5038,N_4611,N_4193);
nor U5039 (N_5039,N_4111,N_4916);
or U5040 (N_5040,N_4623,N_4940);
or U5041 (N_5041,N_4463,N_4780);
nor U5042 (N_5042,N_4797,N_4977);
or U5043 (N_5043,N_4299,N_4117);
nand U5044 (N_5044,N_4722,N_4494);
nand U5045 (N_5045,N_4754,N_4931);
nor U5046 (N_5046,N_4328,N_4106);
nand U5047 (N_5047,N_4075,N_4973);
and U5048 (N_5048,N_4851,N_4732);
or U5049 (N_5049,N_4114,N_4358);
nand U5050 (N_5050,N_4581,N_4063);
nor U5051 (N_5051,N_4034,N_4515);
nand U5052 (N_5052,N_4168,N_4011);
nand U5053 (N_5053,N_4101,N_4192);
nor U5054 (N_5054,N_4639,N_4454);
xnor U5055 (N_5055,N_4149,N_4550);
nand U5056 (N_5056,N_4897,N_4486);
nand U5057 (N_5057,N_4187,N_4043);
or U5058 (N_5058,N_4790,N_4451);
and U5059 (N_5059,N_4025,N_4327);
and U5060 (N_5060,N_4881,N_4846);
or U5061 (N_5061,N_4155,N_4690);
nand U5062 (N_5062,N_4428,N_4177);
or U5063 (N_5063,N_4332,N_4092);
or U5064 (N_5064,N_4439,N_4694);
nor U5065 (N_5065,N_4042,N_4932);
nand U5066 (N_5066,N_4033,N_4934);
nor U5067 (N_5067,N_4194,N_4930);
nand U5068 (N_5068,N_4745,N_4396);
and U5069 (N_5069,N_4402,N_4012);
nor U5070 (N_5070,N_4359,N_4131);
xor U5071 (N_5071,N_4340,N_4132);
nand U5072 (N_5072,N_4958,N_4984);
nor U5073 (N_5073,N_4369,N_4264);
nand U5074 (N_5074,N_4862,N_4799);
and U5075 (N_5075,N_4174,N_4507);
nand U5076 (N_5076,N_4180,N_4764);
nor U5077 (N_5077,N_4109,N_4344);
nand U5078 (N_5078,N_4160,N_4250);
and U5079 (N_5079,N_4350,N_4374);
nor U5080 (N_5080,N_4724,N_4102);
or U5081 (N_5081,N_4049,N_4693);
nor U5082 (N_5082,N_4593,N_4217);
xnor U5083 (N_5083,N_4855,N_4580);
nor U5084 (N_5084,N_4538,N_4470);
nor U5085 (N_5085,N_4774,N_4479);
and U5086 (N_5086,N_4309,N_4165);
and U5087 (N_5087,N_4715,N_4083);
nor U5088 (N_5088,N_4617,N_4378);
and U5089 (N_5089,N_4618,N_4186);
xnor U5090 (N_5090,N_4682,N_4680);
and U5091 (N_5091,N_4364,N_4395);
and U5092 (N_5092,N_4508,N_4471);
and U5093 (N_5093,N_4635,N_4727);
nand U5094 (N_5094,N_4927,N_4438);
nor U5095 (N_5095,N_4053,N_4162);
or U5096 (N_5096,N_4864,N_4016);
and U5097 (N_5097,N_4633,N_4274);
and U5098 (N_5098,N_4979,N_4269);
nor U5099 (N_5099,N_4926,N_4182);
nand U5100 (N_5100,N_4554,N_4295);
xnor U5101 (N_5101,N_4133,N_4630);
nor U5102 (N_5102,N_4949,N_4057);
or U5103 (N_5103,N_4459,N_4139);
and U5104 (N_5104,N_4620,N_4873);
nor U5105 (N_5105,N_4349,N_4301);
nand U5106 (N_5106,N_4052,N_4654);
and U5107 (N_5107,N_4272,N_4073);
nand U5108 (N_5108,N_4152,N_4711);
nand U5109 (N_5109,N_4552,N_4670);
and U5110 (N_5110,N_4730,N_4902);
nand U5111 (N_5111,N_4159,N_4223);
or U5112 (N_5112,N_4579,N_4736);
nand U5113 (N_5113,N_4840,N_4390);
or U5114 (N_5114,N_4681,N_4061);
and U5115 (N_5115,N_4172,N_4282);
and U5116 (N_5116,N_4546,N_4408);
nor U5117 (N_5117,N_4523,N_4235);
nand U5118 (N_5118,N_4688,N_4807);
xnor U5119 (N_5119,N_4339,N_4373);
and U5120 (N_5120,N_4006,N_4310);
and U5121 (N_5121,N_4003,N_4585);
nor U5122 (N_5122,N_4288,N_4820);
or U5123 (N_5123,N_4956,N_4305);
or U5124 (N_5124,N_4353,N_4489);
nor U5125 (N_5125,N_4244,N_4826);
nand U5126 (N_5126,N_4007,N_4885);
or U5127 (N_5127,N_4533,N_4386);
nand U5128 (N_5128,N_4298,N_4341);
and U5129 (N_5129,N_4936,N_4184);
nand U5130 (N_5130,N_4222,N_4800);
and U5131 (N_5131,N_4675,N_4360);
nor U5132 (N_5132,N_4590,N_4525);
or U5133 (N_5133,N_4695,N_4857);
and U5134 (N_5134,N_4994,N_4542);
xor U5135 (N_5135,N_4485,N_4937);
or U5136 (N_5136,N_4683,N_4082);
nand U5137 (N_5137,N_4655,N_4225);
nand U5138 (N_5138,N_4260,N_4998);
nor U5139 (N_5139,N_4241,N_4963);
and U5140 (N_5140,N_4607,N_4959);
or U5141 (N_5141,N_4661,N_4944);
and U5142 (N_5142,N_4608,N_4478);
or U5143 (N_5143,N_4738,N_4975);
and U5144 (N_5144,N_4067,N_4400);
nor U5145 (N_5145,N_4725,N_4041);
or U5146 (N_5146,N_4475,N_4397);
nand U5147 (N_5147,N_4817,N_4208);
or U5148 (N_5148,N_4314,N_4803);
nand U5149 (N_5149,N_4498,N_4472);
nor U5150 (N_5150,N_4572,N_4146);
nand U5151 (N_5151,N_4559,N_4316);
or U5152 (N_5152,N_4154,N_4627);
and U5153 (N_5153,N_4018,N_4509);
xor U5154 (N_5154,N_4822,N_4444);
and U5155 (N_5155,N_4104,N_4816);
or U5156 (N_5156,N_4443,N_4772);
or U5157 (N_5157,N_4920,N_4322);
nand U5158 (N_5158,N_4909,N_4878);
nor U5159 (N_5159,N_4136,N_4346);
and U5160 (N_5160,N_4074,N_4370);
xnor U5161 (N_5161,N_4560,N_4547);
and U5162 (N_5162,N_4591,N_4895);
nor U5163 (N_5163,N_4631,N_4905);
nor U5164 (N_5164,N_4477,N_4115);
or U5165 (N_5165,N_4179,N_4189);
nand U5166 (N_5166,N_4610,N_4548);
nor U5167 (N_5167,N_4896,N_4206);
and U5168 (N_5168,N_4935,N_4423);
and U5169 (N_5169,N_4445,N_4870);
nand U5170 (N_5170,N_4888,N_4535);
and U5171 (N_5171,N_4586,N_4563);
or U5172 (N_5172,N_4048,N_4526);
nand U5173 (N_5173,N_4330,N_4524);
nor U5174 (N_5174,N_4775,N_4708);
and U5175 (N_5175,N_4098,N_4512);
nand U5176 (N_5176,N_4584,N_4245);
nand U5177 (N_5177,N_4704,N_4262);
or U5178 (N_5178,N_4231,N_4796);
nand U5179 (N_5179,N_4466,N_4939);
nand U5180 (N_5180,N_4363,N_4990);
xor U5181 (N_5181,N_4794,N_4137);
or U5182 (N_5182,N_4352,N_4384);
and U5183 (N_5183,N_4992,N_4859);
or U5184 (N_5184,N_4519,N_4424);
nand U5185 (N_5185,N_4326,N_4827);
nand U5186 (N_5186,N_4233,N_4838);
or U5187 (N_5187,N_4672,N_4592);
and U5188 (N_5188,N_4853,N_4457);
nand U5189 (N_5189,N_4306,N_4642);
nand U5190 (N_5190,N_4679,N_4382);
nand U5191 (N_5191,N_4516,N_4410);
or U5192 (N_5192,N_4334,N_4718);
or U5193 (N_5193,N_4839,N_4333);
nand U5194 (N_5194,N_4153,N_4000);
or U5195 (N_5195,N_4664,N_4232);
and U5196 (N_5196,N_4029,N_4294);
nand U5197 (N_5197,N_4786,N_4157);
and U5198 (N_5198,N_4988,N_4687);
or U5199 (N_5199,N_4776,N_4481);
or U5200 (N_5200,N_4125,N_4831);
xnor U5201 (N_5201,N_4270,N_4211);
nand U5202 (N_5202,N_4464,N_4120);
nand U5203 (N_5203,N_4268,N_4996);
and U5204 (N_5204,N_4907,N_4965);
xor U5205 (N_5205,N_4532,N_4910);
nor U5206 (N_5206,N_4957,N_4170);
or U5207 (N_5207,N_4318,N_4414);
and U5208 (N_5208,N_4791,N_4604);
nor U5209 (N_5209,N_4151,N_4781);
or U5210 (N_5210,N_4228,N_4456);
or U5211 (N_5211,N_4976,N_4666);
nor U5212 (N_5212,N_4520,N_4876);
xnor U5213 (N_5213,N_4014,N_4068);
nand U5214 (N_5214,N_4837,N_4452);
and U5215 (N_5215,N_4698,N_4933);
xnor U5216 (N_5216,N_4224,N_4582);
and U5217 (N_5217,N_4758,N_4219);
or U5218 (N_5218,N_4141,N_4094);
or U5219 (N_5219,N_4742,N_4230);
and U5220 (N_5220,N_4178,N_4482);
and U5221 (N_5221,N_4928,N_4026);
and U5222 (N_5222,N_4615,N_4372);
nand U5223 (N_5223,N_4760,N_4238);
nand U5224 (N_5224,N_4551,N_4882);
nand U5225 (N_5225,N_4834,N_4565);
nor U5226 (N_5226,N_4300,N_4336);
or U5227 (N_5227,N_4678,N_4122);
nor U5228 (N_5228,N_4324,N_4804);
nor U5229 (N_5229,N_4024,N_4064);
nor U5230 (N_5230,N_4038,N_4496);
or U5231 (N_5231,N_4573,N_4942);
and U5232 (N_5232,N_4901,N_4951);
and U5233 (N_5233,N_4046,N_4468);
and U5234 (N_5234,N_4719,N_4662);
nor U5235 (N_5235,N_4616,N_4032);
nand U5236 (N_5236,N_4440,N_4304);
xnor U5237 (N_5237,N_4313,N_4773);
and U5238 (N_5238,N_4929,N_4097);
nor U5239 (N_5239,N_4828,N_4571);
or U5240 (N_5240,N_4562,N_4648);
or U5241 (N_5241,N_4970,N_4710);
or U5242 (N_5242,N_4811,N_4134);
and U5243 (N_5243,N_4065,N_4924);
xor U5244 (N_5244,N_4626,N_4124);
and U5245 (N_5245,N_4070,N_4379);
and U5246 (N_5246,N_4214,N_4045);
nand U5247 (N_5247,N_4376,N_4766);
nor U5248 (N_5248,N_4971,N_4530);
and U5249 (N_5249,N_4892,N_4081);
nand U5250 (N_5250,N_4596,N_4394);
nand U5251 (N_5251,N_4487,N_4506);
and U5252 (N_5252,N_4845,N_4432);
and U5253 (N_5253,N_4380,N_4854);
and U5254 (N_5254,N_4389,N_4981);
xnor U5255 (N_5255,N_4634,N_4557);
nor U5256 (N_5256,N_4815,N_4001);
nand U5257 (N_5257,N_4891,N_4598);
nor U5258 (N_5258,N_4700,N_4023);
nand U5259 (N_5259,N_4351,N_4292);
nor U5260 (N_5260,N_4802,N_4455);
nand U5261 (N_5261,N_4069,N_4315);
nor U5262 (N_5262,N_4521,N_4647);
or U5263 (N_5263,N_4713,N_4676);
xnor U5264 (N_5264,N_4798,N_4289);
or U5265 (N_5265,N_4628,N_4656);
xnor U5266 (N_5266,N_4028,N_4792);
and U5267 (N_5267,N_4961,N_4201);
xnor U5268 (N_5268,N_4392,N_4777);
nand U5269 (N_5269,N_4302,N_4952);
nor U5270 (N_5270,N_4446,N_4941);
nor U5271 (N_5271,N_4311,N_4699);
nand U5272 (N_5272,N_4113,N_4866);
nor U5273 (N_5273,N_4801,N_4646);
and U5274 (N_5274,N_4393,N_4740);
nor U5275 (N_5275,N_4312,N_4721);
nor U5276 (N_5276,N_4946,N_4555);
xor U5277 (N_5277,N_4103,N_4993);
xor U5278 (N_5278,N_4900,N_4367);
nor U5279 (N_5279,N_4020,N_4756);
and U5280 (N_5280,N_4255,N_4100);
nor U5281 (N_5281,N_4884,N_4469);
nor U5282 (N_5282,N_4729,N_4112);
nor U5283 (N_5283,N_4986,N_4744);
nor U5284 (N_5284,N_4858,N_4651);
and U5285 (N_5285,N_4769,N_4543);
xor U5286 (N_5286,N_4476,N_4355);
and U5287 (N_5287,N_4009,N_4991);
nor U5288 (N_5288,N_4419,N_4207);
and U5289 (N_5289,N_4517,N_4673);
or U5290 (N_5290,N_4583,N_4945);
or U5291 (N_5291,N_4465,N_4911);
nor U5292 (N_5292,N_4757,N_4079);
nand U5293 (N_5293,N_4062,N_4785);
and U5294 (N_5294,N_4196,N_4566);
nand U5295 (N_5295,N_4943,N_4095);
xnor U5296 (N_5296,N_4441,N_4739);
nand U5297 (N_5297,N_4188,N_4158);
and U5298 (N_5298,N_4733,N_4505);
or U5299 (N_5299,N_4747,N_4321);
nor U5300 (N_5300,N_4706,N_4595);
nand U5301 (N_5301,N_4450,N_4434);
nand U5302 (N_5302,N_4613,N_4612);
nor U5303 (N_5303,N_4874,N_4401);
nand U5304 (N_5304,N_4087,N_4629);
nand U5305 (N_5305,N_4677,N_4577);
xnor U5306 (N_5306,N_4253,N_4665);
nor U5307 (N_5307,N_4644,N_4190);
xnor U5308 (N_5308,N_4671,N_4267);
nand U5309 (N_5309,N_4653,N_4484);
and U5310 (N_5310,N_4019,N_4527);
nand U5311 (N_5311,N_4784,N_4836);
and U5312 (N_5312,N_4867,N_4904);
or U5313 (N_5313,N_4567,N_4422);
and U5314 (N_5314,N_4737,N_4863);
nand U5315 (N_5315,N_4812,N_4513);
nor U5316 (N_5316,N_4242,N_4649);
nand U5317 (N_5317,N_4541,N_4751);
or U5318 (N_5318,N_4287,N_4728);
and U5319 (N_5319,N_4461,N_4967);
xnor U5320 (N_5320,N_4495,N_4183);
xnor U5321 (N_5321,N_4251,N_4788);
or U5322 (N_5322,N_4342,N_4175);
and U5323 (N_5323,N_4166,N_4717);
xnor U5324 (N_5324,N_4108,N_4076);
and U5325 (N_5325,N_4435,N_4528);
and U5326 (N_5326,N_4237,N_4437);
nor U5327 (N_5327,N_4399,N_4142);
nor U5328 (N_5328,N_4331,N_4659);
or U5329 (N_5329,N_4147,N_4712);
and U5330 (N_5330,N_4017,N_4265);
nand U5331 (N_5331,N_4685,N_4813);
nand U5332 (N_5332,N_4347,N_4276);
or U5333 (N_5333,N_4197,N_4254);
nand U5334 (N_5334,N_4212,N_4406);
and U5335 (N_5335,N_4323,N_4899);
and U5336 (N_5336,N_4638,N_4969);
or U5337 (N_5337,N_4286,N_4668);
nor U5338 (N_5338,N_4636,N_4221);
nor U5339 (N_5339,N_4752,N_4808);
nand U5340 (N_5340,N_4413,N_4868);
xor U5341 (N_5341,N_4814,N_4398);
nand U5342 (N_5342,N_4167,N_4303);
or U5343 (N_5343,N_4368,N_4692);
and U5344 (N_5344,N_4830,N_4872);
nor U5345 (N_5345,N_4409,N_4039);
nand U5346 (N_5346,N_4066,N_4497);
nor U5347 (N_5347,N_4105,N_4056);
nand U5348 (N_5348,N_4150,N_4116);
nand U5349 (N_5349,N_4609,N_4492);
and U5350 (N_5350,N_4010,N_4403);
nor U5351 (N_5351,N_4603,N_4914);
nand U5352 (N_5352,N_4720,N_4962);
or U5353 (N_5353,N_4258,N_4156);
or U5354 (N_5354,N_4058,N_4714);
nand U5355 (N_5355,N_4204,N_4987);
and U5356 (N_5356,N_4416,N_4096);
xor U5357 (N_5357,N_4447,N_4915);
and U5358 (N_5358,N_4544,N_4411);
or U5359 (N_5359,N_4849,N_4433);
or U5360 (N_5360,N_4691,N_4138);
and U5361 (N_5361,N_4889,N_4273);
nor U5362 (N_5362,N_4259,N_4343);
nand U5363 (N_5363,N_4602,N_4388);
nand U5364 (N_5364,N_4575,N_4749);
nand U5365 (N_5365,N_4285,N_4119);
nor U5366 (N_5366,N_4240,N_4974);
nor U5367 (N_5367,N_4044,N_4275);
nor U5368 (N_5368,N_4036,N_4835);
nor U5369 (N_5369,N_4589,N_4880);
and U5370 (N_5370,N_4391,N_4199);
or U5371 (N_5371,N_4473,N_4906);
nor U5372 (N_5372,N_4667,N_4144);
and U5373 (N_5373,N_4123,N_4234);
and U5374 (N_5374,N_4085,N_4841);
or U5375 (N_5375,N_4697,N_4545);
nand U5376 (N_5376,N_4261,N_4357);
nand U5377 (N_5377,N_4021,N_4966);
and U5378 (N_5378,N_4143,N_4126);
or U5379 (N_5379,N_4436,N_4249);
and U5380 (N_5380,N_4818,N_4964);
xor U5381 (N_5381,N_4462,N_4252);
xnor U5382 (N_5382,N_4317,N_4918);
nand U5383 (N_5383,N_4985,N_4027);
nor U5384 (N_5384,N_4848,N_4850);
nor U5385 (N_5385,N_4319,N_4365);
nand U5386 (N_5386,N_4236,N_4832);
xnor U5387 (N_5387,N_4809,N_4226);
xnor U5388 (N_5388,N_4361,N_4825);
or U5389 (N_5389,N_4989,N_4405);
and U5390 (N_5390,N_4587,N_4643);
or U5391 (N_5391,N_4674,N_4632);
nor U5392 (N_5392,N_4999,N_4787);
nand U5393 (N_5393,N_4257,N_4789);
nor U5394 (N_5394,N_4093,N_4431);
nor U5395 (N_5395,N_4570,N_4622);
and U5396 (N_5396,N_4503,N_4227);
or U5397 (N_5397,N_4229,N_4290);
and U5398 (N_5398,N_4202,N_4002);
and U5399 (N_5399,N_4099,N_4842);
nand U5400 (N_5400,N_4657,N_4856);
xnor U5401 (N_5401,N_4597,N_4163);
or U5402 (N_5402,N_4894,N_4564);
nand U5403 (N_5403,N_4488,N_4427);
or U5404 (N_5404,N_4381,N_4127);
nand U5405 (N_5405,N_4426,N_4040);
nor U5406 (N_5406,N_4338,N_4430);
or U5407 (N_5407,N_4703,N_4448);
nand U5408 (N_5408,N_4953,N_4795);
and U5409 (N_5409,N_4037,N_4248);
nand U5410 (N_5410,N_4746,N_4191);
and U5411 (N_5411,N_4080,N_4759);
nand U5412 (N_5412,N_4195,N_4574);
nand U5413 (N_5413,N_4216,N_4625);
nor U5414 (N_5414,N_4059,N_4534);
nand U5415 (N_5415,N_4705,N_4919);
nand U5416 (N_5416,N_4741,N_4561);
and U5417 (N_5417,N_4569,N_4778);
or U5418 (N_5418,N_4362,N_4600);
xor U5419 (N_5419,N_4161,N_4031);
nand U5420 (N_5420,N_4013,N_4348);
and U5421 (N_5421,N_4453,N_4686);
nand U5422 (N_5422,N_4844,N_4239);
or U5423 (N_5423,N_4491,N_4504);
nand U5424 (N_5424,N_4601,N_4783);
nor U5425 (N_5425,N_4621,N_4514);
nor U5426 (N_5426,N_4140,N_4950);
xnor U5427 (N_5427,N_4805,N_4421);
or U5428 (N_5428,N_4823,N_4980);
xnor U5429 (N_5429,N_4549,N_4118);
nor U5430 (N_5430,N_4893,N_4824);
xor U5431 (N_5431,N_4743,N_4243);
nor U5432 (N_5432,N_4684,N_4947);
or U5433 (N_5433,N_4806,N_4084);
nand U5434 (N_5434,N_4490,N_4198);
xnor U5435 (N_5435,N_4898,N_4983);
nor U5436 (N_5436,N_4022,N_4442);
nand U5437 (N_5437,N_4768,N_4467);
xor U5438 (N_5438,N_4641,N_4917);
nand U5439 (N_5439,N_4702,N_4877);
and U5440 (N_5440,N_4090,N_4576);
and U5441 (N_5441,N_4474,N_4335);
and U5442 (N_5442,N_4458,N_4529);
nand U5443 (N_5443,N_4922,N_4110);
nor U5444 (N_5444,N_4645,N_4320);
nand U5445 (N_5445,N_4246,N_4129);
or U5446 (N_5446,N_4875,N_4086);
nand U5447 (N_5447,N_4734,N_4556);
nor U5448 (N_5448,N_4871,N_4810);
or U5449 (N_5449,N_4329,N_4181);
and U5450 (N_5450,N_4750,N_4696);
and U5451 (N_5451,N_4782,N_4765);
nand U5452 (N_5452,N_4307,N_4860);
or U5453 (N_5453,N_4955,N_4948);
xnor U5454 (N_5454,N_4055,N_4723);
xor U5455 (N_5455,N_4890,N_4088);
or U5456 (N_5456,N_4978,N_4176);
nand U5457 (N_5457,N_4921,N_4624);
or U5458 (N_5458,N_4171,N_4869);
or U5459 (N_5459,N_4726,N_4833);
nor U5460 (N_5460,N_4540,N_4035);
nand U5461 (N_5461,N_4325,N_4030);
nor U5462 (N_5462,N_4903,N_4982);
or U5463 (N_5463,N_4536,N_4995);
or U5464 (N_5464,N_4510,N_4107);
and U5465 (N_5465,N_4925,N_4407);
nand U5466 (N_5466,N_4256,N_4308);
or U5467 (N_5467,N_4960,N_4660);
and U5468 (N_5468,N_4501,N_4767);
and U5469 (N_5469,N_4640,N_4865);
nor U5470 (N_5470,N_4493,N_4480);
nor U5471 (N_5471,N_4281,N_4483);
nor U5472 (N_5472,N_4337,N_4297);
nor U5473 (N_5473,N_4908,N_4449);
or U5474 (N_5474,N_4005,N_4354);
nand U5475 (N_5475,N_4279,N_4968);
and U5476 (N_5476,N_4412,N_4731);
nor U5477 (N_5477,N_4415,N_4130);
nor U5478 (N_5478,N_4121,N_4669);
or U5479 (N_5479,N_4072,N_4383);
nor U5480 (N_5480,N_4793,N_4886);
nor U5481 (N_5481,N_4771,N_4203);
nor U5482 (N_5482,N_4173,N_4220);
or U5483 (N_5483,N_4185,N_4008);
and U5484 (N_5484,N_4819,N_4843);
nor U5485 (N_5485,N_4748,N_4071);
xor U5486 (N_5486,N_4291,N_4821);
or U5487 (N_5487,N_4938,N_4578);
and U5488 (N_5488,N_4278,N_4847);
and U5489 (N_5489,N_4050,N_4861);
or U5490 (N_5490,N_4689,N_4366);
nor U5491 (N_5491,N_4599,N_4755);
nand U5492 (N_5492,N_4716,N_4518);
nand U5493 (N_5493,N_4200,N_4089);
or U5494 (N_5494,N_4588,N_4169);
or U5495 (N_5495,N_4558,N_4266);
nor U5496 (N_5496,N_4537,N_4164);
nor U5497 (N_5497,N_4852,N_4652);
nor U5498 (N_5498,N_4637,N_4753);
nand U5499 (N_5499,N_4531,N_4284);
xor U5500 (N_5500,N_4266,N_4393);
and U5501 (N_5501,N_4342,N_4391);
xor U5502 (N_5502,N_4655,N_4259);
nand U5503 (N_5503,N_4243,N_4909);
nand U5504 (N_5504,N_4767,N_4349);
xnor U5505 (N_5505,N_4961,N_4545);
nand U5506 (N_5506,N_4348,N_4358);
nor U5507 (N_5507,N_4974,N_4660);
nor U5508 (N_5508,N_4679,N_4748);
nor U5509 (N_5509,N_4326,N_4462);
or U5510 (N_5510,N_4444,N_4363);
and U5511 (N_5511,N_4554,N_4765);
and U5512 (N_5512,N_4870,N_4524);
nor U5513 (N_5513,N_4498,N_4994);
nand U5514 (N_5514,N_4232,N_4954);
nor U5515 (N_5515,N_4706,N_4167);
or U5516 (N_5516,N_4562,N_4229);
xnor U5517 (N_5517,N_4656,N_4704);
xor U5518 (N_5518,N_4587,N_4303);
nor U5519 (N_5519,N_4646,N_4206);
nand U5520 (N_5520,N_4789,N_4904);
or U5521 (N_5521,N_4166,N_4176);
and U5522 (N_5522,N_4109,N_4611);
and U5523 (N_5523,N_4607,N_4168);
nor U5524 (N_5524,N_4937,N_4717);
and U5525 (N_5525,N_4660,N_4781);
or U5526 (N_5526,N_4290,N_4746);
or U5527 (N_5527,N_4561,N_4102);
nor U5528 (N_5528,N_4513,N_4629);
nor U5529 (N_5529,N_4009,N_4226);
nand U5530 (N_5530,N_4929,N_4709);
and U5531 (N_5531,N_4734,N_4109);
and U5532 (N_5532,N_4508,N_4498);
nor U5533 (N_5533,N_4705,N_4075);
xor U5534 (N_5534,N_4256,N_4464);
and U5535 (N_5535,N_4881,N_4495);
and U5536 (N_5536,N_4211,N_4847);
nor U5537 (N_5537,N_4674,N_4899);
nand U5538 (N_5538,N_4634,N_4607);
and U5539 (N_5539,N_4370,N_4389);
or U5540 (N_5540,N_4240,N_4686);
nand U5541 (N_5541,N_4843,N_4864);
or U5542 (N_5542,N_4316,N_4996);
or U5543 (N_5543,N_4187,N_4510);
nor U5544 (N_5544,N_4269,N_4148);
nand U5545 (N_5545,N_4925,N_4229);
nand U5546 (N_5546,N_4173,N_4442);
xnor U5547 (N_5547,N_4840,N_4720);
nand U5548 (N_5548,N_4330,N_4476);
or U5549 (N_5549,N_4009,N_4645);
or U5550 (N_5550,N_4775,N_4629);
and U5551 (N_5551,N_4577,N_4934);
xor U5552 (N_5552,N_4843,N_4141);
or U5553 (N_5553,N_4714,N_4642);
and U5554 (N_5554,N_4651,N_4713);
xnor U5555 (N_5555,N_4173,N_4710);
nor U5556 (N_5556,N_4583,N_4879);
and U5557 (N_5557,N_4685,N_4816);
or U5558 (N_5558,N_4662,N_4219);
nand U5559 (N_5559,N_4502,N_4497);
or U5560 (N_5560,N_4142,N_4577);
or U5561 (N_5561,N_4959,N_4851);
xor U5562 (N_5562,N_4846,N_4823);
nor U5563 (N_5563,N_4960,N_4360);
nor U5564 (N_5564,N_4819,N_4739);
or U5565 (N_5565,N_4527,N_4506);
and U5566 (N_5566,N_4849,N_4012);
or U5567 (N_5567,N_4959,N_4632);
nor U5568 (N_5568,N_4478,N_4827);
or U5569 (N_5569,N_4385,N_4486);
and U5570 (N_5570,N_4478,N_4171);
or U5571 (N_5571,N_4414,N_4263);
nor U5572 (N_5572,N_4429,N_4781);
nand U5573 (N_5573,N_4150,N_4614);
nor U5574 (N_5574,N_4461,N_4755);
and U5575 (N_5575,N_4254,N_4582);
and U5576 (N_5576,N_4467,N_4106);
nor U5577 (N_5577,N_4695,N_4980);
and U5578 (N_5578,N_4703,N_4333);
or U5579 (N_5579,N_4222,N_4970);
or U5580 (N_5580,N_4305,N_4496);
or U5581 (N_5581,N_4309,N_4271);
nand U5582 (N_5582,N_4414,N_4077);
or U5583 (N_5583,N_4696,N_4856);
or U5584 (N_5584,N_4004,N_4990);
and U5585 (N_5585,N_4321,N_4579);
nor U5586 (N_5586,N_4370,N_4263);
or U5587 (N_5587,N_4957,N_4529);
and U5588 (N_5588,N_4935,N_4487);
nor U5589 (N_5589,N_4343,N_4141);
or U5590 (N_5590,N_4676,N_4327);
xor U5591 (N_5591,N_4953,N_4267);
nand U5592 (N_5592,N_4326,N_4861);
or U5593 (N_5593,N_4437,N_4092);
nand U5594 (N_5594,N_4281,N_4256);
and U5595 (N_5595,N_4972,N_4623);
nand U5596 (N_5596,N_4804,N_4906);
and U5597 (N_5597,N_4477,N_4692);
and U5598 (N_5598,N_4250,N_4555);
or U5599 (N_5599,N_4443,N_4489);
or U5600 (N_5600,N_4797,N_4449);
nand U5601 (N_5601,N_4668,N_4966);
and U5602 (N_5602,N_4755,N_4004);
nand U5603 (N_5603,N_4789,N_4218);
or U5604 (N_5604,N_4852,N_4904);
or U5605 (N_5605,N_4895,N_4942);
nor U5606 (N_5606,N_4130,N_4511);
nand U5607 (N_5607,N_4827,N_4112);
or U5608 (N_5608,N_4998,N_4294);
or U5609 (N_5609,N_4959,N_4406);
nand U5610 (N_5610,N_4228,N_4607);
nand U5611 (N_5611,N_4574,N_4607);
nor U5612 (N_5612,N_4547,N_4677);
nand U5613 (N_5613,N_4942,N_4518);
and U5614 (N_5614,N_4251,N_4644);
nand U5615 (N_5615,N_4300,N_4944);
nand U5616 (N_5616,N_4313,N_4664);
and U5617 (N_5617,N_4736,N_4793);
nor U5618 (N_5618,N_4921,N_4933);
or U5619 (N_5619,N_4880,N_4888);
xor U5620 (N_5620,N_4610,N_4087);
xnor U5621 (N_5621,N_4085,N_4126);
nor U5622 (N_5622,N_4095,N_4613);
nor U5623 (N_5623,N_4282,N_4830);
nor U5624 (N_5624,N_4704,N_4689);
nand U5625 (N_5625,N_4266,N_4548);
nor U5626 (N_5626,N_4431,N_4222);
or U5627 (N_5627,N_4829,N_4185);
nor U5628 (N_5628,N_4926,N_4773);
nor U5629 (N_5629,N_4262,N_4844);
and U5630 (N_5630,N_4850,N_4329);
nand U5631 (N_5631,N_4211,N_4524);
nand U5632 (N_5632,N_4211,N_4560);
nand U5633 (N_5633,N_4448,N_4650);
xnor U5634 (N_5634,N_4008,N_4242);
nor U5635 (N_5635,N_4081,N_4197);
or U5636 (N_5636,N_4578,N_4182);
nand U5637 (N_5637,N_4500,N_4767);
nor U5638 (N_5638,N_4207,N_4998);
or U5639 (N_5639,N_4420,N_4367);
and U5640 (N_5640,N_4373,N_4780);
nand U5641 (N_5641,N_4151,N_4465);
nand U5642 (N_5642,N_4389,N_4555);
xor U5643 (N_5643,N_4251,N_4150);
and U5644 (N_5644,N_4272,N_4718);
and U5645 (N_5645,N_4975,N_4449);
or U5646 (N_5646,N_4727,N_4618);
nor U5647 (N_5647,N_4235,N_4850);
nor U5648 (N_5648,N_4713,N_4775);
nand U5649 (N_5649,N_4391,N_4849);
or U5650 (N_5650,N_4077,N_4753);
or U5651 (N_5651,N_4275,N_4884);
nand U5652 (N_5652,N_4501,N_4667);
nor U5653 (N_5653,N_4384,N_4624);
xor U5654 (N_5654,N_4079,N_4342);
nand U5655 (N_5655,N_4628,N_4779);
nand U5656 (N_5656,N_4186,N_4206);
nand U5657 (N_5657,N_4030,N_4625);
nor U5658 (N_5658,N_4647,N_4643);
xor U5659 (N_5659,N_4921,N_4948);
and U5660 (N_5660,N_4751,N_4896);
nor U5661 (N_5661,N_4217,N_4556);
and U5662 (N_5662,N_4818,N_4344);
nand U5663 (N_5663,N_4622,N_4893);
nand U5664 (N_5664,N_4256,N_4517);
or U5665 (N_5665,N_4368,N_4303);
and U5666 (N_5666,N_4839,N_4595);
and U5667 (N_5667,N_4158,N_4394);
nand U5668 (N_5668,N_4107,N_4325);
xnor U5669 (N_5669,N_4590,N_4691);
nor U5670 (N_5670,N_4568,N_4548);
nand U5671 (N_5671,N_4643,N_4624);
or U5672 (N_5672,N_4712,N_4116);
nand U5673 (N_5673,N_4941,N_4082);
and U5674 (N_5674,N_4308,N_4320);
and U5675 (N_5675,N_4799,N_4311);
or U5676 (N_5676,N_4116,N_4299);
nand U5677 (N_5677,N_4628,N_4097);
nor U5678 (N_5678,N_4682,N_4055);
or U5679 (N_5679,N_4829,N_4589);
nand U5680 (N_5680,N_4157,N_4425);
and U5681 (N_5681,N_4483,N_4020);
or U5682 (N_5682,N_4913,N_4835);
and U5683 (N_5683,N_4694,N_4946);
nand U5684 (N_5684,N_4303,N_4718);
nand U5685 (N_5685,N_4581,N_4704);
nand U5686 (N_5686,N_4664,N_4437);
nor U5687 (N_5687,N_4527,N_4500);
xnor U5688 (N_5688,N_4728,N_4531);
nor U5689 (N_5689,N_4289,N_4826);
xnor U5690 (N_5690,N_4862,N_4440);
nor U5691 (N_5691,N_4377,N_4836);
or U5692 (N_5692,N_4520,N_4200);
nor U5693 (N_5693,N_4571,N_4310);
nor U5694 (N_5694,N_4430,N_4273);
nand U5695 (N_5695,N_4444,N_4118);
nor U5696 (N_5696,N_4884,N_4212);
xor U5697 (N_5697,N_4552,N_4577);
and U5698 (N_5698,N_4097,N_4129);
nor U5699 (N_5699,N_4284,N_4538);
and U5700 (N_5700,N_4750,N_4172);
and U5701 (N_5701,N_4767,N_4341);
and U5702 (N_5702,N_4956,N_4563);
and U5703 (N_5703,N_4521,N_4471);
nand U5704 (N_5704,N_4746,N_4714);
and U5705 (N_5705,N_4069,N_4764);
or U5706 (N_5706,N_4833,N_4283);
xor U5707 (N_5707,N_4628,N_4875);
and U5708 (N_5708,N_4443,N_4139);
nand U5709 (N_5709,N_4489,N_4289);
nor U5710 (N_5710,N_4736,N_4200);
xor U5711 (N_5711,N_4107,N_4865);
nor U5712 (N_5712,N_4478,N_4632);
or U5713 (N_5713,N_4253,N_4609);
nor U5714 (N_5714,N_4293,N_4400);
and U5715 (N_5715,N_4705,N_4804);
nor U5716 (N_5716,N_4649,N_4407);
or U5717 (N_5717,N_4979,N_4217);
xnor U5718 (N_5718,N_4109,N_4304);
or U5719 (N_5719,N_4659,N_4903);
nor U5720 (N_5720,N_4641,N_4174);
nand U5721 (N_5721,N_4625,N_4911);
or U5722 (N_5722,N_4208,N_4105);
xor U5723 (N_5723,N_4667,N_4098);
nand U5724 (N_5724,N_4287,N_4435);
or U5725 (N_5725,N_4635,N_4511);
nor U5726 (N_5726,N_4549,N_4700);
nor U5727 (N_5727,N_4325,N_4059);
and U5728 (N_5728,N_4336,N_4600);
nor U5729 (N_5729,N_4699,N_4129);
or U5730 (N_5730,N_4159,N_4201);
nand U5731 (N_5731,N_4105,N_4527);
and U5732 (N_5732,N_4416,N_4642);
and U5733 (N_5733,N_4528,N_4805);
or U5734 (N_5734,N_4874,N_4750);
nor U5735 (N_5735,N_4301,N_4375);
and U5736 (N_5736,N_4808,N_4792);
xor U5737 (N_5737,N_4507,N_4350);
nand U5738 (N_5738,N_4561,N_4782);
nand U5739 (N_5739,N_4159,N_4443);
or U5740 (N_5740,N_4009,N_4247);
nand U5741 (N_5741,N_4544,N_4334);
or U5742 (N_5742,N_4255,N_4592);
and U5743 (N_5743,N_4183,N_4774);
and U5744 (N_5744,N_4111,N_4957);
or U5745 (N_5745,N_4024,N_4975);
or U5746 (N_5746,N_4005,N_4621);
nand U5747 (N_5747,N_4582,N_4612);
nor U5748 (N_5748,N_4273,N_4380);
nor U5749 (N_5749,N_4456,N_4230);
or U5750 (N_5750,N_4819,N_4329);
nand U5751 (N_5751,N_4718,N_4267);
nor U5752 (N_5752,N_4297,N_4173);
nand U5753 (N_5753,N_4020,N_4090);
nor U5754 (N_5754,N_4422,N_4857);
nand U5755 (N_5755,N_4059,N_4335);
xnor U5756 (N_5756,N_4756,N_4400);
and U5757 (N_5757,N_4519,N_4087);
nand U5758 (N_5758,N_4322,N_4922);
nand U5759 (N_5759,N_4015,N_4642);
xnor U5760 (N_5760,N_4532,N_4462);
nand U5761 (N_5761,N_4037,N_4131);
nor U5762 (N_5762,N_4813,N_4462);
nor U5763 (N_5763,N_4370,N_4468);
or U5764 (N_5764,N_4262,N_4034);
xor U5765 (N_5765,N_4965,N_4275);
or U5766 (N_5766,N_4398,N_4301);
and U5767 (N_5767,N_4255,N_4817);
or U5768 (N_5768,N_4852,N_4516);
nand U5769 (N_5769,N_4745,N_4561);
nor U5770 (N_5770,N_4352,N_4238);
nand U5771 (N_5771,N_4832,N_4108);
nor U5772 (N_5772,N_4343,N_4959);
nand U5773 (N_5773,N_4447,N_4504);
and U5774 (N_5774,N_4074,N_4823);
and U5775 (N_5775,N_4684,N_4130);
and U5776 (N_5776,N_4132,N_4222);
nor U5777 (N_5777,N_4931,N_4787);
or U5778 (N_5778,N_4702,N_4041);
or U5779 (N_5779,N_4160,N_4104);
and U5780 (N_5780,N_4509,N_4857);
nor U5781 (N_5781,N_4175,N_4757);
or U5782 (N_5782,N_4233,N_4086);
and U5783 (N_5783,N_4944,N_4144);
nor U5784 (N_5784,N_4552,N_4459);
nand U5785 (N_5785,N_4060,N_4909);
nor U5786 (N_5786,N_4777,N_4631);
and U5787 (N_5787,N_4614,N_4604);
and U5788 (N_5788,N_4258,N_4397);
or U5789 (N_5789,N_4683,N_4084);
nand U5790 (N_5790,N_4621,N_4801);
nand U5791 (N_5791,N_4690,N_4232);
or U5792 (N_5792,N_4737,N_4861);
nor U5793 (N_5793,N_4391,N_4077);
nor U5794 (N_5794,N_4669,N_4906);
xnor U5795 (N_5795,N_4826,N_4936);
nor U5796 (N_5796,N_4816,N_4770);
xnor U5797 (N_5797,N_4410,N_4757);
nor U5798 (N_5798,N_4956,N_4957);
nand U5799 (N_5799,N_4685,N_4937);
nand U5800 (N_5800,N_4232,N_4592);
and U5801 (N_5801,N_4583,N_4927);
nor U5802 (N_5802,N_4741,N_4105);
or U5803 (N_5803,N_4740,N_4727);
nand U5804 (N_5804,N_4408,N_4450);
xor U5805 (N_5805,N_4728,N_4267);
nand U5806 (N_5806,N_4109,N_4122);
nand U5807 (N_5807,N_4298,N_4839);
and U5808 (N_5808,N_4724,N_4424);
nor U5809 (N_5809,N_4510,N_4269);
and U5810 (N_5810,N_4097,N_4952);
nor U5811 (N_5811,N_4730,N_4381);
nand U5812 (N_5812,N_4593,N_4290);
or U5813 (N_5813,N_4828,N_4242);
or U5814 (N_5814,N_4957,N_4206);
nand U5815 (N_5815,N_4760,N_4848);
and U5816 (N_5816,N_4795,N_4917);
and U5817 (N_5817,N_4810,N_4320);
nor U5818 (N_5818,N_4099,N_4602);
and U5819 (N_5819,N_4093,N_4390);
and U5820 (N_5820,N_4022,N_4031);
or U5821 (N_5821,N_4074,N_4639);
xnor U5822 (N_5822,N_4155,N_4086);
and U5823 (N_5823,N_4688,N_4934);
nand U5824 (N_5824,N_4163,N_4289);
and U5825 (N_5825,N_4663,N_4106);
or U5826 (N_5826,N_4635,N_4951);
or U5827 (N_5827,N_4561,N_4556);
and U5828 (N_5828,N_4801,N_4915);
nand U5829 (N_5829,N_4468,N_4604);
or U5830 (N_5830,N_4372,N_4482);
xor U5831 (N_5831,N_4632,N_4533);
or U5832 (N_5832,N_4896,N_4443);
nand U5833 (N_5833,N_4885,N_4830);
and U5834 (N_5834,N_4012,N_4548);
nor U5835 (N_5835,N_4031,N_4610);
nand U5836 (N_5836,N_4570,N_4743);
nand U5837 (N_5837,N_4377,N_4453);
nor U5838 (N_5838,N_4994,N_4053);
nand U5839 (N_5839,N_4719,N_4130);
nand U5840 (N_5840,N_4898,N_4476);
and U5841 (N_5841,N_4262,N_4857);
nor U5842 (N_5842,N_4760,N_4327);
nand U5843 (N_5843,N_4529,N_4668);
or U5844 (N_5844,N_4941,N_4377);
nor U5845 (N_5845,N_4089,N_4306);
nor U5846 (N_5846,N_4755,N_4415);
and U5847 (N_5847,N_4838,N_4121);
nand U5848 (N_5848,N_4219,N_4616);
nor U5849 (N_5849,N_4006,N_4354);
nand U5850 (N_5850,N_4099,N_4193);
nand U5851 (N_5851,N_4463,N_4192);
nand U5852 (N_5852,N_4218,N_4590);
or U5853 (N_5853,N_4349,N_4813);
nor U5854 (N_5854,N_4773,N_4002);
or U5855 (N_5855,N_4033,N_4096);
nand U5856 (N_5856,N_4333,N_4773);
nand U5857 (N_5857,N_4655,N_4409);
xnor U5858 (N_5858,N_4743,N_4185);
nand U5859 (N_5859,N_4583,N_4988);
and U5860 (N_5860,N_4808,N_4052);
and U5861 (N_5861,N_4716,N_4698);
xor U5862 (N_5862,N_4446,N_4320);
or U5863 (N_5863,N_4211,N_4156);
nor U5864 (N_5864,N_4215,N_4958);
nand U5865 (N_5865,N_4557,N_4543);
or U5866 (N_5866,N_4357,N_4905);
or U5867 (N_5867,N_4659,N_4042);
or U5868 (N_5868,N_4968,N_4446);
and U5869 (N_5869,N_4064,N_4515);
or U5870 (N_5870,N_4958,N_4840);
nand U5871 (N_5871,N_4334,N_4654);
xor U5872 (N_5872,N_4553,N_4432);
and U5873 (N_5873,N_4135,N_4512);
or U5874 (N_5874,N_4877,N_4482);
and U5875 (N_5875,N_4384,N_4901);
xor U5876 (N_5876,N_4494,N_4800);
xnor U5877 (N_5877,N_4861,N_4656);
nand U5878 (N_5878,N_4824,N_4073);
or U5879 (N_5879,N_4673,N_4420);
and U5880 (N_5880,N_4715,N_4029);
and U5881 (N_5881,N_4177,N_4681);
xnor U5882 (N_5882,N_4696,N_4697);
nand U5883 (N_5883,N_4988,N_4462);
or U5884 (N_5884,N_4694,N_4318);
or U5885 (N_5885,N_4949,N_4530);
nor U5886 (N_5886,N_4736,N_4498);
and U5887 (N_5887,N_4735,N_4775);
nor U5888 (N_5888,N_4042,N_4810);
or U5889 (N_5889,N_4529,N_4737);
and U5890 (N_5890,N_4859,N_4700);
or U5891 (N_5891,N_4832,N_4967);
nor U5892 (N_5892,N_4607,N_4898);
and U5893 (N_5893,N_4771,N_4667);
nor U5894 (N_5894,N_4730,N_4395);
xor U5895 (N_5895,N_4456,N_4709);
or U5896 (N_5896,N_4116,N_4829);
or U5897 (N_5897,N_4256,N_4958);
nor U5898 (N_5898,N_4728,N_4919);
nand U5899 (N_5899,N_4815,N_4359);
nor U5900 (N_5900,N_4130,N_4586);
nand U5901 (N_5901,N_4487,N_4536);
xnor U5902 (N_5902,N_4932,N_4235);
nor U5903 (N_5903,N_4235,N_4019);
nand U5904 (N_5904,N_4479,N_4835);
nor U5905 (N_5905,N_4381,N_4332);
and U5906 (N_5906,N_4882,N_4954);
or U5907 (N_5907,N_4396,N_4137);
and U5908 (N_5908,N_4466,N_4836);
nor U5909 (N_5909,N_4165,N_4978);
nand U5910 (N_5910,N_4708,N_4556);
nor U5911 (N_5911,N_4981,N_4215);
nor U5912 (N_5912,N_4792,N_4339);
or U5913 (N_5913,N_4335,N_4850);
nand U5914 (N_5914,N_4915,N_4577);
and U5915 (N_5915,N_4256,N_4417);
nand U5916 (N_5916,N_4530,N_4639);
nor U5917 (N_5917,N_4200,N_4994);
and U5918 (N_5918,N_4717,N_4437);
xor U5919 (N_5919,N_4037,N_4686);
or U5920 (N_5920,N_4921,N_4231);
and U5921 (N_5921,N_4911,N_4918);
nand U5922 (N_5922,N_4579,N_4276);
nor U5923 (N_5923,N_4131,N_4450);
xor U5924 (N_5924,N_4907,N_4524);
xnor U5925 (N_5925,N_4177,N_4200);
nand U5926 (N_5926,N_4670,N_4595);
xnor U5927 (N_5927,N_4272,N_4163);
xor U5928 (N_5928,N_4752,N_4352);
or U5929 (N_5929,N_4610,N_4022);
or U5930 (N_5930,N_4973,N_4608);
nand U5931 (N_5931,N_4346,N_4871);
nor U5932 (N_5932,N_4597,N_4278);
xor U5933 (N_5933,N_4231,N_4953);
nor U5934 (N_5934,N_4330,N_4320);
nor U5935 (N_5935,N_4719,N_4514);
or U5936 (N_5936,N_4654,N_4716);
nor U5937 (N_5937,N_4697,N_4743);
nand U5938 (N_5938,N_4473,N_4565);
or U5939 (N_5939,N_4313,N_4027);
xnor U5940 (N_5940,N_4267,N_4096);
xnor U5941 (N_5941,N_4940,N_4965);
or U5942 (N_5942,N_4286,N_4323);
and U5943 (N_5943,N_4552,N_4909);
nor U5944 (N_5944,N_4857,N_4210);
and U5945 (N_5945,N_4524,N_4268);
or U5946 (N_5946,N_4995,N_4752);
nand U5947 (N_5947,N_4756,N_4588);
nor U5948 (N_5948,N_4597,N_4892);
xor U5949 (N_5949,N_4126,N_4173);
nand U5950 (N_5950,N_4019,N_4309);
xnor U5951 (N_5951,N_4866,N_4854);
nand U5952 (N_5952,N_4972,N_4105);
nand U5953 (N_5953,N_4514,N_4958);
nor U5954 (N_5954,N_4009,N_4053);
and U5955 (N_5955,N_4983,N_4552);
nor U5956 (N_5956,N_4015,N_4667);
or U5957 (N_5957,N_4403,N_4530);
or U5958 (N_5958,N_4330,N_4362);
nor U5959 (N_5959,N_4646,N_4812);
nand U5960 (N_5960,N_4421,N_4058);
nand U5961 (N_5961,N_4275,N_4188);
xnor U5962 (N_5962,N_4369,N_4983);
and U5963 (N_5963,N_4611,N_4755);
or U5964 (N_5964,N_4888,N_4815);
nand U5965 (N_5965,N_4094,N_4228);
or U5966 (N_5966,N_4192,N_4583);
and U5967 (N_5967,N_4199,N_4244);
and U5968 (N_5968,N_4077,N_4251);
nor U5969 (N_5969,N_4678,N_4717);
or U5970 (N_5970,N_4088,N_4847);
nor U5971 (N_5971,N_4063,N_4747);
and U5972 (N_5972,N_4206,N_4816);
nand U5973 (N_5973,N_4948,N_4884);
nor U5974 (N_5974,N_4565,N_4008);
and U5975 (N_5975,N_4126,N_4734);
nand U5976 (N_5976,N_4002,N_4697);
or U5977 (N_5977,N_4694,N_4809);
nand U5978 (N_5978,N_4461,N_4262);
or U5979 (N_5979,N_4237,N_4933);
or U5980 (N_5980,N_4523,N_4355);
xor U5981 (N_5981,N_4025,N_4595);
or U5982 (N_5982,N_4291,N_4872);
nor U5983 (N_5983,N_4958,N_4166);
nand U5984 (N_5984,N_4983,N_4188);
nor U5985 (N_5985,N_4557,N_4775);
nand U5986 (N_5986,N_4105,N_4755);
or U5987 (N_5987,N_4229,N_4429);
nor U5988 (N_5988,N_4893,N_4533);
or U5989 (N_5989,N_4442,N_4960);
xnor U5990 (N_5990,N_4746,N_4201);
nand U5991 (N_5991,N_4301,N_4446);
nor U5992 (N_5992,N_4087,N_4854);
and U5993 (N_5993,N_4291,N_4336);
nor U5994 (N_5994,N_4210,N_4435);
nand U5995 (N_5995,N_4662,N_4473);
nor U5996 (N_5996,N_4867,N_4682);
or U5997 (N_5997,N_4835,N_4150);
or U5998 (N_5998,N_4913,N_4669);
nand U5999 (N_5999,N_4022,N_4111);
and U6000 (N_6000,N_5616,N_5702);
and U6001 (N_6001,N_5118,N_5898);
xnor U6002 (N_6002,N_5104,N_5677);
nand U6003 (N_6003,N_5240,N_5599);
and U6004 (N_6004,N_5031,N_5046);
nor U6005 (N_6005,N_5356,N_5224);
and U6006 (N_6006,N_5633,N_5886);
xor U6007 (N_6007,N_5111,N_5050);
and U6008 (N_6008,N_5249,N_5501);
nor U6009 (N_6009,N_5157,N_5239);
or U6010 (N_6010,N_5470,N_5694);
and U6011 (N_6011,N_5437,N_5986);
nor U6012 (N_6012,N_5640,N_5868);
or U6013 (N_6013,N_5361,N_5927);
and U6014 (N_6014,N_5784,N_5330);
nor U6015 (N_6015,N_5357,N_5754);
nand U6016 (N_6016,N_5611,N_5889);
nor U6017 (N_6017,N_5151,N_5965);
or U6018 (N_6018,N_5628,N_5215);
nor U6019 (N_6019,N_5397,N_5475);
nor U6020 (N_6020,N_5099,N_5897);
and U6021 (N_6021,N_5552,N_5041);
and U6022 (N_6022,N_5533,N_5843);
nor U6023 (N_6023,N_5555,N_5894);
nor U6024 (N_6024,N_5167,N_5158);
or U6025 (N_6025,N_5202,N_5557);
and U6026 (N_6026,N_5862,N_5454);
and U6027 (N_6027,N_5053,N_5171);
nand U6028 (N_6028,N_5573,N_5329);
and U6029 (N_6029,N_5918,N_5753);
or U6030 (N_6030,N_5563,N_5386);
or U6031 (N_6031,N_5322,N_5043);
nand U6032 (N_6032,N_5791,N_5458);
nor U6033 (N_6033,N_5728,N_5941);
xor U6034 (N_6034,N_5101,N_5553);
xor U6035 (N_6035,N_5542,N_5078);
or U6036 (N_6036,N_5696,N_5024);
nor U6037 (N_6037,N_5340,N_5960);
nor U6038 (N_6038,N_5816,N_5917);
nor U6039 (N_6039,N_5478,N_5442);
or U6040 (N_6040,N_5451,N_5001);
nor U6041 (N_6041,N_5013,N_5731);
and U6042 (N_6042,N_5097,N_5829);
or U6043 (N_6043,N_5438,N_5381);
or U6044 (N_6044,N_5583,N_5291);
nand U6045 (N_6045,N_5321,N_5551);
nor U6046 (N_6046,N_5536,N_5887);
or U6047 (N_6047,N_5034,N_5310);
xnor U6048 (N_6048,N_5817,N_5492);
nor U6049 (N_6049,N_5068,N_5429);
nand U6050 (N_6050,N_5448,N_5881);
and U6051 (N_6051,N_5845,N_5937);
and U6052 (N_6052,N_5796,N_5439);
nand U6053 (N_6053,N_5016,N_5926);
nand U6054 (N_6054,N_5936,N_5659);
nand U6055 (N_6055,N_5539,N_5124);
nor U6056 (N_6056,N_5679,N_5947);
nand U6057 (N_6057,N_5328,N_5567);
nor U6058 (N_6058,N_5146,N_5258);
or U6059 (N_6059,N_5675,N_5624);
nor U6060 (N_6060,N_5203,N_5564);
nand U6061 (N_6061,N_5874,N_5715);
and U6062 (N_6062,N_5972,N_5142);
and U6063 (N_6063,N_5968,N_5974);
nand U6064 (N_6064,N_5831,N_5395);
nor U6065 (N_6065,N_5314,N_5586);
and U6066 (N_6066,N_5178,N_5656);
nand U6067 (N_6067,N_5362,N_5390);
or U6068 (N_6068,N_5359,N_5004);
nor U6069 (N_6069,N_5699,N_5517);
and U6070 (N_6070,N_5011,N_5821);
nor U6071 (N_6071,N_5313,N_5037);
or U6072 (N_6072,N_5035,N_5513);
nor U6073 (N_6073,N_5168,N_5226);
and U6074 (N_6074,N_5743,N_5132);
nand U6075 (N_6075,N_5893,N_5687);
nand U6076 (N_6076,N_5629,N_5735);
nor U6077 (N_6077,N_5801,N_5776);
nand U6078 (N_6078,N_5062,N_5990);
and U6079 (N_6079,N_5604,N_5741);
nor U6080 (N_6080,N_5307,N_5562);
or U6081 (N_6081,N_5710,N_5277);
nor U6082 (N_6082,N_5814,N_5755);
nand U6083 (N_6083,N_5266,N_5032);
nor U6084 (N_6084,N_5645,N_5189);
nand U6085 (N_6085,N_5254,N_5726);
nand U6086 (N_6086,N_5353,N_5577);
and U6087 (N_6087,N_5080,N_5740);
nor U6088 (N_6088,N_5932,N_5576);
and U6089 (N_6089,N_5485,N_5566);
xor U6090 (N_6090,N_5825,N_5707);
nor U6091 (N_6091,N_5913,N_5649);
xor U6092 (N_6092,N_5026,N_5738);
xor U6093 (N_6093,N_5499,N_5663);
and U6094 (N_6094,N_5444,N_5771);
and U6095 (N_6095,N_5980,N_5514);
or U6096 (N_6096,N_5900,N_5405);
or U6097 (N_6097,N_5655,N_5569);
or U6098 (N_6098,N_5584,N_5159);
nor U6099 (N_6099,N_5391,N_5131);
and U6100 (N_6100,N_5246,N_5790);
and U6101 (N_6101,N_5427,N_5618);
nand U6102 (N_6102,N_5135,N_5371);
nor U6103 (N_6103,N_5884,N_5846);
or U6104 (N_6104,N_5891,N_5931);
and U6105 (N_6105,N_5867,N_5878);
xnor U6106 (N_6106,N_5579,N_5370);
or U6107 (N_6107,N_5372,N_5875);
nor U6108 (N_6108,N_5476,N_5450);
nor U6109 (N_6109,N_5129,N_5176);
nand U6110 (N_6110,N_5150,N_5349);
nor U6111 (N_6111,N_5905,N_5546);
and U6112 (N_6112,N_5612,N_5198);
xnor U6113 (N_6113,N_5615,N_5217);
xnor U6114 (N_6114,N_5109,N_5412);
and U6115 (N_6115,N_5232,N_5081);
and U6116 (N_6116,N_5393,N_5620);
xnor U6117 (N_6117,N_5250,N_5123);
nand U6118 (N_6118,N_5015,N_5786);
nand U6119 (N_6119,N_5651,N_5712);
xor U6120 (N_6120,N_5487,N_5460);
or U6121 (N_6121,N_5082,N_5009);
and U6122 (N_6122,N_5793,N_5300);
xnor U6123 (N_6123,N_5605,N_5510);
nand U6124 (N_6124,N_5603,N_5734);
nor U6125 (N_6125,N_5709,N_5909);
xnor U6126 (N_6126,N_5423,N_5870);
or U6127 (N_6127,N_5907,N_5653);
and U6128 (N_6128,N_5006,N_5410);
nor U6129 (N_6129,N_5367,N_5084);
nand U6130 (N_6130,N_5234,N_5834);
nor U6131 (N_6131,N_5471,N_5140);
or U6132 (N_6132,N_5835,N_5029);
xnor U6133 (N_6133,N_5928,N_5890);
and U6134 (N_6134,N_5019,N_5264);
xnor U6135 (N_6135,N_5772,N_5216);
nand U6136 (N_6136,N_5924,N_5761);
or U6137 (N_6137,N_5148,N_5207);
or U6138 (N_6138,N_5718,N_5064);
nand U6139 (N_6139,N_5079,N_5672);
or U6140 (N_6140,N_5302,N_5727);
nor U6141 (N_6141,N_5156,N_5063);
nand U6142 (N_6142,N_5344,N_5698);
xor U6143 (N_6143,N_5970,N_5650);
nor U6144 (N_6144,N_5145,N_5752);
or U6145 (N_6145,N_5069,N_5363);
nand U6146 (N_6146,N_5664,N_5319);
and U6147 (N_6147,N_5490,N_5484);
and U6148 (N_6148,N_5701,N_5982);
or U6149 (N_6149,N_5509,N_5975);
nand U6150 (N_6150,N_5978,N_5040);
nor U6151 (N_6151,N_5779,N_5425);
nand U6152 (N_6152,N_5840,N_5428);
xnor U6153 (N_6153,N_5892,N_5805);
and U6154 (N_6154,N_5332,N_5822);
nand U6155 (N_6155,N_5126,N_5273);
nand U6156 (N_6156,N_5408,N_5303);
or U6157 (N_6157,N_5348,N_5417);
nand U6158 (N_6158,N_5808,N_5644);
and U6159 (N_6159,N_5299,N_5634);
or U6160 (N_6160,N_5864,N_5309);
or U6161 (N_6161,N_5060,N_5187);
and U6162 (N_6162,N_5318,N_5456);
nand U6163 (N_6163,N_5942,N_5643);
nor U6164 (N_6164,N_5949,N_5981);
xnor U6165 (N_6165,N_5785,N_5022);
and U6166 (N_6166,N_5690,N_5200);
and U6167 (N_6167,N_5521,N_5983);
and U6168 (N_6168,N_5775,N_5759);
nand U6169 (N_6169,N_5383,N_5241);
and U6170 (N_6170,N_5220,N_5899);
nor U6171 (N_6171,N_5935,N_5872);
and U6172 (N_6172,N_5012,N_5057);
or U6173 (N_6173,N_5961,N_5435);
and U6174 (N_6174,N_5789,N_5376);
or U6175 (N_6175,N_5590,N_5338);
or U6176 (N_6176,N_5952,N_5335);
or U6177 (N_6177,N_5033,N_5360);
nor U6178 (N_6178,N_5121,N_5781);
xnor U6179 (N_6179,N_5914,N_5174);
and U6180 (N_6180,N_5951,N_5815);
and U6181 (N_6181,N_5688,N_5638);
or U6182 (N_6182,N_5175,N_5073);
and U6183 (N_6183,N_5792,N_5185);
nor U6184 (N_6184,N_5221,N_5883);
or U6185 (N_6185,N_5795,N_5021);
and U6186 (N_6186,N_5023,N_5496);
nand U6187 (N_6187,N_5895,N_5166);
nand U6188 (N_6188,N_5901,N_5873);
nor U6189 (N_6189,N_5760,N_5325);
or U6190 (N_6190,N_5107,N_5455);
and U6191 (N_6191,N_5570,N_5988);
and U6192 (N_6192,N_5282,N_5744);
and U6193 (N_6193,N_5794,N_5125);
xnor U6194 (N_6194,N_5445,N_5908);
and U6195 (N_6195,N_5642,N_5762);
nor U6196 (N_6196,N_5305,N_5077);
and U6197 (N_6197,N_5333,N_5502);
nand U6198 (N_6198,N_5392,N_5058);
nand U6199 (N_6199,N_5387,N_5963);
and U6200 (N_6200,N_5337,N_5388);
and U6201 (N_6201,N_5312,N_5269);
and U6202 (N_6202,N_5285,N_5306);
nand U6203 (N_6203,N_5186,N_5100);
or U6204 (N_6204,N_5997,N_5172);
or U6205 (N_6205,N_5304,N_5680);
and U6206 (N_6206,N_5674,N_5538);
or U6207 (N_6207,N_5800,N_5912);
nor U6208 (N_6208,N_5658,N_5466);
nor U6209 (N_6209,N_5700,N_5747);
or U6210 (N_6210,N_5290,N_5347);
nand U6211 (N_6211,N_5297,N_5355);
nand U6212 (N_6212,N_5288,N_5153);
nand U6213 (N_6213,N_5112,N_5432);
nor U6214 (N_6214,N_5452,N_5469);
xor U6215 (N_6215,N_5003,N_5052);
and U6216 (N_6216,N_5182,N_5418);
and U6217 (N_6217,N_5110,N_5416);
nor U6218 (N_6218,N_5406,N_5516);
and U6219 (N_6219,N_5411,N_5719);
or U6220 (N_6220,N_5869,N_5681);
or U6221 (N_6221,N_5703,N_5238);
nor U6222 (N_6222,N_5289,N_5190);
nand U6223 (N_6223,N_5293,N_5341);
nor U6224 (N_6224,N_5682,N_5149);
xnor U6225 (N_6225,N_5880,N_5343);
and U6226 (N_6226,N_5839,N_5910);
nor U6227 (N_6227,N_5515,N_5811);
or U6228 (N_6228,N_5902,N_5705);
nand U6229 (N_6229,N_5797,N_5697);
and U6230 (N_6230,N_5691,N_5998);
or U6231 (N_6231,N_5860,N_5859);
xor U6232 (N_6232,N_5739,N_5920);
and U6233 (N_6233,N_5979,N_5858);
nand U6234 (N_6234,N_5844,N_5896);
or U6235 (N_6235,N_5518,N_5463);
nand U6236 (N_6236,N_5144,N_5541);
and U6237 (N_6237,N_5020,N_5228);
or U6238 (N_6238,N_5352,N_5420);
nand U6239 (N_6239,N_5588,N_5279);
nor U6240 (N_6240,N_5520,N_5946);
xnor U6241 (N_6241,N_5768,N_5547);
or U6242 (N_6242,N_5777,N_5637);
nand U6243 (N_6243,N_5377,N_5530);
and U6244 (N_6244,N_5394,N_5652);
xnor U6245 (N_6245,N_5464,N_5559);
nand U6246 (N_6246,N_5262,N_5400);
nor U6247 (N_6247,N_5724,N_5957);
nand U6248 (N_6248,N_5550,N_5977);
nand U6249 (N_6249,N_5414,N_5255);
or U6250 (N_6250,N_5594,N_5678);
nand U6251 (N_6251,N_5147,N_5301);
nor U6252 (N_6252,N_5545,N_5358);
nor U6253 (N_6253,N_5030,N_5136);
xnor U6254 (N_6254,N_5523,N_5204);
nand U6255 (N_6255,N_5237,N_5434);
nand U6256 (N_6256,N_5810,N_5572);
xor U6257 (N_6257,N_5495,N_5162);
and U6258 (N_6258,N_5180,N_5671);
nand U6259 (N_6259,N_5404,N_5067);
nor U6260 (N_6260,N_5736,N_5823);
nand U6261 (N_6261,N_5128,N_5934);
nand U6262 (N_6262,N_5511,N_5602);
or U6263 (N_6263,N_5746,N_5994);
nand U6264 (N_6264,N_5948,N_5007);
or U6265 (N_6265,N_5818,N_5832);
nor U6266 (N_6266,N_5227,N_5861);
and U6267 (N_6267,N_5422,N_5373);
and U6268 (N_6268,N_5733,N_5116);
and U6269 (N_6269,N_5263,N_5048);
nand U6270 (N_6270,N_5526,N_5196);
nor U6271 (N_6271,N_5560,N_5879);
nor U6272 (N_6272,N_5436,N_5945);
nand U6273 (N_6273,N_5850,N_5660);
nand U6274 (N_6274,N_5222,N_5481);
nand U6275 (N_6275,N_5838,N_5231);
nand U6276 (N_6276,N_5529,N_5218);
and U6277 (N_6277,N_5824,N_5243);
and U6278 (N_6278,N_5704,N_5426);
nand U6279 (N_6279,N_5685,N_5378);
and U6280 (N_6280,N_5117,N_5930);
nor U6281 (N_6281,N_5173,N_5851);
nand U6282 (N_6282,N_5483,N_5014);
and U6283 (N_6283,N_5774,N_5010);
nand U6284 (N_6284,N_5334,N_5711);
or U6285 (N_6285,N_5722,N_5364);
xor U6286 (N_6286,N_5969,N_5298);
nand U6287 (N_6287,N_5443,N_5380);
or U6288 (N_6288,N_5491,N_5091);
and U6289 (N_6289,N_5494,N_5595);
nand U6290 (N_6290,N_5863,N_5339);
or U6291 (N_6291,N_5987,N_5326);
or U6292 (N_6292,N_5807,N_5841);
and U6293 (N_6293,N_5745,N_5544);
nand U6294 (N_6294,N_5580,N_5543);
or U6295 (N_6295,N_5002,N_5809);
nand U6296 (N_6296,N_5877,N_5075);
and U6297 (N_6297,N_5923,N_5954);
xor U6298 (N_6298,N_5548,N_5802);
and U6299 (N_6299,N_5489,N_5154);
and U6300 (N_6300,N_5574,N_5384);
or U6301 (N_6301,N_5284,N_5201);
or U6302 (N_6302,N_5155,N_5856);
nor U6303 (N_6303,N_5556,N_5648);
nor U6304 (N_6304,N_5066,N_5331);
or U6305 (N_6305,N_5431,N_5385);
nand U6306 (N_6306,N_5985,N_5209);
xor U6307 (N_6307,N_5071,N_5163);
or U6308 (N_6308,N_5106,N_5783);
nor U6309 (N_6309,N_5625,N_5374);
or U6310 (N_6310,N_5292,N_5143);
nand U6311 (N_6311,N_5197,N_5267);
or U6312 (N_6312,N_5467,N_5916);
and U6313 (N_6313,N_5996,N_5668);
or U6314 (N_6314,N_5631,N_5787);
nor U6315 (N_6315,N_5183,N_5621);
or U6316 (N_6316,N_5641,N_5087);
and U6317 (N_6317,N_5127,N_5092);
nor U6318 (N_6318,N_5827,N_5504);
nor U6319 (N_6319,N_5453,N_5767);
or U6320 (N_6320,N_5959,N_5626);
nand U6321 (N_6321,N_5676,N_5938);
or U6322 (N_6322,N_5535,N_5323);
nor U6323 (N_6323,N_5508,N_5139);
and U6324 (N_6324,N_5480,N_5268);
nand U6325 (N_6325,N_5119,N_5773);
and U6326 (N_6326,N_5316,N_5120);
or U6327 (N_6327,N_5211,N_5472);
and U6328 (N_6328,N_5336,N_5210);
nor U6329 (N_6329,N_5944,N_5468);
nand U6330 (N_6330,N_5000,N_5906);
nor U6331 (N_6331,N_5113,N_5497);
nand U6332 (N_6332,N_5094,N_5474);
nor U6333 (N_6333,N_5413,N_5571);
nand U6334 (N_6334,N_5219,N_5819);
and U6335 (N_6335,N_5717,N_5493);
xnor U6336 (N_6336,N_5966,N_5854);
and U6337 (N_6337,N_5365,N_5537);
nor U6338 (N_6338,N_5191,N_5430);
or U6339 (N_6339,N_5782,N_5421);
nand U6340 (N_6340,N_5257,N_5047);
and U6341 (N_6341,N_5161,N_5804);
nor U6342 (N_6342,N_5177,N_5181);
nand U6343 (N_6343,N_5830,N_5737);
and U6344 (N_6344,N_5654,N_5554);
nand U6345 (N_6345,N_5179,N_5342);
and U6346 (N_6346,N_5382,N_5607);
nor U6347 (N_6347,N_5610,N_5230);
and U6348 (N_6348,N_5477,N_5991);
xnor U6349 (N_6349,N_5852,N_5503);
nor U6350 (N_6350,N_5065,N_5083);
and U6351 (N_6351,N_5379,N_5138);
and U6352 (N_6352,N_5252,N_5366);
and U6353 (N_6353,N_5882,N_5865);
and U6354 (N_6354,N_5630,N_5184);
xor U6355 (N_6355,N_5636,N_5194);
nand U6356 (N_6356,N_5038,N_5457);
and U6357 (N_6357,N_5133,N_5500);
nand U6358 (N_6358,N_5396,N_5272);
xnor U6359 (N_6359,N_5346,N_5617);
xnor U6360 (N_6360,N_5964,N_5730);
and U6361 (N_6361,N_5585,N_5235);
xor U6362 (N_6362,N_5798,N_5488);
nor U6363 (N_6363,N_5122,N_5939);
or U6364 (N_6364,N_5287,N_5956);
nand U6365 (N_6365,N_5670,N_5995);
nand U6366 (N_6366,N_5044,N_5657);
and U6367 (N_6367,N_5540,N_5647);
and U6368 (N_6368,N_5592,N_5929);
nand U6369 (N_6369,N_5866,N_5130);
and U6370 (N_6370,N_5461,N_5749);
and U6371 (N_6371,N_5223,N_5622);
xor U6372 (N_6372,N_5278,N_5212);
nor U6373 (N_6373,N_5857,N_5855);
nand U6374 (N_6374,N_5609,N_5274);
nor U6375 (N_6375,N_5512,N_5849);
nand U6376 (N_6376,N_5669,N_5311);
nand U6377 (N_6377,N_5164,N_5623);
nor U6378 (N_6378,N_5095,N_5440);
and U6379 (N_6379,N_5419,N_5765);
nor U6380 (N_6380,N_5689,N_5565);
nor U6381 (N_6381,N_5528,N_5806);
and U6382 (N_6382,N_5070,N_5449);
nor U6383 (N_6383,N_5345,N_5188);
or U6384 (N_6384,N_5152,N_5465);
or U6385 (N_6385,N_5601,N_5090);
or U6386 (N_6386,N_5085,N_5244);
nand U6387 (N_6387,N_5708,N_5056);
nor U6388 (N_6388,N_5261,N_5283);
xnor U6389 (N_6389,N_5525,N_5921);
nor U6390 (N_6390,N_5940,N_5294);
or U6391 (N_6391,N_5568,N_5137);
and U6392 (N_6392,N_5320,N_5992);
and U6393 (N_6393,N_5253,N_5072);
nand U6394 (N_6394,N_5614,N_5351);
or U6395 (N_6395,N_5732,N_5665);
nor U6396 (N_6396,N_5295,N_5950);
or U6397 (N_6397,N_5758,N_5195);
and U6398 (N_6398,N_5169,N_5589);
nand U6399 (N_6399,N_5208,N_5531);
nor U6400 (N_6400,N_5275,N_5369);
and U6401 (N_6401,N_5225,N_5751);
xor U6402 (N_6402,N_5661,N_5922);
and U6403 (N_6403,N_5441,N_5778);
or U6404 (N_6404,N_5519,N_5317);
nand U6405 (N_6405,N_5459,N_5141);
and U6406 (N_6406,N_5242,N_5742);
or U6407 (N_6407,N_5027,N_5597);
and U6408 (N_6408,N_5098,N_5591);
or U6409 (N_6409,N_5086,N_5606);
and U6410 (N_6410,N_5581,N_5248);
and U6411 (N_6411,N_5770,N_5943);
nor U6412 (N_6412,N_5549,N_5587);
or U6413 (N_6413,N_5600,N_5308);
nand U6414 (N_6414,N_5462,N_5826);
xor U6415 (N_6415,N_5399,N_5876);
nand U6416 (N_6416,N_5558,N_5105);
nor U6417 (N_6417,N_5389,N_5527);
or U6418 (N_6418,N_5270,N_5375);
nand U6419 (N_6419,N_5976,N_5498);
or U6420 (N_6420,N_5482,N_5769);
nor U6421 (N_6421,N_5415,N_5967);
and U6422 (N_6422,N_5061,N_5885);
xnor U6423 (N_6423,N_5666,N_5256);
nand U6424 (N_6424,N_5054,N_5114);
and U6425 (N_6425,N_5473,N_5296);
and U6426 (N_6426,N_5271,N_5059);
nor U6427 (N_6427,N_5055,N_5206);
nand U6428 (N_6428,N_5534,N_5684);
or U6429 (N_6429,N_5608,N_5984);
nand U6430 (N_6430,N_5911,N_5788);
nand U6431 (N_6431,N_5750,N_5108);
or U6432 (N_6432,N_5327,N_5522);
and U6433 (N_6433,N_5259,N_5134);
and U6434 (N_6434,N_5848,N_5532);
nand U6435 (N_6435,N_5280,N_5925);
nand U6436 (N_6436,N_5757,N_5192);
xor U6437 (N_6437,N_5049,N_5233);
nand U6438 (N_6438,N_5089,N_5005);
or U6439 (N_6439,N_5582,N_5074);
nor U6440 (N_6440,N_5613,N_5424);
nor U6441 (N_6441,N_5993,N_5247);
or U6442 (N_6442,N_5017,N_5102);
and U6443 (N_6443,N_5281,N_5729);
nor U6444 (N_6444,N_5088,N_5667);
and U6445 (N_6445,N_5286,N_5368);
nor U6446 (N_6446,N_5407,N_5276);
or U6447 (N_6447,N_5245,N_5524);
or U6448 (N_6448,N_5933,N_5028);
xnor U6449 (N_6449,N_5214,N_5706);
and U6450 (N_6450,N_5695,N_5999);
nand U6451 (N_6451,N_5662,N_5748);
nor U6452 (N_6452,N_5780,N_5433);
nor U6453 (N_6453,N_5446,N_5409);
nor U6454 (N_6454,N_5989,N_5971);
nor U6455 (N_6455,N_5813,N_5836);
and U6456 (N_6456,N_5561,N_5486);
nor U6457 (N_6457,N_5973,N_5903);
or U6458 (N_6458,N_5693,N_5812);
nor U6459 (N_6459,N_5799,N_5213);
nor U6460 (N_6460,N_5402,N_5627);
or U6461 (N_6461,N_5593,N_5842);
xor U6462 (N_6462,N_5958,N_5042);
or U6463 (N_6463,N_5635,N_5051);
or U6464 (N_6464,N_5324,N_5904);
nand U6465 (N_6465,N_5725,N_5193);
or U6466 (N_6466,N_5803,N_5170);
xor U6467 (N_6467,N_5632,N_5847);
or U6468 (N_6468,N_5575,N_5871);
xnor U6469 (N_6469,N_5008,N_5619);
nor U6470 (N_6470,N_5479,N_5837);
nand U6471 (N_6471,N_5763,N_5639);
or U6472 (N_6472,N_5953,N_5756);
nor U6473 (N_6473,N_5714,N_5045);
nor U6474 (N_6474,N_5354,N_5506);
nand U6475 (N_6475,N_5507,N_5447);
or U6476 (N_6476,N_5598,N_5096);
or U6477 (N_6477,N_5915,N_5251);
or U6478 (N_6478,N_5160,N_5716);
nor U6479 (N_6479,N_5403,N_5350);
nor U6480 (N_6480,N_5888,N_5686);
nand U6481 (N_6481,N_5919,N_5076);
and U6482 (N_6482,N_5713,N_5260);
xnor U6483 (N_6483,N_5265,N_5039);
and U6484 (N_6484,N_5018,N_5398);
nand U6485 (N_6485,N_5955,N_5766);
and U6486 (N_6486,N_5025,N_5229);
and U6487 (N_6487,N_5596,N_5692);
or U6488 (N_6488,N_5646,N_5103);
nand U6489 (N_6489,N_5315,N_5205);
nand U6490 (N_6490,N_5165,N_5578);
nor U6491 (N_6491,N_5093,N_5828);
or U6492 (N_6492,N_5236,N_5115);
nor U6493 (N_6493,N_5683,N_5199);
nand U6494 (N_6494,N_5723,N_5505);
nor U6495 (N_6495,N_5833,N_5721);
nor U6496 (N_6496,N_5853,N_5820);
or U6497 (N_6497,N_5036,N_5720);
or U6498 (N_6498,N_5764,N_5401);
nor U6499 (N_6499,N_5673,N_5962);
nor U6500 (N_6500,N_5892,N_5954);
or U6501 (N_6501,N_5014,N_5629);
xor U6502 (N_6502,N_5980,N_5706);
xor U6503 (N_6503,N_5050,N_5849);
nand U6504 (N_6504,N_5621,N_5378);
and U6505 (N_6505,N_5195,N_5074);
and U6506 (N_6506,N_5010,N_5263);
nor U6507 (N_6507,N_5794,N_5530);
nand U6508 (N_6508,N_5121,N_5369);
nand U6509 (N_6509,N_5861,N_5626);
and U6510 (N_6510,N_5581,N_5021);
nor U6511 (N_6511,N_5919,N_5533);
nand U6512 (N_6512,N_5093,N_5789);
nor U6513 (N_6513,N_5366,N_5060);
nand U6514 (N_6514,N_5778,N_5796);
nand U6515 (N_6515,N_5222,N_5435);
nor U6516 (N_6516,N_5549,N_5671);
xor U6517 (N_6517,N_5874,N_5654);
or U6518 (N_6518,N_5358,N_5892);
and U6519 (N_6519,N_5740,N_5636);
nor U6520 (N_6520,N_5518,N_5796);
and U6521 (N_6521,N_5530,N_5464);
xnor U6522 (N_6522,N_5762,N_5167);
nor U6523 (N_6523,N_5673,N_5469);
or U6524 (N_6524,N_5763,N_5105);
nand U6525 (N_6525,N_5697,N_5782);
nor U6526 (N_6526,N_5963,N_5560);
nor U6527 (N_6527,N_5963,N_5491);
nand U6528 (N_6528,N_5855,N_5824);
nand U6529 (N_6529,N_5102,N_5231);
or U6530 (N_6530,N_5235,N_5824);
nand U6531 (N_6531,N_5207,N_5083);
or U6532 (N_6532,N_5270,N_5913);
nand U6533 (N_6533,N_5830,N_5345);
and U6534 (N_6534,N_5122,N_5133);
and U6535 (N_6535,N_5041,N_5171);
nand U6536 (N_6536,N_5709,N_5095);
and U6537 (N_6537,N_5181,N_5544);
xor U6538 (N_6538,N_5418,N_5644);
or U6539 (N_6539,N_5377,N_5264);
xnor U6540 (N_6540,N_5261,N_5859);
or U6541 (N_6541,N_5944,N_5411);
or U6542 (N_6542,N_5475,N_5991);
nand U6543 (N_6543,N_5914,N_5361);
and U6544 (N_6544,N_5084,N_5501);
nor U6545 (N_6545,N_5948,N_5323);
or U6546 (N_6546,N_5409,N_5005);
nand U6547 (N_6547,N_5697,N_5586);
or U6548 (N_6548,N_5672,N_5430);
and U6549 (N_6549,N_5865,N_5801);
and U6550 (N_6550,N_5522,N_5070);
or U6551 (N_6551,N_5041,N_5488);
nand U6552 (N_6552,N_5499,N_5787);
nand U6553 (N_6553,N_5901,N_5093);
and U6554 (N_6554,N_5788,N_5133);
nand U6555 (N_6555,N_5893,N_5674);
and U6556 (N_6556,N_5212,N_5565);
nand U6557 (N_6557,N_5073,N_5576);
nor U6558 (N_6558,N_5504,N_5280);
nand U6559 (N_6559,N_5333,N_5467);
nor U6560 (N_6560,N_5787,N_5594);
nor U6561 (N_6561,N_5479,N_5754);
and U6562 (N_6562,N_5946,N_5774);
xnor U6563 (N_6563,N_5372,N_5706);
xor U6564 (N_6564,N_5871,N_5583);
and U6565 (N_6565,N_5856,N_5346);
nor U6566 (N_6566,N_5804,N_5158);
nor U6567 (N_6567,N_5700,N_5181);
or U6568 (N_6568,N_5290,N_5845);
nor U6569 (N_6569,N_5823,N_5608);
and U6570 (N_6570,N_5536,N_5760);
or U6571 (N_6571,N_5001,N_5980);
nor U6572 (N_6572,N_5949,N_5437);
nand U6573 (N_6573,N_5026,N_5237);
or U6574 (N_6574,N_5540,N_5682);
or U6575 (N_6575,N_5256,N_5466);
and U6576 (N_6576,N_5812,N_5371);
xor U6577 (N_6577,N_5440,N_5137);
nand U6578 (N_6578,N_5174,N_5284);
or U6579 (N_6579,N_5041,N_5566);
and U6580 (N_6580,N_5619,N_5880);
nor U6581 (N_6581,N_5967,N_5954);
nand U6582 (N_6582,N_5684,N_5887);
or U6583 (N_6583,N_5720,N_5566);
xnor U6584 (N_6584,N_5135,N_5898);
xnor U6585 (N_6585,N_5249,N_5931);
or U6586 (N_6586,N_5447,N_5711);
xnor U6587 (N_6587,N_5569,N_5234);
xnor U6588 (N_6588,N_5612,N_5637);
xor U6589 (N_6589,N_5603,N_5126);
xor U6590 (N_6590,N_5315,N_5522);
nor U6591 (N_6591,N_5989,N_5325);
xor U6592 (N_6592,N_5684,N_5035);
or U6593 (N_6593,N_5423,N_5151);
or U6594 (N_6594,N_5312,N_5950);
xor U6595 (N_6595,N_5829,N_5880);
nor U6596 (N_6596,N_5895,N_5369);
or U6597 (N_6597,N_5963,N_5779);
nor U6598 (N_6598,N_5383,N_5913);
and U6599 (N_6599,N_5569,N_5963);
nand U6600 (N_6600,N_5907,N_5298);
or U6601 (N_6601,N_5076,N_5520);
or U6602 (N_6602,N_5845,N_5838);
and U6603 (N_6603,N_5004,N_5174);
nand U6604 (N_6604,N_5339,N_5996);
nand U6605 (N_6605,N_5934,N_5191);
nand U6606 (N_6606,N_5519,N_5479);
or U6607 (N_6607,N_5819,N_5623);
nand U6608 (N_6608,N_5091,N_5484);
and U6609 (N_6609,N_5070,N_5280);
and U6610 (N_6610,N_5402,N_5558);
nand U6611 (N_6611,N_5982,N_5265);
or U6612 (N_6612,N_5904,N_5696);
nor U6613 (N_6613,N_5260,N_5297);
nor U6614 (N_6614,N_5920,N_5393);
or U6615 (N_6615,N_5750,N_5409);
nor U6616 (N_6616,N_5290,N_5364);
nor U6617 (N_6617,N_5875,N_5381);
nand U6618 (N_6618,N_5232,N_5735);
and U6619 (N_6619,N_5695,N_5803);
nor U6620 (N_6620,N_5338,N_5518);
nand U6621 (N_6621,N_5729,N_5466);
and U6622 (N_6622,N_5161,N_5604);
and U6623 (N_6623,N_5466,N_5809);
nand U6624 (N_6624,N_5318,N_5033);
nor U6625 (N_6625,N_5464,N_5015);
and U6626 (N_6626,N_5966,N_5129);
nand U6627 (N_6627,N_5592,N_5890);
nor U6628 (N_6628,N_5040,N_5689);
nor U6629 (N_6629,N_5383,N_5410);
or U6630 (N_6630,N_5407,N_5321);
and U6631 (N_6631,N_5789,N_5424);
nor U6632 (N_6632,N_5324,N_5088);
and U6633 (N_6633,N_5340,N_5006);
xor U6634 (N_6634,N_5353,N_5878);
nor U6635 (N_6635,N_5673,N_5719);
or U6636 (N_6636,N_5186,N_5801);
nor U6637 (N_6637,N_5446,N_5612);
xor U6638 (N_6638,N_5650,N_5504);
and U6639 (N_6639,N_5433,N_5495);
and U6640 (N_6640,N_5804,N_5056);
or U6641 (N_6641,N_5692,N_5980);
xnor U6642 (N_6642,N_5020,N_5730);
and U6643 (N_6643,N_5516,N_5878);
and U6644 (N_6644,N_5967,N_5531);
or U6645 (N_6645,N_5103,N_5974);
and U6646 (N_6646,N_5451,N_5093);
and U6647 (N_6647,N_5727,N_5218);
and U6648 (N_6648,N_5034,N_5942);
and U6649 (N_6649,N_5021,N_5163);
nand U6650 (N_6650,N_5338,N_5165);
nor U6651 (N_6651,N_5536,N_5868);
and U6652 (N_6652,N_5220,N_5715);
xor U6653 (N_6653,N_5723,N_5288);
nor U6654 (N_6654,N_5142,N_5030);
nand U6655 (N_6655,N_5455,N_5117);
or U6656 (N_6656,N_5772,N_5109);
nor U6657 (N_6657,N_5604,N_5981);
and U6658 (N_6658,N_5092,N_5863);
nand U6659 (N_6659,N_5992,N_5335);
nor U6660 (N_6660,N_5986,N_5980);
nand U6661 (N_6661,N_5415,N_5107);
and U6662 (N_6662,N_5893,N_5077);
xor U6663 (N_6663,N_5387,N_5345);
nor U6664 (N_6664,N_5574,N_5434);
and U6665 (N_6665,N_5457,N_5261);
nor U6666 (N_6666,N_5688,N_5365);
nand U6667 (N_6667,N_5410,N_5000);
and U6668 (N_6668,N_5370,N_5881);
nand U6669 (N_6669,N_5341,N_5389);
nand U6670 (N_6670,N_5545,N_5733);
nand U6671 (N_6671,N_5683,N_5871);
or U6672 (N_6672,N_5773,N_5383);
and U6673 (N_6673,N_5049,N_5482);
and U6674 (N_6674,N_5095,N_5142);
nor U6675 (N_6675,N_5029,N_5509);
nand U6676 (N_6676,N_5867,N_5040);
xor U6677 (N_6677,N_5237,N_5178);
and U6678 (N_6678,N_5973,N_5754);
or U6679 (N_6679,N_5637,N_5667);
and U6680 (N_6680,N_5054,N_5112);
nor U6681 (N_6681,N_5653,N_5270);
and U6682 (N_6682,N_5912,N_5297);
and U6683 (N_6683,N_5422,N_5922);
nor U6684 (N_6684,N_5845,N_5141);
and U6685 (N_6685,N_5676,N_5533);
and U6686 (N_6686,N_5351,N_5206);
and U6687 (N_6687,N_5921,N_5504);
or U6688 (N_6688,N_5959,N_5432);
or U6689 (N_6689,N_5813,N_5810);
nand U6690 (N_6690,N_5347,N_5038);
xnor U6691 (N_6691,N_5001,N_5125);
nand U6692 (N_6692,N_5973,N_5704);
nand U6693 (N_6693,N_5687,N_5933);
nor U6694 (N_6694,N_5394,N_5281);
nand U6695 (N_6695,N_5982,N_5461);
or U6696 (N_6696,N_5467,N_5230);
and U6697 (N_6697,N_5206,N_5372);
xnor U6698 (N_6698,N_5924,N_5919);
nor U6699 (N_6699,N_5034,N_5654);
and U6700 (N_6700,N_5625,N_5633);
nor U6701 (N_6701,N_5393,N_5436);
xor U6702 (N_6702,N_5589,N_5427);
xor U6703 (N_6703,N_5453,N_5740);
and U6704 (N_6704,N_5135,N_5919);
nor U6705 (N_6705,N_5829,N_5571);
nand U6706 (N_6706,N_5766,N_5457);
nor U6707 (N_6707,N_5042,N_5809);
nand U6708 (N_6708,N_5536,N_5672);
nor U6709 (N_6709,N_5105,N_5180);
nand U6710 (N_6710,N_5022,N_5104);
and U6711 (N_6711,N_5442,N_5921);
or U6712 (N_6712,N_5115,N_5948);
and U6713 (N_6713,N_5606,N_5186);
nor U6714 (N_6714,N_5314,N_5336);
nor U6715 (N_6715,N_5484,N_5033);
nand U6716 (N_6716,N_5586,N_5796);
nor U6717 (N_6717,N_5219,N_5078);
or U6718 (N_6718,N_5043,N_5426);
nand U6719 (N_6719,N_5248,N_5756);
xor U6720 (N_6720,N_5020,N_5982);
or U6721 (N_6721,N_5646,N_5833);
nand U6722 (N_6722,N_5687,N_5526);
nand U6723 (N_6723,N_5601,N_5777);
and U6724 (N_6724,N_5922,N_5828);
and U6725 (N_6725,N_5054,N_5707);
xor U6726 (N_6726,N_5855,N_5675);
nand U6727 (N_6727,N_5510,N_5021);
nand U6728 (N_6728,N_5411,N_5498);
or U6729 (N_6729,N_5877,N_5978);
xnor U6730 (N_6730,N_5086,N_5985);
nand U6731 (N_6731,N_5717,N_5012);
and U6732 (N_6732,N_5862,N_5894);
or U6733 (N_6733,N_5243,N_5161);
nor U6734 (N_6734,N_5571,N_5855);
nor U6735 (N_6735,N_5949,N_5425);
and U6736 (N_6736,N_5320,N_5810);
nor U6737 (N_6737,N_5663,N_5342);
nand U6738 (N_6738,N_5382,N_5161);
xor U6739 (N_6739,N_5809,N_5402);
or U6740 (N_6740,N_5122,N_5390);
and U6741 (N_6741,N_5705,N_5240);
nand U6742 (N_6742,N_5573,N_5750);
xnor U6743 (N_6743,N_5316,N_5959);
nand U6744 (N_6744,N_5436,N_5682);
nand U6745 (N_6745,N_5539,N_5436);
and U6746 (N_6746,N_5256,N_5794);
and U6747 (N_6747,N_5928,N_5043);
nand U6748 (N_6748,N_5266,N_5866);
nand U6749 (N_6749,N_5459,N_5140);
or U6750 (N_6750,N_5200,N_5781);
xor U6751 (N_6751,N_5699,N_5349);
nand U6752 (N_6752,N_5755,N_5641);
nand U6753 (N_6753,N_5231,N_5959);
and U6754 (N_6754,N_5266,N_5117);
xor U6755 (N_6755,N_5935,N_5226);
nor U6756 (N_6756,N_5551,N_5690);
or U6757 (N_6757,N_5670,N_5669);
and U6758 (N_6758,N_5808,N_5746);
or U6759 (N_6759,N_5830,N_5518);
nor U6760 (N_6760,N_5982,N_5683);
or U6761 (N_6761,N_5232,N_5198);
nor U6762 (N_6762,N_5410,N_5623);
or U6763 (N_6763,N_5502,N_5274);
nor U6764 (N_6764,N_5127,N_5714);
nand U6765 (N_6765,N_5417,N_5284);
nor U6766 (N_6766,N_5461,N_5100);
and U6767 (N_6767,N_5480,N_5251);
nor U6768 (N_6768,N_5669,N_5300);
nand U6769 (N_6769,N_5014,N_5486);
and U6770 (N_6770,N_5663,N_5445);
nand U6771 (N_6771,N_5056,N_5665);
xnor U6772 (N_6772,N_5672,N_5542);
or U6773 (N_6773,N_5785,N_5970);
nand U6774 (N_6774,N_5967,N_5400);
or U6775 (N_6775,N_5293,N_5729);
and U6776 (N_6776,N_5773,N_5811);
nand U6777 (N_6777,N_5759,N_5051);
and U6778 (N_6778,N_5210,N_5181);
nand U6779 (N_6779,N_5857,N_5429);
and U6780 (N_6780,N_5661,N_5897);
xor U6781 (N_6781,N_5661,N_5087);
and U6782 (N_6782,N_5976,N_5085);
or U6783 (N_6783,N_5671,N_5650);
nor U6784 (N_6784,N_5403,N_5827);
nor U6785 (N_6785,N_5164,N_5577);
or U6786 (N_6786,N_5998,N_5400);
nor U6787 (N_6787,N_5268,N_5770);
and U6788 (N_6788,N_5043,N_5291);
nor U6789 (N_6789,N_5052,N_5379);
xnor U6790 (N_6790,N_5283,N_5123);
and U6791 (N_6791,N_5840,N_5983);
nor U6792 (N_6792,N_5258,N_5950);
nand U6793 (N_6793,N_5011,N_5503);
nand U6794 (N_6794,N_5545,N_5461);
or U6795 (N_6795,N_5267,N_5209);
xnor U6796 (N_6796,N_5013,N_5596);
nor U6797 (N_6797,N_5508,N_5705);
or U6798 (N_6798,N_5285,N_5015);
nand U6799 (N_6799,N_5750,N_5213);
and U6800 (N_6800,N_5000,N_5142);
nor U6801 (N_6801,N_5781,N_5645);
nand U6802 (N_6802,N_5383,N_5091);
nand U6803 (N_6803,N_5951,N_5632);
nor U6804 (N_6804,N_5731,N_5609);
or U6805 (N_6805,N_5902,N_5862);
and U6806 (N_6806,N_5478,N_5030);
or U6807 (N_6807,N_5895,N_5926);
or U6808 (N_6808,N_5684,N_5351);
nand U6809 (N_6809,N_5439,N_5299);
and U6810 (N_6810,N_5439,N_5367);
nand U6811 (N_6811,N_5024,N_5743);
and U6812 (N_6812,N_5378,N_5449);
nor U6813 (N_6813,N_5982,N_5589);
and U6814 (N_6814,N_5280,N_5644);
nand U6815 (N_6815,N_5767,N_5371);
nand U6816 (N_6816,N_5482,N_5629);
nand U6817 (N_6817,N_5791,N_5537);
nand U6818 (N_6818,N_5483,N_5555);
and U6819 (N_6819,N_5686,N_5371);
nand U6820 (N_6820,N_5650,N_5688);
nand U6821 (N_6821,N_5221,N_5649);
nand U6822 (N_6822,N_5554,N_5690);
and U6823 (N_6823,N_5560,N_5886);
nor U6824 (N_6824,N_5006,N_5926);
nor U6825 (N_6825,N_5857,N_5549);
nand U6826 (N_6826,N_5759,N_5861);
nand U6827 (N_6827,N_5467,N_5531);
nor U6828 (N_6828,N_5225,N_5368);
nand U6829 (N_6829,N_5157,N_5435);
nor U6830 (N_6830,N_5576,N_5496);
nand U6831 (N_6831,N_5947,N_5609);
and U6832 (N_6832,N_5270,N_5562);
and U6833 (N_6833,N_5085,N_5956);
or U6834 (N_6834,N_5456,N_5887);
nor U6835 (N_6835,N_5837,N_5546);
nor U6836 (N_6836,N_5432,N_5442);
or U6837 (N_6837,N_5074,N_5876);
or U6838 (N_6838,N_5555,N_5553);
nand U6839 (N_6839,N_5267,N_5727);
or U6840 (N_6840,N_5117,N_5791);
and U6841 (N_6841,N_5777,N_5604);
and U6842 (N_6842,N_5747,N_5600);
or U6843 (N_6843,N_5159,N_5693);
nand U6844 (N_6844,N_5698,N_5800);
or U6845 (N_6845,N_5872,N_5441);
or U6846 (N_6846,N_5521,N_5502);
or U6847 (N_6847,N_5558,N_5172);
xnor U6848 (N_6848,N_5391,N_5190);
xnor U6849 (N_6849,N_5701,N_5746);
nor U6850 (N_6850,N_5280,N_5869);
nor U6851 (N_6851,N_5463,N_5820);
nor U6852 (N_6852,N_5636,N_5322);
nand U6853 (N_6853,N_5466,N_5354);
or U6854 (N_6854,N_5382,N_5354);
nand U6855 (N_6855,N_5388,N_5869);
or U6856 (N_6856,N_5920,N_5542);
and U6857 (N_6857,N_5892,N_5198);
or U6858 (N_6858,N_5864,N_5893);
nand U6859 (N_6859,N_5207,N_5892);
and U6860 (N_6860,N_5145,N_5470);
nor U6861 (N_6861,N_5357,N_5373);
nand U6862 (N_6862,N_5194,N_5930);
nor U6863 (N_6863,N_5275,N_5639);
nor U6864 (N_6864,N_5915,N_5375);
or U6865 (N_6865,N_5527,N_5470);
and U6866 (N_6866,N_5493,N_5567);
nor U6867 (N_6867,N_5554,N_5248);
nand U6868 (N_6868,N_5168,N_5325);
xor U6869 (N_6869,N_5665,N_5603);
nand U6870 (N_6870,N_5111,N_5426);
or U6871 (N_6871,N_5238,N_5745);
or U6872 (N_6872,N_5603,N_5875);
nor U6873 (N_6873,N_5911,N_5802);
xnor U6874 (N_6874,N_5578,N_5928);
nor U6875 (N_6875,N_5710,N_5761);
or U6876 (N_6876,N_5840,N_5156);
xnor U6877 (N_6877,N_5605,N_5947);
nand U6878 (N_6878,N_5612,N_5237);
nor U6879 (N_6879,N_5763,N_5782);
or U6880 (N_6880,N_5878,N_5255);
xor U6881 (N_6881,N_5545,N_5414);
xnor U6882 (N_6882,N_5544,N_5058);
nand U6883 (N_6883,N_5143,N_5126);
nand U6884 (N_6884,N_5475,N_5947);
nor U6885 (N_6885,N_5731,N_5675);
and U6886 (N_6886,N_5162,N_5037);
nor U6887 (N_6887,N_5167,N_5739);
nor U6888 (N_6888,N_5343,N_5807);
nor U6889 (N_6889,N_5400,N_5910);
xnor U6890 (N_6890,N_5267,N_5466);
and U6891 (N_6891,N_5317,N_5330);
and U6892 (N_6892,N_5077,N_5265);
xor U6893 (N_6893,N_5911,N_5182);
xnor U6894 (N_6894,N_5980,N_5899);
nand U6895 (N_6895,N_5594,N_5609);
nand U6896 (N_6896,N_5323,N_5963);
and U6897 (N_6897,N_5186,N_5942);
nand U6898 (N_6898,N_5935,N_5673);
nand U6899 (N_6899,N_5028,N_5915);
and U6900 (N_6900,N_5416,N_5713);
or U6901 (N_6901,N_5112,N_5443);
or U6902 (N_6902,N_5793,N_5732);
or U6903 (N_6903,N_5246,N_5411);
nor U6904 (N_6904,N_5173,N_5871);
or U6905 (N_6905,N_5870,N_5833);
or U6906 (N_6906,N_5229,N_5265);
and U6907 (N_6907,N_5887,N_5550);
or U6908 (N_6908,N_5133,N_5223);
nor U6909 (N_6909,N_5496,N_5507);
or U6910 (N_6910,N_5643,N_5214);
or U6911 (N_6911,N_5204,N_5931);
and U6912 (N_6912,N_5950,N_5517);
nand U6913 (N_6913,N_5716,N_5485);
nor U6914 (N_6914,N_5930,N_5849);
and U6915 (N_6915,N_5980,N_5151);
xnor U6916 (N_6916,N_5075,N_5607);
or U6917 (N_6917,N_5797,N_5859);
nand U6918 (N_6918,N_5605,N_5032);
nor U6919 (N_6919,N_5402,N_5123);
nor U6920 (N_6920,N_5703,N_5636);
nand U6921 (N_6921,N_5193,N_5217);
nand U6922 (N_6922,N_5183,N_5718);
nor U6923 (N_6923,N_5812,N_5880);
nor U6924 (N_6924,N_5780,N_5671);
and U6925 (N_6925,N_5339,N_5467);
or U6926 (N_6926,N_5527,N_5973);
or U6927 (N_6927,N_5937,N_5031);
and U6928 (N_6928,N_5342,N_5728);
nand U6929 (N_6929,N_5517,N_5740);
xor U6930 (N_6930,N_5845,N_5411);
and U6931 (N_6931,N_5031,N_5906);
nor U6932 (N_6932,N_5992,N_5494);
or U6933 (N_6933,N_5795,N_5548);
nor U6934 (N_6934,N_5101,N_5323);
xnor U6935 (N_6935,N_5516,N_5446);
nor U6936 (N_6936,N_5243,N_5849);
and U6937 (N_6937,N_5951,N_5557);
or U6938 (N_6938,N_5847,N_5642);
and U6939 (N_6939,N_5949,N_5870);
nand U6940 (N_6940,N_5489,N_5169);
nand U6941 (N_6941,N_5171,N_5819);
or U6942 (N_6942,N_5457,N_5543);
nand U6943 (N_6943,N_5097,N_5672);
nand U6944 (N_6944,N_5704,N_5516);
nor U6945 (N_6945,N_5795,N_5088);
nor U6946 (N_6946,N_5153,N_5599);
and U6947 (N_6947,N_5162,N_5335);
xnor U6948 (N_6948,N_5274,N_5470);
nand U6949 (N_6949,N_5339,N_5086);
xor U6950 (N_6950,N_5258,N_5810);
or U6951 (N_6951,N_5583,N_5129);
xor U6952 (N_6952,N_5996,N_5358);
nand U6953 (N_6953,N_5310,N_5438);
nand U6954 (N_6954,N_5726,N_5833);
or U6955 (N_6955,N_5959,N_5858);
nand U6956 (N_6956,N_5597,N_5111);
or U6957 (N_6957,N_5186,N_5321);
and U6958 (N_6958,N_5487,N_5413);
and U6959 (N_6959,N_5395,N_5047);
nor U6960 (N_6960,N_5118,N_5007);
or U6961 (N_6961,N_5866,N_5967);
xor U6962 (N_6962,N_5475,N_5407);
nor U6963 (N_6963,N_5536,N_5264);
or U6964 (N_6964,N_5557,N_5865);
or U6965 (N_6965,N_5523,N_5119);
or U6966 (N_6966,N_5283,N_5146);
or U6967 (N_6967,N_5304,N_5374);
nor U6968 (N_6968,N_5637,N_5455);
nor U6969 (N_6969,N_5338,N_5686);
and U6970 (N_6970,N_5529,N_5667);
nor U6971 (N_6971,N_5252,N_5039);
or U6972 (N_6972,N_5980,N_5243);
and U6973 (N_6973,N_5189,N_5826);
or U6974 (N_6974,N_5427,N_5181);
nand U6975 (N_6975,N_5440,N_5318);
or U6976 (N_6976,N_5798,N_5008);
nand U6977 (N_6977,N_5742,N_5892);
nand U6978 (N_6978,N_5508,N_5158);
xor U6979 (N_6979,N_5400,N_5125);
nor U6980 (N_6980,N_5247,N_5388);
xor U6981 (N_6981,N_5714,N_5308);
nand U6982 (N_6982,N_5827,N_5277);
nand U6983 (N_6983,N_5607,N_5238);
nor U6984 (N_6984,N_5291,N_5605);
and U6985 (N_6985,N_5754,N_5478);
or U6986 (N_6986,N_5671,N_5892);
and U6987 (N_6987,N_5289,N_5367);
and U6988 (N_6988,N_5050,N_5989);
and U6989 (N_6989,N_5115,N_5187);
nand U6990 (N_6990,N_5142,N_5489);
nor U6991 (N_6991,N_5294,N_5276);
xor U6992 (N_6992,N_5922,N_5638);
nand U6993 (N_6993,N_5337,N_5784);
nand U6994 (N_6994,N_5221,N_5717);
or U6995 (N_6995,N_5332,N_5696);
nand U6996 (N_6996,N_5431,N_5276);
nand U6997 (N_6997,N_5105,N_5244);
nor U6998 (N_6998,N_5217,N_5082);
and U6999 (N_6999,N_5232,N_5880);
nor U7000 (N_7000,N_6928,N_6720);
and U7001 (N_7001,N_6294,N_6416);
or U7002 (N_7002,N_6120,N_6451);
xor U7003 (N_7003,N_6556,N_6484);
and U7004 (N_7004,N_6076,N_6319);
or U7005 (N_7005,N_6941,N_6985);
or U7006 (N_7006,N_6667,N_6645);
and U7007 (N_7007,N_6878,N_6192);
nand U7008 (N_7008,N_6783,N_6988);
or U7009 (N_7009,N_6763,N_6068);
nor U7010 (N_7010,N_6249,N_6333);
and U7011 (N_7011,N_6111,N_6220);
xor U7012 (N_7012,N_6465,N_6526);
nand U7013 (N_7013,N_6108,N_6398);
and U7014 (N_7014,N_6123,N_6149);
or U7015 (N_7015,N_6103,N_6989);
or U7016 (N_7016,N_6277,N_6724);
nand U7017 (N_7017,N_6512,N_6480);
and U7018 (N_7018,N_6019,N_6182);
nor U7019 (N_7019,N_6644,N_6106);
nand U7020 (N_7020,N_6819,N_6658);
nand U7021 (N_7021,N_6976,N_6715);
or U7022 (N_7022,N_6742,N_6848);
xor U7023 (N_7023,N_6893,N_6823);
or U7024 (N_7024,N_6486,N_6891);
nand U7025 (N_7025,N_6650,N_6520);
or U7026 (N_7026,N_6534,N_6402);
nor U7027 (N_7027,N_6730,N_6401);
nor U7028 (N_7028,N_6688,N_6280);
or U7029 (N_7029,N_6359,N_6602);
nor U7030 (N_7030,N_6614,N_6990);
nor U7031 (N_7031,N_6437,N_6394);
nor U7032 (N_7032,N_6139,N_6231);
xor U7033 (N_7033,N_6272,N_6721);
and U7034 (N_7034,N_6306,N_6755);
nor U7035 (N_7035,N_6154,N_6221);
nand U7036 (N_7036,N_6807,N_6489);
or U7037 (N_7037,N_6565,N_6675);
and U7038 (N_7038,N_6919,N_6148);
nand U7039 (N_7039,N_6685,N_6411);
nor U7040 (N_7040,N_6942,N_6922);
nor U7041 (N_7041,N_6168,N_6733);
or U7042 (N_7042,N_6629,N_6442);
or U7043 (N_7043,N_6234,N_6117);
and U7044 (N_7044,N_6744,N_6821);
or U7045 (N_7045,N_6956,N_6379);
nand U7046 (N_7046,N_6438,N_6992);
nand U7047 (N_7047,N_6110,N_6939);
and U7048 (N_7048,N_6900,N_6918);
or U7049 (N_7049,N_6146,N_6176);
nand U7050 (N_7050,N_6767,N_6548);
nand U7051 (N_7051,N_6226,N_6632);
nor U7052 (N_7052,N_6912,N_6916);
nand U7053 (N_7053,N_6395,N_6017);
and U7054 (N_7054,N_6892,N_6274);
nand U7055 (N_7055,N_6591,N_6731);
and U7056 (N_7056,N_6261,N_6251);
nor U7057 (N_7057,N_6032,N_6809);
and U7058 (N_7058,N_6266,N_6498);
nand U7059 (N_7059,N_6085,N_6356);
nor U7060 (N_7060,N_6430,N_6026);
nand U7061 (N_7061,N_6870,N_6612);
nor U7062 (N_7062,N_6346,N_6616);
and U7063 (N_7063,N_6004,N_6608);
or U7064 (N_7064,N_6115,N_6842);
and U7065 (N_7065,N_6392,N_6164);
nand U7066 (N_7066,N_6178,N_6736);
nand U7067 (N_7067,N_6530,N_6672);
nor U7068 (N_7068,N_6296,N_6691);
and U7069 (N_7069,N_6888,N_6641);
nand U7070 (N_7070,N_6194,N_6706);
nand U7071 (N_7071,N_6128,N_6083);
nand U7072 (N_7072,N_6621,N_6069);
nor U7073 (N_7073,N_6122,N_6041);
and U7074 (N_7074,N_6126,N_6061);
and U7075 (N_7075,N_6967,N_6826);
nand U7076 (N_7076,N_6134,N_6332);
and U7077 (N_7077,N_6406,N_6087);
and U7078 (N_7078,N_6105,N_6660);
xor U7079 (N_7079,N_6801,N_6837);
nor U7080 (N_7080,N_6674,N_6639);
xor U7081 (N_7081,N_6160,N_6790);
nor U7082 (N_7082,N_6454,N_6378);
and U7083 (N_7083,N_6439,N_6716);
nor U7084 (N_7084,N_6093,N_6404);
nor U7085 (N_7085,N_6734,N_6517);
and U7086 (N_7086,N_6034,N_6417);
and U7087 (N_7087,N_6940,N_6228);
nand U7088 (N_7088,N_6066,N_6222);
and U7089 (N_7089,N_6422,N_6005);
nand U7090 (N_7090,N_6380,N_6540);
xnor U7091 (N_7091,N_6633,N_6453);
or U7092 (N_7092,N_6092,N_6574);
and U7093 (N_7093,N_6348,N_6758);
nor U7094 (N_7094,N_6230,N_6963);
xnor U7095 (N_7095,N_6329,N_6118);
or U7096 (N_7096,N_6448,N_6338);
xor U7097 (N_7097,N_6046,N_6945);
nor U7098 (N_7098,N_6617,N_6856);
and U7099 (N_7099,N_6622,N_6365);
nand U7100 (N_7100,N_6743,N_6702);
and U7101 (N_7101,N_6682,N_6000);
and U7102 (N_7102,N_6493,N_6711);
and U7103 (N_7103,N_6590,N_6474);
nand U7104 (N_7104,N_6390,N_6838);
or U7105 (N_7105,N_6127,N_6603);
nor U7106 (N_7106,N_6803,N_6132);
nand U7107 (N_7107,N_6213,N_6492);
xor U7108 (N_7108,N_6926,N_6854);
nor U7109 (N_7109,N_6640,N_6693);
nand U7110 (N_7110,N_6152,N_6853);
nand U7111 (N_7111,N_6352,N_6528);
and U7112 (N_7112,N_6491,N_6973);
and U7113 (N_7113,N_6840,N_6423);
nor U7114 (N_7114,N_6031,N_6812);
nand U7115 (N_7115,N_6445,N_6981);
or U7116 (N_7116,N_6172,N_6158);
nor U7117 (N_7117,N_6206,N_6375);
or U7118 (N_7118,N_6415,N_6909);
or U7119 (N_7119,N_6216,N_6186);
nand U7120 (N_7120,N_6499,N_6875);
and U7121 (N_7121,N_6382,N_6147);
and U7122 (N_7122,N_6386,N_6314);
and U7123 (N_7123,N_6174,N_6615);
nor U7124 (N_7124,N_6999,N_6456);
and U7125 (N_7125,N_6930,N_6855);
nand U7126 (N_7126,N_6572,N_6121);
nand U7127 (N_7127,N_6773,N_6690);
nand U7128 (N_7128,N_6156,N_6472);
nand U7129 (N_7129,N_6585,N_6798);
nor U7130 (N_7130,N_6131,N_6412);
nor U7131 (N_7131,N_6424,N_6259);
nand U7132 (N_7132,N_6817,N_6924);
or U7133 (N_7133,N_6481,N_6765);
nor U7134 (N_7134,N_6063,N_6920);
or U7135 (N_7135,N_6543,N_6113);
or U7136 (N_7136,N_6188,N_6421);
nor U7137 (N_7137,N_6897,N_6223);
nor U7138 (N_7138,N_6255,N_6044);
nand U7139 (N_7139,N_6307,N_6908);
or U7140 (N_7140,N_6818,N_6029);
xnor U7141 (N_7141,N_6579,N_6756);
and U7142 (N_7142,N_6661,N_6538);
xor U7143 (N_7143,N_6880,N_6883);
and U7144 (N_7144,N_6712,N_6642);
and U7145 (N_7145,N_6171,N_6604);
nand U7146 (N_7146,N_6566,N_6646);
and U7147 (N_7147,N_6677,N_6657);
xor U7148 (N_7148,N_6845,N_6710);
xnor U7149 (N_7149,N_6052,N_6905);
xor U7150 (N_7150,N_6876,N_6898);
or U7151 (N_7151,N_6678,N_6769);
nor U7152 (N_7152,N_6847,N_6511);
and U7153 (N_7153,N_6894,N_6931);
or U7154 (N_7154,N_6606,N_6982);
nor U7155 (N_7155,N_6822,N_6850);
or U7156 (N_7156,N_6537,N_6064);
or U7157 (N_7157,N_6978,N_6806);
xnor U7158 (N_7158,N_6620,N_6351);
and U7159 (N_7159,N_6205,N_6473);
xnor U7160 (N_7160,N_6835,N_6746);
and U7161 (N_7161,N_6244,N_6977);
and U7162 (N_7162,N_6671,N_6676);
nor U7163 (N_7163,N_6915,N_6596);
or U7164 (N_7164,N_6887,N_6441);
nor U7165 (N_7165,N_6789,N_6839);
nand U7166 (N_7166,N_6488,N_6525);
nor U7167 (N_7167,N_6181,N_6513);
xnor U7168 (N_7168,N_6331,N_6503);
nand U7169 (N_7169,N_6065,N_6409);
nand U7170 (N_7170,N_6387,N_6549);
or U7171 (N_7171,N_6696,N_6198);
and U7172 (N_7172,N_6637,N_6050);
nor U7173 (N_7173,N_6597,N_6270);
and U7174 (N_7174,N_6284,N_6373);
nand U7175 (N_7175,N_6634,N_6080);
or U7176 (N_7176,N_6607,N_6058);
xnor U7177 (N_7177,N_6384,N_6295);
nor U7178 (N_7178,N_6429,N_6844);
or U7179 (N_7179,N_6325,N_6780);
and U7180 (N_7180,N_6166,N_6405);
nand U7181 (N_7181,N_6399,N_6679);
nor U7182 (N_7182,N_6635,N_6729);
xor U7183 (N_7183,N_6910,N_6025);
xnor U7184 (N_7184,N_6955,N_6136);
nor U7185 (N_7185,N_6062,N_6101);
nor U7186 (N_7186,N_6167,N_6015);
nand U7187 (N_7187,N_6655,N_6033);
and U7188 (N_7188,N_6177,N_6313);
nand U7189 (N_7189,N_6771,N_6190);
nor U7190 (N_7190,N_6252,N_6310);
nand U7191 (N_7191,N_6355,N_6628);
nand U7192 (N_7192,N_6072,N_6954);
or U7193 (N_7193,N_6881,N_6775);
and U7194 (N_7194,N_6248,N_6722);
nor U7195 (N_7195,N_6368,N_6383);
or U7196 (N_7196,N_6593,N_6761);
and U7197 (N_7197,N_6197,N_6584);
xor U7198 (N_7198,N_6573,N_6119);
nand U7199 (N_7199,N_6485,N_6779);
nand U7200 (N_7200,N_6539,N_6400);
nand U7201 (N_7201,N_6476,N_6708);
nor U7202 (N_7202,N_6267,N_6408);
and U7203 (N_7203,N_6559,N_6938);
nand U7204 (N_7204,N_6038,N_6449);
and U7205 (N_7205,N_6654,N_6218);
and U7206 (N_7206,N_6890,N_6723);
or U7207 (N_7207,N_6447,N_6247);
nor U7208 (N_7208,N_6774,N_6345);
and U7209 (N_7209,N_6324,N_6011);
and U7210 (N_7210,N_6665,N_6994);
nand U7211 (N_7211,N_6958,N_6263);
xnor U7212 (N_7212,N_6462,N_6626);
xnor U7213 (N_7213,N_6440,N_6300);
or U7214 (N_7214,N_6529,N_6960);
or U7215 (N_7215,N_6500,N_6290);
nand U7216 (N_7216,N_6814,N_6618);
or U7217 (N_7217,N_6811,N_6023);
and U7218 (N_7218,N_6354,N_6185);
nor U7219 (N_7219,N_6291,N_6159);
nor U7220 (N_7220,N_6283,N_6232);
and U7221 (N_7221,N_6991,N_6053);
nor U7222 (N_7222,N_6951,N_6518);
and U7223 (N_7223,N_6464,N_6326);
nand U7224 (N_7224,N_6911,N_6601);
or U7225 (N_7225,N_6824,N_6074);
nand U7226 (N_7226,N_6795,N_6630);
nand U7227 (N_7227,N_6212,N_6145);
nor U7228 (N_7228,N_6141,N_6843);
and U7229 (N_7229,N_6804,N_6670);
nor U7230 (N_7230,N_6010,N_6575);
or U7231 (N_7231,N_6143,N_6446);
nand U7232 (N_7232,N_6563,N_6717);
nand U7233 (N_7233,N_6552,N_6129);
nor U7234 (N_7234,N_6229,N_6577);
nor U7235 (N_7235,N_6479,N_6376);
nor U7236 (N_7236,N_6169,N_6902);
and U7237 (N_7237,N_6664,N_6377);
or U7238 (N_7238,N_6656,N_6070);
or U7239 (N_7239,N_6201,N_6002);
and U7240 (N_7240,N_6980,N_6210);
nor U7241 (N_7241,N_6458,N_6993);
xor U7242 (N_7242,N_6987,N_6582);
or U7243 (N_7243,N_6813,N_6934);
xnor U7244 (N_7244,N_6625,N_6996);
or U7245 (N_7245,N_6768,N_6700);
and U7246 (N_7246,N_6868,N_6865);
nor U7247 (N_7247,N_6998,N_6482);
nand U7248 (N_7248,N_6086,N_6250);
nand U7249 (N_7249,N_6689,N_6704);
and U7250 (N_7250,N_6820,N_6214);
nand U7251 (N_7251,N_6815,N_6873);
or U7252 (N_7252,N_6112,N_6578);
or U7253 (N_7253,N_6753,N_6531);
nand U7254 (N_7254,N_6344,N_6293);
nor U7255 (N_7255,N_6079,N_6653);
nor U7256 (N_7256,N_6834,N_6305);
nand U7257 (N_7257,N_6935,N_6183);
xnor U7258 (N_7258,N_6547,N_6242);
nand U7259 (N_7259,N_6832,N_6673);
xor U7260 (N_7260,N_6288,N_6564);
or U7261 (N_7261,N_6339,N_6098);
nand U7262 (N_7262,N_6372,N_6490);
nor U7263 (N_7263,N_6937,N_6810);
nor U7264 (N_7264,N_6278,N_6757);
and U7265 (N_7265,N_6195,N_6760);
and U7266 (N_7266,N_6580,N_6199);
xnor U7267 (N_7267,N_6235,N_6081);
nand U7268 (N_7268,N_6546,N_6703);
or U7269 (N_7269,N_6858,N_6516);
nand U7270 (N_7270,N_6340,N_6791);
xnor U7271 (N_7271,N_6239,N_6133);
xnor U7272 (N_7272,N_6778,N_6877);
nor U7273 (N_7273,N_6180,N_6289);
or U7274 (N_7274,N_6867,N_6385);
and U7275 (N_7275,N_6965,N_6561);
or U7276 (N_7276,N_6827,N_6505);
or U7277 (N_7277,N_6478,N_6745);
xnor U7278 (N_7278,N_6586,N_6611);
nand U7279 (N_7279,N_6045,N_6107);
and U7280 (N_7280,N_6899,N_6260);
or U7281 (N_7281,N_6397,N_6381);
nor U7282 (N_7282,N_6638,N_6794);
nor U7283 (N_7283,N_6754,N_6833);
nand U7284 (N_7284,N_6797,N_6871);
or U7285 (N_7285,N_6959,N_6496);
nand U7286 (N_7286,N_6619,N_6841);
nor U7287 (N_7287,N_6581,N_6162);
xnor U7288 (N_7288,N_6784,N_6140);
nor U7289 (N_7289,N_6950,N_6627);
or U7290 (N_7290,N_6849,N_6862);
nand U7291 (N_7291,N_6202,N_6320);
nor U7292 (N_7292,N_6388,N_6738);
and U7293 (N_7293,N_6903,N_6191);
nand U7294 (N_7294,N_6013,N_6923);
and U7295 (N_7295,N_6506,N_6455);
and U7296 (N_7296,N_6217,N_6859);
nor U7297 (N_7297,N_6613,N_6321);
and U7298 (N_7298,N_6334,N_6330);
or U7299 (N_7299,N_6589,N_6460);
or U7300 (N_7300,N_6913,N_6109);
and U7301 (N_7301,N_6308,N_6944);
and U7302 (N_7302,N_6090,N_6037);
nor U7303 (N_7303,N_6253,N_6906);
nor U7304 (N_7304,N_6904,N_6957);
nand U7305 (N_7305,N_6649,N_6009);
nor U7306 (N_7306,N_6343,N_6759);
and U7307 (N_7307,N_6886,N_6522);
or U7308 (N_7308,N_6749,N_6137);
and U7309 (N_7309,N_6692,N_6508);
or U7310 (N_7310,N_6555,N_6925);
and U7311 (N_7311,N_6495,N_6135);
and U7312 (N_7312,N_6125,N_6599);
or U7313 (N_7313,N_6802,N_6327);
or U7314 (N_7314,N_6468,N_6747);
or U7315 (N_7315,N_6907,N_6542);
and U7316 (N_7316,N_6636,N_6095);
or U7317 (N_7317,N_6371,N_6816);
xnor U7318 (N_7318,N_6554,N_6788);
nor U7319 (N_7319,N_6825,N_6681);
and U7320 (N_7320,N_6917,N_6510);
nand U7321 (N_7321,N_6161,N_6983);
and U7322 (N_7322,N_6187,N_6457);
and U7323 (N_7323,N_6772,N_6787);
nand U7324 (N_7324,N_6281,N_6874);
nand U7325 (N_7325,N_6557,N_6995);
nor U7326 (N_7326,N_6091,N_6687);
nand U7327 (N_7327,N_6312,N_6078);
nor U7328 (N_7328,N_6610,N_6219);
or U7329 (N_7329,N_6204,N_6021);
nand U7330 (N_7330,N_6471,N_6001);
nor U7331 (N_7331,N_6102,N_6452);
and U7332 (N_7332,N_6241,N_6286);
and U7333 (N_7333,N_6104,N_6830);
nor U7334 (N_7334,N_6100,N_6921);
and U7335 (N_7335,N_6968,N_6777);
nand U7336 (N_7336,N_6740,N_6966);
xnor U7337 (N_7337,N_6089,N_6279);
or U7338 (N_7338,N_6792,N_6576);
nor U7339 (N_7339,N_6831,N_6796);
or U7340 (N_7340,N_6669,N_6144);
or U7341 (N_7341,N_6369,N_6008);
nand U7342 (N_7342,N_6018,N_6298);
or U7343 (N_7343,N_6022,N_6027);
and U7344 (N_7344,N_6433,N_6726);
nor U7345 (N_7345,N_6467,N_6425);
and U7346 (N_7346,N_6268,N_6605);
nand U7347 (N_7347,N_6275,N_6558);
or U7348 (N_7348,N_6567,N_6553);
nor U7349 (N_7349,N_6895,N_6483);
or U7350 (N_7350,N_6391,N_6735);
xnor U7351 (N_7351,N_6861,N_6536);
and U7352 (N_7352,N_6075,N_6972);
nor U7353 (N_7353,N_6668,N_6297);
nand U7354 (N_7354,N_6420,N_6684);
and U7355 (N_7355,N_6914,N_6750);
nand U7356 (N_7356,N_6648,N_6502);
nand U7357 (N_7357,N_6752,N_6969);
and U7358 (N_7358,N_6364,N_6725);
nand U7359 (N_7359,N_6713,N_6043);
and U7360 (N_7360,N_6322,N_6932);
nand U7361 (N_7361,N_6428,N_6737);
and U7362 (N_7362,N_6936,N_6609);
xnor U7363 (N_7363,N_6389,N_6341);
nand U7364 (N_7364,N_6718,N_6138);
xnor U7365 (N_7365,N_6360,N_6975);
or U7366 (N_7366,N_6652,N_6805);
nand U7367 (N_7367,N_6328,N_6056);
and U7368 (N_7368,N_6071,N_6403);
nand U7369 (N_7369,N_6705,N_6246);
and U7370 (N_7370,N_6431,N_6948);
xnor U7371 (N_7371,N_6273,N_6545);
or U7372 (N_7372,N_6042,N_6523);
xor U7373 (N_7373,N_6535,N_6739);
nand U7374 (N_7374,N_6173,N_6997);
nand U7375 (N_7375,N_6367,N_6459);
nor U7376 (N_7376,N_6509,N_6301);
or U7377 (N_7377,N_6786,N_6407);
and U7378 (N_7378,N_6751,N_6882);
nand U7379 (N_7379,N_6550,N_6527);
and U7380 (N_7380,N_6414,N_6209);
nor U7381 (N_7381,N_6155,N_6984);
nor U7382 (N_7382,N_6766,N_6349);
or U7383 (N_7383,N_6477,N_6410);
nand U7384 (N_7384,N_6088,N_6366);
nor U7385 (N_7385,N_6357,N_6240);
or U7386 (N_7386,N_6224,N_6560);
nand U7387 (N_7387,N_6782,N_6949);
nor U7388 (N_7388,N_6470,N_6342);
nand U7389 (N_7389,N_6163,N_6829);
or U7390 (N_7390,N_6588,N_6040);
and U7391 (N_7391,N_6282,N_6828);
nand U7392 (N_7392,N_6036,N_6541);
and U7393 (N_7393,N_6793,N_6764);
nand U7394 (N_7394,N_6570,N_6964);
nor U7395 (N_7395,N_6979,N_6699);
or U7396 (N_7396,N_6686,N_6683);
nand U7397 (N_7397,N_6084,N_6631);
and U7398 (N_7398,N_6698,N_6124);
or U7399 (N_7399,N_6785,N_6624);
or U7400 (N_7400,N_6257,N_6953);
nor U7401 (N_7401,N_6836,N_6741);
or U7402 (N_7402,N_6256,N_6663);
or U7403 (N_7403,N_6592,N_6233);
xnor U7404 (N_7404,N_6189,N_6303);
and U7405 (N_7405,N_6800,N_6494);
or U7406 (N_7406,N_6323,N_6302);
and U7407 (N_7407,N_6889,N_6695);
and U7408 (N_7408,N_6544,N_6879);
or U7409 (N_7409,N_6258,N_6096);
nand U7410 (N_7410,N_6196,N_6732);
nand U7411 (N_7411,N_6851,N_6647);
and U7412 (N_7412,N_6292,N_6562);
nand U7413 (N_7413,N_6150,N_6362);
nor U7414 (N_7414,N_6238,N_6184);
nor U7415 (N_7415,N_6020,N_6507);
and U7416 (N_7416,N_6727,N_6350);
or U7417 (N_7417,N_6370,N_6666);
and U7418 (N_7418,N_6974,N_6947);
or U7419 (N_7419,N_6236,N_6436);
nor U7420 (N_7420,N_6153,N_6943);
or U7421 (N_7421,N_6175,N_6203);
nor U7422 (N_7422,N_6347,N_6872);
and U7423 (N_7423,N_6336,N_6697);
nor U7424 (N_7424,N_6799,N_6927);
and U7425 (N_7425,N_6396,N_6583);
and U7426 (N_7426,N_6073,N_6643);
nand U7427 (N_7427,N_6262,N_6623);
nand U7428 (N_7428,N_6594,N_6287);
nor U7429 (N_7429,N_6335,N_6701);
nand U7430 (N_7430,N_6551,N_6519);
xor U7431 (N_7431,N_6225,N_6532);
and U7432 (N_7432,N_6469,N_6501);
and U7433 (N_7433,N_6237,N_6450);
nand U7434 (N_7434,N_6961,N_6524);
or U7435 (N_7435,N_6374,N_6709);
and U7436 (N_7436,N_6463,N_6047);
nand U7437 (N_7437,N_6028,N_6208);
nor U7438 (N_7438,N_6014,N_6003);
nor U7439 (N_7439,N_6055,N_6598);
or U7440 (N_7440,N_6600,N_6200);
nand U7441 (N_7441,N_6533,N_6016);
and U7442 (N_7442,N_6568,N_6030);
nor U7443 (N_7443,N_6245,N_6846);
and U7444 (N_7444,N_6986,N_6309);
or U7445 (N_7445,N_6060,N_6317);
or U7446 (N_7446,N_6952,N_6432);
nor U7447 (N_7447,N_6170,N_6243);
or U7448 (N_7448,N_6962,N_6413);
or U7449 (N_7449,N_6116,N_6097);
nor U7450 (N_7450,N_6035,N_6179);
nand U7451 (N_7451,N_6933,N_6901);
and U7452 (N_7452,N_6271,N_6215);
or U7453 (N_7453,N_6719,N_6007);
nor U7454 (N_7454,N_6157,N_6130);
nor U7455 (N_7455,N_6866,N_6265);
or U7456 (N_7456,N_6054,N_6207);
xor U7457 (N_7457,N_6569,N_6051);
nor U7458 (N_7458,N_6694,N_6885);
nand U7459 (N_7459,N_6048,N_6728);
nand U7460 (N_7460,N_6094,N_6316);
and U7461 (N_7461,N_6165,N_6662);
and U7462 (N_7462,N_6211,N_6012);
or U7463 (N_7463,N_6067,N_6863);
and U7464 (N_7464,N_6461,N_6318);
xnor U7465 (N_7465,N_6142,N_6714);
nor U7466 (N_7466,N_6418,N_6363);
nor U7467 (N_7467,N_6680,N_6443);
and U7468 (N_7468,N_6515,N_6337);
or U7469 (N_7469,N_6049,N_6361);
or U7470 (N_7470,N_6419,N_6435);
nand U7471 (N_7471,N_6781,N_6466);
or U7472 (N_7472,N_6929,N_6514);
nor U7473 (N_7473,N_6857,N_6864);
and U7474 (N_7474,N_6748,N_6285);
xor U7475 (N_7475,N_6762,N_6776);
xnor U7476 (N_7476,N_6504,N_6151);
nor U7477 (N_7477,N_6039,N_6651);
nor U7478 (N_7478,N_6884,N_6770);
nand U7479 (N_7479,N_6057,N_6860);
nor U7480 (N_7480,N_6315,N_6227);
nand U7481 (N_7481,N_6077,N_6193);
nand U7482 (N_7482,N_6353,N_6299);
xor U7483 (N_7483,N_6082,N_6971);
or U7484 (N_7484,N_6426,N_6444);
and U7485 (N_7485,N_6707,N_6869);
nand U7486 (N_7486,N_6393,N_6571);
or U7487 (N_7487,N_6595,N_6946);
nand U7488 (N_7488,N_6269,N_6497);
nand U7489 (N_7489,N_6114,N_6487);
nor U7490 (N_7490,N_6475,N_6006);
or U7491 (N_7491,N_6521,N_6587);
or U7492 (N_7492,N_6059,N_6434);
nor U7493 (N_7493,N_6024,N_6311);
nand U7494 (N_7494,N_6970,N_6808);
nand U7495 (N_7495,N_6264,N_6276);
and U7496 (N_7496,N_6427,N_6659);
nor U7497 (N_7497,N_6304,N_6099);
and U7498 (N_7498,N_6896,N_6852);
nand U7499 (N_7499,N_6254,N_6358);
nand U7500 (N_7500,N_6829,N_6038);
and U7501 (N_7501,N_6070,N_6173);
and U7502 (N_7502,N_6885,N_6123);
nor U7503 (N_7503,N_6588,N_6913);
or U7504 (N_7504,N_6331,N_6122);
and U7505 (N_7505,N_6377,N_6054);
or U7506 (N_7506,N_6505,N_6826);
or U7507 (N_7507,N_6912,N_6415);
or U7508 (N_7508,N_6370,N_6352);
nor U7509 (N_7509,N_6272,N_6365);
nor U7510 (N_7510,N_6153,N_6194);
nand U7511 (N_7511,N_6270,N_6323);
and U7512 (N_7512,N_6791,N_6970);
xnor U7513 (N_7513,N_6228,N_6399);
and U7514 (N_7514,N_6954,N_6844);
nor U7515 (N_7515,N_6332,N_6138);
nor U7516 (N_7516,N_6549,N_6906);
or U7517 (N_7517,N_6415,N_6391);
nor U7518 (N_7518,N_6738,N_6391);
or U7519 (N_7519,N_6947,N_6216);
and U7520 (N_7520,N_6903,N_6580);
nand U7521 (N_7521,N_6720,N_6756);
and U7522 (N_7522,N_6246,N_6882);
and U7523 (N_7523,N_6866,N_6005);
and U7524 (N_7524,N_6400,N_6201);
nor U7525 (N_7525,N_6336,N_6686);
and U7526 (N_7526,N_6038,N_6781);
nand U7527 (N_7527,N_6664,N_6619);
nand U7528 (N_7528,N_6984,N_6196);
nor U7529 (N_7529,N_6888,N_6764);
nand U7530 (N_7530,N_6116,N_6356);
nor U7531 (N_7531,N_6431,N_6662);
and U7532 (N_7532,N_6439,N_6782);
xnor U7533 (N_7533,N_6788,N_6626);
nor U7534 (N_7534,N_6491,N_6055);
nand U7535 (N_7535,N_6568,N_6582);
or U7536 (N_7536,N_6007,N_6733);
or U7537 (N_7537,N_6698,N_6936);
nor U7538 (N_7538,N_6237,N_6874);
nand U7539 (N_7539,N_6735,N_6063);
nand U7540 (N_7540,N_6183,N_6904);
or U7541 (N_7541,N_6161,N_6067);
nand U7542 (N_7542,N_6089,N_6830);
or U7543 (N_7543,N_6531,N_6725);
and U7544 (N_7544,N_6115,N_6944);
nor U7545 (N_7545,N_6308,N_6402);
and U7546 (N_7546,N_6809,N_6935);
and U7547 (N_7547,N_6198,N_6023);
and U7548 (N_7548,N_6966,N_6394);
xor U7549 (N_7549,N_6229,N_6038);
and U7550 (N_7550,N_6951,N_6880);
and U7551 (N_7551,N_6408,N_6230);
and U7552 (N_7552,N_6059,N_6105);
and U7553 (N_7553,N_6695,N_6427);
and U7554 (N_7554,N_6943,N_6279);
or U7555 (N_7555,N_6188,N_6899);
nand U7556 (N_7556,N_6728,N_6191);
xnor U7557 (N_7557,N_6931,N_6520);
or U7558 (N_7558,N_6159,N_6710);
nand U7559 (N_7559,N_6073,N_6959);
nor U7560 (N_7560,N_6696,N_6865);
or U7561 (N_7561,N_6960,N_6612);
nand U7562 (N_7562,N_6428,N_6270);
nand U7563 (N_7563,N_6808,N_6737);
nand U7564 (N_7564,N_6414,N_6742);
nand U7565 (N_7565,N_6992,N_6988);
or U7566 (N_7566,N_6523,N_6597);
nor U7567 (N_7567,N_6581,N_6896);
or U7568 (N_7568,N_6139,N_6693);
and U7569 (N_7569,N_6008,N_6685);
or U7570 (N_7570,N_6941,N_6682);
nand U7571 (N_7571,N_6564,N_6701);
and U7572 (N_7572,N_6725,N_6453);
nor U7573 (N_7573,N_6098,N_6725);
nor U7574 (N_7574,N_6745,N_6345);
nor U7575 (N_7575,N_6144,N_6818);
or U7576 (N_7576,N_6769,N_6337);
nor U7577 (N_7577,N_6889,N_6984);
or U7578 (N_7578,N_6284,N_6540);
xnor U7579 (N_7579,N_6116,N_6200);
xor U7580 (N_7580,N_6347,N_6514);
xnor U7581 (N_7581,N_6057,N_6759);
and U7582 (N_7582,N_6436,N_6258);
nand U7583 (N_7583,N_6806,N_6847);
nand U7584 (N_7584,N_6726,N_6963);
and U7585 (N_7585,N_6504,N_6212);
nand U7586 (N_7586,N_6853,N_6405);
nand U7587 (N_7587,N_6790,N_6173);
nand U7588 (N_7588,N_6360,N_6279);
nor U7589 (N_7589,N_6114,N_6651);
nand U7590 (N_7590,N_6202,N_6708);
or U7591 (N_7591,N_6312,N_6765);
nand U7592 (N_7592,N_6159,N_6297);
nor U7593 (N_7593,N_6395,N_6789);
and U7594 (N_7594,N_6257,N_6864);
and U7595 (N_7595,N_6072,N_6759);
nor U7596 (N_7596,N_6225,N_6214);
nor U7597 (N_7597,N_6662,N_6617);
or U7598 (N_7598,N_6935,N_6468);
and U7599 (N_7599,N_6893,N_6279);
nand U7600 (N_7600,N_6827,N_6059);
xnor U7601 (N_7601,N_6563,N_6882);
xnor U7602 (N_7602,N_6430,N_6339);
and U7603 (N_7603,N_6012,N_6468);
nand U7604 (N_7604,N_6713,N_6926);
or U7605 (N_7605,N_6341,N_6648);
nor U7606 (N_7606,N_6659,N_6039);
nand U7607 (N_7607,N_6125,N_6458);
nand U7608 (N_7608,N_6016,N_6775);
nand U7609 (N_7609,N_6134,N_6733);
and U7610 (N_7610,N_6045,N_6747);
or U7611 (N_7611,N_6496,N_6100);
nand U7612 (N_7612,N_6458,N_6342);
and U7613 (N_7613,N_6934,N_6746);
or U7614 (N_7614,N_6389,N_6133);
xor U7615 (N_7615,N_6607,N_6513);
and U7616 (N_7616,N_6367,N_6066);
xor U7617 (N_7617,N_6532,N_6510);
or U7618 (N_7618,N_6107,N_6256);
xor U7619 (N_7619,N_6241,N_6221);
nand U7620 (N_7620,N_6759,N_6412);
xnor U7621 (N_7621,N_6191,N_6408);
nor U7622 (N_7622,N_6602,N_6594);
and U7623 (N_7623,N_6570,N_6103);
nand U7624 (N_7624,N_6025,N_6267);
nand U7625 (N_7625,N_6511,N_6764);
or U7626 (N_7626,N_6878,N_6213);
nor U7627 (N_7627,N_6337,N_6073);
and U7628 (N_7628,N_6770,N_6344);
nor U7629 (N_7629,N_6015,N_6506);
nand U7630 (N_7630,N_6373,N_6647);
and U7631 (N_7631,N_6206,N_6322);
xnor U7632 (N_7632,N_6977,N_6405);
or U7633 (N_7633,N_6456,N_6430);
and U7634 (N_7634,N_6962,N_6839);
or U7635 (N_7635,N_6135,N_6711);
nor U7636 (N_7636,N_6560,N_6952);
and U7637 (N_7637,N_6349,N_6549);
or U7638 (N_7638,N_6153,N_6373);
or U7639 (N_7639,N_6393,N_6118);
nand U7640 (N_7640,N_6667,N_6960);
or U7641 (N_7641,N_6478,N_6046);
nor U7642 (N_7642,N_6535,N_6318);
nor U7643 (N_7643,N_6710,N_6431);
and U7644 (N_7644,N_6511,N_6839);
and U7645 (N_7645,N_6509,N_6046);
nor U7646 (N_7646,N_6742,N_6640);
xor U7647 (N_7647,N_6087,N_6383);
nand U7648 (N_7648,N_6757,N_6293);
or U7649 (N_7649,N_6406,N_6299);
and U7650 (N_7650,N_6455,N_6710);
and U7651 (N_7651,N_6265,N_6991);
and U7652 (N_7652,N_6839,N_6542);
and U7653 (N_7653,N_6881,N_6073);
nand U7654 (N_7654,N_6013,N_6170);
xnor U7655 (N_7655,N_6870,N_6717);
or U7656 (N_7656,N_6732,N_6942);
nand U7657 (N_7657,N_6017,N_6050);
or U7658 (N_7658,N_6498,N_6562);
or U7659 (N_7659,N_6936,N_6920);
and U7660 (N_7660,N_6213,N_6234);
and U7661 (N_7661,N_6280,N_6202);
or U7662 (N_7662,N_6925,N_6369);
or U7663 (N_7663,N_6190,N_6957);
xnor U7664 (N_7664,N_6365,N_6754);
nor U7665 (N_7665,N_6731,N_6801);
and U7666 (N_7666,N_6241,N_6507);
nor U7667 (N_7667,N_6202,N_6189);
nand U7668 (N_7668,N_6930,N_6258);
nor U7669 (N_7669,N_6137,N_6994);
and U7670 (N_7670,N_6790,N_6585);
nor U7671 (N_7671,N_6552,N_6456);
and U7672 (N_7672,N_6888,N_6896);
nand U7673 (N_7673,N_6558,N_6761);
or U7674 (N_7674,N_6173,N_6682);
or U7675 (N_7675,N_6326,N_6441);
xor U7676 (N_7676,N_6505,N_6941);
or U7677 (N_7677,N_6361,N_6372);
nor U7678 (N_7678,N_6487,N_6922);
xnor U7679 (N_7679,N_6359,N_6403);
and U7680 (N_7680,N_6340,N_6219);
nand U7681 (N_7681,N_6206,N_6220);
xnor U7682 (N_7682,N_6428,N_6177);
and U7683 (N_7683,N_6800,N_6400);
or U7684 (N_7684,N_6199,N_6814);
and U7685 (N_7685,N_6060,N_6041);
nand U7686 (N_7686,N_6905,N_6389);
or U7687 (N_7687,N_6178,N_6164);
nand U7688 (N_7688,N_6720,N_6694);
nor U7689 (N_7689,N_6026,N_6504);
nor U7690 (N_7690,N_6714,N_6034);
xnor U7691 (N_7691,N_6652,N_6263);
nand U7692 (N_7692,N_6377,N_6986);
nor U7693 (N_7693,N_6626,N_6080);
and U7694 (N_7694,N_6329,N_6215);
and U7695 (N_7695,N_6344,N_6964);
nand U7696 (N_7696,N_6153,N_6713);
and U7697 (N_7697,N_6255,N_6509);
and U7698 (N_7698,N_6842,N_6912);
or U7699 (N_7699,N_6927,N_6187);
and U7700 (N_7700,N_6184,N_6329);
nand U7701 (N_7701,N_6334,N_6854);
or U7702 (N_7702,N_6271,N_6541);
xor U7703 (N_7703,N_6176,N_6173);
and U7704 (N_7704,N_6633,N_6762);
or U7705 (N_7705,N_6203,N_6570);
nand U7706 (N_7706,N_6699,N_6642);
and U7707 (N_7707,N_6416,N_6901);
or U7708 (N_7708,N_6911,N_6753);
or U7709 (N_7709,N_6447,N_6690);
nor U7710 (N_7710,N_6702,N_6901);
nor U7711 (N_7711,N_6439,N_6078);
xnor U7712 (N_7712,N_6693,N_6041);
nor U7713 (N_7713,N_6535,N_6183);
or U7714 (N_7714,N_6221,N_6568);
xor U7715 (N_7715,N_6559,N_6787);
nor U7716 (N_7716,N_6236,N_6835);
nor U7717 (N_7717,N_6744,N_6485);
and U7718 (N_7718,N_6498,N_6478);
nor U7719 (N_7719,N_6703,N_6759);
or U7720 (N_7720,N_6015,N_6293);
and U7721 (N_7721,N_6316,N_6235);
nor U7722 (N_7722,N_6540,N_6024);
and U7723 (N_7723,N_6398,N_6530);
nand U7724 (N_7724,N_6301,N_6112);
and U7725 (N_7725,N_6241,N_6121);
nor U7726 (N_7726,N_6253,N_6303);
nand U7727 (N_7727,N_6949,N_6757);
or U7728 (N_7728,N_6609,N_6342);
nand U7729 (N_7729,N_6268,N_6054);
nand U7730 (N_7730,N_6819,N_6546);
nand U7731 (N_7731,N_6836,N_6977);
xor U7732 (N_7732,N_6277,N_6726);
or U7733 (N_7733,N_6106,N_6832);
or U7734 (N_7734,N_6201,N_6304);
and U7735 (N_7735,N_6043,N_6018);
and U7736 (N_7736,N_6654,N_6769);
nor U7737 (N_7737,N_6723,N_6775);
and U7738 (N_7738,N_6620,N_6590);
and U7739 (N_7739,N_6794,N_6250);
nor U7740 (N_7740,N_6244,N_6170);
or U7741 (N_7741,N_6635,N_6464);
or U7742 (N_7742,N_6729,N_6198);
nor U7743 (N_7743,N_6867,N_6339);
and U7744 (N_7744,N_6231,N_6145);
nor U7745 (N_7745,N_6311,N_6507);
nor U7746 (N_7746,N_6811,N_6439);
or U7747 (N_7747,N_6926,N_6133);
or U7748 (N_7748,N_6055,N_6716);
nand U7749 (N_7749,N_6553,N_6043);
and U7750 (N_7750,N_6577,N_6904);
nor U7751 (N_7751,N_6531,N_6987);
xor U7752 (N_7752,N_6930,N_6705);
and U7753 (N_7753,N_6906,N_6440);
xor U7754 (N_7754,N_6170,N_6192);
or U7755 (N_7755,N_6448,N_6656);
nor U7756 (N_7756,N_6061,N_6746);
nand U7757 (N_7757,N_6817,N_6649);
or U7758 (N_7758,N_6969,N_6799);
and U7759 (N_7759,N_6089,N_6970);
and U7760 (N_7760,N_6804,N_6039);
nor U7761 (N_7761,N_6202,N_6909);
nor U7762 (N_7762,N_6223,N_6691);
nand U7763 (N_7763,N_6098,N_6606);
or U7764 (N_7764,N_6883,N_6252);
or U7765 (N_7765,N_6991,N_6724);
and U7766 (N_7766,N_6008,N_6034);
nor U7767 (N_7767,N_6308,N_6222);
nand U7768 (N_7768,N_6775,N_6357);
and U7769 (N_7769,N_6128,N_6067);
nand U7770 (N_7770,N_6560,N_6015);
and U7771 (N_7771,N_6914,N_6215);
or U7772 (N_7772,N_6163,N_6350);
nand U7773 (N_7773,N_6729,N_6853);
nand U7774 (N_7774,N_6363,N_6227);
or U7775 (N_7775,N_6784,N_6454);
and U7776 (N_7776,N_6640,N_6581);
or U7777 (N_7777,N_6097,N_6458);
or U7778 (N_7778,N_6494,N_6425);
nor U7779 (N_7779,N_6743,N_6302);
and U7780 (N_7780,N_6727,N_6618);
or U7781 (N_7781,N_6593,N_6007);
nor U7782 (N_7782,N_6702,N_6590);
nand U7783 (N_7783,N_6388,N_6453);
nor U7784 (N_7784,N_6730,N_6567);
and U7785 (N_7785,N_6211,N_6161);
nor U7786 (N_7786,N_6915,N_6638);
xnor U7787 (N_7787,N_6504,N_6448);
or U7788 (N_7788,N_6081,N_6757);
or U7789 (N_7789,N_6810,N_6639);
or U7790 (N_7790,N_6850,N_6607);
and U7791 (N_7791,N_6879,N_6802);
and U7792 (N_7792,N_6331,N_6862);
nor U7793 (N_7793,N_6622,N_6219);
nand U7794 (N_7794,N_6776,N_6750);
and U7795 (N_7795,N_6427,N_6472);
or U7796 (N_7796,N_6565,N_6649);
xnor U7797 (N_7797,N_6798,N_6645);
or U7798 (N_7798,N_6776,N_6001);
xnor U7799 (N_7799,N_6676,N_6171);
or U7800 (N_7800,N_6983,N_6240);
nand U7801 (N_7801,N_6232,N_6664);
nand U7802 (N_7802,N_6928,N_6044);
nand U7803 (N_7803,N_6704,N_6409);
and U7804 (N_7804,N_6034,N_6208);
nor U7805 (N_7805,N_6793,N_6356);
or U7806 (N_7806,N_6256,N_6950);
or U7807 (N_7807,N_6694,N_6355);
nand U7808 (N_7808,N_6920,N_6287);
or U7809 (N_7809,N_6482,N_6687);
and U7810 (N_7810,N_6053,N_6250);
nand U7811 (N_7811,N_6580,N_6048);
and U7812 (N_7812,N_6161,N_6343);
nor U7813 (N_7813,N_6813,N_6433);
nor U7814 (N_7814,N_6377,N_6308);
or U7815 (N_7815,N_6954,N_6753);
or U7816 (N_7816,N_6744,N_6531);
and U7817 (N_7817,N_6224,N_6948);
nand U7818 (N_7818,N_6711,N_6124);
and U7819 (N_7819,N_6234,N_6982);
nand U7820 (N_7820,N_6454,N_6624);
and U7821 (N_7821,N_6627,N_6025);
nor U7822 (N_7822,N_6060,N_6254);
nand U7823 (N_7823,N_6089,N_6292);
nor U7824 (N_7824,N_6465,N_6163);
nor U7825 (N_7825,N_6216,N_6404);
or U7826 (N_7826,N_6055,N_6337);
or U7827 (N_7827,N_6770,N_6308);
or U7828 (N_7828,N_6904,N_6436);
and U7829 (N_7829,N_6716,N_6096);
nor U7830 (N_7830,N_6671,N_6341);
and U7831 (N_7831,N_6047,N_6824);
nor U7832 (N_7832,N_6428,N_6695);
and U7833 (N_7833,N_6226,N_6437);
or U7834 (N_7834,N_6882,N_6561);
nand U7835 (N_7835,N_6805,N_6022);
nor U7836 (N_7836,N_6539,N_6323);
or U7837 (N_7837,N_6401,N_6988);
nand U7838 (N_7838,N_6635,N_6741);
xor U7839 (N_7839,N_6309,N_6809);
nand U7840 (N_7840,N_6346,N_6881);
nand U7841 (N_7841,N_6955,N_6171);
nand U7842 (N_7842,N_6575,N_6067);
nor U7843 (N_7843,N_6446,N_6238);
and U7844 (N_7844,N_6729,N_6755);
nor U7845 (N_7845,N_6962,N_6693);
nand U7846 (N_7846,N_6519,N_6082);
nor U7847 (N_7847,N_6727,N_6490);
xnor U7848 (N_7848,N_6908,N_6360);
xnor U7849 (N_7849,N_6393,N_6824);
or U7850 (N_7850,N_6430,N_6057);
nand U7851 (N_7851,N_6540,N_6378);
nor U7852 (N_7852,N_6297,N_6541);
nand U7853 (N_7853,N_6080,N_6414);
nor U7854 (N_7854,N_6439,N_6876);
or U7855 (N_7855,N_6709,N_6237);
xor U7856 (N_7856,N_6493,N_6530);
or U7857 (N_7857,N_6392,N_6456);
xor U7858 (N_7858,N_6322,N_6602);
and U7859 (N_7859,N_6243,N_6336);
nor U7860 (N_7860,N_6464,N_6476);
nor U7861 (N_7861,N_6464,N_6798);
and U7862 (N_7862,N_6638,N_6757);
or U7863 (N_7863,N_6713,N_6335);
or U7864 (N_7864,N_6091,N_6907);
nand U7865 (N_7865,N_6423,N_6816);
xnor U7866 (N_7866,N_6812,N_6717);
xnor U7867 (N_7867,N_6117,N_6143);
and U7868 (N_7868,N_6533,N_6183);
or U7869 (N_7869,N_6474,N_6239);
xor U7870 (N_7870,N_6276,N_6323);
or U7871 (N_7871,N_6603,N_6563);
or U7872 (N_7872,N_6409,N_6812);
and U7873 (N_7873,N_6420,N_6161);
nor U7874 (N_7874,N_6280,N_6374);
nand U7875 (N_7875,N_6191,N_6164);
xnor U7876 (N_7876,N_6154,N_6014);
or U7877 (N_7877,N_6556,N_6168);
nand U7878 (N_7878,N_6334,N_6746);
or U7879 (N_7879,N_6265,N_6877);
or U7880 (N_7880,N_6872,N_6032);
xnor U7881 (N_7881,N_6647,N_6805);
and U7882 (N_7882,N_6598,N_6154);
nor U7883 (N_7883,N_6402,N_6519);
nand U7884 (N_7884,N_6312,N_6472);
xor U7885 (N_7885,N_6430,N_6782);
xnor U7886 (N_7886,N_6629,N_6975);
or U7887 (N_7887,N_6168,N_6051);
and U7888 (N_7888,N_6245,N_6502);
nor U7889 (N_7889,N_6806,N_6097);
nor U7890 (N_7890,N_6911,N_6933);
and U7891 (N_7891,N_6855,N_6591);
or U7892 (N_7892,N_6575,N_6983);
nor U7893 (N_7893,N_6218,N_6145);
nand U7894 (N_7894,N_6132,N_6479);
or U7895 (N_7895,N_6903,N_6675);
and U7896 (N_7896,N_6297,N_6822);
nor U7897 (N_7897,N_6963,N_6020);
nor U7898 (N_7898,N_6024,N_6636);
or U7899 (N_7899,N_6667,N_6742);
and U7900 (N_7900,N_6268,N_6690);
and U7901 (N_7901,N_6773,N_6146);
or U7902 (N_7902,N_6983,N_6559);
nor U7903 (N_7903,N_6385,N_6635);
nor U7904 (N_7904,N_6509,N_6488);
or U7905 (N_7905,N_6775,N_6672);
or U7906 (N_7906,N_6587,N_6394);
nor U7907 (N_7907,N_6338,N_6410);
and U7908 (N_7908,N_6949,N_6589);
nor U7909 (N_7909,N_6130,N_6337);
nand U7910 (N_7910,N_6449,N_6025);
nand U7911 (N_7911,N_6710,N_6099);
nor U7912 (N_7912,N_6347,N_6234);
nor U7913 (N_7913,N_6074,N_6859);
nor U7914 (N_7914,N_6439,N_6933);
or U7915 (N_7915,N_6351,N_6185);
and U7916 (N_7916,N_6152,N_6947);
nor U7917 (N_7917,N_6491,N_6309);
and U7918 (N_7918,N_6701,N_6681);
xnor U7919 (N_7919,N_6818,N_6237);
or U7920 (N_7920,N_6641,N_6385);
nand U7921 (N_7921,N_6035,N_6725);
nor U7922 (N_7922,N_6965,N_6736);
nor U7923 (N_7923,N_6068,N_6244);
and U7924 (N_7924,N_6034,N_6676);
nor U7925 (N_7925,N_6087,N_6450);
nor U7926 (N_7926,N_6136,N_6144);
nand U7927 (N_7927,N_6145,N_6609);
or U7928 (N_7928,N_6812,N_6179);
and U7929 (N_7929,N_6387,N_6112);
or U7930 (N_7930,N_6467,N_6303);
and U7931 (N_7931,N_6770,N_6304);
nand U7932 (N_7932,N_6837,N_6496);
nand U7933 (N_7933,N_6219,N_6859);
and U7934 (N_7934,N_6212,N_6974);
or U7935 (N_7935,N_6059,N_6048);
xnor U7936 (N_7936,N_6866,N_6205);
and U7937 (N_7937,N_6968,N_6585);
and U7938 (N_7938,N_6920,N_6103);
or U7939 (N_7939,N_6125,N_6081);
nor U7940 (N_7940,N_6260,N_6918);
nor U7941 (N_7941,N_6278,N_6994);
or U7942 (N_7942,N_6589,N_6567);
and U7943 (N_7943,N_6753,N_6316);
nor U7944 (N_7944,N_6314,N_6230);
or U7945 (N_7945,N_6117,N_6580);
nand U7946 (N_7946,N_6486,N_6725);
and U7947 (N_7947,N_6963,N_6795);
xor U7948 (N_7948,N_6514,N_6906);
nor U7949 (N_7949,N_6824,N_6363);
nand U7950 (N_7950,N_6444,N_6784);
nand U7951 (N_7951,N_6046,N_6074);
and U7952 (N_7952,N_6300,N_6510);
nor U7953 (N_7953,N_6757,N_6138);
nor U7954 (N_7954,N_6561,N_6025);
and U7955 (N_7955,N_6424,N_6819);
nand U7956 (N_7956,N_6956,N_6534);
and U7957 (N_7957,N_6757,N_6749);
or U7958 (N_7958,N_6637,N_6893);
nor U7959 (N_7959,N_6277,N_6835);
nor U7960 (N_7960,N_6095,N_6421);
nor U7961 (N_7961,N_6651,N_6902);
nand U7962 (N_7962,N_6441,N_6794);
and U7963 (N_7963,N_6283,N_6186);
and U7964 (N_7964,N_6119,N_6019);
and U7965 (N_7965,N_6176,N_6525);
nand U7966 (N_7966,N_6608,N_6416);
and U7967 (N_7967,N_6846,N_6886);
or U7968 (N_7968,N_6645,N_6747);
or U7969 (N_7969,N_6642,N_6125);
and U7970 (N_7970,N_6555,N_6687);
and U7971 (N_7971,N_6534,N_6592);
nor U7972 (N_7972,N_6662,N_6752);
or U7973 (N_7973,N_6496,N_6492);
nor U7974 (N_7974,N_6789,N_6017);
nor U7975 (N_7975,N_6504,N_6377);
xnor U7976 (N_7976,N_6638,N_6504);
xor U7977 (N_7977,N_6192,N_6753);
nand U7978 (N_7978,N_6353,N_6947);
nand U7979 (N_7979,N_6417,N_6777);
and U7980 (N_7980,N_6682,N_6790);
or U7981 (N_7981,N_6882,N_6525);
nand U7982 (N_7982,N_6264,N_6355);
and U7983 (N_7983,N_6126,N_6905);
xor U7984 (N_7984,N_6585,N_6181);
xnor U7985 (N_7985,N_6559,N_6399);
nand U7986 (N_7986,N_6400,N_6766);
nand U7987 (N_7987,N_6545,N_6694);
and U7988 (N_7988,N_6132,N_6465);
and U7989 (N_7989,N_6148,N_6933);
nor U7990 (N_7990,N_6023,N_6572);
and U7991 (N_7991,N_6324,N_6433);
xnor U7992 (N_7992,N_6322,N_6492);
or U7993 (N_7993,N_6064,N_6735);
nor U7994 (N_7994,N_6240,N_6244);
or U7995 (N_7995,N_6595,N_6747);
nor U7996 (N_7996,N_6068,N_6713);
and U7997 (N_7997,N_6220,N_6338);
nand U7998 (N_7998,N_6099,N_6028);
or U7999 (N_7999,N_6574,N_6696);
xnor U8000 (N_8000,N_7732,N_7394);
nand U8001 (N_8001,N_7148,N_7576);
xor U8002 (N_8002,N_7848,N_7475);
nand U8003 (N_8003,N_7736,N_7866);
nor U8004 (N_8004,N_7833,N_7388);
nor U8005 (N_8005,N_7776,N_7215);
nor U8006 (N_8006,N_7991,N_7610);
nand U8007 (N_8007,N_7362,N_7446);
and U8008 (N_8008,N_7862,N_7285);
and U8009 (N_8009,N_7307,N_7262);
and U8010 (N_8010,N_7643,N_7951);
and U8011 (N_8011,N_7675,N_7419);
or U8012 (N_8012,N_7065,N_7810);
nand U8013 (N_8013,N_7832,N_7664);
nand U8014 (N_8014,N_7024,N_7133);
nor U8015 (N_8015,N_7159,N_7054);
and U8016 (N_8016,N_7391,N_7870);
nor U8017 (N_8017,N_7277,N_7886);
xnor U8018 (N_8018,N_7502,N_7924);
and U8019 (N_8019,N_7642,N_7246);
and U8020 (N_8020,N_7235,N_7968);
nor U8021 (N_8021,N_7009,N_7249);
nor U8022 (N_8022,N_7291,N_7772);
nand U8023 (N_8023,N_7724,N_7858);
nand U8024 (N_8024,N_7267,N_7532);
and U8025 (N_8025,N_7960,N_7428);
nand U8026 (N_8026,N_7914,N_7770);
and U8027 (N_8027,N_7925,N_7969);
nor U8028 (N_8028,N_7090,N_7700);
nor U8029 (N_8029,N_7197,N_7136);
nand U8030 (N_8030,N_7091,N_7041);
or U8031 (N_8031,N_7898,N_7385);
and U8032 (N_8032,N_7907,N_7341);
and U8033 (N_8033,N_7158,N_7651);
nand U8034 (N_8034,N_7245,N_7494);
and U8035 (N_8035,N_7224,N_7276);
nor U8036 (N_8036,N_7712,N_7800);
xor U8037 (N_8037,N_7515,N_7392);
nor U8038 (N_8038,N_7230,N_7613);
nand U8039 (N_8039,N_7584,N_7941);
nor U8040 (N_8040,N_7587,N_7533);
nor U8041 (N_8041,N_7284,N_7372);
and U8042 (N_8042,N_7873,N_7134);
nor U8043 (N_8043,N_7817,N_7104);
or U8044 (N_8044,N_7145,N_7513);
or U8045 (N_8045,N_7489,N_7176);
and U8046 (N_8046,N_7186,N_7835);
xnor U8047 (N_8047,N_7420,N_7320);
nor U8048 (N_8048,N_7668,N_7624);
and U8049 (N_8049,N_7363,N_7043);
nand U8050 (N_8050,N_7930,N_7807);
or U8051 (N_8051,N_7495,N_7926);
nand U8052 (N_8052,N_7250,N_7892);
nand U8053 (N_8053,N_7872,N_7342);
and U8054 (N_8054,N_7824,N_7188);
nor U8055 (N_8055,N_7260,N_7693);
nand U8056 (N_8056,N_7863,N_7756);
nand U8057 (N_8057,N_7726,N_7424);
and U8058 (N_8058,N_7283,N_7354);
nor U8059 (N_8059,N_7324,N_7961);
and U8060 (N_8060,N_7711,N_7366);
or U8061 (N_8061,N_7801,N_7149);
and U8062 (N_8062,N_7375,N_7384);
nor U8063 (N_8063,N_7055,N_7326);
nor U8064 (N_8064,N_7378,N_7931);
or U8065 (N_8065,N_7628,N_7938);
or U8066 (N_8066,N_7713,N_7293);
or U8067 (N_8067,N_7615,N_7070);
and U8068 (N_8068,N_7803,N_7808);
or U8069 (N_8069,N_7258,N_7737);
and U8070 (N_8070,N_7414,N_7356);
or U8071 (N_8071,N_7944,N_7020);
nor U8072 (N_8072,N_7316,N_7539);
and U8073 (N_8073,N_7202,N_7791);
nand U8074 (N_8074,N_7237,N_7074);
and U8075 (N_8075,N_7228,N_7820);
or U8076 (N_8076,N_7590,N_7006);
or U8077 (N_8077,N_7787,N_7595);
and U8078 (N_8078,N_7196,N_7303);
nand U8079 (N_8079,N_7256,N_7233);
and U8080 (N_8080,N_7195,N_7698);
and U8081 (N_8081,N_7146,N_7184);
nand U8082 (N_8082,N_7002,N_7995);
or U8083 (N_8083,N_7085,N_7236);
or U8084 (N_8084,N_7340,N_7058);
nand U8085 (N_8085,N_7525,N_7554);
nor U8086 (N_8086,N_7157,N_7095);
or U8087 (N_8087,N_7973,N_7234);
xor U8088 (N_8088,N_7804,N_7517);
or U8089 (N_8089,N_7868,N_7555);
or U8090 (N_8090,N_7600,N_7903);
nand U8091 (N_8091,N_7888,N_7871);
and U8092 (N_8092,N_7653,N_7945);
or U8093 (N_8093,N_7131,N_7809);
xnor U8094 (N_8094,N_7435,N_7198);
or U8095 (N_8095,N_7534,N_7257);
nor U8096 (N_8096,N_7942,N_7305);
or U8097 (N_8097,N_7448,N_7847);
and U8098 (N_8098,N_7825,N_7383);
nand U8099 (N_8099,N_7415,N_7916);
xor U8100 (N_8100,N_7500,N_7255);
nor U8101 (N_8101,N_7141,N_7730);
or U8102 (N_8102,N_7781,N_7727);
or U8103 (N_8103,N_7143,N_7223);
nor U8104 (N_8104,N_7193,N_7789);
nor U8105 (N_8105,N_7814,N_7981);
and U8106 (N_8106,N_7492,N_7985);
nor U8107 (N_8107,N_7472,N_7597);
nand U8108 (N_8108,N_7395,N_7618);
or U8109 (N_8109,N_7497,N_7519);
nor U8110 (N_8110,N_7718,N_7839);
or U8111 (N_8111,N_7469,N_7231);
nor U8112 (N_8112,N_7763,N_7268);
or U8113 (N_8113,N_7336,N_7221);
nand U8114 (N_8114,N_7204,N_7742);
or U8115 (N_8115,N_7792,N_7701);
nor U8116 (N_8116,N_7880,N_7550);
nor U8117 (N_8117,N_7069,N_7488);
and U8118 (N_8118,N_7765,N_7456);
xnor U8119 (N_8119,N_7666,N_7442);
and U8120 (N_8120,N_7607,N_7844);
xnor U8121 (N_8121,N_7449,N_7752);
or U8122 (N_8122,N_7251,N_7072);
nand U8123 (N_8123,N_7986,N_7879);
or U8124 (N_8124,N_7567,N_7764);
or U8125 (N_8125,N_7130,N_7429);
nor U8126 (N_8126,N_7466,N_7487);
nor U8127 (N_8127,N_7688,N_7746);
nor U8128 (N_8128,N_7563,N_7694);
and U8129 (N_8129,N_7658,N_7843);
xnor U8130 (N_8130,N_7178,N_7958);
and U8131 (N_8131,N_7891,N_7016);
and U8132 (N_8132,N_7030,N_7670);
nor U8133 (N_8133,N_7450,N_7845);
nand U8134 (N_8134,N_7473,N_7387);
or U8135 (N_8135,N_7767,N_7505);
nand U8136 (N_8136,N_7908,N_7549);
nand U8137 (N_8137,N_7300,N_7779);
and U8138 (N_8138,N_7214,N_7686);
xor U8139 (N_8139,N_7913,N_7678);
nand U8140 (N_8140,N_7876,N_7691);
or U8141 (N_8141,N_7846,N_7882);
nand U8142 (N_8142,N_7496,N_7725);
xor U8143 (N_8143,N_7747,N_7963);
xor U8144 (N_8144,N_7373,N_7103);
xnor U8145 (N_8145,N_7122,N_7327);
and U8146 (N_8146,N_7606,N_7582);
and U8147 (N_8147,N_7482,N_7167);
or U8148 (N_8148,N_7116,N_7194);
nor U8149 (N_8149,N_7271,N_7912);
nand U8150 (N_8150,N_7865,N_7875);
nand U8151 (N_8151,N_7967,N_7071);
and U8152 (N_8152,N_7463,N_7950);
xnor U8153 (N_8153,N_7138,N_7954);
and U8154 (N_8154,N_7162,N_7884);
nor U8155 (N_8155,N_7783,N_7971);
nor U8156 (N_8156,N_7589,N_7042);
or U8157 (N_8157,N_7001,N_7035);
and U8158 (N_8158,N_7286,N_7546);
or U8159 (N_8159,N_7522,N_7743);
nor U8160 (N_8160,N_7761,N_7634);
nor U8161 (N_8161,N_7766,N_7979);
or U8162 (N_8162,N_7485,N_7717);
nor U8163 (N_8163,N_7460,N_7626);
and U8164 (N_8164,N_7859,N_7636);
or U8165 (N_8165,N_7272,N_7218);
xor U8166 (N_8166,N_7568,N_7076);
xor U8167 (N_8167,N_7470,N_7282);
or U8168 (N_8168,N_7706,N_7937);
and U8169 (N_8169,N_7335,N_7580);
or U8170 (N_8170,N_7721,N_7079);
xnor U8171 (N_8171,N_7412,N_7436);
or U8172 (N_8172,N_7003,N_7240);
nand U8173 (N_8173,N_7239,N_7569);
nor U8174 (N_8174,N_7855,N_7955);
nand U8175 (N_8175,N_7050,N_7380);
xnor U8176 (N_8176,N_7238,N_7023);
nand U8177 (N_8177,N_7592,N_7685);
nor U8178 (N_8178,N_7083,N_7894);
and U8179 (N_8179,N_7113,N_7199);
nor U8180 (N_8180,N_7577,N_7683);
xor U8181 (N_8181,N_7611,N_7667);
nor U8182 (N_8182,N_7975,N_7451);
and U8183 (N_8183,N_7118,N_7308);
and U8184 (N_8184,N_7206,N_7353);
and U8185 (N_8185,N_7080,N_7357);
and U8186 (N_8186,N_7132,N_7108);
nor U8187 (N_8187,N_7096,N_7337);
nor U8188 (N_8188,N_7768,N_7889);
nand U8189 (N_8189,N_7039,N_7571);
nor U8190 (N_8190,N_7749,N_7536);
nand U8191 (N_8191,N_7989,N_7754);
xnor U8192 (N_8192,N_7465,N_7430);
nand U8193 (N_8193,N_7144,N_7547);
nand U8194 (N_8194,N_7773,N_7521);
xor U8195 (N_8195,N_7397,N_7213);
nand U8196 (N_8196,N_7757,N_7129);
xor U8197 (N_8197,N_7759,N_7821);
or U8198 (N_8198,N_7735,N_7661);
and U8199 (N_8199,N_7738,N_7540);
and U8200 (N_8200,N_7811,N_7867);
or U8201 (N_8201,N_7431,N_7140);
and U8202 (N_8202,N_7795,N_7191);
nor U8203 (N_8203,N_7333,N_7229);
nor U8204 (N_8204,N_7998,N_7852);
nand U8205 (N_8205,N_7007,N_7922);
or U8206 (N_8206,N_7032,N_7834);
nand U8207 (N_8207,N_7175,N_7544);
and U8208 (N_8208,N_7849,N_7081);
nand U8209 (N_8209,N_7689,N_7920);
nand U8210 (N_8210,N_7687,N_7541);
nor U8211 (N_8211,N_7874,N_7974);
nand U8212 (N_8212,N_7780,N_7232);
or U8213 (N_8213,N_7659,N_7574);
or U8214 (N_8214,N_7641,N_7192);
nor U8215 (N_8215,N_7205,N_7509);
and U8216 (N_8216,N_7287,N_7984);
nand U8217 (N_8217,N_7004,N_7671);
nand U8218 (N_8218,N_7531,N_7796);
or U8219 (N_8219,N_7407,N_7656);
and U8220 (N_8220,N_7921,N_7445);
nand U8221 (N_8221,N_7220,N_7021);
xnor U8222 (N_8222,N_7806,N_7125);
xor U8223 (N_8223,N_7200,N_7947);
nand U8224 (N_8224,N_7343,N_7785);
nand U8225 (N_8225,N_7734,N_7802);
nand U8226 (N_8226,N_7790,N_7181);
nor U8227 (N_8227,N_7943,N_7347);
nand U8228 (N_8228,N_7105,N_7665);
nand U8229 (N_8229,N_7011,N_7705);
or U8230 (N_8230,N_7616,N_7164);
or U8231 (N_8231,N_7581,N_7417);
and U8232 (N_8232,N_7591,N_7923);
nand U8233 (N_8233,N_7608,N_7264);
or U8234 (N_8234,N_7278,N_7025);
or U8235 (N_8235,N_7422,N_7621);
and U8236 (N_8236,N_7895,N_7579);
or U8237 (N_8237,N_7012,N_7681);
nand U8238 (N_8238,N_7421,N_7432);
nor U8239 (N_8239,N_7088,N_7940);
nand U8240 (N_8240,N_7915,N_7329);
nand U8241 (N_8241,N_7457,N_7117);
nor U8242 (N_8242,N_7827,N_7740);
nor U8243 (N_8243,N_7067,N_7322);
xor U8244 (N_8244,N_7498,N_7605);
nor U8245 (N_8245,N_7084,N_7325);
nor U8246 (N_8246,N_7917,N_7508);
nand U8247 (N_8247,N_7161,N_7174);
nand U8248 (N_8248,N_7203,N_7837);
nand U8249 (N_8249,N_7309,N_7682);
and U8250 (N_8250,N_7952,N_7400);
and U8251 (N_8251,N_7729,N_7298);
and U8252 (N_8252,N_7086,N_7160);
nand U8253 (N_8253,N_7062,N_7910);
and U8254 (N_8254,N_7578,N_7553);
or U8255 (N_8255,N_7216,N_7406);
nor U8256 (N_8256,N_7813,N_7114);
nor U8257 (N_8257,N_7993,N_7861);
and U8258 (N_8258,N_7402,N_7112);
xor U8259 (N_8259,N_7321,N_7896);
nor U8260 (N_8260,N_7120,N_7631);
nor U8261 (N_8261,N_7877,N_7017);
nor U8262 (N_8262,N_7075,N_7155);
xnor U8263 (N_8263,N_7269,N_7939);
nor U8264 (N_8264,N_7511,N_7655);
nor U8265 (N_8265,N_7652,N_7295);
or U8266 (N_8266,N_7543,N_7663);
nor U8267 (N_8267,N_7883,N_7040);
or U8268 (N_8268,N_7123,N_7959);
or U8269 (N_8269,N_7438,N_7212);
and U8270 (N_8270,N_7404,N_7819);
nand U8271 (N_8271,N_7454,N_7990);
nand U8272 (N_8272,N_7733,N_7797);
or U8273 (N_8273,N_7098,N_7029);
nor U8274 (N_8274,N_7588,N_7570);
nand U8275 (N_8275,N_7119,N_7654);
xnor U8276 (N_8276,N_7137,N_7049);
nand U8277 (N_8277,N_7516,N_7169);
xor U8278 (N_8278,N_7949,N_7619);
and U8279 (N_8279,N_7933,N_7368);
nor U8280 (N_8280,N_7537,N_7464);
or U8281 (N_8281,N_7599,N_7398);
nor U8282 (N_8282,N_7339,N_7530);
and U8283 (N_8283,N_7296,N_7440);
nand U8284 (N_8284,N_7370,N_7315);
or U8285 (N_8285,N_7453,N_7673);
nand U8286 (N_8286,N_7173,N_7980);
or U8287 (N_8287,N_7805,N_7902);
or U8288 (N_8288,N_7856,N_7279);
xnor U8289 (N_8289,N_7857,N_7786);
nand U8290 (N_8290,N_7106,N_7187);
nand U8291 (N_8291,N_7163,N_7183);
or U8292 (N_8292,N_7270,N_7719);
or U8293 (N_8293,N_7031,N_7242);
and U8294 (N_8294,N_7566,N_7152);
nor U8295 (N_8295,N_7423,N_7679);
xnor U8296 (N_8296,N_7649,N_7828);
and U8297 (N_8297,N_7771,N_7982);
and U8298 (N_8298,N_7330,N_7087);
xor U8299 (N_8299,N_7927,N_7082);
or U8300 (N_8300,N_7593,N_7853);
nor U8301 (N_8301,N_7812,N_7491);
nor U8302 (N_8302,N_7935,N_7099);
or U8303 (N_8303,N_7503,N_7248);
or U8304 (N_8304,N_7999,N_7382);
and U8305 (N_8305,N_7983,N_7227);
xnor U8306 (N_8306,N_7709,N_7153);
and U8307 (N_8307,N_7838,N_7794);
nand U8308 (N_8308,N_7901,N_7244);
and U8309 (N_8309,N_7179,N_7313);
and U8310 (N_8310,N_7288,N_7323);
nor U8311 (N_8311,N_7364,N_7762);
nor U8312 (N_8312,N_7778,N_7374);
nand U8313 (N_8313,N_7028,N_7946);
and U8314 (N_8314,N_7022,N_7210);
or U8315 (N_8315,N_7033,N_7078);
nor U8316 (N_8316,N_7350,N_7317);
nor U8317 (N_8317,N_7758,N_7647);
and U8318 (N_8318,N_7168,N_7714);
and U8319 (N_8319,N_7064,N_7750);
nor U8320 (N_8320,N_7052,N_7189);
xor U8321 (N_8321,N_7760,N_7005);
or U8322 (N_8322,N_7623,N_7273);
and U8323 (N_8323,N_7110,N_7841);
nor U8324 (N_8324,N_7166,N_7369);
nor U8325 (N_8325,N_7299,N_7128);
or U8326 (N_8326,N_7319,N_7826);
nor U8327 (N_8327,N_7425,N_7474);
or U8328 (N_8328,N_7351,N_7657);
nand U8329 (N_8329,N_7561,N_7089);
and U8330 (N_8330,N_7816,N_7545);
nand U8331 (N_8331,N_7622,N_7094);
nand U8332 (N_8332,N_7471,N_7126);
or U8333 (N_8333,N_7992,N_7037);
nand U8334 (N_8334,N_7290,N_7068);
nor U8335 (N_8335,N_7275,N_7928);
nor U8336 (N_8336,N_7602,N_7782);
xnor U8337 (N_8337,N_7798,N_7565);
or U8338 (N_8338,N_7753,N_7409);
xor U8339 (N_8339,N_7976,N_7527);
nand U8340 (N_8340,N_7410,N_7962);
or U8341 (N_8341,N_7170,N_7000);
xor U8342 (N_8342,N_7073,N_7552);
xor U8343 (N_8343,N_7524,N_7411);
or U8344 (N_8344,N_7484,N_7829);
xnor U8345 (N_8345,N_7426,N_7015);
and U8346 (N_8346,N_7887,N_7906);
nand U8347 (N_8347,N_7609,N_7514);
or U8348 (N_8348,N_7107,N_7815);
or U8349 (N_8349,N_7281,N_7632);
and U8350 (N_8350,N_7177,N_7535);
nor U8351 (N_8351,N_7692,N_7121);
xnor U8352 (N_8352,N_7185,N_7728);
or U8353 (N_8353,N_7027,N_7851);
and U8354 (N_8354,N_7919,N_7306);
nand U8355 (N_8355,N_7953,N_7784);
and U8356 (N_8356,N_7217,N_7965);
nand U8357 (N_8357,N_7247,N_7115);
xor U8358 (N_8358,N_7066,N_7154);
and U8359 (N_8359,N_7386,N_7408);
nor U8360 (N_8360,N_7551,N_7201);
or U8361 (N_8361,N_7777,N_7367);
nor U8362 (N_8362,N_7501,N_7696);
nand U8363 (N_8363,N_7289,N_7697);
nand U8364 (N_8364,N_7932,N_7612);
nor U8365 (N_8365,N_7207,N_7057);
and U8366 (N_8366,N_7433,N_7956);
or U8367 (N_8367,N_7528,N_7707);
xnor U8368 (N_8368,N_7878,N_7292);
nand U8369 (N_8369,N_7562,N_7627);
nand U8370 (N_8370,N_7462,N_7948);
and U8371 (N_8371,N_7936,N_7437);
xor U8372 (N_8372,N_7416,N_7645);
and U8373 (N_8373,N_7723,N_7047);
or U8374 (N_8374,N_7477,N_7625);
nand U8375 (N_8375,N_7741,N_7261);
nand U8376 (N_8376,N_7265,N_7225);
nor U8377 (N_8377,N_7629,N_7156);
or U8378 (N_8378,N_7662,N_7389);
and U8379 (N_8379,N_7499,N_7830);
and U8380 (N_8380,N_7427,N_7648);
and U8381 (N_8381,N_7311,N_7312);
or U8382 (N_8382,N_7253,N_7523);
and U8383 (N_8383,N_7051,N_7358);
nor U8384 (N_8384,N_7934,N_7904);
and U8385 (N_8385,N_7480,N_7842);
xor U8386 (N_8386,N_7010,N_7987);
nand U8387 (N_8387,N_7695,N_7211);
xor U8388 (N_8388,N_7441,N_7840);
or U8389 (N_8389,N_7572,N_7413);
and U8390 (N_8390,N_7594,N_7241);
and U8391 (N_8391,N_7646,N_7614);
nand U8392 (N_8392,N_7483,N_7360);
or U8393 (N_8393,N_7059,N_7102);
or U8394 (N_8394,N_7994,N_7703);
or U8395 (N_8395,N_7063,N_7135);
nand U8396 (N_8396,N_7836,N_7854);
nor U8397 (N_8397,N_7966,N_7053);
and U8398 (N_8398,N_7061,N_7359);
nor U8399 (N_8399,N_7092,N_7142);
and U8400 (N_8400,N_7044,N_7510);
nand U8401 (N_8401,N_7997,N_7434);
nor U8402 (N_8402,N_7556,N_7467);
nor U8403 (N_8403,N_7294,N_7644);
nor U8404 (N_8404,N_7575,N_7056);
or U8405 (N_8405,N_7560,N_7722);
or U8406 (N_8406,N_7109,N_7259);
and U8407 (N_8407,N_7310,N_7060);
nor U8408 (N_8408,N_7222,N_7365);
xor U8409 (N_8409,N_7893,N_7799);
nand U8410 (N_8410,N_7638,N_7101);
and U8411 (N_8411,N_7900,N_7744);
nor U8412 (N_8412,N_7371,N_7093);
nor U8413 (N_8413,N_7748,N_7447);
or U8414 (N_8414,N_7390,N_7332);
or U8415 (N_8415,N_7604,N_7669);
and U8416 (N_8416,N_7818,N_7280);
and U8417 (N_8417,N_7909,N_7672);
and U8418 (N_8418,N_7396,N_7559);
and U8419 (N_8419,N_7823,N_7972);
nor U8420 (N_8420,N_7171,N_7637);
or U8421 (N_8421,N_7755,N_7254);
and U8422 (N_8422,N_7716,N_7338);
xnor U8423 (N_8423,N_7557,N_7504);
or U8424 (N_8424,N_7702,N_7209);
nor U8425 (N_8425,N_7585,N_7690);
or U8426 (N_8426,N_7564,N_7476);
nand U8427 (N_8427,N_7850,N_7352);
or U8428 (N_8428,N_7831,N_7529);
or U8429 (N_8429,N_7208,N_7334);
and U8430 (N_8430,N_7348,N_7788);
and U8431 (N_8431,N_7150,N_7520);
nor U8432 (N_8432,N_7019,N_7077);
nand U8433 (N_8433,N_7481,N_7182);
or U8434 (N_8434,N_7680,N_7708);
and U8435 (N_8435,N_7190,N_7458);
and U8436 (N_8436,N_7598,N_7318);
nand U8437 (N_8437,N_7046,N_7774);
nand U8438 (N_8438,N_7172,N_7538);
nand U8439 (N_8439,N_7486,N_7822);
xnor U8440 (N_8440,N_7376,N_7978);
nor U8441 (N_8441,N_7964,N_7860);
nor U8442 (N_8442,N_7452,N_7684);
nor U8443 (N_8443,N_7361,N_7301);
xnor U8444 (N_8444,N_7124,N_7548);
nor U8445 (N_8445,N_7468,N_7165);
and U8446 (N_8446,N_7869,N_7911);
and U8447 (N_8447,N_7731,N_7111);
nand U8448 (N_8448,N_7676,N_7018);
nor U8449 (N_8449,N_7418,N_7518);
or U8450 (N_8450,N_7704,N_7633);
nor U8451 (N_8451,N_7897,N_7266);
nor U8452 (N_8452,N_7793,N_7328);
nand U8453 (N_8453,N_7100,N_7881);
nor U8454 (N_8454,N_7699,N_7304);
or U8455 (N_8455,N_7885,N_7596);
nand U8456 (N_8456,N_7443,N_7674);
xnor U8457 (N_8457,N_7439,N_7478);
and U8458 (N_8458,N_7640,N_7769);
or U8459 (N_8459,N_7639,N_7660);
or U8460 (N_8460,N_7558,N_7890);
xnor U8461 (N_8461,N_7127,N_7745);
or U8462 (N_8462,N_7379,N_7377);
and U8463 (N_8463,N_7048,N_7314);
nor U8464 (N_8464,N_7461,N_7506);
nand U8465 (N_8465,N_7617,N_7929);
nor U8466 (N_8466,N_7526,N_7635);
or U8467 (N_8467,N_7399,N_7775);
or U8468 (N_8468,N_7180,N_7710);
and U8469 (N_8469,N_7344,N_7226);
nor U8470 (N_8470,N_7274,N_7401);
xor U8471 (N_8471,N_7346,N_7996);
nand U8472 (N_8472,N_7355,N_7542);
nand U8473 (N_8473,N_7252,N_7970);
nand U8474 (N_8474,N_7650,N_7493);
nand U8475 (N_8475,N_7403,N_7620);
nand U8476 (N_8476,N_7345,N_7720);
and U8477 (N_8477,N_7583,N_7455);
or U8478 (N_8478,N_7302,N_7034);
nor U8479 (N_8479,N_7097,N_7038);
and U8480 (N_8480,N_7899,N_7751);
nor U8481 (N_8481,N_7263,N_7918);
nor U8482 (N_8482,N_7603,N_7139);
or U8483 (N_8483,N_7512,N_7008);
xor U8484 (N_8484,N_7715,N_7444);
nor U8485 (N_8485,N_7147,N_7014);
or U8486 (N_8486,N_7036,N_7630);
and U8487 (N_8487,N_7349,N_7507);
nor U8488 (N_8488,N_7393,N_7573);
or U8489 (N_8489,N_7739,N_7219);
or U8490 (N_8490,N_7586,N_7013);
nor U8491 (N_8491,N_7479,N_7381);
or U8492 (N_8492,N_7677,N_7977);
nor U8493 (N_8493,N_7490,N_7243);
or U8494 (N_8494,N_7957,N_7601);
nor U8495 (N_8495,N_7905,N_7151);
nor U8496 (N_8496,N_7297,N_7459);
nor U8497 (N_8497,N_7026,N_7045);
or U8498 (N_8498,N_7864,N_7331);
or U8499 (N_8499,N_7405,N_7988);
nand U8500 (N_8500,N_7840,N_7139);
nand U8501 (N_8501,N_7075,N_7080);
nor U8502 (N_8502,N_7469,N_7555);
nand U8503 (N_8503,N_7058,N_7955);
nand U8504 (N_8504,N_7295,N_7354);
or U8505 (N_8505,N_7531,N_7749);
nand U8506 (N_8506,N_7322,N_7201);
or U8507 (N_8507,N_7101,N_7747);
xor U8508 (N_8508,N_7067,N_7834);
and U8509 (N_8509,N_7337,N_7439);
nor U8510 (N_8510,N_7372,N_7811);
nand U8511 (N_8511,N_7285,N_7246);
and U8512 (N_8512,N_7446,N_7255);
and U8513 (N_8513,N_7210,N_7850);
nand U8514 (N_8514,N_7831,N_7795);
or U8515 (N_8515,N_7720,N_7798);
nor U8516 (N_8516,N_7104,N_7237);
nand U8517 (N_8517,N_7610,N_7682);
nor U8518 (N_8518,N_7024,N_7402);
nor U8519 (N_8519,N_7105,N_7190);
and U8520 (N_8520,N_7070,N_7952);
or U8521 (N_8521,N_7843,N_7801);
nand U8522 (N_8522,N_7602,N_7957);
nand U8523 (N_8523,N_7227,N_7047);
or U8524 (N_8524,N_7200,N_7062);
nor U8525 (N_8525,N_7143,N_7898);
or U8526 (N_8526,N_7321,N_7114);
xor U8527 (N_8527,N_7124,N_7842);
and U8528 (N_8528,N_7550,N_7292);
and U8529 (N_8529,N_7003,N_7504);
or U8530 (N_8530,N_7080,N_7104);
and U8531 (N_8531,N_7766,N_7383);
and U8532 (N_8532,N_7885,N_7276);
or U8533 (N_8533,N_7704,N_7385);
and U8534 (N_8534,N_7137,N_7655);
or U8535 (N_8535,N_7043,N_7477);
nor U8536 (N_8536,N_7910,N_7662);
or U8537 (N_8537,N_7023,N_7840);
nor U8538 (N_8538,N_7121,N_7063);
nor U8539 (N_8539,N_7617,N_7393);
nor U8540 (N_8540,N_7381,N_7260);
or U8541 (N_8541,N_7451,N_7128);
nand U8542 (N_8542,N_7758,N_7184);
or U8543 (N_8543,N_7254,N_7352);
nor U8544 (N_8544,N_7189,N_7362);
nand U8545 (N_8545,N_7494,N_7398);
or U8546 (N_8546,N_7436,N_7292);
or U8547 (N_8547,N_7212,N_7579);
or U8548 (N_8548,N_7947,N_7732);
nand U8549 (N_8549,N_7637,N_7389);
and U8550 (N_8550,N_7414,N_7438);
and U8551 (N_8551,N_7708,N_7831);
nor U8552 (N_8552,N_7199,N_7520);
nand U8553 (N_8553,N_7234,N_7974);
nor U8554 (N_8554,N_7075,N_7091);
xor U8555 (N_8555,N_7117,N_7605);
and U8556 (N_8556,N_7294,N_7395);
or U8557 (N_8557,N_7592,N_7837);
nand U8558 (N_8558,N_7697,N_7342);
or U8559 (N_8559,N_7433,N_7538);
nor U8560 (N_8560,N_7046,N_7085);
nor U8561 (N_8561,N_7713,N_7770);
or U8562 (N_8562,N_7551,N_7902);
and U8563 (N_8563,N_7368,N_7244);
nor U8564 (N_8564,N_7297,N_7783);
nand U8565 (N_8565,N_7266,N_7759);
nor U8566 (N_8566,N_7107,N_7198);
or U8567 (N_8567,N_7133,N_7606);
and U8568 (N_8568,N_7167,N_7268);
nor U8569 (N_8569,N_7000,N_7679);
or U8570 (N_8570,N_7063,N_7097);
xnor U8571 (N_8571,N_7250,N_7101);
xor U8572 (N_8572,N_7077,N_7365);
and U8573 (N_8573,N_7352,N_7608);
nand U8574 (N_8574,N_7149,N_7748);
nor U8575 (N_8575,N_7498,N_7019);
or U8576 (N_8576,N_7734,N_7530);
nor U8577 (N_8577,N_7670,N_7191);
nand U8578 (N_8578,N_7707,N_7992);
nor U8579 (N_8579,N_7791,N_7934);
nor U8580 (N_8580,N_7686,N_7651);
nand U8581 (N_8581,N_7424,N_7574);
or U8582 (N_8582,N_7605,N_7857);
and U8583 (N_8583,N_7505,N_7820);
or U8584 (N_8584,N_7778,N_7433);
or U8585 (N_8585,N_7540,N_7881);
nand U8586 (N_8586,N_7785,N_7255);
nand U8587 (N_8587,N_7232,N_7680);
and U8588 (N_8588,N_7863,N_7622);
nor U8589 (N_8589,N_7376,N_7689);
nor U8590 (N_8590,N_7183,N_7083);
and U8591 (N_8591,N_7695,N_7561);
nor U8592 (N_8592,N_7774,N_7494);
and U8593 (N_8593,N_7673,N_7691);
nor U8594 (N_8594,N_7854,N_7005);
nand U8595 (N_8595,N_7709,N_7115);
nor U8596 (N_8596,N_7683,N_7504);
and U8597 (N_8597,N_7655,N_7547);
nand U8598 (N_8598,N_7548,N_7902);
xor U8599 (N_8599,N_7350,N_7744);
and U8600 (N_8600,N_7224,N_7961);
or U8601 (N_8601,N_7026,N_7609);
and U8602 (N_8602,N_7705,N_7728);
xor U8603 (N_8603,N_7318,N_7505);
nor U8604 (N_8604,N_7414,N_7627);
and U8605 (N_8605,N_7560,N_7510);
nor U8606 (N_8606,N_7660,N_7900);
xnor U8607 (N_8607,N_7395,N_7840);
and U8608 (N_8608,N_7675,N_7104);
nand U8609 (N_8609,N_7964,N_7398);
or U8610 (N_8610,N_7896,N_7606);
or U8611 (N_8611,N_7203,N_7927);
nor U8612 (N_8612,N_7568,N_7499);
and U8613 (N_8613,N_7365,N_7150);
nor U8614 (N_8614,N_7701,N_7564);
or U8615 (N_8615,N_7409,N_7084);
nor U8616 (N_8616,N_7826,N_7764);
and U8617 (N_8617,N_7293,N_7367);
nand U8618 (N_8618,N_7345,N_7375);
or U8619 (N_8619,N_7243,N_7578);
and U8620 (N_8620,N_7067,N_7932);
and U8621 (N_8621,N_7549,N_7137);
nor U8622 (N_8622,N_7321,N_7673);
nand U8623 (N_8623,N_7407,N_7013);
and U8624 (N_8624,N_7028,N_7992);
and U8625 (N_8625,N_7327,N_7387);
and U8626 (N_8626,N_7659,N_7258);
xor U8627 (N_8627,N_7515,N_7126);
or U8628 (N_8628,N_7074,N_7558);
or U8629 (N_8629,N_7770,N_7716);
xnor U8630 (N_8630,N_7584,N_7913);
xor U8631 (N_8631,N_7708,N_7872);
or U8632 (N_8632,N_7142,N_7584);
nand U8633 (N_8633,N_7079,N_7688);
nand U8634 (N_8634,N_7216,N_7822);
nor U8635 (N_8635,N_7980,N_7012);
nand U8636 (N_8636,N_7375,N_7436);
nand U8637 (N_8637,N_7066,N_7987);
nand U8638 (N_8638,N_7893,N_7836);
nand U8639 (N_8639,N_7602,N_7549);
nor U8640 (N_8640,N_7350,N_7793);
and U8641 (N_8641,N_7692,N_7338);
or U8642 (N_8642,N_7722,N_7484);
xnor U8643 (N_8643,N_7930,N_7544);
and U8644 (N_8644,N_7619,N_7082);
and U8645 (N_8645,N_7386,N_7908);
nand U8646 (N_8646,N_7141,N_7737);
nand U8647 (N_8647,N_7824,N_7929);
and U8648 (N_8648,N_7695,N_7518);
nand U8649 (N_8649,N_7282,N_7550);
and U8650 (N_8650,N_7874,N_7093);
or U8651 (N_8651,N_7708,N_7710);
or U8652 (N_8652,N_7378,N_7385);
and U8653 (N_8653,N_7436,N_7972);
nand U8654 (N_8654,N_7957,N_7164);
and U8655 (N_8655,N_7011,N_7058);
and U8656 (N_8656,N_7263,N_7144);
nand U8657 (N_8657,N_7958,N_7131);
and U8658 (N_8658,N_7483,N_7803);
and U8659 (N_8659,N_7527,N_7891);
nand U8660 (N_8660,N_7112,N_7990);
and U8661 (N_8661,N_7768,N_7460);
or U8662 (N_8662,N_7237,N_7532);
or U8663 (N_8663,N_7852,N_7315);
nor U8664 (N_8664,N_7711,N_7932);
and U8665 (N_8665,N_7413,N_7759);
nor U8666 (N_8666,N_7488,N_7380);
or U8667 (N_8667,N_7748,N_7566);
or U8668 (N_8668,N_7821,N_7950);
xor U8669 (N_8669,N_7072,N_7460);
and U8670 (N_8670,N_7131,N_7551);
or U8671 (N_8671,N_7466,N_7791);
or U8672 (N_8672,N_7946,N_7779);
nor U8673 (N_8673,N_7128,N_7671);
and U8674 (N_8674,N_7477,N_7200);
xor U8675 (N_8675,N_7741,N_7526);
xor U8676 (N_8676,N_7612,N_7260);
and U8677 (N_8677,N_7021,N_7669);
nand U8678 (N_8678,N_7359,N_7737);
nand U8679 (N_8679,N_7639,N_7129);
and U8680 (N_8680,N_7021,N_7877);
nand U8681 (N_8681,N_7287,N_7752);
or U8682 (N_8682,N_7781,N_7038);
nand U8683 (N_8683,N_7921,N_7765);
nor U8684 (N_8684,N_7050,N_7792);
and U8685 (N_8685,N_7370,N_7544);
and U8686 (N_8686,N_7688,N_7942);
nand U8687 (N_8687,N_7760,N_7676);
nor U8688 (N_8688,N_7687,N_7155);
xnor U8689 (N_8689,N_7612,N_7510);
nor U8690 (N_8690,N_7437,N_7840);
xnor U8691 (N_8691,N_7194,N_7365);
nor U8692 (N_8692,N_7908,N_7813);
nor U8693 (N_8693,N_7178,N_7760);
nand U8694 (N_8694,N_7052,N_7219);
xor U8695 (N_8695,N_7399,N_7453);
xor U8696 (N_8696,N_7602,N_7276);
and U8697 (N_8697,N_7060,N_7597);
nand U8698 (N_8698,N_7631,N_7383);
nor U8699 (N_8699,N_7174,N_7084);
xnor U8700 (N_8700,N_7728,N_7891);
or U8701 (N_8701,N_7536,N_7751);
or U8702 (N_8702,N_7939,N_7898);
xor U8703 (N_8703,N_7571,N_7606);
or U8704 (N_8704,N_7300,N_7577);
or U8705 (N_8705,N_7017,N_7099);
xor U8706 (N_8706,N_7793,N_7587);
or U8707 (N_8707,N_7226,N_7363);
or U8708 (N_8708,N_7918,N_7345);
and U8709 (N_8709,N_7286,N_7986);
or U8710 (N_8710,N_7997,N_7726);
nor U8711 (N_8711,N_7144,N_7082);
and U8712 (N_8712,N_7311,N_7764);
and U8713 (N_8713,N_7507,N_7320);
nor U8714 (N_8714,N_7085,N_7507);
and U8715 (N_8715,N_7814,N_7071);
and U8716 (N_8716,N_7754,N_7746);
nand U8717 (N_8717,N_7168,N_7486);
nor U8718 (N_8718,N_7059,N_7067);
nand U8719 (N_8719,N_7847,N_7836);
or U8720 (N_8720,N_7901,N_7882);
or U8721 (N_8721,N_7240,N_7375);
nor U8722 (N_8722,N_7547,N_7509);
and U8723 (N_8723,N_7807,N_7629);
and U8724 (N_8724,N_7791,N_7672);
nor U8725 (N_8725,N_7086,N_7028);
or U8726 (N_8726,N_7017,N_7227);
nand U8727 (N_8727,N_7576,N_7677);
and U8728 (N_8728,N_7937,N_7861);
nor U8729 (N_8729,N_7377,N_7358);
xor U8730 (N_8730,N_7515,N_7685);
and U8731 (N_8731,N_7899,N_7873);
nand U8732 (N_8732,N_7860,N_7765);
and U8733 (N_8733,N_7785,N_7760);
and U8734 (N_8734,N_7271,N_7221);
xor U8735 (N_8735,N_7332,N_7450);
and U8736 (N_8736,N_7726,N_7577);
or U8737 (N_8737,N_7763,N_7029);
nor U8738 (N_8738,N_7275,N_7828);
nand U8739 (N_8739,N_7086,N_7521);
nand U8740 (N_8740,N_7271,N_7565);
or U8741 (N_8741,N_7788,N_7544);
nor U8742 (N_8742,N_7760,N_7734);
nor U8743 (N_8743,N_7654,N_7812);
and U8744 (N_8744,N_7630,N_7513);
nand U8745 (N_8745,N_7761,N_7259);
and U8746 (N_8746,N_7774,N_7362);
nand U8747 (N_8747,N_7972,N_7990);
nor U8748 (N_8748,N_7599,N_7696);
or U8749 (N_8749,N_7837,N_7186);
xnor U8750 (N_8750,N_7130,N_7443);
nor U8751 (N_8751,N_7647,N_7098);
nand U8752 (N_8752,N_7914,N_7038);
nand U8753 (N_8753,N_7448,N_7110);
nand U8754 (N_8754,N_7492,N_7499);
nand U8755 (N_8755,N_7563,N_7900);
nand U8756 (N_8756,N_7568,N_7578);
nor U8757 (N_8757,N_7740,N_7140);
nor U8758 (N_8758,N_7108,N_7702);
xor U8759 (N_8759,N_7674,N_7425);
or U8760 (N_8760,N_7916,N_7682);
or U8761 (N_8761,N_7779,N_7242);
xnor U8762 (N_8762,N_7631,N_7414);
and U8763 (N_8763,N_7397,N_7810);
and U8764 (N_8764,N_7201,N_7204);
nor U8765 (N_8765,N_7469,N_7405);
nand U8766 (N_8766,N_7642,N_7203);
nand U8767 (N_8767,N_7968,N_7642);
or U8768 (N_8768,N_7909,N_7728);
or U8769 (N_8769,N_7083,N_7801);
xor U8770 (N_8770,N_7480,N_7604);
nor U8771 (N_8771,N_7570,N_7660);
or U8772 (N_8772,N_7902,N_7294);
and U8773 (N_8773,N_7200,N_7961);
nand U8774 (N_8774,N_7846,N_7210);
nand U8775 (N_8775,N_7943,N_7174);
xor U8776 (N_8776,N_7536,N_7490);
xor U8777 (N_8777,N_7344,N_7420);
xor U8778 (N_8778,N_7570,N_7398);
nand U8779 (N_8779,N_7610,N_7079);
nand U8780 (N_8780,N_7091,N_7244);
or U8781 (N_8781,N_7121,N_7497);
or U8782 (N_8782,N_7419,N_7245);
and U8783 (N_8783,N_7961,N_7519);
xnor U8784 (N_8784,N_7020,N_7478);
or U8785 (N_8785,N_7424,N_7094);
nor U8786 (N_8786,N_7488,N_7942);
nor U8787 (N_8787,N_7714,N_7853);
or U8788 (N_8788,N_7418,N_7917);
nand U8789 (N_8789,N_7729,N_7328);
nor U8790 (N_8790,N_7780,N_7954);
nor U8791 (N_8791,N_7778,N_7035);
or U8792 (N_8792,N_7272,N_7298);
and U8793 (N_8793,N_7793,N_7434);
and U8794 (N_8794,N_7294,N_7365);
or U8795 (N_8795,N_7367,N_7883);
and U8796 (N_8796,N_7958,N_7875);
and U8797 (N_8797,N_7103,N_7008);
or U8798 (N_8798,N_7227,N_7446);
nand U8799 (N_8799,N_7186,N_7432);
nor U8800 (N_8800,N_7991,N_7330);
or U8801 (N_8801,N_7367,N_7578);
nor U8802 (N_8802,N_7311,N_7361);
nand U8803 (N_8803,N_7733,N_7619);
xnor U8804 (N_8804,N_7880,N_7336);
nand U8805 (N_8805,N_7880,N_7132);
and U8806 (N_8806,N_7120,N_7337);
nor U8807 (N_8807,N_7923,N_7879);
nor U8808 (N_8808,N_7923,N_7406);
and U8809 (N_8809,N_7976,N_7628);
or U8810 (N_8810,N_7008,N_7445);
or U8811 (N_8811,N_7174,N_7507);
xor U8812 (N_8812,N_7995,N_7546);
nand U8813 (N_8813,N_7847,N_7215);
xnor U8814 (N_8814,N_7085,N_7479);
and U8815 (N_8815,N_7496,N_7657);
nand U8816 (N_8816,N_7261,N_7467);
nand U8817 (N_8817,N_7993,N_7943);
and U8818 (N_8818,N_7119,N_7171);
nand U8819 (N_8819,N_7041,N_7175);
xnor U8820 (N_8820,N_7848,N_7880);
and U8821 (N_8821,N_7470,N_7608);
nand U8822 (N_8822,N_7087,N_7546);
nor U8823 (N_8823,N_7342,N_7344);
or U8824 (N_8824,N_7542,N_7790);
and U8825 (N_8825,N_7124,N_7103);
or U8826 (N_8826,N_7638,N_7231);
and U8827 (N_8827,N_7854,N_7443);
nor U8828 (N_8828,N_7486,N_7332);
nor U8829 (N_8829,N_7516,N_7170);
nand U8830 (N_8830,N_7273,N_7227);
nand U8831 (N_8831,N_7706,N_7408);
and U8832 (N_8832,N_7395,N_7580);
nand U8833 (N_8833,N_7107,N_7774);
nor U8834 (N_8834,N_7532,N_7205);
xor U8835 (N_8835,N_7422,N_7706);
nand U8836 (N_8836,N_7846,N_7059);
nand U8837 (N_8837,N_7196,N_7524);
or U8838 (N_8838,N_7359,N_7240);
or U8839 (N_8839,N_7315,N_7205);
nor U8840 (N_8840,N_7243,N_7205);
and U8841 (N_8841,N_7206,N_7843);
and U8842 (N_8842,N_7866,N_7157);
nand U8843 (N_8843,N_7524,N_7699);
nand U8844 (N_8844,N_7696,N_7950);
nor U8845 (N_8845,N_7180,N_7591);
nor U8846 (N_8846,N_7196,N_7373);
or U8847 (N_8847,N_7155,N_7467);
or U8848 (N_8848,N_7606,N_7390);
or U8849 (N_8849,N_7261,N_7944);
nand U8850 (N_8850,N_7785,N_7249);
or U8851 (N_8851,N_7979,N_7359);
nand U8852 (N_8852,N_7382,N_7823);
nor U8853 (N_8853,N_7947,N_7495);
or U8854 (N_8854,N_7830,N_7652);
xor U8855 (N_8855,N_7152,N_7193);
or U8856 (N_8856,N_7800,N_7784);
and U8857 (N_8857,N_7617,N_7421);
nand U8858 (N_8858,N_7050,N_7647);
or U8859 (N_8859,N_7200,N_7329);
xnor U8860 (N_8860,N_7320,N_7347);
xnor U8861 (N_8861,N_7158,N_7522);
or U8862 (N_8862,N_7107,N_7068);
nand U8863 (N_8863,N_7026,N_7502);
nand U8864 (N_8864,N_7105,N_7677);
and U8865 (N_8865,N_7574,N_7136);
nand U8866 (N_8866,N_7952,N_7198);
or U8867 (N_8867,N_7763,N_7809);
nor U8868 (N_8868,N_7594,N_7544);
nand U8869 (N_8869,N_7461,N_7325);
nor U8870 (N_8870,N_7789,N_7935);
nand U8871 (N_8871,N_7723,N_7557);
xor U8872 (N_8872,N_7257,N_7719);
and U8873 (N_8873,N_7261,N_7531);
or U8874 (N_8874,N_7185,N_7505);
or U8875 (N_8875,N_7929,N_7372);
and U8876 (N_8876,N_7380,N_7068);
nor U8877 (N_8877,N_7930,N_7469);
nor U8878 (N_8878,N_7955,N_7536);
nand U8879 (N_8879,N_7197,N_7857);
and U8880 (N_8880,N_7807,N_7780);
and U8881 (N_8881,N_7910,N_7760);
or U8882 (N_8882,N_7248,N_7163);
and U8883 (N_8883,N_7008,N_7853);
xor U8884 (N_8884,N_7410,N_7382);
nand U8885 (N_8885,N_7468,N_7756);
and U8886 (N_8886,N_7872,N_7152);
nand U8887 (N_8887,N_7025,N_7508);
nor U8888 (N_8888,N_7256,N_7630);
and U8889 (N_8889,N_7175,N_7080);
nor U8890 (N_8890,N_7211,N_7054);
and U8891 (N_8891,N_7116,N_7853);
and U8892 (N_8892,N_7118,N_7943);
xor U8893 (N_8893,N_7406,N_7391);
nor U8894 (N_8894,N_7514,N_7967);
nand U8895 (N_8895,N_7841,N_7396);
and U8896 (N_8896,N_7430,N_7087);
or U8897 (N_8897,N_7243,N_7066);
and U8898 (N_8898,N_7584,N_7837);
nand U8899 (N_8899,N_7280,N_7690);
and U8900 (N_8900,N_7129,N_7763);
xor U8901 (N_8901,N_7176,N_7271);
or U8902 (N_8902,N_7972,N_7124);
or U8903 (N_8903,N_7504,N_7529);
nor U8904 (N_8904,N_7044,N_7479);
nand U8905 (N_8905,N_7958,N_7848);
nor U8906 (N_8906,N_7727,N_7855);
nor U8907 (N_8907,N_7947,N_7636);
nand U8908 (N_8908,N_7335,N_7946);
or U8909 (N_8909,N_7868,N_7846);
or U8910 (N_8910,N_7841,N_7399);
and U8911 (N_8911,N_7971,N_7605);
nand U8912 (N_8912,N_7969,N_7000);
nand U8913 (N_8913,N_7637,N_7999);
nor U8914 (N_8914,N_7537,N_7098);
nor U8915 (N_8915,N_7714,N_7765);
nor U8916 (N_8916,N_7562,N_7709);
xor U8917 (N_8917,N_7186,N_7901);
nand U8918 (N_8918,N_7259,N_7084);
and U8919 (N_8919,N_7121,N_7304);
nor U8920 (N_8920,N_7210,N_7196);
and U8921 (N_8921,N_7692,N_7218);
or U8922 (N_8922,N_7047,N_7659);
and U8923 (N_8923,N_7732,N_7091);
and U8924 (N_8924,N_7601,N_7648);
nor U8925 (N_8925,N_7344,N_7053);
or U8926 (N_8926,N_7407,N_7780);
nor U8927 (N_8927,N_7900,N_7528);
nand U8928 (N_8928,N_7722,N_7692);
and U8929 (N_8929,N_7161,N_7989);
nand U8930 (N_8930,N_7847,N_7254);
nand U8931 (N_8931,N_7769,N_7054);
nor U8932 (N_8932,N_7681,N_7319);
nor U8933 (N_8933,N_7266,N_7545);
nor U8934 (N_8934,N_7735,N_7756);
or U8935 (N_8935,N_7887,N_7324);
or U8936 (N_8936,N_7783,N_7989);
and U8937 (N_8937,N_7241,N_7207);
nor U8938 (N_8938,N_7789,N_7927);
nand U8939 (N_8939,N_7395,N_7280);
nand U8940 (N_8940,N_7926,N_7786);
and U8941 (N_8941,N_7995,N_7821);
and U8942 (N_8942,N_7349,N_7263);
nand U8943 (N_8943,N_7022,N_7316);
or U8944 (N_8944,N_7202,N_7255);
nor U8945 (N_8945,N_7885,N_7837);
nor U8946 (N_8946,N_7901,N_7255);
xnor U8947 (N_8947,N_7066,N_7519);
or U8948 (N_8948,N_7413,N_7126);
xor U8949 (N_8949,N_7948,N_7818);
and U8950 (N_8950,N_7170,N_7837);
or U8951 (N_8951,N_7610,N_7882);
nand U8952 (N_8952,N_7217,N_7782);
xnor U8953 (N_8953,N_7368,N_7239);
nor U8954 (N_8954,N_7924,N_7969);
nor U8955 (N_8955,N_7166,N_7324);
nand U8956 (N_8956,N_7455,N_7023);
or U8957 (N_8957,N_7243,N_7051);
and U8958 (N_8958,N_7847,N_7344);
or U8959 (N_8959,N_7639,N_7488);
xor U8960 (N_8960,N_7305,N_7200);
nand U8961 (N_8961,N_7598,N_7615);
nor U8962 (N_8962,N_7015,N_7874);
xor U8963 (N_8963,N_7362,N_7271);
nand U8964 (N_8964,N_7019,N_7048);
nand U8965 (N_8965,N_7558,N_7672);
nand U8966 (N_8966,N_7745,N_7704);
nor U8967 (N_8967,N_7831,N_7333);
nand U8968 (N_8968,N_7711,N_7098);
nor U8969 (N_8969,N_7270,N_7089);
nor U8970 (N_8970,N_7788,N_7961);
or U8971 (N_8971,N_7541,N_7652);
xor U8972 (N_8972,N_7463,N_7764);
nor U8973 (N_8973,N_7439,N_7049);
xnor U8974 (N_8974,N_7759,N_7225);
or U8975 (N_8975,N_7438,N_7553);
nor U8976 (N_8976,N_7892,N_7008);
nor U8977 (N_8977,N_7418,N_7894);
nand U8978 (N_8978,N_7426,N_7837);
xor U8979 (N_8979,N_7949,N_7247);
nand U8980 (N_8980,N_7015,N_7574);
xor U8981 (N_8981,N_7757,N_7666);
nor U8982 (N_8982,N_7997,N_7224);
nor U8983 (N_8983,N_7710,N_7817);
xnor U8984 (N_8984,N_7328,N_7080);
or U8985 (N_8985,N_7072,N_7223);
nor U8986 (N_8986,N_7228,N_7968);
or U8987 (N_8987,N_7330,N_7001);
and U8988 (N_8988,N_7135,N_7662);
nor U8989 (N_8989,N_7518,N_7640);
or U8990 (N_8990,N_7752,N_7317);
nor U8991 (N_8991,N_7139,N_7914);
or U8992 (N_8992,N_7953,N_7507);
and U8993 (N_8993,N_7833,N_7984);
nor U8994 (N_8994,N_7945,N_7716);
nand U8995 (N_8995,N_7379,N_7620);
or U8996 (N_8996,N_7913,N_7843);
or U8997 (N_8997,N_7463,N_7944);
nand U8998 (N_8998,N_7716,N_7145);
and U8999 (N_8999,N_7039,N_7721);
xnor U9000 (N_9000,N_8261,N_8382);
or U9001 (N_9001,N_8876,N_8226);
nor U9002 (N_9002,N_8600,N_8545);
and U9003 (N_9003,N_8137,N_8059);
nor U9004 (N_9004,N_8171,N_8399);
or U9005 (N_9005,N_8459,N_8042);
nor U9006 (N_9006,N_8515,N_8864);
xor U9007 (N_9007,N_8756,N_8945);
and U9008 (N_9008,N_8832,N_8190);
and U9009 (N_9009,N_8041,N_8485);
nand U9010 (N_9010,N_8166,N_8011);
nand U9011 (N_9011,N_8427,N_8500);
or U9012 (N_9012,N_8622,N_8280);
nor U9013 (N_9013,N_8238,N_8804);
and U9014 (N_9014,N_8263,N_8414);
nand U9015 (N_9015,N_8157,N_8722);
nor U9016 (N_9016,N_8122,N_8257);
nand U9017 (N_9017,N_8734,N_8281);
nor U9018 (N_9018,N_8327,N_8110);
and U9019 (N_9019,N_8540,N_8249);
nor U9020 (N_9020,N_8282,N_8401);
nand U9021 (N_9021,N_8017,N_8848);
or U9022 (N_9022,N_8986,N_8429);
nor U9023 (N_9023,N_8297,N_8340);
nand U9024 (N_9024,N_8370,N_8254);
or U9025 (N_9025,N_8172,N_8589);
nor U9026 (N_9026,N_8532,N_8809);
or U9027 (N_9027,N_8480,N_8939);
xor U9028 (N_9028,N_8522,N_8849);
nor U9029 (N_9029,N_8964,N_8646);
xnor U9030 (N_9030,N_8884,N_8363);
and U9031 (N_9031,N_8347,N_8434);
nand U9032 (N_9032,N_8073,N_8180);
xnor U9033 (N_9033,N_8898,N_8174);
or U9034 (N_9034,N_8627,N_8307);
or U9035 (N_9035,N_8103,N_8360);
or U9036 (N_9036,N_8634,N_8109);
and U9037 (N_9037,N_8018,N_8503);
xor U9038 (N_9038,N_8924,N_8711);
nand U9039 (N_9039,N_8854,N_8529);
and U9040 (N_9040,N_8558,N_8486);
nand U9041 (N_9041,N_8335,N_8315);
nand U9042 (N_9042,N_8195,N_8246);
xnor U9043 (N_9043,N_8816,N_8877);
nand U9044 (N_9044,N_8979,N_8375);
and U9045 (N_9045,N_8141,N_8426);
and U9046 (N_9046,N_8184,N_8085);
nor U9047 (N_9047,N_8683,N_8151);
nand U9048 (N_9048,N_8905,N_8996);
and U9049 (N_9049,N_8436,N_8610);
nor U9050 (N_9050,N_8016,N_8200);
or U9051 (N_9051,N_8690,N_8806);
xnor U9052 (N_9052,N_8118,N_8520);
or U9053 (N_9053,N_8078,N_8973);
nor U9054 (N_9054,N_8243,N_8299);
or U9055 (N_9055,N_8869,N_8620);
and U9056 (N_9056,N_8328,N_8681);
nand U9057 (N_9057,N_8564,N_8423);
xnor U9058 (N_9058,N_8717,N_8855);
or U9059 (N_9059,N_8484,N_8213);
or U9060 (N_9060,N_8206,N_8946);
nand U9061 (N_9061,N_8087,N_8398);
nor U9062 (N_9062,N_8597,N_8612);
xor U9063 (N_9063,N_8794,N_8111);
nor U9064 (N_9064,N_8439,N_8999);
xor U9065 (N_9065,N_8552,N_8630);
nor U9066 (N_9066,N_8736,N_8167);
nand U9067 (N_9067,N_8866,N_8588);
or U9068 (N_9068,N_8223,N_8329);
nor U9069 (N_9069,N_8727,N_8914);
nand U9070 (N_9070,N_8374,N_8005);
nand U9071 (N_9071,N_8472,N_8685);
or U9072 (N_9072,N_8779,N_8661);
or U9073 (N_9073,N_8859,N_8478);
nor U9074 (N_9074,N_8696,N_8183);
xor U9075 (N_9075,N_8524,N_8663);
and U9076 (N_9076,N_8063,N_8325);
nand U9077 (N_9077,N_8628,N_8695);
xnor U9078 (N_9078,N_8265,N_8697);
xor U9079 (N_9079,N_8189,N_8290);
or U9080 (N_9080,N_8050,N_8553);
nand U9081 (N_9081,N_8292,N_8186);
nand U9082 (N_9082,N_8992,N_8908);
nand U9083 (N_9083,N_8693,N_8850);
or U9084 (N_9084,N_8601,N_8729);
and U9085 (N_9085,N_8833,N_8134);
nand U9086 (N_9086,N_8680,N_8421);
nand U9087 (N_9087,N_8231,N_8258);
nor U9088 (N_9088,N_8049,N_8527);
nand U9089 (N_9089,N_8533,N_8959);
or U9090 (N_9090,N_8870,N_8193);
nand U9091 (N_9091,N_8512,N_8772);
and U9092 (N_9092,N_8494,N_8787);
nand U9093 (N_9093,N_8062,N_8726);
or U9094 (N_9094,N_8581,N_8428);
xnor U9095 (N_9095,N_8481,N_8438);
nand U9096 (N_9096,N_8507,N_8926);
nand U9097 (N_9097,N_8210,N_8626);
nand U9098 (N_9098,N_8922,N_8740);
nor U9099 (N_9099,N_8778,N_8351);
or U9100 (N_9100,N_8766,N_8081);
nand U9101 (N_9101,N_8917,N_8514);
and U9102 (N_9102,N_8700,N_8077);
and U9103 (N_9103,N_8170,N_8287);
nor U9104 (N_9104,N_8310,N_8294);
nand U9105 (N_9105,N_8827,N_8036);
and U9106 (N_9106,N_8803,N_8882);
nand U9107 (N_9107,N_8929,N_8356);
and U9108 (N_9108,N_8668,N_8955);
nand U9109 (N_9109,N_8493,N_8599);
nor U9110 (N_9110,N_8055,N_8921);
or U9111 (N_9111,N_8829,N_8400);
nor U9112 (N_9112,N_8760,N_8000);
nand U9113 (N_9113,N_8857,N_8487);
xor U9114 (N_9114,N_8357,N_8152);
nand U9115 (N_9115,N_8079,N_8225);
and U9116 (N_9116,N_8143,N_8311);
nand U9117 (N_9117,N_8277,N_8637);
nor U9118 (N_9118,N_8332,N_8821);
and U9119 (N_9119,N_8703,N_8314);
nor U9120 (N_9120,N_8918,N_8064);
and U9121 (N_9121,N_8271,N_8161);
nor U9122 (N_9122,N_8913,N_8121);
and U9123 (N_9123,N_8535,N_8296);
nand U9124 (N_9124,N_8348,N_8021);
nor U9125 (N_9125,N_8024,N_8454);
nand U9126 (N_9126,N_8495,N_8568);
or U9127 (N_9127,N_8925,N_8526);
nand U9128 (N_9128,N_8679,N_8739);
and U9129 (N_9129,N_8384,N_8886);
nor U9130 (N_9130,N_8108,N_8006);
xnor U9131 (N_9131,N_8227,N_8082);
or U9132 (N_9132,N_8587,N_8355);
and U9133 (N_9133,N_8878,N_8293);
and U9134 (N_9134,N_8684,N_8364);
nor U9135 (N_9135,N_8025,N_8272);
xor U9136 (N_9136,N_8040,N_8798);
nand U9137 (N_9137,N_8754,N_8026);
or U9138 (N_9138,N_8844,N_8657);
nor U9139 (N_9139,N_8031,N_8842);
or U9140 (N_9140,N_8102,N_8268);
nor U9141 (N_9141,N_8592,N_8274);
and U9142 (N_9142,N_8447,N_8686);
nand U9143 (N_9143,N_8219,N_8819);
xor U9144 (N_9144,N_8361,N_8306);
nand U9145 (N_9145,N_8702,N_8642);
nor U9146 (N_9146,N_8010,N_8138);
or U9147 (N_9147,N_8467,N_8463);
or U9148 (N_9148,N_8030,N_8738);
nand U9149 (N_9149,N_8699,N_8892);
and U9150 (N_9150,N_8653,N_8659);
nand U9151 (N_9151,N_8719,N_8625);
nor U9152 (N_9152,N_8070,N_8337);
and U9153 (N_9153,N_8903,N_8951);
or U9154 (N_9154,N_8129,N_8093);
or U9155 (N_9155,N_8741,N_8388);
nor U9156 (N_9156,N_8578,N_8267);
and U9157 (N_9157,N_8196,N_8631);
xnor U9158 (N_9158,N_8713,N_8320);
or U9159 (N_9159,N_8856,N_8199);
nor U9160 (N_9160,N_8912,N_8731);
or U9161 (N_9161,N_8723,N_8674);
nand U9162 (N_9162,N_8156,N_8163);
nand U9163 (N_9163,N_8165,N_8053);
nor U9164 (N_9164,N_8765,N_8004);
and U9165 (N_9165,N_8369,N_8120);
or U9166 (N_9166,N_8385,N_8594);
nand U9167 (N_9167,N_8034,N_8839);
or U9168 (N_9168,N_8843,N_8119);
and U9169 (N_9169,N_8732,N_8403);
nor U9170 (N_9170,N_8966,N_8720);
xor U9171 (N_9171,N_8896,N_8830);
nor U9172 (N_9172,N_8339,N_8919);
xor U9173 (N_9173,N_8473,N_8577);
or U9174 (N_9174,N_8058,N_8264);
nand U9175 (N_9175,N_8932,N_8396);
xor U9176 (N_9176,N_8636,N_8669);
nor U9177 (N_9177,N_8840,N_8618);
nand U9178 (N_9178,N_8198,N_8813);
nand U9179 (N_9179,N_8409,N_8682);
and U9180 (N_9180,N_8323,N_8373);
nor U9181 (N_9181,N_8776,N_8621);
nor U9182 (N_9182,N_8446,N_8981);
nor U9183 (N_9183,N_8104,N_8688);
and U9184 (N_9184,N_8284,N_8963);
or U9185 (N_9185,N_8549,N_8145);
nor U9186 (N_9186,N_8786,N_8393);
nand U9187 (N_9187,N_8784,N_8013);
nor U9188 (N_9188,N_8752,N_8433);
or U9189 (N_9189,N_8479,N_8379);
nor U9190 (N_9190,N_8458,N_8221);
nor U9191 (N_9191,N_8389,N_8229);
nor U9192 (N_9192,N_8415,N_8107);
nand U9193 (N_9193,N_8838,N_8825);
nor U9194 (N_9194,N_8550,N_8205);
and U9195 (N_9195,N_8617,N_8037);
and U9196 (N_9196,N_8974,N_8262);
nand U9197 (N_9197,N_8574,N_8344);
nand U9198 (N_9198,N_8606,N_8451);
and U9199 (N_9199,N_8442,N_8075);
nor U9200 (N_9200,N_8633,N_8716);
nor U9201 (N_9201,N_8420,N_8216);
nand U9202 (N_9202,N_8289,N_8969);
and U9203 (N_9203,N_8020,N_8498);
nor U9204 (N_9204,N_8312,N_8687);
nand U9205 (N_9205,N_8065,N_8569);
and U9206 (N_9206,N_8022,N_8132);
and U9207 (N_9207,N_8678,N_8902);
and U9208 (N_9208,N_8441,N_8091);
or U9209 (N_9209,N_8150,N_8097);
and U9210 (N_9210,N_8283,N_8531);
and U9211 (N_9211,N_8188,N_8660);
xnor U9212 (N_9212,N_8126,N_8613);
xnor U9213 (N_9213,N_8256,N_8831);
xnor U9214 (N_9214,N_8247,N_8962);
nand U9215 (N_9215,N_8303,N_8185);
nand U9216 (N_9216,N_8380,N_8362);
nand U9217 (N_9217,N_8865,N_8977);
nor U9218 (N_9218,N_8906,N_8985);
or U9219 (N_9219,N_8432,N_8288);
and U9220 (N_9220,N_8395,N_8012);
nand U9221 (N_9221,N_8858,N_8169);
or U9222 (N_9222,N_8704,N_8565);
and U9223 (N_9223,N_8639,N_8582);
nor U9224 (N_9224,N_8950,N_8341);
or U9225 (N_9225,N_8513,N_8390);
and U9226 (N_9226,N_8412,N_8546);
and U9227 (N_9227,N_8954,N_8192);
and U9228 (N_9228,N_8602,N_8098);
and U9229 (N_9229,N_8497,N_8818);
or U9230 (N_9230,N_8934,N_8159);
and U9231 (N_9231,N_8894,N_8116);
or U9232 (N_9232,N_8260,N_8506);
nand U9233 (N_9233,N_8080,N_8240);
nand U9234 (N_9234,N_8795,N_8106);
and U9235 (N_9235,N_8496,N_8972);
or U9236 (N_9236,N_8182,N_8570);
nor U9237 (N_9237,N_8321,N_8523);
and U9238 (N_9238,N_8092,N_8608);
nand U9239 (N_9239,N_8381,N_8591);
xor U9240 (N_9240,N_8793,N_8655);
or U9241 (N_9241,N_8504,N_8881);
nand U9242 (N_9242,N_8450,N_8233);
or U9243 (N_9243,N_8730,N_8468);
nand U9244 (N_9244,N_8510,N_8861);
and U9245 (N_9245,N_8354,N_8490);
nand U9246 (N_9246,N_8953,N_8105);
nor U9247 (N_9247,N_8237,N_8907);
or U9248 (N_9248,N_8774,N_8001);
and U9249 (N_9249,N_8769,N_8534);
nand U9250 (N_9250,N_8853,N_8689);
and U9251 (N_9251,N_8476,N_8828);
nand U9252 (N_9252,N_8002,N_8714);
xor U9253 (N_9253,N_8757,N_8957);
nand U9254 (N_9254,N_8125,N_8147);
nor U9255 (N_9255,N_8241,N_8649);
and U9256 (N_9256,N_8931,N_8043);
and U9257 (N_9257,N_8367,N_8135);
xor U9258 (N_9258,N_8672,N_8291);
and U9259 (N_9259,N_8692,N_8658);
xor U9260 (N_9260,N_8457,N_8194);
xnor U9261 (N_9261,N_8099,N_8837);
and U9262 (N_9262,N_8557,N_8643);
nor U9263 (N_9263,N_8242,N_8470);
nor U9264 (N_9264,N_8269,N_8815);
nand U9265 (N_9265,N_8960,N_8449);
nand U9266 (N_9266,N_8807,N_8285);
nand U9267 (N_9267,N_8895,N_8780);
nor U9268 (N_9268,N_8645,N_8236);
nor U9269 (N_9269,N_8768,N_8667);
and U9270 (N_9270,N_8234,N_8923);
or U9271 (N_9271,N_8090,N_8547);
xnor U9272 (N_9272,N_8154,N_8418);
or U9273 (N_9273,N_8517,N_8245);
or U9274 (N_9274,N_8595,N_8317);
or U9275 (N_9275,N_8061,N_8750);
nand U9276 (N_9276,N_8862,N_8224);
xnor U9277 (N_9277,N_8847,N_8140);
nand U9278 (N_9278,N_8875,N_8650);
nand U9279 (N_9279,N_8286,N_8761);
and U9280 (N_9280,N_8253,N_8202);
and U9281 (N_9281,N_8177,N_8007);
and U9282 (N_9282,N_8812,N_8980);
nand U9283 (N_9283,N_8179,N_8580);
nor U9284 (N_9284,N_8089,N_8252);
nor U9285 (N_9285,N_8841,N_8901);
xnor U9286 (N_9286,N_8128,N_8644);
xnor U9287 (N_9287,N_8456,N_8845);
and U9288 (N_9288,N_8475,N_8067);
and U9289 (N_9289,N_8027,N_8573);
nand U9290 (N_9290,N_8763,N_8383);
nor U9291 (N_9291,N_8676,N_8176);
or U9292 (N_9292,N_8300,N_8805);
nor U9293 (N_9293,N_8397,N_8791);
nand U9294 (N_9294,N_8425,N_8516);
and U9295 (N_9295,N_8100,N_8997);
xor U9296 (N_9296,N_8709,N_8318);
and U9297 (N_9297,N_8057,N_8915);
nand U9298 (N_9298,N_8160,N_8941);
or U9299 (N_9299,N_8215,N_8590);
nor U9300 (N_9300,N_8958,N_8583);
and U9301 (N_9301,N_8008,N_8899);
or U9302 (N_9302,N_8114,N_8651);
or U9303 (N_9303,N_8753,N_8789);
and U9304 (N_9304,N_8343,N_8993);
xor U9305 (N_9305,N_8619,N_8910);
or U9306 (N_9306,N_8788,N_8302);
and U9307 (N_9307,N_8987,N_8708);
nand U9308 (N_9308,N_8086,N_8469);
or U9309 (N_9309,N_8989,N_8153);
xor U9310 (N_9310,N_8054,N_8652);
xnor U9311 (N_9311,N_8244,N_8604);
or U9312 (N_9312,N_8142,N_8800);
and U9313 (N_9313,N_8824,N_8598);
nor U9314 (N_9314,N_8411,N_8746);
and U9315 (N_9315,N_8773,N_8220);
and U9316 (N_9316,N_8255,N_8047);
nor U9317 (N_9317,N_8874,N_8408);
xor U9318 (N_9318,N_8424,N_8266);
nor U9319 (N_9319,N_8440,N_8453);
nor U9320 (N_9320,N_8489,N_8820);
or U9321 (N_9321,N_8419,N_8422);
xor U9322 (N_9322,N_8701,N_8691);
nor U9323 (N_9323,N_8248,N_8968);
or U9324 (N_9324,N_8326,N_8095);
nor U9325 (N_9325,N_8209,N_8175);
nand U9326 (N_9326,N_8967,N_8782);
nand U9327 (N_9327,N_8930,N_8920);
nor U9328 (N_9328,N_8561,N_8197);
xor U9329 (N_9329,N_8448,N_8541);
xnor U9330 (N_9330,N_8671,N_8836);
nor U9331 (N_9331,N_8330,N_8528);
nand U9332 (N_9332,N_8543,N_8066);
xor U9333 (N_9333,N_8144,N_8888);
xnor U9334 (N_9334,N_8304,N_8413);
or U9335 (N_9335,N_8358,N_8554);
nor U9336 (N_9336,N_8365,N_8983);
nor U9337 (N_9337,N_8217,N_8952);
nor U9338 (N_9338,N_8431,N_8771);
and U9339 (N_9339,N_8797,N_8083);
nand U9340 (N_9340,N_8947,N_8576);
xnor U9341 (N_9341,N_8149,N_8635);
or U9342 (N_9342,N_8571,N_8046);
and U9343 (N_9343,N_8715,N_8662);
or U9344 (N_9344,N_8251,N_8823);
nor U9345 (N_9345,N_8904,N_8916);
or U9346 (N_9346,N_8308,N_8101);
nor U9347 (N_9347,N_8410,N_8596);
xnor U9348 (N_9348,N_8508,N_8405);
nand U9349 (N_9349,N_8279,N_8712);
or U9350 (N_9350,N_8530,N_8810);
xor U9351 (N_9351,N_8935,N_8937);
and U9352 (N_9352,N_8607,N_8052);
or U9353 (N_9353,N_8994,N_8605);
nor U9354 (N_9354,N_8511,N_8563);
nor U9355 (N_9355,N_8970,N_8749);
nand U9356 (N_9356,N_8259,N_8991);
xnor U9357 (N_9357,N_8088,N_8614);
xor U9358 (N_9358,N_8965,N_8278);
or U9359 (N_9359,N_8044,N_8759);
xnor U9360 (N_9360,N_8499,N_8665);
and U9361 (N_9361,N_8214,N_8725);
and U9362 (N_9362,N_8368,N_8204);
nand U9363 (N_9363,N_8477,N_8474);
or U9364 (N_9364,N_8444,N_8270);
xnor U9365 (N_9365,N_8136,N_8584);
and U9366 (N_9366,N_8465,N_8112);
and U9367 (N_9367,N_8035,N_8208);
or U9368 (N_9368,N_8933,N_8938);
nand U9369 (N_9369,N_8352,N_8298);
or U9370 (N_9370,N_8801,N_8664);
xor U9371 (N_9371,N_8559,N_8033);
nor U9372 (N_9372,N_8316,N_8232);
xnor U9373 (N_9373,N_8911,N_8377);
or U9374 (N_9374,N_8871,N_8045);
or U9375 (N_9375,N_8212,N_8386);
or U9376 (N_9376,N_8982,N_8751);
nand U9377 (N_9377,N_8603,N_8928);
or U9378 (N_9378,N_8562,N_8015);
nand U9379 (N_9379,N_8975,N_8071);
nor U9380 (N_9380,N_8984,N_8538);
nor U9381 (N_9381,N_8747,N_8029);
nand U9382 (N_9382,N_8471,N_8301);
nor U9383 (N_9383,N_8406,N_8346);
nand U9384 (N_9384,N_8319,N_8191);
and U9385 (N_9385,N_8014,N_8131);
nor U9386 (N_9386,N_8133,N_8366);
and U9387 (N_9387,N_8452,N_8623);
nor U9388 (N_9388,N_8767,N_8048);
nand U9389 (N_9389,N_8525,N_8735);
or U9390 (N_9390,N_8228,N_8654);
nand U9391 (N_9391,N_8371,N_8742);
or U9392 (N_9392,N_8796,N_8218);
xnor U9393 (N_9393,N_8437,N_8814);
nand U9394 (N_9394,N_8867,N_8537);
nor U9395 (N_9395,N_8158,N_8944);
nand U9396 (N_9396,N_8758,N_8548);
nor U9397 (N_9397,N_8491,N_8187);
and U9398 (N_9398,N_8295,N_8976);
and U9399 (N_9399,N_8893,N_8462);
nor U9400 (N_9400,N_8863,N_8338);
and U9401 (N_9401,N_8394,N_8404);
and U9402 (N_9402,N_8518,N_8705);
xor U9403 (N_9403,N_8971,N_8019);
nand U9404 (N_9404,N_8333,N_8909);
nand U9405 (N_9405,N_8350,N_8127);
nor U9406 (N_9406,N_8488,N_8168);
nor U9407 (N_9407,N_8275,N_8790);
nand U9408 (N_9408,N_8885,N_8178);
xor U9409 (N_9409,N_8706,N_8609);
xor U9410 (N_9410,N_8748,N_8505);
and U9411 (N_9411,N_8900,N_8762);
and U9412 (N_9412,N_8586,N_8094);
and U9413 (N_9413,N_8276,N_8113);
xor U9414 (N_9414,N_8961,N_8808);
and U9415 (N_9415,N_8579,N_8336);
nand U9416 (N_9416,N_8978,N_8309);
nor U9417 (N_9417,N_8811,N_8852);
or U9418 (N_9418,N_8359,N_8416);
nand U9419 (N_9419,N_8028,N_8694);
and U9420 (N_9420,N_8641,N_8943);
nand U9421 (N_9421,N_8542,N_8076);
and U9422 (N_9422,N_8211,N_8781);
or U9423 (N_9423,N_8860,N_8764);
nor U9424 (N_9424,N_8826,N_8755);
nand U9425 (N_9425,N_8555,N_8956);
nand U9426 (N_9426,N_8455,N_8124);
nand U9427 (N_9427,N_8201,N_8743);
nand U9428 (N_9428,N_8733,N_8164);
nand U9429 (N_9429,N_8544,N_8353);
nor U9430 (N_9430,N_8203,N_8873);
nand U9431 (N_9431,N_8273,N_8936);
or U9432 (N_9432,N_8521,N_8567);
or U9433 (N_9433,N_8988,N_8677);
and U9434 (N_9434,N_8927,N_8482);
nor U9435 (N_9435,N_8949,N_8995);
xnor U9436 (N_9436,N_8376,N_8430);
xor U9437 (N_9437,N_8670,N_8775);
nand U9438 (N_9438,N_8009,N_8799);
nand U9439 (N_9439,N_8560,N_8407);
or U9440 (N_9440,N_8536,N_8069);
nor U9441 (N_9441,N_8624,N_8575);
or U9442 (N_9442,N_8728,N_8435);
or U9443 (N_9443,N_8744,N_8585);
and U9444 (N_9444,N_8003,N_8834);
and U9445 (N_9445,N_8445,N_8032);
xor U9446 (N_9446,N_8207,N_8239);
and U9447 (N_9447,N_8509,N_8222);
nor U9448 (N_9448,N_8890,N_8777);
and U9449 (N_9449,N_8466,N_8391);
or U9450 (N_9450,N_8673,N_8710);
nand U9451 (N_9451,N_8460,N_8334);
nand U9452 (N_9452,N_8770,N_8173);
xnor U9453 (N_9453,N_8785,N_8392);
or U9454 (N_9454,N_8130,N_8123);
nor U9455 (N_9455,N_8638,N_8675);
or U9456 (N_9456,N_8056,N_8868);
nand U9457 (N_9457,N_8155,N_8698);
xnor U9458 (N_9458,N_8707,N_8802);
or U9459 (N_9459,N_8887,N_8942);
nand U9460 (N_9460,N_8074,N_8551);
and U9461 (N_9461,N_8593,N_8656);
nand U9462 (N_9462,N_8060,N_8897);
xnor U9463 (N_9463,N_8872,N_8648);
and U9464 (N_9464,N_8324,N_8068);
xor U9465 (N_9465,N_8084,N_8117);
and U9466 (N_9466,N_8322,N_8162);
or U9467 (N_9467,N_8566,N_8611);
nand U9468 (N_9468,N_8940,N_8879);
xor U9469 (N_9469,N_8443,N_8880);
xor U9470 (N_9470,N_8783,N_8737);
or U9471 (N_9471,N_8666,N_8072);
nand U9472 (N_9472,N_8115,N_8250);
nor U9473 (N_9473,N_8349,N_8313);
nor U9474 (N_9474,N_8039,N_8615);
nor U9475 (N_9475,N_8023,N_8331);
nor U9476 (N_9476,N_8822,N_8718);
nand U9477 (N_9477,N_8148,N_8724);
or U9478 (N_9478,N_8891,N_8835);
nand U9479 (N_9479,N_8181,N_8461);
nand U9480 (N_9480,N_8556,N_8502);
nand U9481 (N_9481,N_8632,N_8230);
nor U9482 (N_9482,N_8519,N_8402);
xor U9483 (N_9483,N_8851,N_8235);
xnor U9484 (N_9484,N_8305,N_8889);
nand U9485 (N_9485,N_8721,N_8745);
xor U9486 (N_9486,N_8817,N_8038);
and U9487 (N_9487,N_8572,N_8629);
nand U9488 (N_9488,N_8616,N_8464);
xor U9489 (N_9489,N_8342,N_8387);
or U9490 (N_9490,N_8051,N_8345);
nand U9491 (N_9491,N_8146,N_8372);
nor U9492 (N_9492,N_8417,N_8483);
and U9493 (N_9493,N_8492,N_8990);
or U9494 (N_9494,N_8378,N_8139);
nand U9495 (N_9495,N_8539,N_8883);
nor U9496 (N_9496,N_8998,N_8846);
xnor U9497 (N_9497,N_8647,N_8096);
nand U9498 (N_9498,N_8792,N_8501);
nor U9499 (N_9499,N_8948,N_8640);
nor U9500 (N_9500,N_8868,N_8477);
nor U9501 (N_9501,N_8265,N_8026);
and U9502 (N_9502,N_8086,N_8775);
nand U9503 (N_9503,N_8858,N_8363);
nand U9504 (N_9504,N_8615,N_8380);
and U9505 (N_9505,N_8698,N_8058);
or U9506 (N_9506,N_8565,N_8876);
and U9507 (N_9507,N_8659,N_8439);
nand U9508 (N_9508,N_8254,N_8288);
or U9509 (N_9509,N_8146,N_8289);
xor U9510 (N_9510,N_8222,N_8469);
nor U9511 (N_9511,N_8360,N_8886);
and U9512 (N_9512,N_8153,N_8413);
or U9513 (N_9513,N_8064,N_8514);
or U9514 (N_9514,N_8959,N_8080);
or U9515 (N_9515,N_8441,N_8128);
or U9516 (N_9516,N_8969,N_8221);
nand U9517 (N_9517,N_8771,N_8216);
and U9518 (N_9518,N_8550,N_8957);
nand U9519 (N_9519,N_8011,N_8959);
or U9520 (N_9520,N_8672,N_8964);
nor U9521 (N_9521,N_8864,N_8724);
and U9522 (N_9522,N_8002,N_8623);
xnor U9523 (N_9523,N_8106,N_8232);
nor U9524 (N_9524,N_8640,N_8465);
nand U9525 (N_9525,N_8252,N_8734);
nor U9526 (N_9526,N_8484,N_8777);
and U9527 (N_9527,N_8780,N_8705);
and U9528 (N_9528,N_8711,N_8970);
nor U9529 (N_9529,N_8508,N_8149);
nor U9530 (N_9530,N_8200,N_8724);
and U9531 (N_9531,N_8324,N_8688);
nor U9532 (N_9532,N_8569,N_8494);
nor U9533 (N_9533,N_8073,N_8297);
nand U9534 (N_9534,N_8523,N_8880);
nand U9535 (N_9535,N_8378,N_8946);
nand U9536 (N_9536,N_8416,N_8368);
and U9537 (N_9537,N_8662,N_8523);
or U9538 (N_9538,N_8048,N_8938);
and U9539 (N_9539,N_8292,N_8246);
or U9540 (N_9540,N_8938,N_8922);
nor U9541 (N_9541,N_8887,N_8847);
and U9542 (N_9542,N_8925,N_8998);
or U9543 (N_9543,N_8553,N_8439);
xor U9544 (N_9544,N_8883,N_8670);
or U9545 (N_9545,N_8893,N_8912);
and U9546 (N_9546,N_8197,N_8533);
and U9547 (N_9547,N_8412,N_8230);
or U9548 (N_9548,N_8878,N_8206);
or U9549 (N_9549,N_8438,N_8839);
or U9550 (N_9550,N_8362,N_8364);
nor U9551 (N_9551,N_8702,N_8845);
nor U9552 (N_9552,N_8039,N_8069);
and U9553 (N_9553,N_8721,N_8431);
or U9554 (N_9554,N_8629,N_8707);
nand U9555 (N_9555,N_8131,N_8247);
nor U9556 (N_9556,N_8983,N_8366);
or U9557 (N_9557,N_8731,N_8179);
nand U9558 (N_9558,N_8849,N_8173);
and U9559 (N_9559,N_8042,N_8152);
nand U9560 (N_9560,N_8355,N_8756);
nor U9561 (N_9561,N_8196,N_8607);
nand U9562 (N_9562,N_8631,N_8201);
and U9563 (N_9563,N_8467,N_8021);
nand U9564 (N_9564,N_8065,N_8250);
and U9565 (N_9565,N_8598,N_8024);
nand U9566 (N_9566,N_8657,N_8635);
nand U9567 (N_9567,N_8570,N_8711);
or U9568 (N_9568,N_8089,N_8114);
nand U9569 (N_9569,N_8694,N_8310);
or U9570 (N_9570,N_8543,N_8680);
nor U9571 (N_9571,N_8342,N_8270);
xor U9572 (N_9572,N_8436,N_8051);
nand U9573 (N_9573,N_8037,N_8041);
or U9574 (N_9574,N_8801,N_8689);
xor U9575 (N_9575,N_8649,N_8722);
nor U9576 (N_9576,N_8508,N_8072);
nand U9577 (N_9577,N_8257,N_8046);
and U9578 (N_9578,N_8754,N_8417);
nor U9579 (N_9579,N_8095,N_8750);
nor U9580 (N_9580,N_8262,N_8004);
nand U9581 (N_9581,N_8897,N_8357);
xnor U9582 (N_9582,N_8567,N_8148);
or U9583 (N_9583,N_8466,N_8272);
xnor U9584 (N_9584,N_8005,N_8538);
nor U9585 (N_9585,N_8712,N_8349);
or U9586 (N_9586,N_8373,N_8444);
nor U9587 (N_9587,N_8524,N_8315);
nor U9588 (N_9588,N_8805,N_8144);
or U9589 (N_9589,N_8243,N_8102);
and U9590 (N_9590,N_8806,N_8595);
nand U9591 (N_9591,N_8431,N_8777);
and U9592 (N_9592,N_8487,N_8744);
xnor U9593 (N_9593,N_8247,N_8398);
nor U9594 (N_9594,N_8964,N_8506);
nor U9595 (N_9595,N_8184,N_8066);
nand U9596 (N_9596,N_8317,N_8325);
or U9597 (N_9597,N_8138,N_8165);
nand U9598 (N_9598,N_8726,N_8271);
nand U9599 (N_9599,N_8413,N_8930);
nand U9600 (N_9600,N_8148,N_8444);
nor U9601 (N_9601,N_8287,N_8700);
nand U9602 (N_9602,N_8441,N_8078);
nor U9603 (N_9603,N_8469,N_8596);
and U9604 (N_9604,N_8814,N_8611);
and U9605 (N_9605,N_8865,N_8741);
and U9606 (N_9606,N_8463,N_8741);
xnor U9607 (N_9607,N_8124,N_8652);
nor U9608 (N_9608,N_8700,N_8861);
nand U9609 (N_9609,N_8106,N_8739);
nor U9610 (N_9610,N_8970,N_8892);
and U9611 (N_9611,N_8977,N_8077);
nand U9612 (N_9612,N_8624,N_8517);
nor U9613 (N_9613,N_8474,N_8765);
nor U9614 (N_9614,N_8910,N_8545);
xor U9615 (N_9615,N_8725,N_8668);
and U9616 (N_9616,N_8500,N_8825);
nand U9617 (N_9617,N_8542,N_8818);
nand U9618 (N_9618,N_8076,N_8530);
and U9619 (N_9619,N_8366,N_8180);
or U9620 (N_9620,N_8156,N_8218);
nor U9621 (N_9621,N_8539,N_8178);
and U9622 (N_9622,N_8148,N_8737);
nor U9623 (N_9623,N_8155,N_8638);
nand U9624 (N_9624,N_8041,N_8152);
and U9625 (N_9625,N_8813,N_8298);
nor U9626 (N_9626,N_8327,N_8254);
nor U9627 (N_9627,N_8993,N_8723);
nor U9628 (N_9628,N_8553,N_8249);
or U9629 (N_9629,N_8588,N_8089);
and U9630 (N_9630,N_8121,N_8438);
nand U9631 (N_9631,N_8501,N_8908);
or U9632 (N_9632,N_8526,N_8926);
and U9633 (N_9633,N_8804,N_8475);
or U9634 (N_9634,N_8018,N_8263);
or U9635 (N_9635,N_8721,N_8459);
or U9636 (N_9636,N_8955,N_8276);
nor U9637 (N_9637,N_8435,N_8495);
or U9638 (N_9638,N_8756,N_8831);
or U9639 (N_9639,N_8918,N_8928);
and U9640 (N_9640,N_8569,N_8042);
nor U9641 (N_9641,N_8462,N_8953);
nor U9642 (N_9642,N_8378,N_8502);
nand U9643 (N_9643,N_8052,N_8366);
nor U9644 (N_9644,N_8056,N_8124);
nor U9645 (N_9645,N_8214,N_8171);
and U9646 (N_9646,N_8045,N_8617);
and U9647 (N_9647,N_8096,N_8453);
or U9648 (N_9648,N_8059,N_8923);
and U9649 (N_9649,N_8932,N_8077);
nand U9650 (N_9650,N_8676,N_8904);
nor U9651 (N_9651,N_8734,N_8183);
or U9652 (N_9652,N_8976,N_8109);
or U9653 (N_9653,N_8277,N_8627);
nand U9654 (N_9654,N_8863,N_8913);
nor U9655 (N_9655,N_8440,N_8185);
nand U9656 (N_9656,N_8248,N_8009);
and U9657 (N_9657,N_8312,N_8268);
xnor U9658 (N_9658,N_8141,N_8194);
or U9659 (N_9659,N_8692,N_8905);
nor U9660 (N_9660,N_8493,N_8624);
nand U9661 (N_9661,N_8216,N_8128);
nand U9662 (N_9662,N_8721,N_8738);
and U9663 (N_9663,N_8439,N_8648);
or U9664 (N_9664,N_8525,N_8140);
xnor U9665 (N_9665,N_8078,N_8594);
and U9666 (N_9666,N_8509,N_8130);
or U9667 (N_9667,N_8681,N_8391);
nor U9668 (N_9668,N_8116,N_8323);
nor U9669 (N_9669,N_8414,N_8494);
nor U9670 (N_9670,N_8481,N_8560);
xor U9671 (N_9671,N_8744,N_8650);
nand U9672 (N_9672,N_8375,N_8370);
or U9673 (N_9673,N_8079,N_8961);
nor U9674 (N_9674,N_8136,N_8108);
nand U9675 (N_9675,N_8687,N_8546);
or U9676 (N_9676,N_8340,N_8747);
or U9677 (N_9677,N_8915,N_8313);
nand U9678 (N_9678,N_8948,N_8821);
and U9679 (N_9679,N_8495,N_8211);
xnor U9680 (N_9680,N_8146,N_8432);
nor U9681 (N_9681,N_8495,N_8779);
or U9682 (N_9682,N_8696,N_8044);
or U9683 (N_9683,N_8559,N_8543);
nand U9684 (N_9684,N_8387,N_8378);
nor U9685 (N_9685,N_8191,N_8970);
xnor U9686 (N_9686,N_8913,N_8064);
nand U9687 (N_9687,N_8722,N_8549);
nor U9688 (N_9688,N_8992,N_8216);
nor U9689 (N_9689,N_8115,N_8461);
or U9690 (N_9690,N_8093,N_8556);
or U9691 (N_9691,N_8984,N_8099);
nand U9692 (N_9692,N_8425,N_8707);
or U9693 (N_9693,N_8898,N_8398);
or U9694 (N_9694,N_8474,N_8317);
or U9695 (N_9695,N_8172,N_8566);
nand U9696 (N_9696,N_8238,N_8261);
nor U9697 (N_9697,N_8833,N_8717);
nand U9698 (N_9698,N_8817,N_8144);
and U9699 (N_9699,N_8778,N_8720);
and U9700 (N_9700,N_8104,N_8843);
and U9701 (N_9701,N_8618,N_8366);
nand U9702 (N_9702,N_8654,N_8421);
or U9703 (N_9703,N_8122,N_8914);
xor U9704 (N_9704,N_8997,N_8298);
or U9705 (N_9705,N_8224,N_8668);
and U9706 (N_9706,N_8223,N_8120);
nor U9707 (N_9707,N_8901,N_8713);
nand U9708 (N_9708,N_8788,N_8621);
or U9709 (N_9709,N_8599,N_8964);
xor U9710 (N_9710,N_8413,N_8465);
or U9711 (N_9711,N_8130,N_8589);
nor U9712 (N_9712,N_8215,N_8122);
or U9713 (N_9713,N_8921,N_8283);
and U9714 (N_9714,N_8603,N_8707);
and U9715 (N_9715,N_8501,N_8139);
and U9716 (N_9716,N_8631,N_8683);
nand U9717 (N_9717,N_8402,N_8977);
or U9718 (N_9718,N_8687,N_8624);
or U9719 (N_9719,N_8670,N_8459);
nor U9720 (N_9720,N_8766,N_8975);
nor U9721 (N_9721,N_8853,N_8229);
xor U9722 (N_9722,N_8128,N_8163);
xnor U9723 (N_9723,N_8312,N_8062);
nor U9724 (N_9724,N_8957,N_8444);
nand U9725 (N_9725,N_8447,N_8182);
nand U9726 (N_9726,N_8221,N_8157);
nor U9727 (N_9727,N_8488,N_8241);
and U9728 (N_9728,N_8791,N_8916);
or U9729 (N_9729,N_8322,N_8170);
nor U9730 (N_9730,N_8919,N_8235);
nor U9731 (N_9731,N_8946,N_8032);
nor U9732 (N_9732,N_8863,N_8337);
or U9733 (N_9733,N_8032,N_8088);
or U9734 (N_9734,N_8912,N_8220);
or U9735 (N_9735,N_8845,N_8354);
nand U9736 (N_9736,N_8630,N_8356);
nand U9737 (N_9737,N_8631,N_8221);
and U9738 (N_9738,N_8397,N_8741);
or U9739 (N_9739,N_8417,N_8562);
nor U9740 (N_9740,N_8962,N_8480);
or U9741 (N_9741,N_8566,N_8000);
or U9742 (N_9742,N_8639,N_8642);
nor U9743 (N_9743,N_8053,N_8870);
nor U9744 (N_9744,N_8006,N_8887);
or U9745 (N_9745,N_8351,N_8030);
nor U9746 (N_9746,N_8182,N_8500);
nor U9747 (N_9747,N_8810,N_8850);
nor U9748 (N_9748,N_8002,N_8046);
nand U9749 (N_9749,N_8759,N_8395);
nor U9750 (N_9750,N_8866,N_8537);
or U9751 (N_9751,N_8929,N_8248);
nand U9752 (N_9752,N_8837,N_8855);
or U9753 (N_9753,N_8707,N_8805);
and U9754 (N_9754,N_8058,N_8502);
or U9755 (N_9755,N_8046,N_8480);
nand U9756 (N_9756,N_8355,N_8482);
nand U9757 (N_9757,N_8707,N_8667);
xnor U9758 (N_9758,N_8917,N_8644);
and U9759 (N_9759,N_8521,N_8849);
or U9760 (N_9760,N_8993,N_8772);
nor U9761 (N_9761,N_8307,N_8353);
nand U9762 (N_9762,N_8212,N_8959);
and U9763 (N_9763,N_8964,N_8747);
or U9764 (N_9764,N_8923,N_8657);
nand U9765 (N_9765,N_8285,N_8936);
nor U9766 (N_9766,N_8282,N_8725);
nand U9767 (N_9767,N_8044,N_8730);
xor U9768 (N_9768,N_8452,N_8700);
or U9769 (N_9769,N_8379,N_8242);
or U9770 (N_9770,N_8805,N_8538);
nor U9771 (N_9771,N_8635,N_8603);
nor U9772 (N_9772,N_8888,N_8576);
and U9773 (N_9773,N_8536,N_8060);
nand U9774 (N_9774,N_8572,N_8103);
xnor U9775 (N_9775,N_8869,N_8731);
and U9776 (N_9776,N_8802,N_8491);
or U9777 (N_9777,N_8631,N_8064);
or U9778 (N_9778,N_8744,N_8649);
or U9779 (N_9779,N_8796,N_8013);
nor U9780 (N_9780,N_8726,N_8296);
nand U9781 (N_9781,N_8114,N_8261);
and U9782 (N_9782,N_8548,N_8679);
nor U9783 (N_9783,N_8818,N_8450);
nand U9784 (N_9784,N_8368,N_8840);
nand U9785 (N_9785,N_8798,N_8836);
nor U9786 (N_9786,N_8028,N_8656);
nor U9787 (N_9787,N_8266,N_8478);
nand U9788 (N_9788,N_8306,N_8507);
or U9789 (N_9789,N_8882,N_8188);
nor U9790 (N_9790,N_8892,N_8315);
nand U9791 (N_9791,N_8497,N_8803);
nor U9792 (N_9792,N_8954,N_8174);
or U9793 (N_9793,N_8768,N_8211);
nor U9794 (N_9794,N_8244,N_8211);
xnor U9795 (N_9795,N_8813,N_8946);
and U9796 (N_9796,N_8518,N_8961);
or U9797 (N_9797,N_8907,N_8410);
nor U9798 (N_9798,N_8818,N_8649);
or U9799 (N_9799,N_8403,N_8494);
nand U9800 (N_9800,N_8253,N_8411);
nor U9801 (N_9801,N_8386,N_8223);
and U9802 (N_9802,N_8168,N_8864);
and U9803 (N_9803,N_8176,N_8184);
and U9804 (N_9804,N_8453,N_8831);
xor U9805 (N_9805,N_8096,N_8147);
and U9806 (N_9806,N_8737,N_8948);
xnor U9807 (N_9807,N_8313,N_8710);
nor U9808 (N_9808,N_8236,N_8992);
nand U9809 (N_9809,N_8432,N_8613);
nand U9810 (N_9810,N_8011,N_8224);
nand U9811 (N_9811,N_8820,N_8347);
nand U9812 (N_9812,N_8400,N_8391);
or U9813 (N_9813,N_8752,N_8195);
nand U9814 (N_9814,N_8830,N_8280);
nand U9815 (N_9815,N_8016,N_8236);
nand U9816 (N_9816,N_8386,N_8533);
xor U9817 (N_9817,N_8000,N_8491);
nand U9818 (N_9818,N_8789,N_8882);
nor U9819 (N_9819,N_8219,N_8424);
nand U9820 (N_9820,N_8129,N_8292);
nand U9821 (N_9821,N_8664,N_8304);
and U9822 (N_9822,N_8736,N_8894);
nand U9823 (N_9823,N_8092,N_8775);
and U9824 (N_9824,N_8738,N_8417);
nor U9825 (N_9825,N_8392,N_8288);
and U9826 (N_9826,N_8415,N_8607);
and U9827 (N_9827,N_8794,N_8668);
and U9828 (N_9828,N_8197,N_8482);
or U9829 (N_9829,N_8898,N_8276);
or U9830 (N_9830,N_8492,N_8878);
nor U9831 (N_9831,N_8768,N_8969);
and U9832 (N_9832,N_8242,N_8343);
or U9833 (N_9833,N_8195,N_8311);
nand U9834 (N_9834,N_8126,N_8474);
nor U9835 (N_9835,N_8312,N_8704);
nor U9836 (N_9836,N_8088,N_8702);
and U9837 (N_9837,N_8426,N_8270);
nand U9838 (N_9838,N_8553,N_8590);
xnor U9839 (N_9839,N_8012,N_8528);
nor U9840 (N_9840,N_8338,N_8109);
nor U9841 (N_9841,N_8173,N_8818);
and U9842 (N_9842,N_8202,N_8845);
nand U9843 (N_9843,N_8274,N_8393);
or U9844 (N_9844,N_8642,N_8326);
nand U9845 (N_9845,N_8439,N_8134);
nor U9846 (N_9846,N_8960,N_8645);
nor U9847 (N_9847,N_8138,N_8843);
and U9848 (N_9848,N_8247,N_8582);
and U9849 (N_9849,N_8541,N_8576);
and U9850 (N_9850,N_8487,N_8452);
or U9851 (N_9851,N_8098,N_8154);
nand U9852 (N_9852,N_8419,N_8297);
or U9853 (N_9853,N_8384,N_8905);
and U9854 (N_9854,N_8938,N_8059);
nand U9855 (N_9855,N_8784,N_8572);
or U9856 (N_9856,N_8612,N_8684);
or U9857 (N_9857,N_8754,N_8678);
nand U9858 (N_9858,N_8288,N_8206);
or U9859 (N_9859,N_8208,N_8268);
nand U9860 (N_9860,N_8973,N_8351);
and U9861 (N_9861,N_8122,N_8348);
and U9862 (N_9862,N_8279,N_8921);
and U9863 (N_9863,N_8507,N_8736);
nand U9864 (N_9864,N_8946,N_8518);
or U9865 (N_9865,N_8094,N_8723);
or U9866 (N_9866,N_8195,N_8998);
nand U9867 (N_9867,N_8404,N_8047);
nor U9868 (N_9868,N_8946,N_8341);
nor U9869 (N_9869,N_8651,N_8561);
and U9870 (N_9870,N_8820,N_8952);
and U9871 (N_9871,N_8371,N_8663);
xor U9872 (N_9872,N_8796,N_8678);
nor U9873 (N_9873,N_8882,N_8475);
xor U9874 (N_9874,N_8946,N_8173);
and U9875 (N_9875,N_8033,N_8158);
nand U9876 (N_9876,N_8752,N_8079);
nand U9877 (N_9877,N_8836,N_8114);
or U9878 (N_9878,N_8164,N_8749);
and U9879 (N_9879,N_8658,N_8300);
and U9880 (N_9880,N_8732,N_8952);
nor U9881 (N_9881,N_8897,N_8054);
xnor U9882 (N_9882,N_8051,N_8815);
and U9883 (N_9883,N_8420,N_8448);
and U9884 (N_9884,N_8006,N_8649);
nor U9885 (N_9885,N_8323,N_8789);
nor U9886 (N_9886,N_8114,N_8258);
nand U9887 (N_9887,N_8083,N_8321);
and U9888 (N_9888,N_8225,N_8944);
nand U9889 (N_9889,N_8767,N_8230);
nand U9890 (N_9890,N_8210,N_8097);
nor U9891 (N_9891,N_8617,N_8325);
nor U9892 (N_9892,N_8704,N_8316);
and U9893 (N_9893,N_8785,N_8273);
nand U9894 (N_9894,N_8028,N_8109);
or U9895 (N_9895,N_8756,N_8692);
nand U9896 (N_9896,N_8756,N_8588);
nand U9897 (N_9897,N_8994,N_8418);
and U9898 (N_9898,N_8693,N_8351);
nand U9899 (N_9899,N_8056,N_8038);
or U9900 (N_9900,N_8498,N_8155);
nor U9901 (N_9901,N_8366,N_8607);
or U9902 (N_9902,N_8025,N_8164);
or U9903 (N_9903,N_8862,N_8784);
and U9904 (N_9904,N_8027,N_8270);
nor U9905 (N_9905,N_8112,N_8503);
xor U9906 (N_9906,N_8106,N_8488);
nor U9907 (N_9907,N_8416,N_8070);
or U9908 (N_9908,N_8110,N_8485);
and U9909 (N_9909,N_8109,N_8631);
and U9910 (N_9910,N_8976,N_8409);
nor U9911 (N_9911,N_8857,N_8258);
or U9912 (N_9912,N_8710,N_8908);
nor U9913 (N_9913,N_8355,N_8508);
xnor U9914 (N_9914,N_8741,N_8825);
or U9915 (N_9915,N_8865,N_8742);
xnor U9916 (N_9916,N_8929,N_8496);
and U9917 (N_9917,N_8622,N_8994);
nor U9918 (N_9918,N_8390,N_8378);
or U9919 (N_9919,N_8913,N_8085);
nand U9920 (N_9920,N_8671,N_8894);
nand U9921 (N_9921,N_8403,N_8054);
and U9922 (N_9922,N_8594,N_8154);
xnor U9923 (N_9923,N_8449,N_8308);
nand U9924 (N_9924,N_8411,N_8987);
and U9925 (N_9925,N_8735,N_8172);
nand U9926 (N_9926,N_8569,N_8625);
and U9927 (N_9927,N_8937,N_8936);
and U9928 (N_9928,N_8128,N_8973);
nand U9929 (N_9929,N_8242,N_8797);
nor U9930 (N_9930,N_8365,N_8692);
nor U9931 (N_9931,N_8967,N_8641);
or U9932 (N_9932,N_8325,N_8926);
and U9933 (N_9933,N_8350,N_8564);
and U9934 (N_9934,N_8491,N_8242);
xnor U9935 (N_9935,N_8094,N_8030);
nand U9936 (N_9936,N_8342,N_8895);
or U9937 (N_9937,N_8074,N_8901);
nand U9938 (N_9938,N_8796,N_8422);
nand U9939 (N_9939,N_8969,N_8215);
and U9940 (N_9940,N_8268,N_8798);
nand U9941 (N_9941,N_8425,N_8713);
and U9942 (N_9942,N_8779,N_8446);
and U9943 (N_9943,N_8656,N_8142);
nor U9944 (N_9944,N_8223,N_8359);
nand U9945 (N_9945,N_8355,N_8497);
or U9946 (N_9946,N_8195,N_8624);
and U9947 (N_9947,N_8770,N_8735);
or U9948 (N_9948,N_8000,N_8972);
nor U9949 (N_9949,N_8946,N_8392);
xnor U9950 (N_9950,N_8565,N_8538);
and U9951 (N_9951,N_8417,N_8449);
and U9952 (N_9952,N_8971,N_8390);
and U9953 (N_9953,N_8658,N_8860);
nor U9954 (N_9954,N_8031,N_8608);
and U9955 (N_9955,N_8415,N_8779);
nand U9956 (N_9956,N_8108,N_8629);
or U9957 (N_9957,N_8533,N_8651);
or U9958 (N_9958,N_8329,N_8058);
or U9959 (N_9959,N_8940,N_8703);
or U9960 (N_9960,N_8932,N_8222);
nand U9961 (N_9961,N_8420,N_8531);
nor U9962 (N_9962,N_8184,N_8637);
nand U9963 (N_9963,N_8394,N_8015);
or U9964 (N_9964,N_8887,N_8891);
nor U9965 (N_9965,N_8063,N_8231);
and U9966 (N_9966,N_8241,N_8139);
nor U9967 (N_9967,N_8361,N_8991);
xor U9968 (N_9968,N_8672,N_8534);
nand U9969 (N_9969,N_8617,N_8808);
nand U9970 (N_9970,N_8126,N_8660);
nand U9971 (N_9971,N_8287,N_8486);
nor U9972 (N_9972,N_8829,N_8520);
nand U9973 (N_9973,N_8143,N_8711);
nand U9974 (N_9974,N_8462,N_8626);
nor U9975 (N_9975,N_8988,N_8146);
nand U9976 (N_9976,N_8009,N_8051);
xnor U9977 (N_9977,N_8913,N_8625);
nand U9978 (N_9978,N_8789,N_8144);
or U9979 (N_9979,N_8455,N_8475);
nor U9980 (N_9980,N_8626,N_8867);
or U9981 (N_9981,N_8895,N_8877);
nand U9982 (N_9982,N_8635,N_8547);
and U9983 (N_9983,N_8236,N_8949);
nand U9984 (N_9984,N_8160,N_8204);
xor U9985 (N_9985,N_8633,N_8774);
nor U9986 (N_9986,N_8635,N_8110);
or U9987 (N_9987,N_8245,N_8987);
nand U9988 (N_9988,N_8812,N_8154);
nor U9989 (N_9989,N_8714,N_8973);
or U9990 (N_9990,N_8312,N_8102);
nor U9991 (N_9991,N_8180,N_8410);
nand U9992 (N_9992,N_8528,N_8464);
nand U9993 (N_9993,N_8460,N_8303);
or U9994 (N_9994,N_8925,N_8708);
nand U9995 (N_9995,N_8986,N_8251);
nand U9996 (N_9996,N_8633,N_8927);
nand U9997 (N_9997,N_8387,N_8058);
or U9998 (N_9998,N_8093,N_8324);
or U9999 (N_9999,N_8296,N_8004);
or UO_0 (O_0,N_9938,N_9659);
nor UO_1 (O_1,N_9974,N_9109);
or UO_2 (O_2,N_9627,N_9143);
or UO_3 (O_3,N_9475,N_9604);
or UO_4 (O_4,N_9149,N_9590);
nand UO_5 (O_5,N_9963,N_9424);
nand UO_6 (O_6,N_9298,N_9207);
nor UO_7 (O_7,N_9849,N_9618);
and UO_8 (O_8,N_9168,N_9610);
or UO_9 (O_9,N_9321,N_9570);
and UO_10 (O_10,N_9024,N_9259);
xor UO_11 (O_11,N_9546,N_9383);
xnor UO_12 (O_12,N_9529,N_9930);
nor UO_13 (O_13,N_9134,N_9809);
and UO_14 (O_14,N_9851,N_9791);
nor UO_15 (O_15,N_9885,N_9036);
nand UO_16 (O_16,N_9421,N_9380);
and UO_17 (O_17,N_9758,N_9234);
and UO_18 (O_18,N_9718,N_9931);
and UO_19 (O_19,N_9883,N_9429);
nor UO_20 (O_20,N_9446,N_9281);
nand UO_21 (O_21,N_9169,N_9616);
and UO_22 (O_22,N_9348,N_9318);
and UO_23 (O_23,N_9991,N_9669);
nor UO_24 (O_24,N_9064,N_9801);
xor UO_25 (O_25,N_9743,N_9932);
nor UO_26 (O_26,N_9273,N_9910);
nor UO_27 (O_27,N_9629,N_9969);
or UO_28 (O_28,N_9994,N_9263);
or UO_29 (O_29,N_9157,N_9470);
or UO_30 (O_30,N_9903,N_9844);
nor UO_31 (O_31,N_9527,N_9017);
nor UO_32 (O_32,N_9648,N_9120);
xnor UO_33 (O_33,N_9661,N_9432);
xnor UO_34 (O_34,N_9807,N_9401);
nand UO_35 (O_35,N_9044,N_9006);
nand UO_36 (O_36,N_9127,N_9637);
or UO_37 (O_37,N_9272,N_9726);
nor UO_38 (O_38,N_9768,N_9238);
and UO_39 (O_39,N_9331,N_9685);
and UO_40 (O_40,N_9247,N_9598);
nor UO_41 (O_41,N_9816,N_9116);
nor UO_42 (O_42,N_9735,N_9536);
or UO_43 (O_43,N_9206,N_9955);
xor UO_44 (O_44,N_9379,N_9093);
nor UO_45 (O_45,N_9395,N_9534);
or UO_46 (O_46,N_9047,N_9454);
or UO_47 (O_47,N_9684,N_9130);
or UO_48 (O_48,N_9069,N_9192);
nor UO_49 (O_49,N_9804,N_9524);
xor UO_50 (O_50,N_9092,N_9794);
nor UO_51 (O_51,N_9004,N_9893);
and UO_52 (O_52,N_9439,N_9222);
or UO_53 (O_53,N_9276,N_9205);
or UO_54 (O_54,N_9811,N_9753);
and UO_55 (O_55,N_9392,N_9232);
nor UO_56 (O_56,N_9566,N_9463);
or UO_57 (O_57,N_9803,N_9547);
nand UO_58 (O_58,N_9900,N_9191);
nand UO_59 (O_59,N_9246,N_9831);
or UO_60 (O_60,N_9407,N_9688);
or UO_61 (O_61,N_9625,N_9808);
or UO_62 (O_62,N_9389,N_9950);
or UO_63 (O_63,N_9320,N_9757);
nand UO_64 (O_64,N_9196,N_9738);
and UO_65 (O_65,N_9133,N_9488);
and UO_66 (O_66,N_9698,N_9022);
and UO_67 (O_67,N_9484,N_9248);
nand UO_68 (O_68,N_9382,N_9179);
nor UO_69 (O_69,N_9736,N_9881);
nand UO_70 (O_70,N_9655,N_9282);
and UO_71 (O_71,N_9198,N_9864);
nand UO_72 (O_72,N_9554,N_9819);
nand UO_73 (O_73,N_9433,N_9613);
nand UO_74 (O_74,N_9345,N_9194);
xnor UO_75 (O_75,N_9100,N_9413);
or UO_76 (O_76,N_9430,N_9761);
nor UO_77 (O_77,N_9905,N_9227);
nor UO_78 (O_78,N_9099,N_9894);
nor UO_79 (O_79,N_9887,N_9557);
nor UO_80 (O_80,N_9663,N_9142);
nand UO_81 (O_81,N_9215,N_9280);
nand UO_82 (O_82,N_9593,N_9465);
or UO_83 (O_83,N_9519,N_9285);
and UO_84 (O_84,N_9654,N_9474);
nor UO_85 (O_85,N_9733,N_9986);
xor UO_86 (O_86,N_9747,N_9362);
nand UO_87 (O_87,N_9843,N_9633);
nand UO_88 (O_88,N_9029,N_9140);
or UO_89 (O_89,N_9967,N_9602);
nand UO_90 (O_90,N_9845,N_9094);
nor UO_91 (O_91,N_9796,N_9213);
nand UO_92 (O_92,N_9390,N_9649);
nor UO_93 (O_93,N_9652,N_9533);
nand UO_94 (O_94,N_9152,N_9219);
nand UO_95 (O_95,N_9256,N_9328);
or UO_96 (O_96,N_9708,N_9115);
nor UO_97 (O_97,N_9104,N_9060);
nand UO_98 (O_98,N_9119,N_9783);
and UO_99 (O_99,N_9568,N_9224);
and UO_100 (O_100,N_9335,N_9946);
and UO_101 (O_101,N_9854,N_9707);
and UO_102 (O_102,N_9396,N_9358);
xnor UO_103 (O_103,N_9971,N_9990);
nor UO_104 (O_104,N_9098,N_9691);
and UO_105 (O_105,N_9371,N_9672);
or UO_106 (O_106,N_9692,N_9287);
and UO_107 (O_107,N_9216,N_9283);
nor UO_108 (O_108,N_9765,N_9599);
nand UO_109 (O_109,N_9727,N_9666);
nand UO_110 (O_110,N_9680,N_9428);
nor UO_111 (O_111,N_9049,N_9875);
xor UO_112 (O_112,N_9309,N_9585);
or UO_113 (O_113,N_9630,N_9861);
or UO_114 (O_114,N_9010,N_9609);
or UO_115 (O_115,N_9715,N_9805);
nor UO_116 (O_116,N_9769,N_9138);
and UO_117 (O_117,N_9236,N_9072);
nand UO_118 (O_118,N_9467,N_9787);
and UO_119 (O_119,N_9916,N_9958);
or UO_120 (O_120,N_9068,N_9552);
xor UO_121 (O_121,N_9079,N_9520);
xor UO_122 (O_122,N_9813,N_9989);
or UO_123 (O_123,N_9908,N_9890);
nor UO_124 (O_124,N_9458,N_9344);
nor UO_125 (O_125,N_9589,N_9001);
and UO_126 (O_126,N_9487,N_9151);
nand UO_127 (O_127,N_9173,N_9944);
and UO_128 (O_128,N_9180,N_9834);
nor UO_129 (O_129,N_9026,N_9634);
or UO_130 (O_130,N_9776,N_9514);
nor UO_131 (O_131,N_9499,N_9928);
or UO_132 (O_132,N_9640,N_9110);
and UO_133 (O_133,N_9300,N_9830);
or UO_134 (O_134,N_9435,N_9892);
nand UO_135 (O_135,N_9306,N_9737);
or UO_136 (O_136,N_9876,N_9538);
or UO_137 (O_137,N_9444,N_9373);
and UO_138 (O_138,N_9644,N_9954);
or UO_139 (O_139,N_9150,N_9048);
or UO_140 (O_140,N_9495,N_9440);
and UO_141 (O_141,N_9919,N_9218);
and UO_142 (O_142,N_9906,N_9132);
nor UO_143 (O_143,N_9752,N_9453);
or UO_144 (O_144,N_9178,N_9709);
nand UO_145 (O_145,N_9159,N_9711);
nand UO_146 (O_146,N_9891,N_9667);
nor UO_147 (O_147,N_9107,N_9106);
nor UO_148 (O_148,N_9292,N_9089);
and UO_149 (O_149,N_9387,N_9720);
nor UO_150 (O_150,N_9869,N_9350);
nor UO_151 (O_151,N_9645,N_9368);
xnor UO_152 (O_152,N_9375,N_9673);
nand UO_153 (O_153,N_9491,N_9541);
or UO_154 (O_154,N_9310,N_9087);
nand UO_155 (O_155,N_9393,N_9793);
or UO_156 (O_156,N_9105,N_9493);
and UO_157 (O_157,N_9122,N_9330);
nor UO_158 (O_158,N_9795,N_9798);
and UO_159 (O_159,N_9199,N_9785);
xnor UO_160 (O_160,N_9459,N_9391);
xor UO_161 (O_161,N_9983,N_9777);
or UO_162 (O_162,N_9638,N_9927);
nand UO_163 (O_163,N_9739,N_9347);
and UO_164 (O_164,N_9114,N_9307);
nor UO_165 (O_165,N_9647,N_9681);
xor UO_166 (O_166,N_9510,N_9355);
and UO_167 (O_167,N_9577,N_9278);
and UO_168 (O_168,N_9741,N_9126);
or UO_169 (O_169,N_9690,N_9066);
xnor UO_170 (O_170,N_9865,N_9003);
nand UO_171 (O_171,N_9102,N_9405);
xnor UO_172 (O_172,N_9624,N_9055);
and UO_173 (O_173,N_9501,N_9964);
xor UO_174 (O_174,N_9472,N_9270);
or UO_175 (O_175,N_9118,N_9592);
or UO_176 (O_176,N_9981,N_9399);
nor UO_177 (O_177,N_9154,N_9235);
nand UO_178 (O_178,N_9548,N_9935);
nor UO_179 (O_179,N_9351,N_9337);
nand UO_180 (O_180,N_9483,N_9223);
xor UO_181 (O_181,N_9365,N_9515);
nand UO_182 (O_182,N_9978,N_9852);
or UO_183 (O_183,N_9188,N_9045);
xor UO_184 (O_184,N_9177,N_9160);
and UO_185 (O_185,N_9023,N_9131);
xor UO_186 (O_186,N_9578,N_9124);
nor UO_187 (O_187,N_9556,N_9790);
and UO_188 (O_188,N_9305,N_9677);
nand UO_189 (O_189,N_9972,N_9564);
nor UO_190 (O_190,N_9586,N_9897);
nand UO_191 (O_191,N_9918,N_9961);
or UO_192 (O_192,N_9540,N_9823);
nand UO_193 (O_193,N_9810,N_9418);
or UO_194 (O_194,N_9423,N_9940);
and UO_195 (O_195,N_9740,N_9988);
nand UO_196 (O_196,N_9880,N_9898);
and UO_197 (O_197,N_9144,N_9657);
and UO_198 (O_198,N_9689,N_9101);
and UO_199 (O_199,N_9855,N_9075);
and UO_200 (O_200,N_9388,N_9301);
nand UO_201 (O_201,N_9296,N_9749);
and UO_202 (O_202,N_9806,N_9706);
and UO_203 (O_203,N_9063,N_9748);
xnor UO_204 (O_204,N_9203,N_9859);
nor UO_205 (O_205,N_9195,N_9770);
nand UO_206 (O_206,N_9056,N_9125);
nand UO_207 (O_207,N_9032,N_9694);
nand UO_208 (O_208,N_9999,N_9080);
and UO_209 (O_209,N_9582,N_9584);
nor UO_210 (O_210,N_9754,N_9966);
or UO_211 (O_211,N_9204,N_9703);
xnor UO_212 (O_212,N_9477,N_9948);
nand UO_213 (O_213,N_9530,N_9286);
or UO_214 (O_214,N_9512,N_9266);
xor UO_215 (O_215,N_9612,N_9426);
and UO_216 (O_216,N_9136,N_9090);
or UO_217 (O_217,N_9818,N_9549);
and UO_218 (O_218,N_9265,N_9658);
nor UO_219 (O_219,N_9028,N_9394);
xnor UO_220 (O_220,N_9000,N_9705);
xnor UO_221 (O_221,N_9619,N_9051);
or UO_222 (O_222,N_9034,N_9614);
nand UO_223 (O_223,N_9926,N_9052);
or UO_224 (O_224,N_9678,N_9033);
nand UO_225 (O_225,N_9366,N_9464);
or UO_226 (O_226,N_9863,N_9868);
nor UO_227 (O_227,N_9683,N_9998);
and UO_228 (O_228,N_9088,N_9268);
nor UO_229 (O_229,N_9412,N_9302);
and UO_230 (O_230,N_9895,N_9294);
nor UO_231 (O_231,N_9921,N_9532);
nand UO_232 (O_232,N_9323,N_9084);
and UO_233 (O_233,N_9836,N_9386);
nor UO_234 (O_234,N_9731,N_9710);
nand UO_235 (O_235,N_9511,N_9535);
nor UO_236 (O_236,N_9313,N_9824);
nand UO_237 (O_237,N_9874,N_9257);
or UO_238 (O_238,N_9112,N_9187);
nand UO_239 (O_239,N_9628,N_9042);
nor UO_240 (O_240,N_9171,N_9817);
and UO_241 (O_241,N_9077,N_9409);
xnor UO_242 (O_242,N_9841,N_9901);
nand UO_243 (O_243,N_9742,N_9065);
nand UO_244 (O_244,N_9481,N_9277);
nor UO_245 (O_245,N_9274,N_9580);
nor UO_246 (O_246,N_9882,N_9976);
nand UO_247 (O_247,N_9226,N_9860);
nand UO_248 (O_248,N_9837,N_9631);
and UO_249 (O_249,N_9997,N_9025);
and UO_250 (O_250,N_9704,N_9443);
nand UO_251 (O_251,N_9018,N_9732);
or UO_252 (O_252,N_9528,N_9670);
and UO_253 (O_253,N_9719,N_9632);
or UO_254 (O_254,N_9623,N_9922);
or UO_255 (O_255,N_9786,N_9867);
nor UO_256 (O_256,N_9031,N_9550);
and UO_257 (O_257,N_9091,N_9996);
nand UO_258 (O_258,N_9987,N_9596);
and UO_259 (O_259,N_9293,N_9588);
xnor UO_260 (O_260,N_9660,N_9039);
or UO_261 (O_261,N_9304,N_9279);
nor UO_262 (O_262,N_9057,N_9146);
or UO_263 (O_263,N_9494,N_9815);
nor UO_264 (O_264,N_9531,N_9078);
and UO_265 (O_265,N_9832,N_9923);
or UO_266 (O_266,N_9889,N_9427);
nor UO_267 (O_267,N_9664,N_9622);
nor UO_268 (O_268,N_9252,N_9436);
or UO_269 (O_269,N_9594,N_9076);
xor UO_270 (O_270,N_9925,N_9856);
or UO_271 (O_271,N_9573,N_9097);
nor UO_272 (O_272,N_9015,N_9264);
nand UO_273 (O_273,N_9408,N_9829);
or UO_274 (O_274,N_9471,N_9716);
nor UO_275 (O_275,N_9936,N_9486);
or UO_276 (O_276,N_9158,N_9209);
xor UO_277 (O_277,N_9043,N_9163);
nor UO_278 (O_278,N_9186,N_9788);
or UO_279 (O_279,N_9929,N_9384);
and UO_280 (O_280,N_9575,N_9404);
nor UO_281 (O_281,N_9516,N_9979);
nor UO_282 (O_282,N_9242,N_9434);
nor UO_283 (O_283,N_9261,N_9041);
nand UO_284 (O_284,N_9642,N_9466);
and UO_285 (O_285,N_9431,N_9643);
nor UO_286 (O_286,N_9447,N_9668);
nand UO_287 (O_287,N_9046,N_9489);
and UO_288 (O_288,N_9942,N_9696);
nor UO_289 (O_289,N_9952,N_9081);
xor UO_290 (O_290,N_9343,N_9067);
or UO_291 (O_291,N_9909,N_9975);
and UO_292 (O_292,N_9469,N_9878);
or UO_293 (O_293,N_9956,N_9544);
or UO_294 (O_294,N_9326,N_9848);
nor UO_295 (O_295,N_9579,N_9904);
nor UO_296 (O_296,N_9385,N_9462);
nand UO_297 (O_297,N_9581,N_9461);
nand UO_298 (O_298,N_9085,N_9812);
and UO_299 (O_299,N_9237,N_9840);
or UO_300 (O_300,N_9962,N_9912);
or UO_301 (O_301,N_9086,N_9289);
or UO_302 (O_302,N_9369,N_9576);
and UO_303 (O_303,N_9117,N_9712);
nor UO_304 (O_304,N_9083,N_9784);
nand UO_305 (O_305,N_9312,N_9509);
and UO_306 (O_306,N_9230,N_9062);
or UO_307 (O_307,N_9574,N_9951);
or UO_308 (O_308,N_9839,N_9513);
and UO_309 (O_309,N_9949,N_9751);
nor UO_310 (O_310,N_9190,N_9240);
or UO_311 (O_311,N_9103,N_9821);
and UO_312 (O_312,N_9934,N_9479);
nor UO_313 (O_313,N_9792,N_9697);
and UO_314 (O_314,N_9400,N_9175);
or UO_315 (O_315,N_9311,N_9721);
or UO_316 (O_316,N_9492,N_9773);
xnor UO_317 (O_317,N_9148,N_9445);
and UO_318 (O_318,N_9377,N_9525);
nor UO_319 (O_319,N_9181,N_9258);
and UO_320 (O_320,N_9641,N_9676);
or UO_321 (O_321,N_9021,N_9496);
or UO_322 (O_322,N_9059,N_9886);
nand UO_323 (O_323,N_9202,N_9896);
nand UO_324 (O_324,N_9702,N_9162);
and UO_325 (O_325,N_9053,N_9452);
or UO_326 (O_326,N_9241,N_9772);
nor UO_327 (O_327,N_9338,N_9621);
nand UO_328 (O_328,N_9601,N_9071);
nor UO_329 (O_329,N_9555,N_9866);
and UO_330 (O_330,N_9771,N_9014);
or UO_331 (O_331,N_9724,N_9482);
xor UO_332 (O_332,N_9425,N_9953);
xnor UO_333 (O_333,N_9030,N_9070);
and UO_334 (O_334,N_9485,N_9317);
nand UO_335 (O_335,N_9503,N_9517);
and UO_336 (O_336,N_9322,N_9789);
nand UO_337 (O_337,N_9255,N_9959);
nand UO_338 (O_338,N_9438,N_9591);
or UO_339 (O_339,N_9411,N_9123);
nor UO_340 (O_340,N_9340,N_9381);
nor UO_341 (O_341,N_9500,N_9723);
or UO_342 (O_342,N_9835,N_9450);
or UO_343 (O_343,N_9879,N_9497);
nand UO_344 (O_344,N_9559,N_9185);
and UO_345 (O_345,N_9675,N_9838);
nand UO_346 (O_346,N_9490,N_9239);
xnor UO_347 (O_347,N_9376,N_9973);
or UO_348 (O_348,N_9308,N_9161);
nor UO_349 (O_349,N_9888,N_9135);
nand UO_350 (O_350,N_9468,N_9137);
nand UO_351 (O_351,N_9802,N_9508);
or UO_352 (O_352,N_9750,N_9560);
nor UO_353 (O_353,N_9367,N_9016);
nor UO_354 (O_354,N_9410,N_9937);
nand UO_355 (O_355,N_9853,N_9040);
and UO_356 (O_356,N_9332,N_9558);
nor UO_357 (O_357,N_9542,N_9378);
nor UO_358 (O_358,N_9374,N_9406);
nand UO_359 (O_359,N_9319,N_9920);
nand UO_360 (O_360,N_9422,N_9651);
xnor UO_361 (O_361,N_9924,N_9457);
nand UO_362 (O_362,N_9626,N_9267);
nand UO_363 (O_363,N_9775,N_9361);
and UO_364 (O_364,N_9857,N_9299);
or UO_365 (O_365,N_9221,N_9870);
nand UO_366 (O_366,N_9744,N_9128);
nand UO_367 (O_367,N_9800,N_9420);
and UO_368 (O_368,N_9288,N_9250);
and UO_369 (O_369,N_9569,N_9526);
and UO_370 (O_370,N_9722,N_9725);
nand UO_371 (O_371,N_9774,N_9201);
nor UO_372 (O_372,N_9013,N_9518);
nor UO_373 (O_373,N_9172,N_9600);
nor UO_374 (O_374,N_9460,N_9419);
xnor UO_375 (O_375,N_9507,N_9605);
or UO_376 (O_376,N_9871,N_9957);
and UO_377 (O_377,N_9011,N_9695);
nand UO_378 (O_378,N_9760,N_9231);
nand UO_379 (O_379,N_9417,N_9814);
or UO_380 (O_380,N_9746,N_9797);
and UO_381 (O_381,N_9603,N_9767);
and UO_382 (O_382,N_9403,N_9756);
and UO_383 (O_383,N_9873,N_9139);
or UO_384 (O_384,N_9545,N_9448);
nor UO_385 (O_385,N_9073,N_9650);
or UO_386 (O_386,N_9007,N_9363);
nor UO_387 (O_387,N_9714,N_9686);
or UO_388 (O_388,N_9617,N_9597);
and UO_389 (O_389,N_9553,N_9314);
and UO_390 (O_390,N_9701,N_9189);
nor UO_391 (O_391,N_9842,N_9176);
nand UO_392 (O_392,N_9762,N_9325);
and UO_393 (O_393,N_9595,N_9303);
nor UO_394 (O_394,N_9269,N_9228);
and UO_395 (O_395,N_9220,N_9850);
and UO_396 (O_396,N_9476,N_9939);
nand UO_397 (O_397,N_9012,N_9780);
nand UO_398 (O_398,N_9037,N_9193);
nand UO_399 (O_399,N_9164,N_9565);
nor UO_400 (O_400,N_9061,N_9416);
xor UO_401 (O_401,N_9297,N_9153);
nor UO_402 (O_402,N_9970,N_9349);
nand UO_403 (O_403,N_9341,N_9523);
xor UO_404 (O_404,N_9437,N_9357);
nand UO_405 (O_405,N_9020,N_9415);
xnor UO_406 (O_406,N_9782,N_9372);
or UO_407 (O_407,N_9096,N_9449);
or UO_408 (O_408,N_9182,N_9933);
and UO_409 (O_409,N_9442,N_9402);
nor UO_410 (O_410,N_9473,N_9284);
or UO_411 (O_411,N_9915,N_9095);
or UO_412 (O_412,N_9346,N_9945);
nor UO_413 (O_413,N_9167,N_9778);
and UO_414 (O_414,N_9561,N_9271);
or UO_415 (O_415,N_9606,N_9397);
or UO_416 (O_416,N_9730,N_9211);
or UO_417 (O_417,N_9478,N_9262);
and UO_418 (O_418,N_9862,N_9847);
nor UO_419 (O_419,N_9414,N_9984);
or UO_420 (O_420,N_9911,N_9764);
and UO_421 (O_421,N_9249,N_9572);
nor UO_422 (O_422,N_9229,N_9295);
and UO_423 (O_423,N_9941,N_9208);
or UO_424 (O_424,N_9662,N_9155);
and UO_425 (O_425,N_9822,N_9364);
nand UO_426 (O_426,N_9693,N_9826);
nand UO_427 (O_427,N_9342,N_9985);
or UO_428 (O_428,N_9441,N_9074);
or UO_429 (O_429,N_9129,N_9166);
nor UO_430 (O_430,N_9245,N_9009);
nand UO_431 (O_431,N_9354,N_9339);
nand UO_432 (O_432,N_9872,N_9563);
and UO_433 (O_433,N_9111,N_9827);
nor UO_434 (O_434,N_9197,N_9145);
nor UO_435 (O_435,N_9899,N_9759);
and UO_436 (O_436,N_9779,N_9451);
nand UO_437 (O_437,N_9551,N_9543);
nor UO_438 (O_438,N_9562,N_9914);
or UO_439 (O_439,N_9646,N_9699);
xor UO_440 (O_440,N_9333,N_9260);
and UO_441 (O_441,N_9968,N_9156);
nand UO_442 (O_442,N_9522,N_9960);
xor UO_443 (O_443,N_9636,N_9687);
nand UO_444 (O_444,N_9058,N_9992);
or UO_445 (O_445,N_9352,N_9682);
or UO_446 (O_446,N_9700,N_9665);
nand UO_447 (O_447,N_9587,N_9583);
xnor UO_448 (O_448,N_9502,N_9980);
or UO_449 (O_449,N_9456,N_9141);
or UO_450 (O_450,N_9253,N_9027);
nand UO_451 (O_451,N_9877,N_9054);
nand UO_452 (O_452,N_9917,N_9828);
nand UO_453 (O_453,N_9212,N_9327);
nand UO_454 (O_454,N_9728,N_9275);
nand UO_455 (O_455,N_9539,N_9982);
nand UO_456 (O_456,N_9336,N_9965);
and UO_457 (O_457,N_9121,N_9745);
and UO_458 (O_458,N_9005,N_9356);
or UO_459 (O_459,N_9315,N_9902);
and UO_460 (O_460,N_9833,N_9884);
nand UO_461 (O_461,N_9567,N_9907);
nor UO_462 (O_462,N_9002,N_9506);
and UO_463 (O_463,N_9244,N_9329);
xor UO_464 (O_464,N_9147,N_9184);
nand UO_465 (O_465,N_9038,N_9316);
and UO_466 (O_466,N_9225,N_9113);
or UO_467 (O_467,N_9635,N_9995);
and UO_468 (O_468,N_9008,N_9480);
nor UO_469 (O_469,N_9656,N_9679);
nand UO_470 (O_470,N_9200,N_9183);
nor UO_471 (O_471,N_9537,N_9825);
and UO_472 (O_472,N_9734,N_9165);
xnor UO_473 (O_473,N_9653,N_9639);
nand UO_474 (O_474,N_9243,N_9370);
nor UO_475 (O_475,N_9251,N_9050);
nand UO_476 (O_476,N_9170,N_9359);
or UO_477 (O_477,N_9214,N_9611);
or UO_478 (O_478,N_9455,N_9082);
or UO_479 (O_479,N_9846,N_9608);
nor UO_480 (O_480,N_9521,N_9353);
or UO_481 (O_481,N_9674,N_9498);
and UO_482 (O_482,N_9108,N_9019);
xor UO_483 (O_483,N_9505,N_9713);
nand UO_484 (O_484,N_9571,N_9799);
or UO_485 (O_485,N_9820,N_9291);
or UO_486 (O_486,N_9360,N_9781);
nand UO_487 (O_487,N_9324,N_9504);
or UO_488 (O_488,N_9174,N_9398);
nor UO_489 (O_489,N_9766,N_9254);
and UO_490 (O_490,N_9217,N_9913);
xor UO_491 (O_491,N_9755,N_9858);
or UO_492 (O_492,N_9607,N_9943);
nor UO_493 (O_493,N_9615,N_9977);
nor UO_494 (O_494,N_9717,N_9334);
and UO_495 (O_495,N_9233,N_9763);
and UO_496 (O_496,N_9035,N_9671);
nor UO_497 (O_497,N_9729,N_9290);
nand UO_498 (O_498,N_9210,N_9947);
nand UO_499 (O_499,N_9620,N_9993);
nand UO_500 (O_500,N_9935,N_9977);
or UO_501 (O_501,N_9719,N_9524);
nand UO_502 (O_502,N_9692,N_9991);
and UO_503 (O_503,N_9248,N_9216);
nor UO_504 (O_504,N_9338,N_9987);
xor UO_505 (O_505,N_9121,N_9184);
nor UO_506 (O_506,N_9575,N_9741);
nor UO_507 (O_507,N_9760,N_9433);
and UO_508 (O_508,N_9278,N_9701);
and UO_509 (O_509,N_9211,N_9134);
nand UO_510 (O_510,N_9524,N_9861);
or UO_511 (O_511,N_9887,N_9990);
nand UO_512 (O_512,N_9777,N_9717);
and UO_513 (O_513,N_9075,N_9370);
nor UO_514 (O_514,N_9064,N_9402);
and UO_515 (O_515,N_9469,N_9558);
nand UO_516 (O_516,N_9910,N_9847);
or UO_517 (O_517,N_9550,N_9294);
and UO_518 (O_518,N_9392,N_9480);
nand UO_519 (O_519,N_9556,N_9375);
and UO_520 (O_520,N_9226,N_9289);
nor UO_521 (O_521,N_9328,N_9280);
nor UO_522 (O_522,N_9124,N_9906);
and UO_523 (O_523,N_9810,N_9935);
or UO_524 (O_524,N_9944,N_9516);
or UO_525 (O_525,N_9638,N_9254);
xor UO_526 (O_526,N_9665,N_9642);
and UO_527 (O_527,N_9653,N_9762);
nand UO_528 (O_528,N_9712,N_9312);
or UO_529 (O_529,N_9134,N_9515);
nand UO_530 (O_530,N_9859,N_9601);
nor UO_531 (O_531,N_9482,N_9879);
and UO_532 (O_532,N_9897,N_9065);
and UO_533 (O_533,N_9743,N_9491);
nor UO_534 (O_534,N_9693,N_9380);
or UO_535 (O_535,N_9324,N_9633);
nand UO_536 (O_536,N_9164,N_9119);
or UO_537 (O_537,N_9448,N_9544);
and UO_538 (O_538,N_9583,N_9977);
and UO_539 (O_539,N_9122,N_9782);
and UO_540 (O_540,N_9382,N_9209);
xnor UO_541 (O_541,N_9297,N_9457);
nand UO_542 (O_542,N_9523,N_9247);
or UO_543 (O_543,N_9561,N_9269);
xnor UO_544 (O_544,N_9655,N_9089);
xnor UO_545 (O_545,N_9362,N_9020);
or UO_546 (O_546,N_9244,N_9254);
nand UO_547 (O_547,N_9582,N_9943);
or UO_548 (O_548,N_9754,N_9685);
nor UO_549 (O_549,N_9588,N_9663);
nand UO_550 (O_550,N_9209,N_9038);
or UO_551 (O_551,N_9414,N_9663);
and UO_552 (O_552,N_9667,N_9258);
nor UO_553 (O_553,N_9883,N_9965);
and UO_554 (O_554,N_9651,N_9226);
or UO_555 (O_555,N_9229,N_9207);
nor UO_556 (O_556,N_9303,N_9042);
nor UO_557 (O_557,N_9715,N_9469);
and UO_558 (O_558,N_9336,N_9873);
or UO_559 (O_559,N_9267,N_9144);
nand UO_560 (O_560,N_9533,N_9944);
or UO_561 (O_561,N_9465,N_9926);
nor UO_562 (O_562,N_9139,N_9144);
nor UO_563 (O_563,N_9668,N_9458);
nor UO_564 (O_564,N_9909,N_9928);
nand UO_565 (O_565,N_9766,N_9047);
and UO_566 (O_566,N_9477,N_9930);
or UO_567 (O_567,N_9692,N_9704);
nand UO_568 (O_568,N_9933,N_9240);
nand UO_569 (O_569,N_9049,N_9509);
or UO_570 (O_570,N_9637,N_9191);
nor UO_571 (O_571,N_9409,N_9841);
nor UO_572 (O_572,N_9458,N_9348);
nand UO_573 (O_573,N_9003,N_9777);
or UO_574 (O_574,N_9059,N_9260);
xor UO_575 (O_575,N_9886,N_9389);
nand UO_576 (O_576,N_9381,N_9365);
nand UO_577 (O_577,N_9454,N_9210);
nor UO_578 (O_578,N_9616,N_9984);
nand UO_579 (O_579,N_9439,N_9658);
or UO_580 (O_580,N_9965,N_9726);
or UO_581 (O_581,N_9751,N_9673);
nand UO_582 (O_582,N_9645,N_9650);
or UO_583 (O_583,N_9609,N_9961);
nand UO_584 (O_584,N_9439,N_9883);
nor UO_585 (O_585,N_9591,N_9685);
nand UO_586 (O_586,N_9430,N_9214);
xor UO_587 (O_587,N_9502,N_9231);
or UO_588 (O_588,N_9291,N_9581);
and UO_589 (O_589,N_9182,N_9976);
and UO_590 (O_590,N_9308,N_9645);
nand UO_591 (O_591,N_9207,N_9209);
and UO_592 (O_592,N_9300,N_9071);
and UO_593 (O_593,N_9076,N_9027);
nand UO_594 (O_594,N_9814,N_9382);
nor UO_595 (O_595,N_9123,N_9091);
nand UO_596 (O_596,N_9344,N_9884);
and UO_597 (O_597,N_9351,N_9655);
nor UO_598 (O_598,N_9575,N_9302);
nand UO_599 (O_599,N_9507,N_9536);
nor UO_600 (O_600,N_9696,N_9888);
nor UO_601 (O_601,N_9599,N_9554);
or UO_602 (O_602,N_9107,N_9490);
nor UO_603 (O_603,N_9071,N_9716);
or UO_604 (O_604,N_9047,N_9212);
nor UO_605 (O_605,N_9235,N_9571);
and UO_606 (O_606,N_9036,N_9472);
and UO_607 (O_607,N_9701,N_9729);
nand UO_608 (O_608,N_9942,N_9244);
and UO_609 (O_609,N_9579,N_9248);
nor UO_610 (O_610,N_9720,N_9945);
nand UO_611 (O_611,N_9936,N_9571);
nand UO_612 (O_612,N_9886,N_9725);
or UO_613 (O_613,N_9356,N_9300);
or UO_614 (O_614,N_9585,N_9228);
nand UO_615 (O_615,N_9049,N_9508);
or UO_616 (O_616,N_9796,N_9355);
nand UO_617 (O_617,N_9821,N_9531);
xnor UO_618 (O_618,N_9453,N_9909);
nor UO_619 (O_619,N_9635,N_9676);
xnor UO_620 (O_620,N_9427,N_9364);
nor UO_621 (O_621,N_9143,N_9025);
or UO_622 (O_622,N_9470,N_9660);
or UO_623 (O_623,N_9841,N_9306);
xnor UO_624 (O_624,N_9613,N_9512);
and UO_625 (O_625,N_9288,N_9370);
nor UO_626 (O_626,N_9112,N_9858);
nor UO_627 (O_627,N_9478,N_9647);
nor UO_628 (O_628,N_9494,N_9697);
and UO_629 (O_629,N_9426,N_9845);
nor UO_630 (O_630,N_9460,N_9381);
nor UO_631 (O_631,N_9874,N_9997);
and UO_632 (O_632,N_9667,N_9467);
nand UO_633 (O_633,N_9271,N_9293);
or UO_634 (O_634,N_9160,N_9753);
or UO_635 (O_635,N_9808,N_9410);
nor UO_636 (O_636,N_9841,N_9759);
nor UO_637 (O_637,N_9750,N_9562);
nand UO_638 (O_638,N_9836,N_9888);
nor UO_639 (O_639,N_9831,N_9360);
or UO_640 (O_640,N_9153,N_9563);
or UO_641 (O_641,N_9267,N_9598);
xor UO_642 (O_642,N_9659,N_9900);
and UO_643 (O_643,N_9961,N_9915);
or UO_644 (O_644,N_9541,N_9266);
and UO_645 (O_645,N_9244,N_9819);
or UO_646 (O_646,N_9103,N_9498);
and UO_647 (O_647,N_9264,N_9571);
xor UO_648 (O_648,N_9527,N_9943);
or UO_649 (O_649,N_9901,N_9530);
nand UO_650 (O_650,N_9898,N_9377);
nand UO_651 (O_651,N_9128,N_9177);
nor UO_652 (O_652,N_9488,N_9567);
nand UO_653 (O_653,N_9896,N_9237);
and UO_654 (O_654,N_9791,N_9142);
nand UO_655 (O_655,N_9812,N_9746);
nor UO_656 (O_656,N_9150,N_9889);
or UO_657 (O_657,N_9542,N_9330);
nor UO_658 (O_658,N_9958,N_9105);
nor UO_659 (O_659,N_9166,N_9065);
and UO_660 (O_660,N_9384,N_9555);
and UO_661 (O_661,N_9807,N_9978);
nor UO_662 (O_662,N_9824,N_9343);
or UO_663 (O_663,N_9528,N_9425);
nand UO_664 (O_664,N_9383,N_9714);
nand UO_665 (O_665,N_9205,N_9398);
or UO_666 (O_666,N_9720,N_9866);
or UO_667 (O_667,N_9614,N_9456);
nor UO_668 (O_668,N_9036,N_9313);
or UO_669 (O_669,N_9254,N_9523);
nand UO_670 (O_670,N_9901,N_9169);
or UO_671 (O_671,N_9317,N_9866);
nand UO_672 (O_672,N_9671,N_9085);
nand UO_673 (O_673,N_9875,N_9187);
nor UO_674 (O_674,N_9751,N_9281);
nor UO_675 (O_675,N_9284,N_9329);
nor UO_676 (O_676,N_9133,N_9013);
or UO_677 (O_677,N_9113,N_9583);
or UO_678 (O_678,N_9530,N_9663);
and UO_679 (O_679,N_9656,N_9721);
or UO_680 (O_680,N_9669,N_9012);
and UO_681 (O_681,N_9913,N_9581);
or UO_682 (O_682,N_9363,N_9297);
xnor UO_683 (O_683,N_9960,N_9805);
and UO_684 (O_684,N_9259,N_9029);
and UO_685 (O_685,N_9329,N_9728);
xor UO_686 (O_686,N_9299,N_9811);
nor UO_687 (O_687,N_9077,N_9260);
and UO_688 (O_688,N_9522,N_9558);
nor UO_689 (O_689,N_9514,N_9507);
or UO_690 (O_690,N_9039,N_9686);
nor UO_691 (O_691,N_9112,N_9267);
or UO_692 (O_692,N_9225,N_9071);
or UO_693 (O_693,N_9859,N_9239);
nand UO_694 (O_694,N_9865,N_9451);
or UO_695 (O_695,N_9971,N_9758);
nand UO_696 (O_696,N_9883,N_9623);
nand UO_697 (O_697,N_9582,N_9459);
nor UO_698 (O_698,N_9488,N_9787);
or UO_699 (O_699,N_9891,N_9353);
and UO_700 (O_700,N_9459,N_9617);
nand UO_701 (O_701,N_9340,N_9977);
and UO_702 (O_702,N_9065,N_9962);
nand UO_703 (O_703,N_9249,N_9263);
or UO_704 (O_704,N_9450,N_9521);
nor UO_705 (O_705,N_9187,N_9180);
nor UO_706 (O_706,N_9534,N_9258);
and UO_707 (O_707,N_9879,N_9597);
nor UO_708 (O_708,N_9223,N_9376);
and UO_709 (O_709,N_9342,N_9138);
xor UO_710 (O_710,N_9395,N_9276);
and UO_711 (O_711,N_9664,N_9850);
nor UO_712 (O_712,N_9583,N_9827);
or UO_713 (O_713,N_9565,N_9652);
and UO_714 (O_714,N_9876,N_9132);
xnor UO_715 (O_715,N_9566,N_9232);
and UO_716 (O_716,N_9800,N_9801);
nor UO_717 (O_717,N_9060,N_9390);
nor UO_718 (O_718,N_9705,N_9106);
nor UO_719 (O_719,N_9994,N_9810);
or UO_720 (O_720,N_9305,N_9321);
nand UO_721 (O_721,N_9506,N_9618);
xor UO_722 (O_722,N_9885,N_9121);
nand UO_723 (O_723,N_9832,N_9598);
nor UO_724 (O_724,N_9049,N_9811);
or UO_725 (O_725,N_9814,N_9752);
nor UO_726 (O_726,N_9618,N_9665);
or UO_727 (O_727,N_9597,N_9902);
or UO_728 (O_728,N_9214,N_9646);
nor UO_729 (O_729,N_9170,N_9915);
nand UO_730 (O_730,N_9422,N_9582);
xor UO_731 (O_731,N_9833,N_9406);
nand UO_732 (O_732,N_9267,N_9330);
and UO_733 (O_733,N_9516,N_9785);
nand UO_734 (O_734,N_9587,N_9927);
nand UO_735 (O_735,N_9727,N_9757);
nor UO_736 (O_736,N_9723,N_9606);
nor UO_737 (O_737,N_9559,N_9337);
nand UO_738 (O_738,N_9478,N_9082);
nor UO_739 (O_739,N_9502,N_9785);
nor UO_740 (O_740,N_9783,N_9318);
nand UO_741 (O_741,N_9153,N_9195);
and UO_742 (O_742,N_9240,N_9103);
and UO_743 (O_743,N_9111,N_9833);
and UO_744 (O_744,N_9399,N_9694);
nor UO_745 (O_745,N_9813,N_9675);
or UO_746 (O_746,N_9499,N_9644);
or UO_747 (O_747,N_9609,N_9193);
or UO_748 (O_748,N_9077,N_9212);
and UO_749 (O_749,N_9775,N_9566);
nor UO_750 (O_750,N_9126,N_9706);
nand UO_751 (O_751,N_9377,N_9048);
xnor UO_752 (O_752,N_9451,N_9605);
nor UO_753 (O_753,N_9784,N_9793);
or UO_754 (O_754,N_9222,N_9349);
nand UO_755 (O_755,N_9765,N_9664);
or UO_756 (O_756,N_9522,N_9986);
and UO_757 (O_757,N_9464,N_9382);
and UO_758 (O_758,N_9775,N_9393);
nand UO_759 (O_759,N_9329,N_9918);
and UO_760 (O_760,N_9615,N_9025);
or UO_761 (O_761,N_9375,N_9659);
nor UO_762 (O_762,N_9544,N_9241);
nor UO_763 (O_763,N_9044,N_9052);
nand UO_764 (O_764,N_9717,N_9249);
nand UO_765 (O_765,N_9822,N_9709);
and UO_766 (O_766,N_9887,N_9117);
and UO_767 (O_767,N_9250,N_9925);
nand UO_768 (O_768,N_9493,N_9220);
or UO_769 (O_769,N_9584,N_9603);
nand UO_770 (O_770,N_9134,N_9176);
nor UO_771 (O_771,N_9957,N_9595);
and UO_772 (O_772,N_9119,N_9299);
nor UO_773 (O_773,N_9598,N_9187);
nand UO_774 (O_774,N_9809,N_9748);
xor UO_775 (O_775,N_9665,N_9490);
nand UO_776 (O_776,N_9027,N_9167);
nand UO_777 (O_777,N_9023,N_9092);
and UO_778 (O_778,N_9634,N_9932);
or UO_779 (O_779,N_9527,N_9224);
or UO_780 (O_780,N_9338,N_9394);
and UO_781 (O_781,N_9612,N_9032);
or UO_782 (O_782,N_9575,N_9440);
nand UO_783 (O_783,N_9136,N_9511);
nand UO_784 (O_784,N_9337,N_9215);
and UO_785 (O_785,N_9479,N_9437);
nor UO_786 (O_786,N_9308,N_9371);
nand UO_787 (O_787,N_9451,N_9328);
xor UO_788 (O_788,N_9664,N_9120);
nand UO_789 (O_789,N_9421,N_9238);
nand UO_790 (O_790,N_9742,N_9593);
and UO_791 (O_791,N_9272,N_9125);
nand UO_792 (O_792,N_9656,N_9014);
and UO_793 (O_793,N_9192,N_9984);
nand UO_794 (O_794,N_9673,N_9353);
nand UO_795 (O_795,N_9996,N_9922);
nand UO_796 (O_796,N_9777,N_9838);
and UO_797 (O_797,N_9176,N_9654);
nand UO_798 (O_798,N_9290,N_9637);
or UO_799 (O_799,N_9941,N_9186);
xnor UO_800 (O_800,N_9926,N_9898);
nand UO_801 (O_801,N_9577,N_9914);
and UO_802 (O_802,N_9838,N_9509);
and UO_803 (O_803,N_9369,N_9551);
or UO_804 (O_804,N_9888,N_9584);
nand UO_805 (O_805,N_9182,N_9185);
nand UO_806 (O_806,N_9165,N_9250);
nor UO_807 (O_807,N_9251,N_9912);
or UO_808 (O_808,N_9059,N_9797);
or UO_809 (O_809,N_9323,N_9047);
and UO_810 (O_810,N_9055,N_9466);
nor UO_811 (O_811,N_9642,N_9421);
or UO_812 (O_812,N_9682,N_9822);
nor UO_813 (O_813,N_9840,N_9637);
and UO_814 (O_814,N_9977,N_9459);
and UO_815 (O_815,N_9132,N_9416);
nor UO_816 (O_816,N_9578,N_9532);
and UO_817 (O_817,N_9503,N_9303);
nor UO_818 (O_818,N_9441,N_9886);
and UO_819 (O_819,N_9028,N_9503);
nand UO_820 (O_820,N_9698,N_9724);
nor UO_821 (O_821,N_9097,N_9172);
nand UO_822 (O_822,N_9216,N_9580);
nor UO_823 (O_823,N_9783,N_9293);
and UO_824 (O_824,N_9628,N_9614);
nor UO_825 (O_825,N_9276,N_9594);
nor UO_826 (O_826,N_9353,N_9279);
nand UO_827 (O_827,N_9785,N_9706);
or UO_828 (O_828,N_9042,N_9348);
nor UO_829 (O_829,N_9817,N_9077);
and UO_830 (O_830,N_9506,N_9757);
or UO_831 (O_831,N_9965,N_9125);
or UO_832 (O_832,N_9435,N_9200);
xor UO_833 (O_833,N_9426,N_9287);
nor UO_834 (O_834,N_9307,N_9988);
and UO_835 (O_835,N_9904,N_9660);
or UO_836 (O_836,N_9220,N_9318);
nand UO_837 (O_837,N_9885,N_9058);
xnor UO_838 (O_838,N_9128,N_9884);
nor UO_839 (O_839,N_9047,N_9748);
nand UO_840 (O_840,N_9362,N_9985);
and UO_841 (O_841,N_9725,N_9753);
and UO_842 (O_842,N_9878,N_9857);
and UO_843 (O_843,N_9954,N_9741);
xor UO_844 (O_844,N_9329,N_9644);
nor UO_845 (O_845,N_9221,N_9712);
nor UO_846 (O_846,N_9991,N_9601);
nand UO_847 (O_847,N_9446,N_9952);
and UO_848 (O_848,N_9293,N_9865);
nor UO_849 (O_849,N_9674,N_9119);
nor UO_850 (O_850,N_9212,N_9129);
nor UO_851 (O_851,N_9267,N_9592);
or UO_852 (O_852,N_9589,N_9402);
and UO_853 (O_853,N_9038,N_9531);
and UO_854 (O_854,N_9587,N_9519);
nand UO_855 (O_855,N_9748,N_9964);
and UO_856 (O_856,N_9785,N_9133);
or UO_857 (O_857,N_9695,N_9676);
and UO_858 (O_858,N_9331,N_9817);
nor UO_859 (O_859,N_9465,N_9380);
nand UO_860 (O_860,N_9752,N_9008);
nor UO_861 (O_861,N_9230,N_9457);
nand UO_862 (O_862,N_9632,N_9856);
nand UO_863 (O_863,N_9005,N_9179);
nand UO_864 (O_864,N_9773,N_9928);
nor UO_865 (O_865,N_9387,N_9455);
and UO_866 (O_866,N_9030,N_9172);
or UO_867 (O_867,N_9137,N_9984);
nor UO_868 (O_868,N_9493,N_9956);
and UO_869 (O_869,N_9566,N_9373);
or UO_870 (O_870,N_9173,N_9100);
or UO_871 (O_871,N_9660,N_9913);
and UO_872 (O_872,N_9202,N_9997);
and UO_873 (O_873,N_9204,N_9580);
nand UO_874 (O_874,N_9000,N_9393);
nor UO_875 (O_875,N_9510,N_9018);
and UO_876 (O_876,N_9029,N_9811);
or UO_877 (O_877,N_9708,N_9698);
xor UO_878 (O_878,N_9124,N_9779);
or UO_879 (O_879,N_9174,N_9820);
nand UO_880 (O_880,N_9911,N_9650);
nor UO_881 (O_881,N_9720,N_9643);
and UO_882 (O_882,N_9329,N_9669);
and UO_883 (O_883,N_9386,N_9399);
nand UO_884 (O_884,N_9480,N_9084);
and UO_885 (O_885,N_9520,N_9292);
or UO_886 (O_886,N_9551,N_9250);
nand UO_887 (O_887,N_9915,N_9281);
or UO_888 (O_888,N_9011,N_9221);
and UO_889 (O_889,N_9056,N_9001);
or UO_890 (O_890,N_9447,N_9223);
nor UO_891 (O_891,N_9776,N_9792);
or UO_892 (O_892,N_9603,N_9563);
nand UO_893 (O_893,N_9281,N_9934);
nor UO_894 (O_894,N_9244,N_9216);
xnor UO_895 (O_895,N_9423,N_9425);
nor UO_896 (O_896,N_9394,N_9263);
nand UO_897 (O_897,N_9429,N_9289);
nor UO_898 (O_898,N_9149,N_9600);
and UO_899 (O_899,N_9378,N_9758);
or UO_900 (O_900,N_9353,N_9976);
or UO_901 (O_901,N_9262,N_9814);
nand UO_902 (O_902,N_9122,N_9074);
and UO_903 (O_903,N_9948,N_9249);
and UO_904 (O_904,N_9324,N_9241);
nand UO_905 (O_905,N_9606,N_9527);
xor UO_906 (O_906,N_9887,N_9531);
and UO_907 (O_907,N_9489,N_9153);
nor UO_908 (O_908,N_9888,N_9456);
nor UO_909 (O_909,N_9691,N_9591);
or UO_910 (O_910,N_9860,N_9976);
nor UO_911 (O_911,N_9976,N_9079);
xnor UO_912 (O_912,N_9576,N_9824);
nor UO_913 (O_913,N_9392,N_9159);
nand UO_914 (O_914,N_9680,N_9057);
nand UO_915 (O_915,N_9960,N_9135);
or UO_916 (O_916,N_9186,N_9285);
nand UO_917 (O_917,N_9937,N_9094);
or UO_918 (O_918,N_9337,N_9532);
or UO_919 (O_919,N_9854,N_9627);
or UO_920 (O_920,N_9682,N_9440);
and UO_921 (O_921,N_9703,N_9652);
or UO_922 (O_922,N_9571,N_9848);
nor UO_923 (O_923,N_9339,N_9362);
xnor UO_924 (O_924,N_9406,N_9540);
nand UO_925 (O_925,N_9360,N_9037);
xnor UO_926 (O_926,N_9582,N_9913);
or UO_927 (O_927,N_9347,N_9261);
xnor UO_928 (O_928,N_9591,N_9241);
and UO_929 (O_929,N_9373,N_9656);
and UO_930 (O_930,N_9923,N_9348);
nor UO_931 (O_931,N_9654,N_9513);
nor UO_932 (O_932,N_9490,N_9232);
or UO_933 (O_933,N_9660,N_9952);
or UO_934 (O_934,N_9066,N_9993);
and UO_935 (O_935,N_9179,N_9181);
and UO_936 (O_936,N_9357,N_9825);
and UO_937 (O_937,N_9159,N_9549);
or UO_938 (O_938,N_9306,N_9988);
nand UO_939 (O_939,N_9760,N_9169);
and UO_940 (O_940,N_9255,N_9586);
nand UO_941 (O_941,N_9544,N_9170);
nor UO_942 (O_942,N_9267,N_9507);
and UO_943 (O_943,N_9864,N_9179);
and UO_944 (O_944,N_9671,N_9247);
nor UO_945 (O_945,N_9625,N_9539);
and UO_946 (O_946,N_9370,N_9303);
or UO_947 (O_947,N_9943,N_9977);
or UO_948 (O_948,N_9225,N_9924);
nor UO_949 (O_949,N_9500,N_9161);
nand UO_950 (O_950,N_9730,N_9980);
or UO_951 (O_951,N_9279,N_9023);
nand UO_952 (O_952,N_9214,N_9890);
and UO_953 (O_953,N_9360,N_9966);
nor UO_954 (O_954,N_9538,N_9758);
or UO_955 (O_955,N_9986,N_9285);
and UO_956 (O_956,N_9612,N_9009);
and UO_957 (O_957,N_9828,N_9997);
and UO_958 (O_958,N_9028,N_9326);
or UO_959 (O_959,N_9336,N_9433);
or UO_960 (O_960,N_9653,N_9966);
or UO_961 (O_961,N_9842,N_9773);
xor UO_962 (O_962,N_9448,N_9092);
nor UO_963 (O_963,N_9084,N_9972);
or UO_964 (O_964,N_9740,N_9477);
and UO_965 (O_965,N_9011,N_9968);
xnor UO_966 (O_966,N_9928,N_9228);
or UO_967 (O_967,N_9645,N_9099);
and UO_968 (O_968,N_9561,N_9332);
nand UO_969 (O_969,N_9094,N_9119);
nand UO_970 (O_970,N_9920,N_9115);
and UO_971 (O_971,N_9403,N_9624);
xnor UO_972 (O_972,N_9366,N_9501);
and UO_973 (O_973,N_9685,N_9846);
or UO_974 (O_974,N_9040,N_9802);
and UO_975 (O_975,N_9463,N_9280);
or UO_976 (O_976,N_9196,N_9464);
xor UO_977 (O_977,N_9467,N_9922);
or UO_978 (O_978,N_9017,N_9326);
nand UO_979 (O_979,N_9899,N_9986);
nor UO_980 (O_980,N_9538,N_9879);
or UO_981 (O_981,N_9328,N_9024);
or UO_982 (O_982,N_9236,N_9551);
and UO_983 (O_983,N_9996,N_9931);
or UO_984 (O_984,N_9791,N_9981);
xor UO_985 (O_985,N_9441,N_9463);
nand UO_986 (O_986,N_9636,N_9989);
nand UO_987 (O_987,N_9832,N_9489);
nand UO_988 (O_988,N_9265,N_9055);
xnor UO_989 (O_989,N_9052,N_9347);
nor UO_990 (O_990,N_9658,N_9145);
nor UO_991 (O_991,N_9740,N_9124);
or UO_992 (O_992,N_9632,N_9295);
nand UO_993 (O_993,N_9114,N_9019);
xnor UO_994 (O_994,N_9440,N_9744);
nand UO_995 (O_995,N_9429,N_9928);
or UO_996 (O_996,N_9305,N_9436);
and UO_997 (O_997,N_9031,N_9770);
nor UO_998 (O_998,N_9054,N_9065);
xor UO_999 (O_999,N_9692,N_9215);
nor UO_1000 (O_1000,N_9774,N_9739);
xnor UO_1001 (O_1001,N_9843,N_9063);
nand UO_1002 (O_1002,N_9080,N_9075);
or UO_1003 (O_1003,N_9948,N_9246);
nor UO_1004 (O_1004,N_9225,N_9697);
or UO_1005 (O_1005,N_9146,N_9461);
or UO_1006 (O_1006,N_9392,N_9089);
xor UO_1007 (O_1007,N_9538,N_9353);
or UO_1008 (O_1008,N_9278,N_9200);
nand UO_1009 (O_1009,N_9753,N_9346);
or UO_1010 (O_1010,N_9012,N_9390);
and UO_1011 (O_1011,N_9752,N_9604);
xnor UO_1012 (O_1012,N_9786,N_9637);
or UO_1013 (O_1013,N_9420,N_9240);
or UO_1014 (O_1014,N_9621,N_9663);
nor UO_1015 (O_1015,N_9551,N_9726);
nand UO_1016 (O_1016,N_9115,N_9722);
xor UO_1017 (O_1017,N_9320,N_9278);
nor UO_1018 (O_1018,N_9228,N_9938);
nand UO_1019 (O_1019,N_9952,N_9717);
nand UO_1020 (O_1020,N_9912,N_9458);
and UO_1021 (O_1021,N_9705,N_9382);
or UO_1022 (O_1022,N_9345,N_9994);
and UO_1023 (O_1023,N_9770,N_9441);
nand UO_1024 (O_1024,N_9899,N_9430);
nor UO_1025 (O_1025,N_9256,N_9097);
and UO_1026 (O_1026,N_9912,N_9476);
or UO_1027 (O_1027,N_9253,N_9418);
nand UO_1028 (O_1028,N_9804,N_9185);
nor UO_1029 (O_1029,N_9086,N_9069);
nand UO_1030 (O_1030,N_9611,N_9261);
or UO_1031 (O_1031,N_9962,N_9605);
and UO_1032 (O_1032,N_9574,N_9968);
and UO_1033 (O_1033,N_9009,N_9281);
and UO_1034 (O_1034,N_9055,N_9209);
nand UO_1035 (O_1035,N_9962,N_9293);
nand UO_1036 (O_1036,N_9134,N_9531);
and UO_1037 (O_1037,N_9331,N_9021);
and UO_1038 (O_1038,N_9159,N_9307);
nand UO_1039 (O_1039,N_9257,N_9611);
nand UO_1040 (O_1040,N_9736,N_9232);
and UO_1041 (O_1041,N_9717,N_9744);
nor UO_1042 (O_1042,N_9025,N_9501);
or UO_1043 (O_1043,N_9930,N_9918);
or UO_1044 (O_1044,N_9274,N_9641);
xnor UO_1045 (O_1045,N_9774,N_9938);
nor UO_1046 (O_1046,N_9068,N_9668);
or UO_1047 (O_1047,N_9894,N_9853);
or UO_1048 (O_1048,N_9125,N_9831);
or UO_1049 (O_1049,N_9315,N_9352);
nor UO_1050 (O_1050,N_9784,N_9835);
nor UO_1051 (O_1051,N_9810,N_9102);
or UO_1052 (O_1052,N_9393,N_9678);
nand UO_1053 (O_1053,N_9353,N_9351);
and UO_1054 (O_1054,N_9028,N_9932);
nor UO_1055 (O_1055,N_9171,N_9322);
or UO_1056 (O_1056,N_9464,N_9503);
nand UO_1057 (O_1057,N_9987,N_9913);
or UO_1058 (O_1058,N_9004,N_9227);
nand UO_1059 (O_1059,N_9975,N_9369);
or UO_1060 (O_1060,N_9623,N_9448);
nor UO_1061 (O_1061,N_9208,N_9122);
nand UO_1062 (O_1062,N_9788,N_9400);
and UO_1063 (O_1063,N_9958,N_9357);
nand UO_1064 (O_1064,N_9658,N_9555);
and UO_1065 (O_1065,N_9752,N_9095);
nor UO_1066 (O_1066,N_9915,N_9535);
and UO_1067 (O_1067,N_9761,N_9023);
and UO_1068 (O_1068,N_9259,N_9397);
nor UO_1069 (O_1069,N_9716,N_9068);
or UO_1070 (O_1070,N_9153,N_9579);
or UO_1071 (O_1071,N_9217,N_9442);
and UO_1072 (O_1072,N_9119,N_9290);
and UO_1073 (O_1073,N_9493,N_9341);
or UO_1074 (O_1074,N_9841,N_9890);
or UO_1075 (O_1075,N_9313,N_9026);
and UO_1076 (O_1076,N_9598,N_9720);
and UO_1077 (O_1077,N_9462,N_9688);
and UO_1078 (O_1078,N_9702,N_9085);
or UO_1079 (O_1079,N_9282,N_9875);
xor UO_1080 (O_1080,N_9655,N_9938);
nor UO_1081 (O_1081,N_9925,N_9332);
and UO_1082 (O_1082,N_9224,N_9592);
nand UO_1083 (O_1083,N_9105,N_9712);
nor UO_1084 (O_1084,N_9763,N_9118);
nand UO_1085 (O_1085,N_9467,N_9871);
nand UO_1086 (O_1086,N_9363,N_9251);
xnor UO_1087 (O_1087,N_9926,N_9612);
and UO_1088 (O_1088,N_9028,N_9077);
nor UO_1089 (O_1089,N_9569,N_9071);
nand UO_1090 (O_1090,N_9899,N_9649);
and UO_1091 (O_1091,N_9217,N_9925);
or UO_1092 (O_1092,N_9711,N_9684);
nor UO_1093 (O_1093,N_9853,N_9486);
nand UO_1094 (O_1094,N_9287,N_9202);
and UO_1095 (O_1095,N_9395,N_9425);
nor UO_1096 (O_1096,N_9608,N_9549);
nand UO_1097 (O_1097,N_9970,N_9530);
and UO_1098 (O_1098,N_9590,N_9705);
and UO_1099 (O_1099,N_9206,N_9551);
or UO_1100 (O_1100,N_9685,N_9351);
or UO_1101 (O_1101,N_9369,N_9948);
nand UO_1102 (O_1102,N_9528,N_9822);
nand UO_1103 (O_1103,N_9733,N_9597);
nand UO_1104 (O_1104,N_9714,N_9101);
or UO_1105 (O_1105,N_9232,N_9048);
xnor UO_1106 (O_1106,N_9179,N_9720);
nor UO_1107 (O_1107,N_9488,N_9209);
or UO_1108 (O_1108,N_9340,N_9625);
and UO_1109 (O_1109,N_9490,N_9547);
or UO_1110 (O_1110,N_9789,N_9479);
or UO_1111 (O_1111,N_9262,N_9901);
nor UO_1112 (O_1112,N_9319,N_9077);
nand UO_1113 (O_1113,N_9464,N_9022);
and UO_1114 (O_1114,N_9864,N_9852);
and UO_1115 (O_1115,N_9999,N_9231);
or UO_1116 (O_1116,N_9040,N_9018);
nand UO_1117 (O_1117,N_9591,N_9487);
and UO_1118 (O_1118,N_9376,N_9321);
nand UO_1119 (O_1119,N_9828,N_9273);
or UO_1120 (O_1120,N_9140,N_9891);
or UO_1121 (O_1121,N_9484,N_9256);
xnor UO_1122 (O_1122,N_9903,N_9397);
nor UO_1123 (O_1123,N_9290,N_9515);
and UO_1124 (O_1124,N_9246,N_9508);
nand UO_1125 (O_1125,N_9182,N_9415);
nor UO_1126 (O_1126,N_9008,N_9565);
and UO_1127 (O_1127,N_9046,N_9833);
or UO_1128 (O_1128,N_9067,N_9511);
or UO_1129 (O_1129,N_9474,N_9523);
or UO_1130 (O_1130,N_9241,N_9848);
nand UO_1131 (O_1131,N_9807,N_9671);
nor UO_1132 (O_1132,N_9456,N_9044);
nor UO_1133 (O_1133,N_9176,N_9318);
nor UO_1134 (O_1134,N_9698,N_9131);
nor UO_1135 (O_1135,N_9940,N_9988);
nor UO_1136 (O_1136,N_9036,N_9121);
nor UO_1137 (O_1137,N_9328,N_9788);
nand UO_1138 (O_1138,N_9252,N_9167);
nor UO_1139 (O_1139,N_9163,N_9931);
nand UO_1140 (O_1140,N_9808,N_9197);
and UO_1141 (O_1141,N_9913,N_9453);
and UO_1142 (O_1142,N_9077,N_9058);
nand UO_1143 (O_1143,N_9854,N_9431);
nor UO_1144 (O_1144,N_9882,N_9483);
or UO_1145 (O_1145,N_9573,N_9811);
nor UO_1146 (O_1146,N_9086,N_9088);
xor UO_1147 (O_1147,N_9433,N_9437);
and UO_1148 (O_1148,N_9817,N_9280);
nor UO_1149 (O_1149,N_9258,N_9368);
nor UO_1150 (O_1150,N_9698,N_9192);
nand UO_1151 (O_1151,N_9519,N_9491);
and UO_1152 (O_1152,N_9167,N_9327);
nand UO_1153 (O_1153,N_9443,N_9890);
nand UO_1154 (O_1154,N_9816,N_9075);
nand UO_1155 (O_1155,N_9899,N_9938);
and UO_1156 (O_1156,N_9440,N_9625);
or UO_1157 (O_1157,N_9712,N_9196);
xnor UO_1158 (O_1158,N_9948,N_9544);
nand UO_1159 (O_1159,N_9966,N_9769);
nand UO_1160 (O_1160,N_9664,N_9293);
nand UO_1161 (O_1161,N_9737,N_9076);
nor UO_1162 (O_1162,N_9265,N_9593);
or UO_1163 (O_1163,N_9053,N_9097);
nand UO_1164 (O_1164,N_9547,N_9689);
nand UO_1165 (O_1165,N_9935,N_9096);
xnor UO_1166 (O_1166,N_9695,N_9395);
nor UO_1167 (O_1167,N_9792,N_9417);
or UO_1168 (O_1168,N_9464,N_9226);
nor UO_1169 (O_1169,N_9263,N_9137);
nor UO_1170 (O_1170,N_9143,N_9257);
or UO_1171 (O_1171,N_9027,N_9860);
nor UO_1172 (O_1172,N_9498,N_9106);
or UO_1173 (O_1173,N_9339,N_9389);
nor UO_1174 (O_1174,N_9954,N_9228);
nand UO_1175 (O_1175,N_9706,N_9027);
nand UO_1176 (O_1176,N_9288,N_9100);
or UO_1177 (O_1177,N_9221,N_9781);
or UO_1178 (O_1178,N_9032,N_9678);
nand UO_1179 (O_1179,N_9143,N_9118);
or UO_1180 (O_1180,N_9702,N_9990);
and UO_1181 (O_1181,N_9904,N_9539);
nor UO_1182 (O_1182,N_9815,N_9935);
nor UO_1183 (O_1183,N_9785,N_9536);
or UO_1184 (O_1184,N_9809,N_9634);
xnor UO_1185 (O_1185,N_9393,N_9782);
nor UO_1186 (O_1186,N_9474,N_9695);
and UO_1187 (O_1187,N_9805,N_9305);
nand UO_1188 (O_1188,N_9813,N_9966);
nor UO_1189 (O_1189,N_9280,N_9708);
nor UO_1190 (O_1190,N_9608,N_9423);
nor UO_1191 (O_1191,N_9017,N_9028);
and UO_1192 (O_1192,N_9292,N_9251);
or UO_1193 (O_1193,N_9537,N_9736);
or UO_1194 (O_1194,N_9744,N_9389);
and UO_1195 (O_1195,N_9011,N_9767);
and UO_1196 (O_1196,N_9213,N_9741);
xnor UO_1197 (O_1197,N_9884,N_9174);
or UO_1198 (O_1198,N_9403,N_9148);
nor UO_1199 (O_1199,N_9502,N_9565);
and UO_1200 (O_1200,N_9291,N_9838);
nor UO_1201 (O_1201,N_9401,N_9227);
or UO_1202 (O_1202,N_9473,N_9505);
xor UO_1203 (O_1203,N_9874,N_9643);
nand UO_1204 (O_1204,N_9289,N_9643);
nand UO_1205 (O_1205,N_9823,N_9959);
nor UO_1206 (O_1206,N_9447,N_9050);
nand UO_1207 (O_1207,N_9270,N_9870);
nor UO_1208 (O_1208,N_9342,N_9667);
nor UO_1209 (O_1209,N_9925,N_9509);
nand UO_1210 (O_1210,N_9077,N_9486);
or UO_1211 (O_1211,N_9586,N_9946);
or UO_1212 (O_1212,N_9807,N_9501);
or UO_1213 (O_1213,N_9428,N_9448);
and UO_1214 (O_1214,N_9045,N_9626);
nor UO_1215 (O_1215,N_9222,N_9477);
or UO_1216 (O_1216,N_9921,N_9327);
nor UO_1217 (O_1217,N_9257,N_9540);
nor UO_1218 (O_1218,N_9504,N_9542);
xnor UO_1219 (O_1219,N_9808,N_9684);
and UO_1220 (O_1220,N_9127,N_9311);
nor UO_1221 (O_1221,N_9089,N_9447);
xor UO_1222 (O_1222,N_9886,N_9873);
or UO_1223 (O_1223,N_9048,N_9251);
nor UO_1224 (O_1224,N_9671,N_9762);
nor UO_1225 (O_1225,N_9497,N_9095);
nand UO_1226 (O_1226,N_9854,N_9619);
or UO_1227 (O_1227,N_9699,N_9961);
nor UO_1228 (O_1228,N_9904,N_9179);
nor UO_1229 (O_1229,N_9907,N_9015);
nor UO_1230 (O_1230,N_9522,N_9268);
and UO_1231 (O_1231,N_9338,N_9845);
nor UO_1232 (O_1232,N_9888,N_9018);
nor UO_1233 (O_1233,N_9969,N_9433);
nor UO_1234 (O_1234,N_9258,N_9909);
nand UO_1235 (O_1235,N_9971,N_9935);
nor UO_1236 (O_1236,N_9982,N_9650);
and UO_1237 (O_1237,N_9211,N_9426);
and UO_1238 (O_1238,N_9147,N_9849);
nand UO_1239 (O_1239,N_9458,N_9860);
and UO_1240 (O_1240,N_9342,N_9528);
or UO_1241 (O_1241,N_9469,N_9103);
nand UO_1242 (O_1242,N_9826,N_9983);
nor UO_1243 (O_1243,N_9752,N_9953);
nor UO_1244 (O_1244,N_9269,N_9643);
xor UO_1245 (O_1245,N_9921,N_9287);
and UO_1246 (O_1246,N_9869,N_9956);
nor UO_1247 (O_1247,N_9944,N_9539);
nor UO_1248 (O_1248,N_9068,N_9108);
nor UO_1249 (O_1249,N_9150,N_9303);
and UO_1250 (O_1250,N_9443,N_9882);
nand UO_1251 (O_1251,N_9727,N_9927);
nand UO_1252 (O_1252,N_9068,N_9959);
nor UO_1253 (O_1253,N_9652,N_9415);
or UO_1254 (O_1254,N_9219,N_9942);
nand UO_1255 (O_1255,N_9993,N_9720);
nand UO_1256 (O_1256,N_9637,N_9043);
and UO_1257 (O_1257,N_9820,N_9669);
and UO_1258 (O_1258,N_9054,N_9947);
xnor UO_1259 (O_1259,N_9850,N_9287);
nor UO_1260 (O_1260,N_9585,N_9296);
nand UO_1261 (O_1261,N_9723,N_9215);
nor UO_1262 (O_1262,N_9582,N_9000);
nor UO_1263 (O_1263,N_9707,N_9899);
nand UO_1264 (O_1264,N_9711,N_9382);
and UO_1265 (O_1265,N_9638,N_9026);
nor UO_1266 (O_1266,N_9863,N_9034);
nor UO_1267 (O_1267,N_9064,N_9217);
nand UO_1268 (O_1268,N_9508,N_9252);
and UO_1269 (O_1269,N_9599,N_9924);
xor UO_1270 (O_1270,N_9923,N_9674);
nor UO_1271 (O_1271,N_9202,N_9820);
or UO_1272 (O_1272,N_9743,N_9908);
and UO_1273 (O_1273,N_9534,N_9087);
or UO_1274 (O_1274,N_9796,N_9016);
nand UO_1275 (O_1275,N_9715,N_9451);
nor UO_1276 (O_1276,N_9906,N_9130);
nand UO_1277 (O_1277,N_9439,N_9871);
and UO_1278 (O_1278,N_9728,N_9509);
nor UO_1279 (O_1279,N_9217,N_9879);
nand UO_1280 (O_1280,N_9494,N_9674);
or UO_1281 (O_1281,N_9026,N_9490);
nor UO_1282 (O_1282,N_9134,N_9078);
and UO_1283 (O_1283,N_9156,N_9554);
nor UO_1284 (O_1284,N_9333,N_9159);
nor UO_1285 (O_1285,N_9746,N_9436);
or UO_1286 (O_1286,N_9957,N_9210);
nand UO_1287 (O_1287,N_9095,N_9983);
and UO_1288 (O_1288,N_9431,N_9218);
and UO_1289 (O_1289,N_9882,N_9972);
or UO_1290 (O_1290,N_9957,N_9126);
nor UO_1291 (O_1291,N_9014,N_9411);
or UO_1292 (O_1292,N_9076,N_9253);
or UO_1293 (O_1293,N_9770,N_9382);
xnor UO_1294 (O_1294,N_9568,N_9672);
or UO_1295 (O_1295,N_9119,N_9023);
nor UO_1296 (O_1296,N_9426,N_9133);
nor UO_1297 (O_1297,N_9723,N_9849);
and UO_1298 (O_1298,N_9677,N_9292);
xor UO_1299 (O_1299,N_9546,N_9931);
or UO_1300 (O_1300,N_9738,N_9874);
nor UO_1301 (O_1301,N_9357,N_9844);
nor UO_1302 (O_1302,N_9573,N_9804);
nor UO_1303 (O_1303,N_9443,N_9364);
nand UO_1304 (O_1304,N_9436,N_9680);
nand UO_1305 (O_1305,N_9128,N_9345);
xor UO_1306 (O_1306,N_9018,N_9775);
and UO_1307 (O_1307,N_9075,N_9635);
nor UO_1308 (O_1308,N_9017,N_9044);
nand UO_1309 (O_1309,N_9843,N_9269);
or UO_1310 (O_1310,N_9361,N_9939);
or UO_1311 (O_1311,N_9705,N_9038);
and UO_1312 (O_1312,N_9481,N_9442);
nor UO_1313 (O_1313,N_9518,N_9728);
nand UO_1314 (O_1314,N_9423,N_9817);
nor UO_1315 (O_1315,N_9043,N_9479);
nor UO_1316 (O_1316,N_9250,N_9900);
xor UO_1317 (O_1317,N_9022,N_9057);
nor UO_1318 (O_1318,N_9113,N_9663);
and UO_1319 (O_1319,N_9851,N_9381);
and UO_1320 (O_1320,N_9257,N_9300);
and UO_1321 (O_1321,N_9608,N_9852);
and UO_1322 (O_1322,N_9099,N_9238);
xor UO_1323 (O_1323,N_9334,N_9656);
xnor UO_1324 (O_1324,N_9619,N_9768);
and UO_1325 (O_1325,N_9981,N_9587);
nand UO_1326 (O_1326,N_9965,N_9526);
and UO_1327 (O_1327,N_9861,N_9130);
nor UO_1328 (O_1328,N_9956,N_9203);
and UO_1329 (O_1329,N_9206,N_9850);
xnor UO_1330 (O_1330,N_9381,N_9482);
nand UO_1331 (O_1331,N_9591,N_9195);
or UO_1332 (O_1332,N_9460,N_9751);
xnor UO_1333 (O_1333,N_9617,N_9660);
and UO_1334 (O_1334,N_9781,N_9249);
nor UO_1335 (O_1335,N_9750,N_9461);
or UO_1336 (O_1336,N_9337,N_9974);
and UO_1337 (O_1337,N_9392,N_9371);
and UO_1338 (O_1338,N_9655,N_9241);
nand UO_1339 (O_1339,N_9589,N_9083);
or UO_1340 (O_1340,N_9164,N_9341);
and UO_1341 (O_1341,N_9686,N_9826);
nand UO_1342 (O_1342,N_9182,N_9117);
nand UO_1343 (O_1343,N_9618,N_9478);
nor UO_1344 (O_1344,N_9149,N_9989);
nand UO_1345 (O_1345,N_9717,N_9871);
and UO_1346 (O_1346,N_9070,N_9708);
and UO_1347 (O_1347,N_9607,N_9539);
nand UO_1348 (O_1348,N_9323,N_9134);
nand UO_1349 (O_1349,N_9848,N_9559);
nor UO_1350 (O_1350,N_9059,N_9402);
or UO_1351 (O_1351,N_9667,N_9452);
nand UO_1352 (O_1352,N_9869,N_9588);
or UO_1353 (O_1353,N_9784,N_9995);
nor UO_1354 (O_1354,N_9960,N_9735);
nand UO_1355 (O_1355,N_9183,N_9810);
nand UO_1356 (O_1356,N_9581,N_9009);
xnor UO_1357 (O_1357,N_9906,N_9044);
xor UO_1358 (O_1358,N_9990,N_9001);
nor UO_1359 (O_1359,N_9847,N_9909);
xor UO_1360 (O_1360,N_9718,N_9732);
and UO_1361 (O_1361,N_9830,N_9337);
and UO_1362 (O_1362,N_9848,N_9836);
nand UO_1363 (O_1363,N_9022,N_9456);
or UO_1364 (O_1364,N_9080,N_9684);
xor UO_1365 (O_1365,N_9483,N_9349);
nor UO_1366 (O_1366,N_9980,N_9280);
nand UO_1367 (O_1367,N_9783,N_9939);
nand UO_1368 (O_1368,N_9820,N_9924);
and UO_1369 (O_1369,N_9438,N_9636);
nand UO_1370 (O_1370,N_9303,N_9510);
nor UO_1371 (O_1371,N_9072,N_9029);
nor UO_1372 (O_1372,N_9980,N_9918);
nor UO_1373 (O_1373,N_9253,N_9516);
or UO_1374 (O_1374,N_9601,N_9644);
nor UO_1375 (O_1375,N_9824,N_9572);
nor UO_1376 (O_1376,N_9953,N_9324);
nor UO_1377 (O_1377,N_9064,N_9904);
or UO_1378 (O_1378,N_9171,N_9279);
xor UO_1379 (O_1379,N_9185,N_9038);
nor UO_1380 (O_1380,N_9874,N_9758);
xnor UO_1381 (O_1381,N_9136,N_9939);
nand UO_1382 (O_1382,N_9332,N_9441);
and UO_1383 (O_1383,N_9694,N_9277);
xor UO_1384 (O_1384,N_9922,N_9921);
xor UO_1385 (O_1385,N_9242,N_9714);
and UO_1386 (O_1386,N_9876,N_9010);
nand UO_1387 (O_1387,N_9156,N_9909);
nand UO_1388 (O_1388,N_9665,N_9339);
and UO_1389 (O_1389,N_9619,N_9542);
nand UO_1390 (O_1390,N_9527,N_9561);
and UO_1391 (O_1391,N_9931,N_9274);
nand UO_1392 (O_1392,N_9687,N_9198);
and UO_1393 (O_1393,N_9421,N_9955);
nand UO_1394 (O_1394,N_9773,N_9146);
nor UO_1395 (O_1395,N_9426,N_9206);
nand UO_1396 (O_1396,N_9141,N_9923);
nand UO_1397 (O_1397,N_9414,N_9431);
nor UO_1398 (O_1398,N_9827,N_9312);
nand UO_1399 (O_1399,N_9020,N_9969);
nor UO_1400 (O_1400,N_9794,N_9933);
and UO_1401 (O_1401,N_9615,N_9256);
or UO_1402 (O_1402,N_9154,N_9028);
and UO_1403 (O_1403,N_9913,N_9333);
or UO_1404 (O_1404,N_9162,N_9243);
nand UO_1405 (O_1405,N_9618,N_9453);
and UO_1406 (O_1406,N_9981,N_9470);
and UO_1407 (O_1407,N_9577,N_9034);
xor UO_1408 (O_1408,N_9330,N_9877);
nor UO_1409 (O_1409,N_9413,N_9492);
nand UO_1410 (O_1410,N_9308,N_9629);
or UO_1411 (O_1411,N_9722,N_9914);
and UO_1412 (O_1412,N_9126,N_9705);
nand UO_1413 (O_1413,N_9698,N_9500);
and UO_1414 (O_1414,N_9236,N_9738);
nor UO_1415 (O_1415,N_9940,N_9458);
and UO_1416 (O_1416,N_9064,N_9294);
nand UO_1417 (O_1417,N_9227,N_9820);
nand UO_1418 (O_1418,N_9888,N_9260);
xor UO_1419 (O_1419,N_9387,N_9272);
xor UO_1420 (O_1420,N_9262,N_9799);
or UO_1421 (O_1421,N_9764,N_9312);
and UO_1422 (O_1422,N_9790,N_9347);
nand UO_1423 (O_1423,N_9062,N_9994);
nand UO_1424 (O_1424,N_9944,N_9011);
and UO_1425 (O_1425,N_9590,N_9594);
and UO_1426 (O_1426,N_9270,N_9934);
or UO_1427 (O_1427,N_9968,N_9339);
xnor UO_1428 (O_1428,N_9565,N_9538);
nor UO_1429 (O_1429,N_9122,N_9002);
and UO_1430 (O_1430,N_9690,N_9976);
nand UO_1431 (O_1431,N_9865,N_9308);
nor UO_1432 (O_1432,N_9824,N_9003);
nor UO_1433 (O_1433,N_9248,N_9980);
nor UO_1434 (O_1434,N_9309,N_9829);
nand UO_1435 (O_1435,N_9517,N_9143);
nor UO_1436 (O_1436,N_9692,N_9211);
nand UO_1437 (O_1437,N_9532,N_9811);
and UO_1438 (O_1438,N_9846,N_9241);
nor UO_1439 (O_1439,N_9977,N_9576);
xor UO_1440 (O_1440,N_9113,N_9356);
nor UO_1441 (O_1441,N_9257,N_9310);
nand UO_1442 (O_1442,N_9502,N_9507);
and UO_1443 (O_1443,N_9992,N_9789);
and UO_1444 (O_1444,N_9137,N_9194);
xnor UO_1445 (O_1445,N_9756,N_9180);
or UO_1446 (O_1446,N_9222,N_9512);
nor UO_1447 (O_1447,N_9953,N_9731);
nor UO_1448 (O_1448,N_9814,N_9906);
nor UO_1449 (O_1449,N_9655,N_9209);
or UO_1450 (O_1450,N_9546,N_9080);
nand UO_1451 (O_1451,N_9448,N_9838);
nor UO_1452 (O_1452,N_9419,N_9048);
nand UO_1453 (O_1453,N_9132,N_9117);
or UO_1454 (O_1454,N_9566,N_9803);
or UO_1455 (O_1455,N_9162,N_9722);
and UO_1456 (O_1456,N_9300,N_9395);
nand UO_1457 (O_1457,N_9877,N_9217);
nand UO_1458 (O_1458,N_9707,N_9790);
nor UO_1459 (O_1459,N_9551,N_9294);
nand UO_1460 (O_1460,N_9285,N_9838);
xnor UO_1461 (O_1461,N_9151,N_9736);
xnor UO_1462 (O_1462,N_9545,N_9059);
nor UO_1463 (O_1463,N_9548,N_9167);
nor UO_1464 (O_1464,N_9924,N_9098);
nand UO_1465 (O_1465,N_9445,N_9174);
nand UO_1466 (O_1466,N_9722,N_9986);
nand UO_1467 (O_1467,N_9026,N_9043);
nand UO_1468 (O_1468,N_9961,N_9850);
and UO_1469 (O_1469,N_9640,N_9998);
nor UO_1470 (O_1470,N_9488,N_9779);
or UO_1471 (O_1471,N_9126,N_9731);
and UO_1472 (O_1472,N_9170,N_9968);
or UO_1473 (O_1473,N_9302,N_9608);
and UO_1474 (O_1474,N_9887,N_9088);
xnor UO_1475 (O_1475,N_9964,N_9424);
or UO_1476 (O_1476,N_9738,N_9026);
or UO_1477 (O_1477,N_9675,N_9310);
xor UO_1478 (O_1478,N_9582,N_9349);
nand UO_1479 (O_1479,N_9257,N_9813);
nor UO_1480 (O_1480,N_9116,N_9559);
nor UO_1481 (O_1481,N_9920,N_9881);
or UO_1482 (O_1482,N_9451,N_9765);
nand UO_1483 (O_1483,N_9615,N_9892);
xor UO_1484 (O_1484,N_9545,N_9690);
or UO_1485 (O_1485,N_9490,N_9283);
or UO_1486 (O_1486,N_9588,N_9284);
or UO_1487 (O_1487,N_9271,N_9692);
and UO_1488 (O_1488,N_9037,N_9938);
and UO_1489 (O_1489,N_9279,N_9893);
or UO_1490 (O_1490,N_9511,N_9541);
nor UO_1491 (O_1491,N_9219,N_9770);
nor UO_1492 (O_1492,N_9657,N_9089);
and UO_1493 (O_1493,N_9673,N_9956);
or UO_1494 (O_1494,N_9283,N_9503);
or UO_1495 (O_1495,N_9037,N_9109);
or UO_1496 (O_1496,N_9333,N_9234);
nor UO_1497 (O_1497,N_9132,N_9096);
xnor UO_1498 (O_1498,N_9084,N_9767);
nor UO_1499 (O_1499,N_9679,N_9152);
endmodule