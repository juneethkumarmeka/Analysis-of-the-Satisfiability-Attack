module basic_500_3000_500_15_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_219,In_416);
xor U1 (N_1,In_371,In_124);
nor U2 (N_2,In_201,In_100);
or U3 (N_3,In_482,In_128);
nor U4 (N_4,In_208,In_277);
and U5 (N_5,In_391,In_260);
nand U6 (N_6,In_339,In_424);
or U7 (N_7,In_334,In_417);
and U8 (N_8,In_419,In_269);
xnor U9 (N_9,In_303,In_394);
nor U10 (N_10,In_93,In_484);
and U11 (N_11,In_478,In_18);
nor U12 (N_12,In_171,In_400);
nand U13 (N_13,In_425,In_249);
xor U14 (N_14,In_163,In_407);
and U15 (N_15,In_215,In_69);
and U16 (N_16,In_200,In_228);
nor U17 (N_17,In_483,In_396);
and U18 (N_18,In_42,In_57);
nand U19 (N_19,In_469,In_19);
and U20 (N_20,In_265,In_467);
or U21 (N_21,In_236,In_241);
and U22 (N_22,In_49,In_178);
nand U23 (N_23,In_248,In_452);
nand U24 (N_24,In_133,In_488);
nor U25 (N_25,In_312,In_86);
xor U26 (N_26,In_109,In_14);
and U27 (N_27,In_287,In_311);
nor U28 (N_28,In_496,In_186);
xor U29 (N_29,In_237,In_43);
xnor U30 (N_30,In_121,In_472);
or U31 (N_31,In_390,In_7);
xnor U32 (N_32,In_380,In_24);
xnor U33 (N_33,In_62,In_113);
nand U34 (N_34,In_214,In_91);
and U35 (N_35,In_145,In_261);
nand U36 (N_36,In_354,In_232);
nand U37 (N_37,In_479,In_205);
and U38 (N_38,In_358,In_310);
nand U39 (N_39,In_323,In_130);
and U40 (N_40,In_92,In_392);
nand U41 (N_41,In_460,In_383);
nor U42 (N_42,In_397,In_209);
and U43 (N_43,In_0,In_111);
nand U44 (N_44,In_393,In_387);
or U45 (N_45,In_17,In_430);
nor U46 (N_46,In_435,In_78);
and U47 (N_47,In_363,In_247);
or U48 (N_48,In_355,In_122);
xnor U49 (N_49,In_444,In_262);
nor U50 (N_50,In_218,In_436);
nand U51 (N_51,In_448,In_26);
nand U52 (N_52,In_487,In_217);
or U53 (N_53,In_70,In_67);
nor U54 (N_54,In_333,In_348);
xor U55 (N_55,In_212,In_153);
nor U56 (N_56,In_254,In_96);
nor U57 (N_57,In_377,In_8);
xor U58 (N_58,In_114,In_389);
or U59 (N_59,In_41,In_313);
nand U60 (N_60,In_495,In_328);
and U61 (N_61,In_188,In_319);
xnor U62 (N_62,In_224,In_335);
nand U63 (N_63,In_330,In_169);
xor U64 (N_64,In_280,In_149);
nor U65 (N_65,In_192,In_183);
or U66 (N_66,In_221,In_185);
xor U67 (N_67,In_30,In_85);
nor U68 (N_68,In_88,In_459);
nand U69 (N_69,In_369,In_252);
or U70 (N_70,In_167,In_83);
and U71 (N_71,In_464,In_320);
xnor U72 (N_72,In_256,In_471);
nand U73 (N_73,In_61,In_158);
nand U74 (N_74,In_284,In_184);
or U75 (N_75,In_204,In_53);
xnor U76 (N_76,In_21,In_47);
xnor U77 (N_77,In_272,In_152);
xor U78 (N_78,In_409,In_31);
or U79 (N_79,In_292,In_118);
and U80 (N_80,In_197,In_54);
nor U81 (N_81,In_90,In_418);
nor U82 (N_82,In_9,In_338);
nand U83 (N_83,In_125,In_266);
and U84 (N_84,In_162,In_202);
nand U85 (N_85,In_33,In_3);
nor U86 (N_86,In_422,In_140);
and U87 (N_87,In_139,In_71);
xor U88 (N_88,In_456,In_494);
xor U89 (N_89,In_365,In_263);
nand U90 (N_90,In_300,In_443);
nand U91 (N_91,In_28,In_58);
nor U92 (N_92,In_246,In_203);
nor U93 (N_93,In_108,In_147);
xor U94 (N_94,In_485,In_6);
or U95 (N_95,In_274,In_308);
nand U96 (N_96,In_326,In_412);
and U97 (N_97,In_293,In_322);
or U98 (N_98,In_314,In_89);
xnor U99 (N_99,In_492,In_229);
xnor U100 (N_100,In_198,In_259);
and U101 (N_101,In_361,In_136);
nand U102 (N_102,In_127,In_131);
xor U103 (N_103,In_283,In_276);
xor U104 (N_104,In_65,In_156);
nor U105 (N_105,In_1,In_309);
or U106 (N_106,In_376,In_220);
xor U107 (N_107,In_325,In_110);
nand U108 (N_108,In_141,In_350);
nor U109 (N_109,In_150,In_196);
xnor U110 (N_110,In_135,In_170);
and U111 (N_111,In_332,In_279);
xor U112 (N_112,In_429,In_63);
nand U113 (N_113,In_123,In_480);
nand U114 (N_114,In_102,In_51);
nand U115 (N_115,In_231,In_275);
and U116 (N_116,In_404,In_362);
nand U117 (N_117,In_45,In_420);
nand U118 (N_118,In_98,In_405);
nor U119 (N_119,In_81,In_164);
nor U120 (N_120,In_427,In_129);
xor U121 (N_121,In_367,In_455);
nor U122 (N_122,In_336,In_445);
xor U123 (N_123,In_306,In_37);
or U124 (N_124,In_281,In_408);
and U125 (N_125,In_120,In_402);
xor U126 (N_126,In_352,In_449);
or U127 (N_127,In_321,In_301);
xor U128 (N_128,In_395,In_79);
and U129 (N_129,In_453,In_16);
nand U130 (N_130,In_59,In_52);
nor U131 (N_131,In_75,In_193);
xnor U132 (N_132,In_490,In_251);
nor U133 (N_133,In_257,In_493);
or U134 (N_134,In_375,In_77);
xnor U135 (N_135,In_34,In_182);
and U136 (N_136,In_11,In_491);
or U137 (N_137,In_398,In_366);
xnor U138 (N_138,In_25,In_437);
xor U139 (N_139,In_433,In_465);
or U140 (N_140,In_142,In_337);
and U141 (N_141,In_466,In_373);
or U142 (N_142,In_50,In_97);
xor U143 (N_143,In_116,In_32);
xnor U144 (N_144,In_438,In_174);
nand U145 (N_145,In_76,In_39);
xnor U146 (N_146,In_225,In_144);
nand U147 (N_147,In_357,In_137);
nor U148 (N_148,In_415,In_381);
and U149 (N_149,In_173,In_372);
nand U150 (N_150,In_329,In_382);
xor U151 (N_151,In_233,In_119);
nor U152 (N_152,In_187,In_5);
xnor U153 (N_153,In_27,In_454);
nor U154 (N_154,In_195,In_44);
nor U155 (N_155,In_294,In_457);
and U156 (N_156,In_344,In_399);
xor U157 (N_157,In_160,In_264);
nand U158 (N_158,In_99,In_177);
or U159 (N_159,In_489,In_331);
and U160 (N_160,In_349,In_370);
nor U161 (N_161,In_305,In_179);
nor U162 (N_162,In_48,In_406);
nor U163 (N_163,In_106,In_72);
xnor U164 (N_164,In_166,In_288);
xor U165 (N_165,In_290,In_413);
xor U166 (N_166,In_181,In_286);
nor U167 (N_167,In_298,In_296);
nor U168 (N_168,In_403,In_268);
nand U169 (N_169,In_428,In_38);
or U170 (N_170,In_35,In_258);
and U171 (N_171,In_473,In_213);
nand U172 (N_172,In_64,In_346);
nand U173 (N_173,In_15,In_84);
nor U174 (N_174,In_476,In_388);
nand U175 (N_175,In_463,In_324);
nor U176 (N_176,In_176,In_60);
xor U177 (N_177,In_107,In_384);
nand U178 (N_178,In_240,In_230);
nor U179 (N_179,In_441,In_12);
or U180 (N_180,In_22,In_80);
xnor U181 (N_181,In_235,In_447);
nor U182 (N_182,In_56,In_359);
nor U183 (N_183,In_253,In_434);
nand U184 (N_184,In_289,In_104);
nand U185 (N_185,In_304,In_4);
nor U186 (N_186,In_112,In_317);
nor U187 (N_187,In_87,In_159);
nor U188 (N_188,In_411,In_55);
xor U189 (N_189,In_341,In_73);
or U190 (N_190,In_23,In_285);
and U191 (N_191,In_343,In_401);
xnor U192 (N_192,In_295,In_497);
nand U193 (N_193,In_134,In_297);
and U194 (N_194,In_29,In_327);
xnor U195 (N_195,In_345,In_481);
nand U196 (N_196,In_442,In_316);
nor U197 (N_197,In_347,In_82);
xor U198 (N_198,In_199,In_175);
nand U199 (N_199,In_191,In_103);
nor U200 (N_200,N_22,N_91);
and U201 (N_201,N_142,N_199);
xor U202 (N_202,N_51,In_271);
nor U203 (N_203,N_43,In_94);
nand U204 (N_204,In_440,N_143);
nand U205 (N_205,N_170,N_118);
and U206 (N_206,In_172,In_273);
nor U207 (N_207,In_499,In_475);
nor U208 (N_208,N_144,In_207);
and U209 (N_209,N_181,N_8);
and U210 (N_210,N_50,In_374);
or U211 (N_211,N_96,N_150);
xnor U212 (N_212,N_17,In_210);
nand U213 (N_213,In_66,In_216);
nor U214 (N_214,In_368,N_28);
nor U215 (N_215,In_117,N_115);
nand U216 (N_216,N_134,N_110);
xor U217 (N_217,In_46,In_244);
or U218 (N_218,N_80,In_386);
and U219 (N_219,N_139,In_356);
nor U220 (N_220,N_78,N_158);
xnor U221 (N_221,N_145,N_123);
and U222 (N_222,In_155,N_178);
or U223 (N_223,In_2,N_183);
and U224 (N_224,In_138,N_193);
or U225 (N_225,In_161,N_186);
nand U226 (N_226,N_55,N_168);
and U227 (N_227,N_32,N_133);
xnor U228 (N_228,N_138,In_105);
nor U229 (N_229,N_14,In_364);
nor U230 (N_230,In_378,In_245);
or U231 (N_231,In_431,N_74);
xnor U232 (N_232,N_0,N_73);
and U233 (N_233,N_2,N_26);
nand U234 (N_234,N_154,N_47);
and U235 (N_235,N_173,N_169);
and U236 (N_236,N_12,N_40);
nor U237 (N_237,N_182,In_146);
xnor U238 (N_238,N_58,N_48);
nand U239 (N_239,N_180,In_379);
nand U240 (N_240,N_97,In_238);
xor U241 (N_241,N_135,N_108);
xnor U242 (N_242,In_126,N_29);
and U243 (N_243,In_474,In_189);
and U244 (N_244,N_87,In_426);
nor U245 (N_245,N_167,N_100);
and U246 (N_246,In_458,In_291);
or U247 (N_247,In_462,In_450);
and U248 (N_248,N_69,In_239);
xnor U249 (N_249,N_84,In_410);
and U250 (N_250,N_191,N_41);
nand U251 (N_251,N_157,N_4);
nor U252 (N_252,N_165,N_116);
nand U253 (N_253,N_57,In_180);
nand U254 (N_254,N_136,N_103);
and U255 (N_255,N_141,N_131);
nor U256 (N_256,N_6,In_477);
xor U257 (N_257,N_52,N_76);
nand U258 (N_258,N_152,N_90);
nand U259 (N_259,N_149,N_35);
nand U260 (N_260,N_95,In_385);
nand U261 (N_261,N_146,N_153);
nor U262 (N_262,N_163,N_162);
or U263 (N_263,In_165,N_75);
nor U264 (N_264,N_147,In_414);
and U265 (N_265,N_175,In_168);
and U266 (N_266,N_30,In_154);
or U267 (N_267,N_189,N_121);
xor U268 (N_268,N_194,In_40);
nor U269 (N_269,In_315,N_132);
and U270 (N_270,In_13,N_85);
or U271 (N_271,N_20,N_45);
nand U272 (N_272,In_223,N_11);
nand U273 (N_273,In_95,N_187);
or U274 (N_274,In_340,In_461);
and U275 (N_275,N_124,N_81);
or U276 (N_276,In_446,N_60);
and U277 (N_277,N_198,In_211);
nor U278 (N_278,N_125,N_59);
or U279 (N_279,N_195,N_172);
and U280 (N_280,In_318,N_127);
xor U281 (N_281,In_432,In_74);
nand U282 (N_282,In_353,N_19);
and U283 (N_283,N_161,N_86);
nand U284 (N_284,N_185,In_470);
or U285 (N_285,N_126,In_143);
and U286 (N_286,In_148,In_151);
or U287 (N_287,N_56,In_190);
nand U288 (N_288,N_179,N_24);
nor U289 (N_289,In_278,In_242);
nand U290 (N_290,N_9,N_106);
nand U291 (N_291,N_18,N_122);
nor U292 (N_292,In_360,N_1);
xor U293 (N_293,N_105,N_176);
nor U294 (N_294,N_174,In_20);
and U295 (N_295,N_160,N_155);
or U296 (N_296,N_104,N_190);
xnor U297 (N_297,N_62,N_89);
xor U298 (N_298,N_7,N_71);
nor U299 (N_299,N_49,N_88);
and U300 (N_300,In_243,N_21);
nor U301 (N_301,N_171,In_234);
or U302 (N_302,N_114,N_102);
and U303 (N_303,N_101,In_194);
nor U304 (N_304,In_222,In_351);
and U305 (N_305,In_302,In_68);
nor U306 (N_306,In_227,N_3);
or U307 (N_307,N_111,N_113);
and U308 (N_308,N_151,In_451);
nor U309 (N_309,N_129,N_82);
nor U310 (N_310,N_166,In_10);
xnor U311 (N_311,In_270,In_36);
nand U312 (N_312,N_23,N_63);
nand U313 (N_313,N_46,N_148);
or U314 (N_314,N_83,N_112);
xor U315 (N_315,In_226,N_34);
xnor U316 (N_316,N_5,In_423);
nand U317 (N_317,N_156,In_307);
nand U318 (N_318,N_39,N_192);
and U319 (N_319,N_196,In_439);
nor U320 (N_320,N_130,N_70);
xor U321 (N_321,N_184,N_27);
nand U322 (N_322,In_342,In_267);
or U323 (N_323,N_119,N_25);
nand U324 (N_324,N_107,In_421);
and U325 (N_325,In_157,N_93);
nand U326 (N_326,N_37,N_54);
or U327 (N_327,N_77,N_61);
xnor U328 (N_328,N_42,N_38);
nor U329 (N_329,N_177,N_66);
xnor U330 (N_330,In_255,N_117);
nor U331 (N_331,N_164,N_64);
nor U332 (N_332,N_120,N_140);
nor U333 (N_333,In_498,In_486);
xnor U334 (N_334,N_99,N_16);
nand U335 (N_335,In_101,N_68);
nand U336 (N_336,N_79,N_137);
or U337 (N_337,In_299,N_31);
and U338 (N_338,In_132,N_53);
or U339 (N_339,N_128,N_92);
or U340 (N_340,In_282,N_65);
nor U341 (N_341,In_250,N_44);
nor U342 (N_342,N_94,N_72);
xor U343 (N_343,N_33,N_188);
xnor U344 (N_344,In_468,N_13);
xor U345 (N_345,N_109,N_159);
nor U346 (N_346,In_206,N_10);
xor U347 (N_347,N_15,N_67);
nor U348 (N_348,N_36,In_115);
and U349 (N_349,N_197,N_98);
nor U350 (N_350,N_183,N_20);
xor U351 (N_351,In_498,N_11);
nor U352 (N_352,In_154,N_32);
or U353 (N_353,In_226,N_180);
nand U354 (N_354,In_126,N_44);
nand U355 (N_355,N_181,N_158);
nor U356 (N_356,In_146,N_107);
and U357 (N_357,N_118,N_31);
xnor U358 (N_358,In_227,In_157);
xor U359 (N_359,N_18,In_132);
or U360 (N_360,In_351,N_104);
and U361 (N_361,N_122,N_24);
nor U362 (N_362,N_163,In_364);
and U363 (N_363,N_163,In_95);
nor U364 (N_364,N_181,N_70);
and U365 (N_365,N_83,In_291);
nand U366 (N_366,In_95,N_154);
nand U367 (N_367,N_7,N_142);
xor U368 (N_368,N_104,N_3);
or U369 (N_369,N_28,In_216);
and U370 (N_370,N_122,N_162);
and U371 (N_371,N_10,N_171);
nor U372 (N_372,In_74,In_385);
nor U373 (N_373,N_42,N_55);
xnor U374 (N_374,N_84,In_477);
or U375 (N_375,N_116,N_22);
xnor U376 (N_376,N_39,In_216);
nor U377 (N_377,N_5,In_20);
xnor U378 (N_378,In_234,In_227);
xor U379 (N_379,N_84,N_96);
nand U380 (N_380,N_125,N_100);
or U381 (N_381,N_75,N_162);
nor U382 (N_382,N_26,N_114);
or U383 (N_383,N_163,N_190);
nor U384 (N_384,N_199,N_195);
and U385 (N_385,N_64,N_84);
nand U386 (N_386,N_6,In_161);
nor U387 (N_387,In_273,In_10);
or U388 (N_388,N_103,N_112);
xnor U389 (N_389,N_14,N_143);
or U390 (N_390,N_82,N_173);
or U391 (N_391,N_133,N_139);
nand U392 (N_392,In_342,N_154);
nand U393 (N_393,N_14,N_46);
nor U394 (N_394,In_282,In_474);
and U395 (N_395,N_163,N_75);
nand U396 (N_396,N_199,In_222);
nor U397 (N_397,N_28,In_318);
xor U398 (N_398,In_126,N_9);
or U399 (N_399,N_98,N_69);
and U400 (N_400,N_321,N_259);
nand U401 (N_401,N_232,N_227);
nand U402 (N_402,N_255,N_308);
xnor U403 (N_403,N_280,N_339);
or U404 (N_404,N_384,N_303);
nand U405 (N_405,N_353,N_230);
nor U406 (N_406,N_225,N_299);
or U407 (N_407,N_285,N_296);
and U408 (N_408,N_291,N_302);
and U409 (N_409,N_206,N_346);
nor U410 (N_410,N_392,N_389);
nor U411 (N_411,N_390,N_354);
or U412 (N_412,N_385,N_279);
nand U413 (N_413,N_231,N_342);
and U414 (N_414,N_309,N_314);
nand U415 (N_415,N_377,N_345);
or U416 (N_416,N_359,N_239);
and U417 (N_417,N_203,N_347);
nand U418 (N_418,N_387,N_257);
or U419 (N_419,N_240,N_262);
nand U420 (N_420,N_341,N_229);
nor U421 (N_421,N_266,N_357);
and U422 (N_422,N_290,N_307);
nand U423 (N_423,N_256,N_252);
nor U424 (N_424,N_331,N_287);
nand U425 (N_425,N_355,N_216);
nand U426 (N_426,N_275,N_368);
or U427 (N_427,N_284,N_222);
nor U428 (N_428,N_329,N_361);
nor U429 (N_429,N_282,N_319);
xnor U430 (N_430,N_265,N_327);
nand U431 (N_431,N_322,N_212);
xor U432 (N_432,N_236,N_218);
xnor U433 (N_433,N_318,N_379);
and U434 (N_434,N_317,N_298);
or U435 (N_435,N_343,N_270);
and U436 (N_436,N_253,N_395);
nand U437 (N_437,N_245,N_242);
or U438 (N_438,N_383,N_363);
and U439 (N_439,N_350,N_250);
or U440 (N_440,N_348,N_382);
nor U441 (N_441,N_247,N_202);
xor U442 (N_442,N_393,N_233);
nand U443 (N_443,N_249,N_278);
xnor U444 (N_444,N_378,N_267);
or U445 (N_445,N_221,N_365);
nor U446 (N_446,N_316,N_208);
nand U447 (N_447,N_237,N_367);
and U448 (N_448,N_351,N_224);
or U449 (N_449,N_215,N_205);
and U450 (N_450,N_333,N_332);
or U451 (N_451,N_288,N_399);
and U452 (N_452,N_328,N_235);
xnor U453 (N_453,N_300,N_293);
nor U454 (N_454,N_209,N_323);
nand U455 (N_455,N_281,N_356);
xnor U456 (N_456,N_268,N_243);
nand U457 (N_457,N_373,N_277);
xnor U458 (N_458,N_213,N_201);
nor U459 (N_459,N_364,N_254);
xnor U460 (N_460,N_394,N_386);
nor U461 (N_461,N_210,N_334);
nor U462 (N_462,N_220,N_305);
nand U463 (N_463,N_313,N_234);
xnor U464 (N_464,N_217,N_228);
nand U465 (N_465,N_274,N_369);
and U466 (N_466,N_310,N_204);
nor U467 (N_467,N_397,N_312);
and U468 (N_468,N_349,N_375);
nand U469 (N_469,N_258,N_286);
nor U470 (N_470,N_238,N_264);
xor U471 (N_471,N_396,N_295);
and U472 (N_472,N_251,N_372);
xnor U473 (N_473,N_362,N_226);
nand U474 (N_474,N_304,N_260);
xnor U475 (N_475,N_297,N_223);
xor U476 (N_476,N_371,N_219);
or U477 (N_477,N_338,N_360);
or U478 (N_478,N_330,N_292);
and U479 (N_479,N_211,N_276);
nor U480 (N_480,N_374,N_271);
and U481 (N_481,N_241,N_388);
and U482 (N_482,N_306,N_263);
nand U483 (N_483,N_320,N_261);
or U484 (N_484,N_336,N_283);
and U485 (N_485,N_337,N_358);
xor U486 (N_486,N_246,N_335);
nand U487 (N_487,N_391,N_324);
xor U488 (N_488,N_207,N_366);
nor U489 (N_489,N_248,N_294);
xnor U490 (N_490,N_315,N_200);
and U491 (N_491,N_344,N_376);
xor U492 (N_492,N_272,N_370);
and U493 (N_493,N_273,N_289);
xor U494 (N_494,N_352,N_214);
or U495 (N_495,N_380,N_326);
xor U496 (N_496,N_311,N_340);
nor U497 (N_497,N_325,N_398);
xor U498 (N_498,N_381,N_301);
nand U499 (N_499,N_244,N_269);
xnor U500 (N_500,N_345,N_216);
nand U501 (N_501,N_299,N_252);
and U502 (N_502,N_399,N_205);
xor U503 (N_503,N_317,N_258);
and U504 (N_504,N_272,N_232);
xnor U505 (N_505,N_374,N_392);
nand U506 (N_506,N_295,N_298);
nand U507 (N_507,N_265,N_354);
xnor U508 (N_508,N_274,N_287);
nor U509 (N_509,N_292,N_399);
nor U510 (N_510,N_395,N_307);
nand U511 (N_511,N_247,N_330);
and U512 (N_512,N_287,N_311);
or U513 (N_513,N_380,N_339);
nor U514 (N_514,N_301,N_309);
nand U515 (N_515,N_221,N_278);
nand U516 (N_516,N_333,N_328);
and U517 (N_517,N_319,N_216);
nand U518 (N_518,N_381,N_226);
nand U519 (N_519,N_362,N_209);
nand U520 (N_520,N_304,N_310);
nor U521 (N_521,N_242,N_212);
xnor U522 (N_522,N_223,N_279);
nor U523 (N_523,N_231,N_279);
xor U524 (N_524,N_350,N_212);
or U525 (N_525,N_279,N_245);
and U526 (N_526,N_381,N_319);
and U527 (N_527,N_248,N_262);
or U528 (N_528,N_239,N_218);
xnor U529 (N_529,N_232,N_335);
xor U530 (N_530,N_331,N_225);
and U531 (N_531,N_378,N_262);
xnor U532 (N_532,N_307,N_331);
nor U533 (N_533,N_221,N_292);
and U534 (N_534,N_291,N_398);
or U535 (N_535,N_347,N_228);
xnor U536 (N_536,N_310,N_330);
xor U537 (N_537,N_222,N_203);
xnor U538 (N_538,N_313,N_265);
nand U539 (N_539,N_351,N_269);
nor U540 (N_540,N_222,N_295);
and U541 (N_541,N_311,N_351);
and U542 (N_542,N_302,N_230);
nand U543 (N_543,N_225,N_248);
nor U544 (N_544,N_207,N_324);
and U545 (N_545,N_258,N_343);
or U546 (N_546,N_257,N_394);
nand U547 (N_547,N_207,N_241);
xor U548 (N_548,N_256,N_241);
xnor U549 (N_549,N_385,N_384);
or U550 (N_550,N_325,N_217);
nand U551 (N_551,N_294,N_374);
nand U552 (N_552,N_273,N_262);
nor U553 (N_553,N_355,N_282);
nor U554 (N_554,N_211,N_239);
or U555 (N_555,N_277,N_316);
and U556 (N_556,N_249,N_207);
xor U557 (N_557,N_271,N_357);
nand U558 (N_558,N_293,N_341);
xnor U559 (N_559,N_382,N_309);
nand U560 (N_560,N_303,N_239);
nor U561 (N_561,N_365,N_271);
nand U562 (N_562,N_321,N_373);
or U563 (N_563,N_294,N_240);
nand U564 (N_564,N_301,N_245);
or U565 (N_565,N_263,N_222);
xor U566 (N_566,N_396,N_315);
and U567 (N_567,N_235,N_204);
nor U568 (N_568,N_316,N_263);
nand U569 (N_569,N_224,N_209);
nor U570 (N_570,N_302,N_286);
and U571 (N_571,N_329,N_253);
nand U572 (N_572,N_235,N_258);
and U573 (N_573,N_249,N_280);
or U574 (N_574,N_333,N_242);
xnor U575 (N_575,N_257,N_292);
xor U576 (N_576,N_357,N_390);
nor U577 (N_577,N_225,N_339);
nor U578 (N_578,N_204,N_361);
or U579 (N_579,N_235,N_342);
nand U580 (N_580,N_267,N_337);
or U581 (N_581,N_288,N_275);
and U582 (N_582,N_315,N_341);
nand U583 (N_583,N_391,N_268);
xnor U584 (N_584,N_326,N_288);
nand U585 (N_585,N_271,N_339);
nand U586 (N_586,N_299,N_333);
nor U587 (N_587,N_262,N_395);
xor U588 (N_588,N_295,N_398);
nand U589 (N_589,N_252,N_381);
nand U590 (N_590,N_266,N_231);
xnor U591 (N_591,N_210,N_298);
or U592 (N_592,N_281,N_293);
nand U593 (N_593,N_349,N_348);
xor U594 (N_594,N_331,N_234);
or U595 (N_595,N_275,N_258);
and U596 (N_596,N_213,N_281);
nor U597 (N_597,N_302,N_379);
and U598 (N_598,N_343,N_377);
or U599 (N_599,N_341,N_340);
xor U600 (N_600,N_561,N_451);
or U601 (N_601,N_588,N_463);
and U602 (N_602,N_470,N_578);
nand U603 (N_603,N_536,N_453);
or U604 (N_604,N_527,N_583);
xor U605 (N_605,N_417,N_446);
nand U606 (N_606,N_425,N_493);
nand U607 (N_607,N_540,N_550);
nor U608 (N_608,N_564,N_500);
xor U609 (N_609,N_598,N_418);
xor U610 (N_610,N_434,N_538);
and U611 (N_611,N_520,N_459);
and U612 (N_612,N_537,N_531);
or U613 (N_613,N_497,N_482);
or U614 (N_614,N_568,N_424);
nand U615 (N_615,N_580,N_433);
nand U616 (N_616,N_579,N_414);
nand U617 (N_617,N_480,N_530);
or U618 (N_618,N_510,N_552);
or U619 (N_619,N_545,N_539);
and U620 (N_620,N_413,N_526);
or U621 (N_621,N_515,N_448);
and U622 (N_622,N_542,N_548);
xor U623 (N_623,N_554,N_491);
or U624 (N_624,N_428,N_421);
or U625 (N_625,N_533,N_507);
nand U626 (N_626,N_443,N_441);
xor U627 (N_627,N_590,N_522);
nand U628 (N_628,N_592,N_562);
or U629 (N_629,N_513,N_437);
and U630 (N_630,N_400,N_514);
nor U631 (N_631,N_436,N_573);
and U632 (N_632,N_456,N_535);
nor U633 (N_633,N_547,N_460);
and U634 (N_634,N_486,N_401);
and U635 (N_635,N_442,N_420);
or U636 (N_636,N_532,N_474);
nor U637 (N_637,N_560,N_586);
nand U638 (N_638,N_449,N_521);
nand U639 (N_639,N_557,N_431);
xor U640 (N_640,N_485,N_412);
xnor U641 (N_641,N_574,N_423);
or U642 (N_642,N_458,N_426);
nor U643 (N_643,N_517,N_498);
xnor U644 (N_644,N_454,N_439);
xnor U645 (N_645,N_508,N_455);
nor U646 (N_646,N_571,N_438);
nand U647 (N_647,N_501,N_489);
xnor U648 (N_648,N_499,N_492);
nand U649 (N_649,N_525,N_406);
xnor U650 (N_650,N_402,N_587);
xor U651 (N_651,N_502,N_558);
and U652 (N_652,N_551,N_445);
and U653 (N_653,N_567,N_468);
nor U654 (N_654,N_496,N_503);
or U655 (N_655,N_565,N_559);
nand U656 (N_656,N_519,N_511);
and U657 (N_657,N_473,N_435);
nand U658 (N_658,N_410,N_415);
and U659 (N_659,N_528,N_516);
nand U660 (N_660,N_440,N_505);
nor U661 (N_661,N_490,N_541);
and U662 (N_662,N_484,N_509);
or U663 (N_663,N_582,N_553);
nand U664 (N_664,N_405,N_512);
nor U665 (N_665,N_429,N_591);
nor U666 (N_666,N_506,N_403);
xnor U667 (N_667,N_452,N_581);
and U668 (N_668,N_476,N_596);
nor U669 (N_669,N_518,N_466);
xor U670 (N_670,N_404,N_523);
and U671 (N_671,N_467,N_427);
nor U672 (N_672,N_444,N_543);
xor U673 (N_673,N_407,N_461);
xnor U674 (N_674,N_462,N_494);
nor U675 (N_675,N_487,N_585);
and U676 (N_676,N_471,N_469);
nand U677 (N_677,N_483,N_544);
nor U678 (N_678,N_563,N_430);
and U679 (N_679,N_475,N_464);
xor U680 (N_680,N_450,N_478);
nor U681 (N_681,N_595,N_411);
and U682 (N_682,N_419,N_422);
xor U683 (N_683,N_546,N_416);
xor U684 (N_684,N_566,N_529);
nor U685 (N_685,N_488,N_593);
nand U686 (N_686,N_569,N_481);
xnor U687 (N_687,N_577,N_447);
nor U688 (N_688,N_594,N_570);
or U689 (N_689,N_576,N_556);
xnor U690 (N_690,N_584,N_599);
xor U691 (N_691,N_479,N_465);
or U692 (N_692,N_597,N_495);
or U693 (N_693,N_555,N_408);
and U694 (N_694,N_589,N_524);
xor U695 (N_695,N_534,N_409);
and U696 (N_696,N_572,N_432);
xnor U697 (N_697,N_549,N_575);
xnor U698 (N_698,N_504,N_472);
and U699 (N_699,N_457,N_477);
and U700 (N_700,N_461,N_423);
nand U701 (N_701,N_541,N_497);
or U702 (N_702,N_427,N_420);
xor U703 (N_703,N_577,N_441);
and U704 (N_704,N_529,N_563);
nor U705 (N_705,N_473,N_503);
nand U706 (N_706,N_536,N_407);
xor U707 (N_707,N_526,N_513);
xnor U708 (N_708,N_482,N_472);
and U709 (N_709,N_572,N_478);
nor U710 (N_710,N_518,N_581);
xnor U711 (N_711,N_403,N_474);
and U712 (N_712,N_586,N_585);
and U713 (N_713,N_488,N_407);
nor U714 (N_714,N_454,N_404);
nand U715 (N_715,N_513,N_510);
nand U716 (N_716,N_446,N_551);
xnor U717 (N_717,N_517,N_509);
or U718 (N_718,N_476,N_517);
and U719 (N_719,N_538,N_473);
xnor U720 (N_720,N_412,N_500);
nand U721 (N_721,N_466,N_573);
nand U722 (N_722,N_546,N_571);
nor U723 (N_723,N_556,N_541);
xor U724 (N_724,N_433,N_471);
xnor U725 (N_725,N_438,N_504);
nor U726 (N_726,N_520,N_530);
nor U727 (N_727,N_479,N_444);
and U728 (N_728,N_425,N_449);
nand U729 (N_729,N_491,N_498);
nand U730 (N_730,N_573,N_413);
nand U731 (N_731,N_527,N_531);
or U732 (N_732,N_584,N_548);
and U733 (N_733,N_537,N_477);
nor U734 (N_734,N_589,N_469);
xor U735 (N_735,N_519,N_477);
nor U736 (N_736,N_525,N_561);
xor U737 (N_737,N_523,N_584);
xor U738 (N_738,N_540,N_592);
nor U739 (N_739,N_509,N_587);
xor U740 (N_740,N_599,N_445);
nand U741 (N_741,N_440,N_483);
or U742 (N_742,N_531,N_562);
xor U743 (N_743,N_470,N_408);
and U744 (N_744,N_461,N_538);
and U745 (N_745,N_506,N_546);
nand U746 (N_746,N_592,N_426);
or U747 (N_747,N_543,N_589);
or U748 (N_748,N_524,N_485);
or U749 (N_749,N_440,N_422);
nor U750 (N_750,N_527,N_405);
nor U751 (N_751,N_575,N_495);
or U752 (N_752,N_472,N_515);
and U753 (N_753,N_586,N_420);
or U754 (N_754,N_426,N_410);
xnor U755 (N_755,N_422,N_481);
and U756 (N_756,N_554,N_438);
nand U757 (N_757,N_555,N_403);
and U758 (N_758,N_521,N_498);
xnor U759 (N_759,N_552,N_593);
nand U760 (N_760,N_577,N_599);
or U761 (N_761,N_516,N_581);
nor U762 (N_762,N_421,N_510);
nand U763 (N_763,N_488,N_554);
or U764 (N_764,N_480,N_586);
nand U765 (N_765,N_484,N_500);
nor U766 (N_766,N_542,N_496);
and U767 (N_767,N_422,N_520);
and U768 (N_768,N_462,N_491);
nand U769 (N_769,N_429,N_572);
and U770 (N_770,N_545,N_478);
xor U771 (N_771,N_582,N_528);
xor U772 (N_772,N_409,N_450);
nor U773 (N_773,N_473,N_471);
nor U774 (N_774,N_591,N_468);
or U775 (N_775,N_525,N_526);
nand U776 (N_776,N_543,N_439);
nand U777 (N_777,N_483,N_433);
or U778 (N_778,N_464,N_597);
and U779 (N_779,N_541,N_414);
or U780 (N_780,N_592,N_424);
xnor U781 (N_781,N_510,N_582);
xnor U782 (N_782,N_431,N_495);
nor U783 (N_783,N_418,N_442);
nor U784 (N_784,N_543,N_538);
nand U785 (N_785,N_449,N_480);
nor U786 (N_786,N_571,N_464);
and U787 (N_787,N_480,N_524);
and U788 (N_788,N_447,N_544);
and U789 (N_789,N_486,N_523);
xnor U790 (N_790,N_587,N_564);
nand U791 (N_791,N_578,N_459);
nand U792 (N_792,N_501,N_571);
xor U793 (N_793,N_412,N_514);
nor U794 (N_794,N_573,N_452);
nor U795 (N_795,N_585,N_516);
or U796 (N_796,N_569,N_525);
nand U797 (N_797,N_536,N_513);
or U798 (N_798,N_475,N_555);
or U799 (N_799,N_563,N_552);
or U800 (N_800,N_721,N_760);
nand U801 (N_801,N_707,N_787);
or U802 (N_802,N_746,N_713);
or U803 (N_803,N_688,N_774);
or U804 (N_804,N_708,N_745);
and U805 (N_805,N_653,N_648);
nand U806 (N_806,N_665,N_710);
xor U807 (N_807,N_635,N_777);
nand U808 (N_808,N_643,N_634);
nor U809 (N_809,N_767,N_678);
nand U810 (N_810,N_766,N_797);
and U811 (N_811,N_646,N_703);
or U812 (N_812,N_748,N_613);
nor U813 (N_813,N_671,N_786);
and U814 (N_814,N_758,N_605);
nor U815 (N_815,N_723,N_728);
nand U816 (N_816,N_675,N_655);
nor U817 (N_817,N_725,N_649);
nor U818 (N_818,N_765,N_658);
or U819 (N_819,N_689,N_631);
nor U820 (N_820,N_693,N_743);
and U821 (N_821,N_684,N_733);
nand U822 (N_822,N_661,N_638);
xnor U823 (N_823,N_657,N_781);
nand U824 (N_824,N_764,N_736);
xor U825 (N_825,N_735,N_785);
nor U826 (N_826,N_718,N_604);
nand U827 (N_827,N_667,N_670);
xnor U828 (N_828,N_647,N_633);
nand U829 (N_829,N_744,N_669);
xnor U830 (N_830,N_600,N_716);
and U831 (N_831,N_753,N_796);
and U832 (N_832,N_612,N_637);
nor U833 (N_833,N_697,N_666);
and U834 (N_834,N_754,N_630);
nor U835 (N_835,N_795,N_662);
or U836 (N_836,N_762,N_724);
or U837 (N_837,N_621,N_792);
nand U838 (N_838,N_783,N_639);
xnor U839 (N_839,N_717,N_695);
nand U840 (N_840,N_629,N_676);
xnor U841 (N_841,N_645,N_626);
or U842 (N_842,N_627,N_782);
xor U843 (N_843,N_650,N_619);
and U844 (N_844,N_642,N_757);
xor U845 (N_845,N_720,N_778);
nor U846 (N_846,N_779,N_614);
nand U847 (N_847,N_660,N_674);
or U848 (N_848,N_691,N_739);
nor U849 (N_849,N_794,N_668);
xor U850 (N_850,N_664,N_673);
nor U851 (N_851,N_776,N_722);
xor U852 (N_852,N_750,N_756);
or U853 (N_853,N_609,N_768);
xnor U854 (N_854,N_652,N_732);
and U855 (N_855,N_628,N_700);
xnor U856 (N_856,N_632,N_715);
xnor U857 (N_857,N_611,N_687);
and U858 (N_858,N_771,N_624);
or U859 (N_859,N_686,N_706);
nor U860 (N_860,N_636,N_784);
and U861 (N_861,N_663,N_726);
nand U862 (N_862,N_789,N_698);
nor U863 (N_863,N_730,N_702);
and U864 (N_864,N_615,N_699);
and U865 (N_865,N_677,N_780);
xor U866 (N_866,N_690,N_749);
nor U867 (N_867,N_682,N_618);
xor U868 (N_868,N_759,N_775);
xnor U869 (N_869,N_681,N_685);
and U870 (N_870,N_719,N_602);
nand U871 (N_871,N_773,N_731);
nand U872 (N_872,N_763,N_601);
nor U873 (N_873,N_798,N_606);
nand U874 (N_874,N_701,N_656);
and U875 (N_875,N_694,N_747);
or U876 (N_876,N_622,N_625);
or U877 (N_877,N_696,N_799);
or U878 (N_878,N_623,N_752);
nor U879 (N_879,N_729,N_737);
nand U880 (N_880,N_692,N_620);
xor U881 (N_881,N_704,N_603);
xnor U882 (N_882,N_680,N_640);
xor U883 (N_883,N_644,N_616);
or U884 (N_884,N_709,N_714);
or U885 (N_885,N_654,N_641);
and U886 (N_886,N_651,N_610);
nor U887 (N_887,N_761,N_617);
nor U888 (N_888,N_741,N_734);
nand U889 (N_889,N_751,N_742);
nor U890 (N_890,N_790,N_683);
or U891 (N_891,N_672,N_727);
and U892 (N_892,N_755,N_705);
or U893 (N_893,N_607,N_788);
or U894 (N_894,N_791,N_679);
xor U895 (N_895,N_711,N_772);
or U896 (N_896,N_659,N_793);
or U897 (N_897,N_712,N_738);
nand U898 (N_898,N_770,N_769);
nand U899 (N_899,N_740,N_608);
or U900 (N_900,N_642,N_756);
xor U901 (N_901,N_615,N_726);
nand U902 (N_902,N_720,N_791);
nand U903 (N_903,N_668,N_648);
xor U904 (N_904,N_744,N_617);
xnor U905 (N_905,N_705,N_796);
or U906 (N_906,N_706,N_711);
nor U907 (N_907,N_794,N_647);
nand U908 (N_908,N_701,N_721);
or U909 (N_909,N_785,N_645);
or U910 (N_910,N_642,N_703);
nand U911 (N_911,N_635,N_747);
nor U912 (N_912,N_740,N_683);
nor U913 (N_913,N_611,N_681);
xor U914 (N_914,N_704,N_623);
xnor U915 (N_915,N_723,N_617);
nor U916 (N_916,N_619,N_793);
or U917 (N_917,N_622,N_652);
nor U918 (N_918,N_645,N_784);
nand U919 (N_919,N_647,N_780);
nand U920 (N_920,N_608,N_741);
nor U921 (N_921,N_758,N_723);
or U922 (N_922,N_697,N_649);
nor U923 (N_923,N_695,N_739);
nand U924 (N_924,N_647,N_782);
xnor U925 (N_925,N_705,N_611);
or U926 (N_926,N_783,N_660);
or U927 (N_927,N_723,N_648);
nand U928 (N_928,N_652,N_734);
nor U929 (N_929,N_735,N_644);
and U930 (N_930,N_741,N_748);
or U931 (N_931,N_628,N_726);
nand U932 (N_932,N_655,N_649);
and U933 (N_933,N_763,N_728);
and U934 (N_934,N_608,N_633);
xnor U935 (N_935,N_677,N_720);
or U936 (N_936,N_646,N_765);
or U937 (N_937,N_651,N_775);
nor U938 (N_938,N_662,N_723);
xnor U939 (N_939,N_631,N_668);
xnor U940 (N_940,N_759,N_735);
or U941 (N_941,N_710,N_739);
and U942 (N_942,N_795,N_606);
and U943 (N_943,N_743,N_762);
nand U944 (N_944,N_684,N_703);
nor U945 (N_945,N_793,N_658);
or U946 (N_946,N_751,N_776);
nor U947 (N_947,N_762,N_623);
or U948 (N_948,N_747,N_706);
nand U949 (N_949,N_670,N_638);
xor U950 (N_950,N_637,N_672);
nor U951 (N_951,N_702,N_671);
and U952 (N_952,N_684,N_736);
nand U953 (N_953,N_617,N_604);
and U954 (N_954,N_650,N_699);
nand U955 (N_955,N_643,N_752);
xnor U956 (N_956,N_615,N_697);
nand U957 (N_957,N_749,N_694);
and U958 (N_958,N_645,N_755);
and U959 (N_959,N_769,N_632);
or U960 (N_960,N_661,N_632);
nand U961 (N_961,N_677,N_688);
nand U962 (N_962,N_656,N_616);
nand U963 (N_963,N_733,N_683);
nand U964 (N_964,N_795,N_639);
or U965 (N_965,N_762,N_778);
or U966 (N_966,N_728,N_652);
nand U967 (N_967,N_756,N_738);
nor U968 (N_968,N_698,N_685);
or U969 (N_969,N_604,N_751);
nand U970 (N_970,N_643,N_798);
and U971 (N_971,N_732,N_786);
nor U972 (N_972,N_622,N_769);
nand U973 (N_973,N_607,N_702);
and U974 (N_974,N_742,N_668);
xor U975 (N_975,N_772,N_652);
and U976 (N_976,N_738,N_628);
nor U977 (N_977,N_797,N_779);
xnor U978 (N_978,N_643,N_677);
nand U979 (N_979,N_641,N_728);
nand U980 (N_980,N_731,N_681);
xor U981 (N_981,N_741,N_721);
and U982 (N_982,N_737,N_799);
xor U983 (N_983,N_623,N_650);
and U984 (N_984,N_611,N_762);
nor U985 (N_985,N_628,N_604);
and U986 (N_986,N_618,N_748);
and U987 (N_987,N_707,N_612);
or U988 (N_988,N_768,N_724);
nand U989 (N_989,N_792,N_667);
xor U990 (N_990,N_601,N_643);
nor U991 (N_991,N_655,N_710);
nand U992 (N_992,N_781,N_642);
and U993 (N_993,N_763,N_600);
nor U994 (N_994,N_776,N_744);
nor U995 (N_995,N_785,N_657);
or U996 (N_996,N_627,N_640);
nand U997 (N_997,N_603,N_785);
xor U998 (N_998,N_638,N_630);
or U999 (N_999,N_776,N_657);
xnor U1000 (N_1000,N_830,N_956);
xnor U1001 (N_1001,N_825,N_966);
and U1002 (N_1002,N_884,N_813);
nor U1003 (N_1003,N_987,N_991);
nand U1004 (N_1004,N_858,N_839);
and U1005 (N_1005,N_871,N_897);
nand U1006 (N_1006,N_856,N_806);
nand U1007 (N_1007,N_873,N_885);
or U1008 (N_1008,N_931,N_978);
nand U1009 (N_1009,N_879,N_900);
nor U1010 (N_1010,N_828,N_805);
xnor U1011 (N_1011,N_802,N_822);
and U1012 (N_1012,N_855,N_886);
nor U1013 (N_1013,N_851,N_928);
nor U1014 (N_1014,N_870,N_914);
and U1015 (N_1015,N_869,N_906);
nand U1016 (N_1016,N_949,N_860);
or U1017 (N_1017,N_846,N_843);
nand U1018 (N_1018,N_877,N_980);
and U1019 (N_1019,N_927,N_974);
xor U1020 (N_1020,N_863,N_904);
and U1021 (N_1021,N_852,N_959);
and U1022 (N_1022,N_896,N_887);
and U1023 (N_1023,N_936,N_926);
xor U1024 (N_1024,N_821,N_849);
nor U1025 (N_1025,N_901,N_819);
xor U1026 (N_1026,N_973,N_976);
xnor U1027 (N_1027,N_890,N_984);
nand U1028 (N_1028,N_985,N_874);
nor U1029 (N_1029,N_932,N_841);
and U1030 (N_1030,N_803,N_918);
nor U1031 (N_1031,N_883,N_840);
nand U1032 (N_1032,N_996,N_923);
nand U1033 (N_1033,N_809,N_969);
or U1034 (N_1034,N_810,N_958);
and U1035 (N_1035,N_834,N_895);
nand U1036 (N_1036,N_977,N_971);
nor U1037 (N_1037,N_820,N_917);
xnor U1038 (N_1038,N_951,N_903);
xnor U1039 (N_1039,N_935,N_850);
or U1040 (N_1040,N_800,N_939);
nor U1041 (N_1041,N_947,N_981);
or U1042 (N_1042,N_934,N_905);
and U1043 (N_1043,N_911,N_964);
and U1044 (N_1044,N_866,N_993);
or U1045 (N_1045,N_963,N_992);
nor U1046 (N_1046,N_893,N_845);
nor U1047 (N_1047,N_990,N_831);
or U1048 (N_1048,N_999,N_954);
xor U1049 (N_1049,N_952,N_994);
or U1050 (N_1050,N_943,N_930);
or U1051 (N_1051,N_922,N_837);
or U1052 (N_1052,N_909,N_946);
nand U1053 (N_1053,N_962,N_907);
xnor U1054 (N_1054,N_836,N_889);
nand U1055 (N_1055,N_875,N_986);
nand U1056 (N_1056,N_913,N_832);
and U1057 (N_1057,N_848,N_835);
nand U1058 (N_1058,N_925,N_957);
nor U1059 (N_1059,N_853,N_876);
xnor U1060 (N_1060,N_908,N_972);
or U1061 (N_1061,N_814,N_892);
nand U1062 (N_1062,N_961,N_812);
nor U1063 (N_1063,N_859,N_968);
and U1064 (N_1064,N_867,N_944);
and U1065 (N_1065,N_967,N_882);
nor U1066 (N_1066,N_941,N_899);
nand U1067 (N_1067,N_833,N_920);
nand U1068 (N_1068,N_854,N_940);
xnor U1069 (N_1069,N_945,N_912);
nor U1070 (N_1070,N_868,N_937);
nand U1071 (N_1071,N_861,N_801);
nor U1072 (N_1072,N_815,N_933);
or U1073 (N_1073,N_826,N_811);
and U1074 (N_1074,N_983,N_818);
nand U1075 (N_1075,N_942,N_919);
nand U1076 (N_1076,N_910,N_998);
nand U1077 (N_1077,N_948,N_921);
or U1078 (N_1078,N_847,N_929);
and U1079 (N_1079,N_807,N_898);
nand U1080 (N_1080,N_808,N_857);
nor U1081 (N_1081,N_995,N_878);
and U1082 (N_1082,N_988,N_997);
or U1083 (N_1083,N_838,N_953);
nand U1084 (N_1084,N_891,N_872);
nand U1085 (N_1085,N_989,N_827);
nor U1086 (N_1086,N_965,N_975);
and U1087 (N_1087,N_864,N_955);
xor U1088 (N_1088,N_842,N_982);
xnor U1089 (N_1089,N_824,N_881);
and U1090 (N_1090,N_829,N_816);
and U1091 (N_1091,N_924,N_970);
or U1092 (N_1092,N_938,N_979);
nor U1093 (N_1093,N_804,N_894);
nand U1094 (N_1094,N_865,N_915);
nor U1095 (N_1095,N_902,N_950);
and U1096 (N_1096,N_880,N_844);
and U1097 (N_1097,N_817,N_823);
nor U1098 (N_1098,N_960,N_888);
nor U1099 (N_1099,N_862,N_916);
nor U1100 (N_1100,N_958,N_887);
xor U1101 (N_1101,N_880,N_887);
xor U1102 (N_1102,N_821,N_990);
nand U1103 (N_1103,N_898,N_995);
xnor U1104 (N_1104,N_907,N_809);
xor U1105 (N_1105,N_909,N_862);
and U1106 (N_1106,N_942,N_811);
xor U1107 (N_1107,N_964,N_849);
and U1108 (N_1108,N_830,N_837);
or U1109 (N_1109,N_809,N_961);
xnor U1110 (N_1110,N_953,N_945);
nor U1111 (N_1111,N_831,N_978);
and U1112 (N_1112,N_828,N_839);
or U1113 (N_1113,N_865,N_892);
nand U1114 (N_1114,N_921,N_900);
and U1115 (N_1115,N_865,N_914);
xnor U1116 (N_1116,N_815,N_943);
or U1117 (N_1117,N_863,N_948);
nor U1118 (N_1118,N_841,N_915);
and U1119 (N_1119,N_810,N_812);
nor U1120 (N_1120,N_847,N_898);
and U1121 (N_1121,N_959,N_819);
xnor U1122 (N_1122,N_894,N_913);
nand U1123 (N_1123,N_934,N_838);
nor U1124 (N_1124,N_940,N_805);
xnor U1125 (N_1125,N_830,N_881);
and U1126 (N_1126,N_885,N_971);
or U1127 (N_1127,N_973,N_925);
nor U1128 (N_1128,N_914,N_907);
or U1129 (N_1129,N_919,N_816);
xor U1130 (N_1130,N_928,N_992);
xor U1131 (N_1131,N_982,N_914);
or U1132 (N_1132,N_832,N_897);
and U1133 (N_1133,N_848,N_823);
nand U1134 (N_1134,N_982,N_981);
xor U1135 (N_1135,N_811,N_916);
nand U1136 (N_1136,N_955,N_943);
and U1137 (N_1137,N_809,N_885);
and U1138 (N_1138,N_848,N_961);
or U1139 (N_1139,N_906,N_850);
and U1140 (N_1140,N_873,N_942);
and U1141 (N_1141,N_966,N_862);
nor U1142 (N_1142,N_832,N_802);
nand U1143 (N_1143,N_855,N_826);
xor U1144 (N_1144,N_967,N_803);
and U1145 (N_1145,N_945,N_989);
nand U1146 (N_1146,N_824,N_982);
nand U1147 (N_1147,N_923,N_924);
nand U1148 (N_1148,N_964,N_821);
nand U1149 (N_1149,N_945,N_902);
and U1150 (N_1150,N_850,N_858);
nand U1151 (N_1151,N_900,N_897);
nor U1152 (N_1152,N_993,N_911);
and U1153 (N_1153,N_989,N_902);
and U1154 (N_1154,N_978,N_820);
nand U1155 (N_1155,N_897,N_966);
and U1156 (N_1156,N_855,N_843);
and U1157 (N_1157,N_956,N_951);
nand U1158 (N_1158,N_947,N_902);
and U1159 (N_1159,N_843,N_907);
xnor U1160 (N_1160,N_804,N_835);
xnor U1161 (N_1161,N_842,N_892);
or U1162 (N_1162,N_839,N_900);
nor U1163 (N_1163,N_975,N_933);
nor U1164 (N_1164,N_888,N_917);
nor U1165 (N_1165,N_934,N_809);
nand U1166 (N_1166,N_953,N_927);
xor U1167 (N_1167,N_995,N_858);
nand U1168 (N_1168,N_910,N_876);
and U1169 (N_1169,N_941,N_975);
or U1170 (N_1170,N_922,N_968);
nand U1171 (N_1171,N_925,N_944);
nor U1172 (N_1172,N_963,N_922);
and U1173 (N_1173,N_920,N_882);
or U1174 (N_1174,N_889,N_891);
and U1175 (N_1175,N_906,N_926);
and U1176 (N_1176,N_971,N_820);
xnor U1177 (N_1177,N_830,N_918);
nand U1178 (N_1178,N_960,N_840);
and U1179 (N_1179,N_965,N_820);
nor U1180 (N_1180,N_941,N_897);
nand U1181 (N_1181,N_926,N_887);
and U1182 (N_1182,N_939,N_935);
or U1183 (N_1183,N_802,N_856);
and U1184 (N_1184,N_928,N_852);
xnor U1185 (N_1185,N_979,N_885);
nand U1186 (N_1186,N_921,N_994);
nor U1187 (N_1187,N_991,N_976);
nand U1188 (N_1188,N_876,N_880);
or U1189 (N_1189,N_993,N_968);
xor U1190 (N_1190,N_935,N_861);
nand U1191 (N_1191,N_839,N_948);
and U1192 (N_1192,N_851,N_925);
xnor U1193 (N_1193,N_879,N_895);
and U1194 (N_1194,N_998,N_832);
nor U1195 (N_1195,N_965,N_913);
and U1196 (N_1196,N_830,N_936);
and U1197 (N_1197,N_807,N_835);
and U1198 (N_1198,N_871,N_920);
or U1199 (N_1199,N_953,N_937);
and U1200 (N_1200,N_1164,N_1079);
or U1201 (N_1201,N_1145,N_1125);
xor U1202 (N_1202,N_1007,N_1151);
and U1203 (N_1203,N_1045,N_1120);
nand U1204 (N_1204,N_1016,N_1115);
xor U1205 (N_1205,N_1185,N_1152);
xor U1206 (N_1206,N_1069,N_1082);
nor U1207 (N_1207,N_1121,N_1157);
nor U1208 (N_1208,N_1170,N_1075);
xnor U1209 (N_1209,N_1021,N_1139);
nand U1210 (N_1210,N_1133,N_1107);
and U1211 (N_1211,N_1055,N_1108);
nand U1212 (N_1212,N_1083,N_1197);
or U1213 (N_1213,N_1070,N_1117);
or U1214 (N_1214,N_1192,N_1030);
nand U1215 (N_1215,N_1028,N_1052);
xor U1216 (N_1216,N_1057,N_1112);
xnor U1217 (N_1217,N_1074,N_1081);
and U1218 (N_1218,N_1095,N_1088);
xnor U1219 (N_1219,N_1061,N_1011);
and U1220 (N_1220,N_1163,N_1009);
xnor U1221 (N_1221,N_1129,N_1029);
nor U1222 (N_1222,N_1172,N_1130);
or U1223 (N_1223,N_1171,N_1160);
and U1224 (N_1224,N_1198,N_1041);
nor U1225 (N_1225,N_1022,N_1187);
nor U1226 (N_1226,N_1182,N_1199);
xor U1227 (N_1227,N_1018,N_1102);
nand U1228 (N_1228,N_1039,N_1140);
nor U1229 (N_1229,N_1058,N_1142);
nor U1230 (N_1230,N_1191,N_1038);
or U1231 (N_1231,N_1091,N_1031);
and U1232 (N_1232,N_1099,N_1060);
xnor U1233 (N_1233,N_1092,N_1054);
and U1234 (N_1234,N_1138,N_1094);
nand U1235 (N_1235,N_1023,N_1050);
nand U1236 (N_1236,N_1017,N_1013);
nand U1237 (N_1237,N_1098,N_1113);
nand U1238 (N_1238,N_1114,N_1096);
and U1239 (N_1239,N_1166,N_1175);
nor U1240 (N_1240,N_1062,N_1150);
nor U1241 (N_1241,N_1004,N_1179);
nor U1242 (N_1242,N_1123,N_1049);
and U1243 (N_1243,N_1040,N_1046);
or U1244 (N_1244,N_1027,N_1181);
xor U1245 (N_1245,N_1002,N_1100);
nor U1246 (N_1246,N_1131,N_1110);
and U1247 (N_1247,N_1090,N_1137);
xor U1248 (N_1248,N_1183,N_1064);
or U1249 (N_1249,N_1159,N_1173);
and U1250 (N_1250,N_1124,N_1006);
nand U1251 (N_1251,N_1126,N_1026);
and U1252 (N_1252,N_1118,N_1167);
nor U1253 (N_1253,N_1056,N_1005);
nand U1254 (N_1254,N_1155,N_1086);
xor U1255 (N_1255,N_1067,N_1084);
and U1256 (N_1256,N_1174,N_1019);
xnor U1257 (N_1257,N_1127,N_1048);
or U1258 (N_1258,N_1196,N_1116);
or U1259 (N_1259,N_1063,N_1105);
or U1260 (N_1260,N_1189,N_1085);
xnor U1261 (N_1261,N_1154,N_1162);
and U1262 (N_1262,N_1015,N_1003);
nor U1263 (N_1263,N_1008,N_1068);
xor U1264 (N_1264,N_1122,N_1193);
nor U1265 (N_1265,N_1106,N_1188);
or U1266 (N_1266,N_1143,N_1073);
nand U1267 (N_1267,N_1077,N_1053);
and U1268 (N_1268,N_1025,N_1044);
nand U1269 (N_1269,N_1000,N_1109);
nand U1270 (N_1270,N_1153,N_1037);
and U1271 (N_1271,N_1161,N_1184);
xor U1272 (N_1272,N_1178,N_1186);
nand U1273 (N_1273,N_1020,N_1156);
and U1274 (N_1274,N_1168,N_1180);
xnor U1275 (N_1275,N_1149,N_1103);
xnor U1276 (N_1276,N_1080,N_1101);
nor U1277 (N_1277,N_1042,N_1071);
nor U1278 (N_1278,N_1035,N_1001);
and U1279 (N_1279,N_1043,N_1034);
nor U1280 (N_1280,N_1104,N_1165);
and U1281 (N_1281,N_1134,N_1047);
or U1282 (N_1282,N_1146,N_1128);
nor U1283 (N_1283,N_1195,N_1097);
nor U1284 (N_1284,N_1014,N_1036);
and U1285 (N_1285,N_1089,N_1141);
and U1286 (N_1286,N_1065,N_1147);
nor U1287 (N_1287,N_1119,N_1093);
and U1288 (N_1288,N_1144,N_1059);
xor U1289 (N_1289,N_1066,N_1072);
or U1290 (N_1290,N_1169,N_1158);
and U1291 (N_1291,N_1136,N_1024);
nor U1292 (N_1292,N_1194,N_1176);
nand U1293 (N_1293,N_1177,N_1190);
nand U1294 (N_1294,N_1051,N_1033);
xor U1295 (N_1295,N_1135,N_1076);
or U1296 (N_1296,N_1087,N_1078);
nor U1297 (N_1297,N_1012,N_1111);
or U1298 (N_1298,N_1032,N_1010);
xor U1299 (N_1299,N_1132,N_1148);
nand U1300 (N_1300,N_1095,N_1086);
or U1301 (N_1301,N_1098,N_1011);
or U1302 (N_1302,N_1164,N_1073);
xnor U1303 (N_1303,N_1027,N_1020);
nor U1304 (N_1304,N_1139,N_1011);
nor U1305 (N_1305,N_1013,N_1029);
nor U1306 (N_1306,N_1025,N_1150);
and U1307 (N_1307,N_1091,N_1032);
nand U1308 (N_1308,N_1043,N_1131);
and U1309 (N_1309,N_1029,N_1028);
and U1310 (N_1310,N_1039,N_1067);
nor U1311 (N_1311,N_1072,N_1075);
or U1312 (N_1312,N_1046,N_1169);
nor U1313 (N_1313,N_1145,N_1191);
nor U1314 (N_1314,N_1110,N_1008);
or U1315 (N_1315,N_1163,N_1008);
nor U1316 (N_1316,N_1050,N_1027);
nand U1317 (N_1317,N_1117,N_1094);
nand U1318 (N_1318,N_1088,N_1163);
and U1319 (N_1319,N_1117,N_1069);
xor U1320 (N_1320,N_1167,N_1100);
or U1321 (N_1321,N_1062,N_1197);
or U1322 (N_1322,N_1091,N_1001);
nand U1323 (N_1323,N_1118,N_1121);
nor U1324 (N_1324,N_1075,N_1177);
nor U1325 (N_1325,N_1039,N_1054);
nor U1326 (N_1326,N_1023,N_1121);
nand U1327 (N_1327,N_1010,N_1151);
xor U1328 (N_1328,N_1058,N_1123);
nor U1329 (N_1329,N_1043,N_1141);
nand U1330 (N_1330,N_1060,N_1165);
or U1331 (N_1331,N_1077,N_1082);
and U1332 (N_1332,N_1114,N_1045);
nor U1333 (N_1333,N_1166,N_1116);
nor U1334 (N_1334,N_1131,N_1096);
and U1335 (N_1335,N_1141,N_1169);
xor U1336 (N_1336,N_1073,N_1027);
and U1337 (N_1337,N_1088,N_1043);
nand U1338 (N_1338,N_1017,N_1185);
nand U1339 (N_1339,N_1030,N_1128);
and U1340 (N_1340,N_1120,N_1000);
or U1341 (N_1341,N_1124,N_1062);
xnor U1342 (N_1342,N_1012,N_1072);
xor U1343 (N_1343,N_1119,N_1050);
nor U1344 (N_1344,N_1039,N_1197);
xnor U1345 (N_1345,N_1151,N_1101);
and U1346 (N_1346,N_1108,N_1092);
nand U1347 (N_1347,N_1050,N_1101);
xnor U1348 (N_1348,N_1173,N_1042);
or U1349 (N_1349,N_1015,N_1030);
or U1350 (N_1350,N_1110,N_1039);
nand U1351 (N_1351,N_1069,N_1109);
nor U1352 (N_1352,N_1022,N_1097);
nand U1353 (N_1353,N_1158,N_1185);
or U1354 (N_1354,N_1138,N_1124);
and U1355 (N_1355,N_1085,N_1067);
xnor U1356 (N_1356,N_1163,N_1143);
nand U1357 (N_1357,N_1148,N_1084);
xor U1358 (N_1358,N_1192,N_1165);
nand U1359 (N_1359,N_1114,N_1079);
and U1360 (N_1360,N_1065,N_1027);
nand U1361 (N_1361,N_1065,N_1018);
or U1362 (N_1362,N_1019,N_1155);
xor U1363 (N_1363,N_1175,N_1102);
xor U1364 (N_1364,N_1153,N_1015);
nand U1365 (N_1365,N_1187,N_1096);
nand U1366 (N_1366,N_1149,N_1014);
xnor U1367 (N_1367,N_1133,N_1007);
xnor U1368 (N_1368,N_1132,N_1164);
and U1369 (N_1369,N_1185,N_1165);
xnor U1370 (N_1370,N_1114,N_1033);
and U1371 (N_1371,N_1171,N_1120);
and U1372 (N_1372,N_1016,N_1052);
nor U1373 (N_1373,N_1121,N_1146);
xnor U1374 (N_1374,N_1109,N_1065);
nand U1375 (N_1375,N_1108,N_1182);
nor U1376 (N_1376,N_1091,N_1123);
and U1377 (N_1377,N_1101,N_1113);
nand U1378 (N_1378,N_1070,N_1198);
and U1379 (N_1379,N_1176,N_1153);
nor U1380 (N_1380,N_1199,N_1093);
and U1381 (N_1381,N_1018,N_1076);
xor U1382 (N_1382,N_1164,N_1161);
xnor U1383 (N_1383,N_1031,N_1056);
xnor U1384 (N_1384,N_1026,N_1003);
xor U1385 (N_1385,N_1143,N_1195);
xnor U1386 (N_1386,N_1156,N_1009);
xor U1387 (N_1387,N_1107,N_1199);
or U1388 (N_1388,N_1051,N_1059);
and U1389 (N_1389,N_1079,N_1166);
or U1390 (N_1390,N_1005,N_1023);
nand U1391 (N_1391,N_1166,N_1170);
or U1392 (N_1392,N_1180,N_1147);
and U1393 (N_1393,N_1175,N_1055);
nand U1394 (N_1394,N_1133,N_1122);
nor U1395 (N_1395,N_1026,N_1143);
and U1396 (N_1396,N_1049,N_1090);
nand U1397 (N_1397,N_1039,N_1123);
nand U1398 (N_1398,N_1044,N_1132);
and U1399 (N_1399,N_1048,N_1059);
and U1400 (N_1400,N_1348,N_1227);
xor U1401 (N_1401,N_1321,N_1328);
or U1402 (N_1402,N_1354,N_1327);
or U1403 (N_1403,N_1363,N_1260);
nor U1404 (N_1404,N_1343,N_1345);
xor U1405 (N_1405,N_1295,N_1281);
nand U1406 (N_1406,N_1293,N_1394);
or U1407 (N_1407,N_1228,N_1296);
and U1408 (N_1408,N_1310,N_1330);
or U1409 (N_1409,N_1332,N_1358);
nor U1410 (N_1410,N_1356,N_1306);
nor U1411 (N_1411,N_1230,N_1371);
or U1412 (N_1412,N_1304,N_1208);
nand U1413 (N_1413,N_1273,N_1253);
nor U1414 (N_1414,N_1312,N_1256);
nand U1415 (N_1415,N_1396,N_1251);
xor U1416 (N_1416,N_1301,N_1391);
xor U1417 (N_1417,N_1382,N_1229);
nand U1418 (N_1418,N_1282,N_1344);
or U1419 (N_1419,N_1302,N_1237);
nand U1420 (N_1420,N_1242,N_1376);
nor U1421 (N_1421,N_1368,N_1323);
xnor U1422 (N_1422,N_1265,N_1210);
nand U1423 (N_1423,N_1387,N_1316);
xor U1424 (N_1424,N_1221,N_1381);
and U1425 (N_1425,N_1209,N_1378);
nor U1426 (N_1426,N_1393,N_1283);
nor U1427 (N_1427,N_1319,N_1211);
xnor U1428 (N_1428,N_1215,N_1335);
nand U1429 (N_1429,N_1369,N_1284);
and U1430 (N_1430,N_1325,N_1231);
nand U1431 (N_1431,N_1373,N_1259);
xor U1432 (N_1432,N_1290,N_1285);
nand U1433 (N_1433,N_1223,N_1362);
nand U1434 (N_1434,N_1297,N_1355);
xnor U1435 (N_1435,N_1204,N_1232);
xor U1436 (N_1436,N_1266,N_1206);
and U1437 (N_1437,N_1276,N_1274);
nor U1438 (N_1438,N_1240,N_1261);
xor U1439 (N_1439,N_1292,N_1257);
or U1440 (N_1440,N_1350,N_1203);
nor U1441 (N_1441,N_1289,N_1226);
nor U1442 (N_1442,N_1225,N_1339);
or U1443 (N_1443,N_1252,N_1275);
nor U1444 (N_1444,N_1380,N_1336);
and U1445 (N_1445,N_1269,N_1311);
xor U1446 (N_1446,N_1217,N_1219);
and U1447 (N_1447,N_1399,N_1234);
nand U1448 (N_1448,N_1334,N_1291);
nand U1449 (N_1449,N_1397,N_1294);
nor U1450 (N_1450,N_1377,N_1201);
xor U1451 (N_1451,N_1392,N_1305);
and U1452 (N_1452,N_1383,N_1338);
or U1453 (N_1453,N_1249,N_1268);
or U1454 (N_1454,N_1353,N_1360);
nor U1455 (N_1455,N_1303,N_1395);
nand U1456 (N_1456,N_1247,N_1386);
nand U1457 (N_1457,N_1244,N_1340);
or U1458 (N_1458,N_1236,N_1320);
xor U1459 (N_1459,N_1389,N_1374);
xnor U1460 (N_1460,N_1213,N_1326);
and U1461 (N_1461,N_1263,N_1390);
nor U1462 (N_1462,N_1309,N_1352);
or U1463 (N_1463,N_1337,N_1216);
or U1464 (N_1464,N_1347,N_1238);
nor U1465 (N_1465,N_1298,N_1388);
nand U1466 (N_1466,N_1280,N_1235);
and U1467 (N_1467,N_1364,N_1342);
xnor U1468 (N_1468,N_1333,N_1384);
xor U1469 (N_1469,N_1288,N_1264);
xor U1470 (N_1470,N_1375,N_1218);
nand U1471 (N_1471,N_1365,N_1341);
and U1472 (N_1472,N_1271,N_1258);
xnor U1473 (N_1473,N_1361,N_1212);
nor U1474 (N_1474,N_1398,N_1262);
xnor U1475 (N_1475,N_1299,N_1254);
nand U1476 (N_1476,N_1222,N_1385);
and U1477 (N_1477,N_1346,N_1308);
and U1478 (N_1478,N_1313,N_1277);
nor U1479 (N_1479,N_1214,N_1307);
or U1480 (N_1480,N_1359,N_1255);
or U1481 (N_1481,N_1287,N_1220);
nor U1482 (N_1482,N_1246,N_1317);
and U1483 (N_1483,N_1366,N_1207);
nand U1484 (N_1484,N_1270,N_1318);
and U1485 (N_1485,N_1286,N_1202);
xor U1486 (N_1486,N_1351,N_1243);
xor U1487 (N_1487,N_1370,N_1279);
nand U1488 (N_1488,N_1372,N_1300);
or U1489 (N_1489,N_1205,N_1329);
or U1490 (N_1490,N_1349,N_1357);
or U1491 (N_1491,N_1267,N_1322);
nor U1492 (N_1492,N_1367,N_1379);
nand U1493 (N_1493,N_1331,N_1314);
nand U1494 (N_1494,N_1200,N_1224);
nand U1495 (N_1495,N_1315,N_1241);
or U1496 (N_1496,N_1239,N_1245);
or U1497 (N_1497,N_1248,N_1272);
xor U1498 (N_1498,N_1324,N_1250);
or U1499 (N_1499,N_1278,N_1233);
or U1500 (N_1500,N_1339,N_1393);
or U1501 (N_1501,N_1370,N_1323);
xor U1502 (N_1502,N_1274,N_1290);
xnor U1503 (N_1503,N_1375,N_1240);
nand U1504 (N_1504,N_1337,N_1206);
or U1505 (N_1505,N_1318,N_1298);
xnor U1506 (N_1506,N_1282,N_1245);
and U1507 (N_1507,N_1376,N_1294);
and U1508 (N_1508,N_1290,N_1252);
or U1509 (N_1509,N_1337,N_1316);
and U1510 (N_1510,N_1381,N_1276);
nor U1511 (N_1511,N_1315,N_1301);
xnor U1512 (N_1512,N_1329,N_1369);
nand U1513 (N_1513,N_1295,N_1270);
and U1514 (N_1514,N_1295,N_1313);
xor U1515 (N_1515,N_1253,N_1321);
nor U1516 (N_1516,N_1384,N_1274);
nor U1517 (N_1517,N_1365,N_1219);
or U1518 (N_1518,N_1334,N_1243);
nor U1519 (N_1519,N_1334,N_1320);
nand U1520 (N_1520,N_1350,N_1337);
nor U1521 (N_1521,N_1387,N_1294);
nand U1522 (N_1522,N_1249,N_1257);
and U1523 (N_1523,N_1395,N_1238);
nor U1524 (N_1524,N_1287,N_1343);
or U1525 (N_1525,N_1354,N_1305);
and U1526 (N_1526,N_1372,N_1329);
and U1527 (N_1527,N_1398,N_1248);
nor U1528 (N_1528,N_1233,N_1323);
and U1529 (N_1529,N_1337,N_1254);
or U1530 (N_1530,N_1200,N_1219);
or U1531 (N_1531,N_1230,N_1213);
nand U1532 (N_1532,N_1322,N_1287);
xnor U1533 (N_1533,N_1218,N_1265);
and U1534 (N_1534,N_1220,N_1369);
nand U1535 (N_1535,N_1287,N_1327);
and U1536 (N_1536,N_1209,N_1327);
nor U1537 (N_1537,N_1296,N_1255);
nor U1538 (N_1538,N_1379,N_1273);
xnor U1539 (N_1539,N_1306,N_1381);
nor U1540 (N_1540,N_1382,N_1220);
nor U1541 (N_1541,N_1385,N_1352);
and U1542 (N_1542,N_1389,N_1324);
nor U1543 (N_1543,N_1370,N_1392);
nand U1544 (N_1544,N_1246,N_1235);
nand U1545 (N_1545,N_1264,N_1388);
nor U1546 (N_1546,N_1235,N_1232);
xor U1547 (N_1547,N_1395,N_1388);
or U1548 (N_1548,N_1388,N_1321);
and U1549 (N_1549,N_1323,N_1263);
and U1550 (N_1550,N_1377,N_1365);
nand U1551 (N_1551,N_1341,N_1285);
or U1552 (N_1552,N_1366,N_1343);
nand U1553 (N_1553,N_1392,N_1302);
nor U1554 (N_1554,N_1373,N_1276);
nor U1555 (N_1555,N_1240,N_1244);
or U1556 (N_1556,N_1322,N_1317);
and U1557 (N_1557,N_1345,N_1246);
nand U1558 (N_1558,N_1387,N_1239);
or U1559 (N_1559,N_1365,N_1396);
nor U1560 (N_1560,N_1253,N_1294);
or U1561 (N_1561,N_1354,N_1377);
xnor U1562 (N_1562,N_1214,N_1266);
nor U1563 (N_1563,N_1394,N_1222);
nor U1564 (N_1564,N_1308,N_1393);
or U1565 (N_1565,N_1241,N_1335);
nand U1566 (N_1566,N_1346,N_1322);
nor U1567 (N_1567,N_1296,N_1322);
nor U1568 (N_1568,N_1315,N_1209);
xor U1569 (N_1569,N_1223,N_1268);
nor U1570 (N_1570,N_1295,N_1310);
or U1571 (N_1571,N_1367,N_1352);
or U1572 (N_1572,N_1294,N_1298);
xnor U1573 (N_1573,N_1205,N_1399);
nand U1574 (N_1574,N_1343,N_1214);
or U1575 (N_1575,N_1351,N_1213);
and U1576 (N_1576,N_1377,N_1266);
xor U1577 (N_1577,N_1372,N_1204);
nor U1578 (N_1578,N_1379,N_1233);
xnor U1579 (N_1579,N_1266,N_1289);
nand U1580 (N_1580,N_1274,N_1263);
or U1581 (N_1581,N_1259,N_1200);
nor U1582 (N_1582,N_1398,N_1329);
and U1583 (N_1583,N_1208,N_1295);
and U1584 (N_1584,N_1255,N_1384);
nand U1585 (N_1585,N_1253,N_1218);
and U1586 (N_1586,N_1395,N_1300);
xor U1587 (N_1587,N_1281,N_1359);
and U1588 (N_1588,N_1268,N_1305);
nand U1589 (N_1589,N_1255,N_1336);
and U1590 (N_1590,N_1353,N_1219);
or U1591 (N_1591,N_1236,N_1394);
or U1592 (N_1592,N_1287,N_1318);
nor U1593 (N_1593,N_1352,N_1259);
xnor U1594 (N_1594,N_1206,N_1317);
xor U1595 (N_1595,N_1299,N_1355);
or U1596 (N_1596,N_1222,N_1305);
and U1597 (N_1597,N_1205,N_1279);
and U1598 (N_1598,N_1275,N_1335);
and U1599 (N_1599,N_1334,N_1322);
or U1600 (N_1600,N_1577,N_1501);
nand U1601 (N_1601,N_1531,N_1520);
or U1602 (N_1602,N_1572,N_1453);
and U1603 (N_1603,N_1443,N_1529);
nor U1604 (N_1604,N_1588,N_1444);
and U1605 (N_1605,N_1543,N_1484);
nor U1606 (N_1606,N_1506,N_1562);
or U1607 (N_1607,N_1412,N_1481);
nor U1608 (N_1608,N_1558,N_1541);
nand U1609 (N_1609,N_1589,N_1440);
or U1610 (N_1610,N_1425,N_1555);
or U1611 (N_1611,N_1441,N_1581);
nand U1612 (N_1612,N_1505,N_1451);
or U1613 (N_1613,N_1573,N_1504);
or U1614 (N_1614,N_1430,N_1512);
or U1615 (N_1615,N_1473,N_1515);
or U1616 (N_1616,N_1466,N_1547);
nor U1617 (N_1617,N_1475,N_1404);
or U1618 (N_1618,N_1542,N_1493);
nand U1619 (N_1619,N_1550,N_1546);
and U1620 (N_1620,N_1421,N_1445);
and U1621 (N_1621,N_1522,N_1486);
nor U1622 (N_1622,N_1594,N_1527);
nor U1623 (N_1623,N_1403,N_1536);
xor U1624 (N_1624,N_1407,N_1449);
and U1625 (N_1625,N_1409,N_1540);
nor U1626 (N_1626,N_1578,N_1530);
nor U1627 (N_1627,N_1569,N_1591);
nor U1628 (N_1628,N_1482,N_1458);
xor U1629 (N_1629,N_1570,N_1513);
xor U1630 (N_1630,N_1593,N_1585);
or U1631 (N_1631,N_1414,N_1438);
xnor U1632 (N_1632,N_1479,N_1496);
xor U1633 (N_1633,N_1582,N_1457);
and U1634 (N_1634,N_1519,N_1433);
nor U1635 (N_1635,N_1495,N_1419);
nor U1636 (N_1636,N_1532,N_1507);
nand U1637 (N_1637,N_1411,N_1420);
xnor U1638 (N_1638,N_1463,N_1521);
and U1639 (N_1639,N_1478,N_1565);
nand U1640 (N_1640,N_1456,N_1423);
and U1641 (N_1641,N_1447,N_1450);
and U1642 (N_1642,N_1491,N_1537);
nor U1643 (N_1643,N_1575,N_1485);
and U1644 (N_1644,N_1410,N_1413);
or U1645 (N_1645,N_1415,N_1592);
or U1646 (N_1646,N_1476,N_1516);
or U1647 (N_1647,N_1597,N_1470);
nor U1648 (N_1648,N_1439,N_1525);
nor U1649 (N_1649,N_1517,N_1535);
nand U1650 (N_1650,N_1406,N_1446);
and U1651 (N_1651,N_1544,N_1472);
nand U1652 (N_1652,N_1469,N_1598);
xnor U1653 (N_1653,N_1499,N_1417);
xor U1654 (N_1654,N_1566,N_1538);
xor U1655 (N_1655,N_1556,N_1452);
nor U1656 (N_1656,N_1477,N_1510);
and U1657 (N_1657,N_1471,N_1432);
and U1658 (N_1658,N_1545,N_1528);
and U1659 (N_1659,N_1400,N_1462);
or U1660 (N_1660,N_1436,N_1431);
and U1661 (N_1661,N_1428,N_1422);
nand U1662 (N_1662,N_1539,N_1559);
or U1663 (N_1663,N_1587,N_1574);
nor U1664 (N_1664,N_1526,N_1560);
nand U1665 (N_1665,N_1596,N_1502);
and U1666 (N_1666,N_1567,N_1568);
nor U1667 (N_1667,N_1474,N_1579);
xnor U1668 (N_1668,N_1563,N_1584);
nand U1669 (N_1669,N_1427,N_1401);
and U1670 (N_1670,N_1498,N_1424);
xnor U1671 (N_1671,N_1599,N_1551);
nand U1672 (N_1672,N_1454,N_1595);
and U1673 (N_1673,N_1590,N_1586);
nor U1674 (N_1674,N_1497,N_1464);
nand U1675 (N_1675,N_1576,N_1549);
and U1676 (N_1676,N_1416,N_1455);
xnor U1677 (N_1677,N_1467,N_1494);
and U1678 (N_1678,N_1554,N_1402);
and U1679 (N_1679,N_1426,N_1487);
nor U1680 (N_1680,N_1489,N_1448);
and U1681 (N_1681,N_1583,N_1459);
xor U1682 (N_1682,N_1533,N_1518);
nand U1683 (N_1683,N_1418,N_1514);
and U1684 (N_1684,N_1523,N_1488);
nor U1685 (N_1685,N_1552,N_1511);
or U1686 (N_1686,N_1500,N_1492);
and U1687 (N_1687,N_1437,N_1405);
nor U1688 (N_1688,N_1553,N_1557);
nand U1689 (N_1689,N_1509,N_1442);
nand U1690 (N_1690,N_1468,N_1429);
xnor U1691 (N_1691,N_1460,N_1503);
nand U1692 (N_1692,N_1465,N_1571);
or U1693 (N_1693,N_1561,N_1435);
nor U1694 (N_1694,N_1408,N_1434);
xnor U1695 (N_1695,N_1548,N_1483);
nand U1696 (N_1696,N_1534,N_1564);
or U1697 (N_1697,N_1524,N_1461);
nor U1698 (N_1698,N_1480,N_1490);
or U1699 (N_1699,N_1580,N_1508);
xnor U1700 (N_1700,N_1461,N_1480);
and U1701 (N_1701,N_1593,N_1519);
xor U1702 (N_1702,N_1474,N_1423);
nand U1703 (N_1703,N_1450,N_1445);
nor U1704 (N_1704,N_1435,N_1508);
and U1705 (N_1705,N_1524,N_1591);
nand U1706 (N_1706,N_1518,N_1402);
nand U1707 (N_1707,N_1403,N_1537);
or U1708 (N_1708,N_1456,N_1440);
or U1709 (N_1709,N_1502,N_1424);
and U1710 (N_1710,N_1450,N_1438);
and U1711 (N_1711,N_1500,N_1450);
and U1712 (N_1712,N_1599,N_1542);
and U1713 (N_1713,N_1553,N_1571);
nand U1714 (N_1714,N_1586,N_1584);
or U1715 (N_1715,N_1492,N_1598);
nand U1716 (N_1716,N_1562,N_1502);
or U1717 (N_1717,N_1568,N_1511);
nand U1718 (N_1718,N_1584,N_1541);
xor U1719 (N_1719,N_1576,N_1470);
nor U1720 (N_1720,N_1454,N_1464);
nor U1721 (N_1721,N_1454,N_1475);
xor U1722 (N_1722,N_1510,N_1437);
nor U1723 (N_1723,N_1417,N_1560);
nor U1724 (N_1724,N_1472,N_1568);
or U1725 (N_1725,N_1484,N_1592);
xnor U1726 (N_1726,N_1575,N_1543);
xor U1727 (N_1727,N_1528,N_1580);
nand U1728 (N_1728,N_1460,N_1567);
nor U1729 (N_1729,N_1510,N_1497);
and U1730 (N_1730,N_1537,N_1420);
or U1731 (N_1731,N_1402,N_1538);
and U1732 (N_1732,N_1452,N_1574);
or U1733 (N_1733,N_1406,N_1558);
and U1734 (N_1734,N_1520,N_1532);
nor U1735 (N_1735,N_1585,N_1457);
and U1736 (N_1736,N_1592,N_1557);
nand U1737 (N_1737,N_1489,N_1410);
or U1738 (N_1738,N_1582,N_1442);
nand U1739 (N_1739,N_1462,N_1587);
and U1740 (N_1740,N_1572,N_1443);
nand U1741 (N_1741,N_1542,N_1545);
nor U1742 (N_1742,N_1597,N_1530);
or U1743 (N_1743,N_1548,N_1512);
xnor U1744 (N_1744,N_1527,N_1588);
nand U1745 (N_1745,N_1580,N_1457);
nor U1746 (N_1746,N_1558,N_1453);
nor U1747 (N_1747,N_1462,N_1497);
or U1748 (N_1748,N_1554,N_1548);
and U1749 (N_1749,N_1422,N_1573);
nand U1750 (N_1750,N_1562,N_1573);
xor U1751 (N_1751,N_1579,N_1505);
nand U1752 (N_1752,N_1400,N_1468);
nor U1753 (N_1753,N_1440,N_1554);
and U1754 (N_1754,N_1414,N_1429);
and U1755 (N_1755,N_1584,N_1507);
or U1756 (N_1756,N_1580,N_1566);
nor U1757 (N_1757,N_1592,N_1423);
nor U1758 (N_1758,N_1574,N_1454);
or U1759 (N_1759,N_1593,N_1555);
nor U1760 (N_1760,N_1452,N_1442);
and U1761 (N_1761,N_1518,N_1482);
nor U1762 (N_1762,N_1415,N_1471);
xnor U1763 (N_1763,N_1479,N_1544);
nor U1764 (N_1764,N_1410,N_1559);
nand U1765 (N_1765,N_1598,N_1540);
nor U1766 (N_1766,N_1500,N_1504);
and U1767 (N_1767,N_1501,N_1427);
nor U1768 (N_1768,N_1553,N_1427);
or U1769 (N_1769,N_1562,N_1530);
xor U1770 (N_1770,N_1570,N_1512);
xor U1771 (N_1771,N_1525,N_1412);
xor U1772 (N_1772,N_1436,N_1503);
or U1773 (N_1773,N_1413,N_1521);
xor U1774 (N_1774,N_1453,N_1596);
or U1775 (N_1775,N_1580,N_1474);
or U1776 (N_1776,N_1409,N_1587);
nand U1777 (N_1777,N_1457,N_1400);
or U1778 (N_1778,N_1571,N_1500);
and U1779 (N_1779,N_1535,N_1471);
or U1780 (N_1780,N_1413,N_1475);
or U1781 (N_1781,N_1401,N_1424);
xor U1782 (N_1782,N_1459,N_1490);
or U1783 (N_1783,N_1453,N_1484);
or U1784 (N_1784,N_1480,N_1550);
nand U1785 (N_1785,N_1495,N_1543);
nor U1786 (N_1786,N_1516,N_1457);
and U1787 (N_1787,N_1427,N_1529);
and U1788 (N_1788,N_1568,N_1486);
and U1789 (N_1789,N_1538,N_1419);
xor U1790 (N_1790,N_1581,N_1552);
nand U1791 (N_1791,N_1546,N_1415);
xor U1792 (N_1792,N_1444,N_1416);
nand U1793 (N_1793,N_1447,N_1566);
nand U1794 (N_1794,N_1565,N_1447);
or U1795 (N_1795,N_1503,N_1522);
xor U1796 (N_1796,N_1558,N_1484);
xor U1797 (N_1797,N_1598,N_1429);
xor U1798 (N_1798,N_1428,N_1413);
and U1799 (N_1799,N_1503,N_1448);
nand U1800 (N_1800,N_1613,N_1696);
or U1801 (N_1801,N_1766,N_1765);
and U1802 (N_1802,N_1683,N_1713);
xnor U1803 (N_1803,N_1620,N_1758);
xor U1804 (N_1804,N_1720,N_1705);
nand U1805 (N_1805,N_1667,N_1690);
xnor U1806 (N_1806,N_1799,N_1733);
nor U1807 (N_1807,N_1751,N_1626);
nor U1808 (N_1808,N_1681,N_1777);
and U1809 (N_1809,N_1749,N_1601);
nor U1810 (N_1810,N_1687,N_1792);
nand U1811 (N_1811,N_1688,N_1776);
xnor U1812 (N_1812,N_1670,N_1628);
or U1813 (N_1813,N_1700,N_1660);
nand U1814 (N_1814,N_1662,N_1711);
and U1815 (N_1815,N_1630,N_1772);
or U1816 (N_1816,N_1656,N_1697);
xnor U1817 (N_1817,N_1605,N_1779);
nor U1818 (N_1818,N_1784,N_1666);
or U1819 (N_1819,N_1695,N_1646);
nor U1820 (N_1820,N_1633,N_1685);
nand U1821 (N_1821,N_1669,N_1638);
and U1822 (N_1822,N_1787,N_1781);
or U1823 (N_1823,N_1657,N_1727);
nand U1824 (N_1824,N_1791,N_1714);
xnor U1825 (N_1825,N_1709,N_1684);
and U1826 (N_1826,N_1736,N_1739);
xnor U1827 (N_1827,N_1724,N_1715);
or U1828 (N_1828,N_1770,N_1769);
or U1829 (N_1829,N_1655,N_1755);
nand U1830 (N_1830,N_1627,N_1742);
nor U1831 (N_1831,N_1671,N_1757);
nor U1832 (N_1832,N_1753,N_1761);
nor U1833 (N_1833,N_1722,N_1623);
xnor U1834 (N_1834,N_1756,N_1686);
or U1835 (N_1835,N_1763,N_1678);
nand U1836 (N_1836,N_1621,N_1796);
or U1837 (N_1837,N_1746,N_1743);
and U1838 (N_1838,N_1704,N_1616);
nand U1839 (N_1839,N_1634,N_1619);
and U1840 (N_1840,N_1728,N_1637);
nor U1841 (N_1841,N_1615,N_1754);
nand U1842 (N_1842,N_1734,N_1618);
and U1843 (N_1843,N_1694,N_1699);
xnor U1844 (N_1844,N_1716,N_1691);
or U1845 (N_1845,N_1760,N_1622);
or U1846 (N_1846,N_1644,N_1710);
or U1847 (N_1847,N_1659,N_1794);
or U1848 (N_1848,N_1707,N_1698);
or U1849 (N_1849,N_1782,N_1617);
xnor U1850 (N_1850,N_1729,N_1653);
or U1851 (N_1851,N_1737,N_1732);
nand U1852 (N_1852,N_1680,N_1606);
or U1853 (N_1853,N_1668,N_1677);
nor U1854 (N_1854,N_1672,N_1611);
nand U1855 (N_1855,N_1730,N_1645);
nand U1856 (N_1856,N_1648,N_1676);
nand U1857 (N_1857,N_1726,N_1786);
or U1858 (N_1858,N_1759,N_1624);
or U1859 (N_1859,N_1798,N_1607);
and U1860 (N_1860,N_1775,N_1712);
nor U1861 (N_1861,N_1767,N_1641);
and U1862 (N_1862,N_1702,N_1738);
xor U1863 (N_1863,N_1762,N_1604);
and U1864 (N_1864,N_1706,N_1647);
or U1865 (N_1865,N_1747,N_1797);
or U1866 (N_1866,N_1740,N_1643);
nand U1867 (N_1867,N_1771,N_1631);
and U1868 (N_1868,N_1674,N_1750);
nand U1869 (N_1869,N_1741,N_1636);
nand U1870 (N_1870,N_1719,N_1793);
or U1871 (N_1871,N_1774,N_1651);
nand U1872 (N_1872,N_1639,N_1723);
nand U1873 (N_1873,N_1752,N_1768);
or U1874 (N_1874,N_1795,N_1612);
nor U1875 (N_1875,N_1679,N_1790);
xnor U1876 (N_1876,N_1783,N_1654);
nor U1877 (N_1877,N_1785,N_1600);
nor U1878 (N_1878,N_1635,N_1778);
nand U1879 (N_1879,N_1652,N_1614);
or U1880 (N_1880,N_1689,N_1673);
and U1881 (N_1881,N_1629,N_1632);
nor U1882 (N_1882,N_1675,N_1650);
xor U1883 (N_1883,N_1764,N_1748);
or U1884 (N_1884,N_1665,N_1708);
xor U1885 (N_1885,N_1701,N_1731);
and U1886 (N_1886,N_1664,N_1640);
nand U1887 (N_1887,N_1745,N_1603);
or U1888 (N_1888,N_1642,N_1780);
and U1889 (N_1889,N_1744,N_1625);
nor U1890 (N_1890,N_1773,N_1658);
nor U1891 (N_1891,N_1649,N_1608);
nand U1892 (N_1892,N_1692,N_1788);
nor U1893 (N_1893,N_1718,N_1661);
and U1894 (N_1894,N_1721,N_1610);
and U1895 (N_1895,N_1789,N_1735);
xnor U1896 (N_1896,N_1602,N_1663);
xnor U1897 (N_1897,N_1725,N_1703);
and U1898 (N_1898,N_1609,N_1682);
xnor U1899 (N_1899,N_1717,N_1693);
nand U1900 (N_1900,N_1772,N_1722);
and U1901 (N_1901,N_1631,N_1686);
or U1902 (N_1902,N_1750,N_1649);
nor U1903 (N_1903,N_1630,N_1739);
and U1904 (N_1904,N_1736,N_1707);
nand U1905 (N_1905,N_1685,N_1700);
nand U1906 (N_1906,N_1787,N_1621);
or U1907 (N_1907,N_1772,N_1728);
xor U1908 (N_1908,N_1738,N_1687);
nor U1909 (N_1909,N_1602,N_1756);
nand U1910 (N_1910,N_1682,N_1728);
nand U1911 (N_1911,N_1644,N_1601);
and U1912 (N_1912,N_1779,N_1614);
xor U1913 (N_1913,N_1676,N_1682);
nand U1914 (N_1914,N_1653,N_1796);
or U1915 (N_1915,N_1797,N_1746);
nand U1916 (N_1916,N_1726,N_1634);
and U1917 (N_1917,N_1798,N_1797);
xor U1918 (N_1918,N_1657,N_1774);
xnor U1919 (N_1919,N_1616,N_1759);
xor U1920 (N_1920,N_1775,N_1692);
nor U1921 (N_1921,N_1620,N_1791);
nand U1922 (N_1922,N_1626,N_1649);
xor U1923 (N_1923,N_1639,N_1631);
and U1924 (N_1924,N_1799,N_1779);
or U1925 (N_1925,N_1636,N_1732);
nor U1926 (N_1926,N_1607,N_1764);
and U1927 (N_1927,N_1617,N_1609);
or U1928 (N_1928,N_1664,N_1787);
and U1929 (N_1929,N_1670,N_1634);
or U1930 (N_1930,N_1740,N_1605);
xor U1931 (N_1931,N_1794,N_1620);
or U1932 (N_1932,N_1661,N_1726);
xor U1933 (N_1933,N_1706,N_1798);
and U1934 (N_1934,N_1799,N_1774);
or U1935 (N_1935,N_1691,N_1777);
and U1936 (N_1936,N_1763,N_1758);
nor U1937 (N_1937,N_1702,N_1785);
and U1938 (N_1938,N_1788,N_1677);
nor U1939 (N_1939,N_1796,N_1752);
and U1940 (N_1940,N_1686,N_1627);
xor U1941 (N_1941,N_1714,N_1676);
xor U1942 (N_1942,N_1687,N_1614);
xor U1943 (N_1943,N_1783,N_1676);
nor U1944 (N_1944,N_1611,N_1668);
nand U1945 (N_1945,N_1651,N_1709);
or U1946 (N_1946,N_1745,N_1607);
and U1947 (N_1947,N_1606,N_1727);
xor U1948 (N_1948,N_1646,N_1788);
and U1949 (N_1949,N_1688,N_1749);
xor U1950 (N_1950,N_1691,N_1737);
or U1951 (N_1951,N_1738,N_1714);
xor U1952 (N_1952,N_1758,N_1694);
nor U1953 (N_1953,N_1734,N_1769);
or U1954 (N_1954,N_1769,N_1676);
nand U1955 (N_1955,N_1654,N_1645);
nor U1956 (N_1956,N_1675,N_1783);
nand U1957 (N_1957,N_1682,N_1651);
and U1958 (N_1958,N_1628,N_1730);
and U1959 (N_1959,N_1612,N_1757);
or U1960 (N_1960,N_1759,N_1708);
and U1961 (N_1961,N_1698,N_1673);
xor U1962 (N_1962,N_1640,N_1618);
nand U1963 (N_1963,N_1646,N_1783);
nand U1964 (N_1964,N_1625,N_1701);
nor U1965 (N_1965,N_1771,N_1666);
nor U1966 (N_1966,N_1627,N_1741);
xnor U1967 (N_1967,N_1627,N_1784);
and U1968 (N_1968,N_1761,N_1702);
xnor U1969 (N_1969,N_1784,N_1651);
nor U1970 (N_1970,N_1654,N_1656);
xor U1971 (N_1971,N_1746,N_1684);
nand U1972 (N_1972,N_1641,N_1691);
or U1973 (N_1973,N_1712,N_1693);
nor U1974 (N_1974,N_1706,N_1620);
nand U1975 (N_1975,N_1664,N_1783);
and U1976 (N_1976,N_1715,N_1705);
and U1977 (N_1977,N_1642,N_1623);
nor U1978 (N_1978,N_1767,N_1664);
nand U1979 (N_1979,N_1785,N_1664);
nand U1980 (N_1980,N_1703,N_1606);
and U1981 (N_1981,N_1691,N_1704);
nor U1982 (N_1982,N_1748,N_1651);
and U1983 (N_1983,N_1689,N_1621);
nand U1984 (N_1984,N_1788,N_1690);
xor U1985 (N_1985,N_1741,N_1689);
nand U1986 (N_1986,N_1752,N_1712);
and U1987 (N_1987,N_1790,N_1777);
nor U1988 (N_1988,N_1714,N_1707);
or U1989 (N_1989,N_1718,N_1799);
xnor U1990 (N_1990,N_1619,N_1605);
and U1991 (N_1991,N_1637,N_1649);
and U1992 (N_1992,N_1611,N_1656);
nor U1993 (N_1993,N_1754,N_1699);
xor U1994 (N_1994,N_1758,N_1713);
xor U1995 (N_1995,N_1766,N_1763);
nor U1996 (N_1996,N_1647,N_1688);
or U1997 (N_1997,N_1664,N_1760);
nand U1998 (N_1998,N_1646,N_1610);
nor U1999 (N_1999,N_1613,N_1671);
nor U2000 (N_2000,N_1817,N_1903);
or U2001 (N_2001,N_1944,N_1839);
and U2002 (N_2002,N_1917,N_1874);
and U2003 (N_2003,N_1900,N_1985);
nand U2004 (N_2004,N_1858,N_1881);
and U2005 (N_2005,N_1921,N_1904);
xnor U2006 (N_2006,N_1989,N_1928);
xor U2007 (N_2007,N_1969,N_1870);
nor U2008 (N_2008,N_1841,N_1914);
or U2009 (N_2009,N_1978,N_1923);
xnor U2010 (N_2010,N_1962,N_1851);
nand U2011 (N_2011,N_1803,N_1860);
xnor U2012 (N_2012,N_1953,N_1902);
nor U2013 (N_2013,N_1849,N_1973);
and U2014 (N_2014,N_1826,N_1875);
nand U2015 (N_2015,N_1886,N_1888);
nand U2016 (N_2016,N_1949,N_1837);
nor U2017 (N_2017,N_1877,N_1807);
xnor U2018 (N_2018,N_1983,N_1979);
nand U2019 (N_2019,N_1905,N_1846);
xnor U2020 (N_2020,N_1899,N_1880);
nor U2021 (N_2021,N_1920,N_1852);
nor U2022 (N_2022,N_1993,N_1943);
xor U2023 (N_2023,N_1857,N_1977);
nor U2024 (N_2024,N_1980,N_1909);
and U2025 (N_2025,N_1862,N_1997);
xnor U2026 (N_2026,N_1891,N_1829);
nor U2027 (N_2027,N_1879,N_1840);
nand U2028 (N_2028,N_1810,N_1935);
and U2029 (N_2029,N_1984,N_1827);
xor U2030 (N_2030,N_1843,N_1883);
xor U2031 (N_2031,N_1863,N_1834);
xor U2032 (N_2032,N_1975,N_1919);
nand U2033 (N_2033,N_1866,N_1882);
or U2034 (N_2034,N_1836,N_1832);
or U2035 (N_2035,N_1824,N_1945);
and U2036 (N_2036,N_1815,N_1897);
and U2037 (N_2037,N_1952,N_1901);
and U2038 (N_2038,N_1936,N_1848);
and U2039 (N_2039,N_1987,N_1964);
nor U2040 (N_2040,N_1842,N_1868);
xnor U2041 (N_2041,N_1820,N_1951);
or U2042 (N_2042,N_1916,N_1976);
nor U2043 (N_2043,N_1992,N_1942);
or U2044 (N_2044,N_1924,N_1999);
nor U2045 (N_2045,N_1885,N_1871);
xor U2046 (N_2046,N_1922,N_1908);
nand U2047 (N_2047,N_1811,N_1889);
nand U2048 (N_2048,N_1938,N_1963);
nor U2049 (N_2049,N_1825,N_1933);
and U2050 (N_2050,N_1828,N_1876);
nand U2051 (N_2051,N_1958,N_1996);
nand U2052 (N_2052,N_1872,N_1910);
or U2053 (N_2053,N_1971,N_1954);
or U2054 (N_2054,N_1847,N_1890);
nand U2055 (N_2055,N_1819,N_1844);
nor U2056 (N_2056,N_1855,N_1995);
nand U2057 (N_2057,N_1966,N_1986);
nor U2058 (N_2058,N_1906,N_1927);
or U2059 (N_2059,N_1925,N_1968);
xor U2060 (N_2060,N_1974,N_1961);
nand U2061 (N_2061,N_1965,N_1895);
or U2062 (N_2062,N_1934,N_1887);
nand U2063 (N_2063,N_1960,N_1854);
nand U2064 (N_2064,N_1896,N_1864);
and U2065 (N_2065,N_1835,N_1816);
or U2066 (N_2066,N_1818,N_1931);
and U2067 (N_2067,N_1937,N_1939);
or U2068 (N_2068,N_1956,N_1821);
or U2069 (N_2069,N_1845,N_1959);
xor U2070 (N_2070,N_1941,N_1981);
and U2071 (N_2071,N_1957,N_1806);
and U2072 (N_2072,N_1893,N_1915);
nand U2073 (N_2073,N_1929,N_1808);
and U2074 (N_2074,N_1946,N_1898);
nand U2075 (N_2075,N_1833,N_1907);
or U2076 (N_2076,N_1918,N_1894);
or U2077 (N_2077,N_1804,N_1991);
xor U2078 (N_2078,N_1912,N_1955);
nand U2079 (N_2079,N_1911,N_1809);
nor U2080 (N_2080,N_1801,N_1913);
or U2081 (N_2081,N_1967,N_1932);
nand U2082 (N_2082,N_1970,N_1800);
or U2083 (N_2083,N_1994,N_1859);
nor U2084 (N_2084,N_1813,N_1823);
nor U2085 (N_2085,N_1950,N_1865);
and U2086 (N_2086,N_1814,N_1873);
nand U2087 (N_2087,N_1831,N_1892);
and U2088 (N_2088,N_1972,N_1990);
xnor U2089 (N_2089,N_1988,N_1850);
and U2090 (N_2090,N_1930,N_1861);
nand U2091 (N_2091,N_1856,N_1926);
and U2092 (N_2092,N_1867,N_1982);
nor U2093 (N_2093,N_1998,N_1940);
xnor U2094 (N_2094,N_1805,N_1838);
nand U2095 (N_2095,N_1853,N_1822);
or U2096 (N_2096,N_1869,N_1812);
nor U2097 (N_2097,N_1878,N_1947);
xor U2098 (N_2098,N_1830,N_1948);
nor U2099 (N_2099,N_1802,N_1884);
and U2100 (N_2100,N_1966,N_1835);
or U2101 (N_2101,N_1939,N_1996);
nor U2102 (N_2102,N_1979,N_1862);
nand U2103 (N_2103,N_1839,N_1994);
nor U2104 (N_2104,N_1831,N_1815);
xor U2105 (N_2105,N_1985,N_1924);
and U2106 (N_2106,N_1857,N_1998);
xor U2107 (N_2107,N_1926,N_1919);
or U2108 (N_2108,N_1970,N_1803);
nand U2109 (N_2109,N_1879,N_1978);
and U2110 (N_2110,N_1902,N_1890);
nand U2111 (N_2111,N_1958,N_1989);
and U2112 (N_2112,N_1889,N_1945);
nor U2113 (N_2113,N_1905,N_1839);
and U2114 (N_2114,N_1866,N_1800);
nand U2115 (N_2115,N_1874,N_1803);
xnor U2116 (N_2116,N_1888,N_1836);
xnor U2117 (N_2117,N_1802,N_1937);
nor U2118 (N_2118,N_1952,N_1976);
or U2119 (N_2119,N_1833,N_1951);
and U2120 (N_2120,N_1916,N_1945);
and U2121 (N_2121,N_1944,N_1860);
nand U2122 (N_2122,N_1853,N_1927);
nor U2123 (N_2123,N_1947,N_1901);
and U2124 (N_2124,N_1957,N_1885);
nor U2125 (N_2125,N_1959,N_1877);
xnor U2126 (N_2126,N_1958,N_1837);
xor U2127 (N_2127,N_1933,N_1938);
or U2128 (N_2128,N_1936,N_1880);
xor U2129 (N_2129,N_1808,N_1853);
or U2130 (N_2130,N_1847,N_1949);
nand U2131 (N_2131,N_1910,N_1893);
and U2132 (N_2132,N_1846,N_1818);
and U2133 (N_2133,N_1981,N_1927);
xnor U2134 (N_2134,N_1931,N_1928);
nor U2135 (N_2135,N_1918,N_1847);
xor U2136 (N_2136,N_1877,N_1858);
and U2137 (N_2137,N_1969,N_1907);
xnor U2138 (N_2138,N_1882,N_1902);
nor U2139 (N_2139,N_1871,N_1979);
nand U2140 (N_2140,N_1916,N_1804);
nor U2141 (N_2141,N_1935,N_1917);
or U2142 (N_2142,N_1964,N_1880);
nand U2143 (N_2143,N_1977,N_1855);
or U2144 (N_2144,N_1953,N_1916);
and U2145 (N_2145,N_1921,N_1811);
and U2146 (N_2146,N_1907,N_1865);
xnor U2147 (N_2147,N_1861,N_1905);
nor U2148 (N_2148,N_1803,N_1944);
and U2149 (N_2149,N_1982,N_1952);
and U2150 (N_2150,N_1933,N_1949);
nand U2151 (N_2151,N_1817,N_1966);
and U2152 (N_2152,N_1933,N_1856);
nand U2153 (N_2153,N_1819,N_1946);
or U2154 (N_2154,N_1964,N_1906);
or U2155 (N_2155,N_1837,N_1923);
nand U2156 (N_2156,N_1946,N_1948);
or U2157 (N_2157,N_1806,N_1856);
nor U2158 (N_2158,N_1844,N_1988);
or U2159 (N_2159,N_1865,N_1973);
nand U2160 (N_2160,N_1933,N_1975);
nor U2161 (N_2161,N_1897,N_1873);
nor U2162 (N_2162,N_1819,N_1869);
xor U2163 (N_2163,N_1936,N_1956);
nor U2164 (N_2164,N_1925,N_1867);
or U2165 (N_2165,N_1827,N_1873);
xnor U2166 (N_2166,N_1929,N_1800);
and U2167 (N_2167,N_1985,N_1908);
nor U2168 (N_2168,N_1853,N_1960);
nand U2169 (N_2169,N_1995,N_1894);
nor U2170 (N_2170,N_1858,N_1984);
or U2171 (N_2171,N_1903,N_1832);
xnor U2172 (N_2172,N_1939,N_1994);
or U2173 (N_2173,N_1875,N_1907);
nand U2174 (N_2174,N_1896,N_1941);
nand U2175 (N_2175,N_1885,N_1931);
and U2176 (N_2176,N_1854,N_1913);
nor U2177 (N_2177,N_1995,N_1931);
and U2178 (N_2178,N_1859,N_1993);
xnor U2179 (N_2179,N_1811,N_1960);
xnor U2180 (N_2180,N_1939,N_1817);
or U2181 (N_2181,N_1823,N_1951);
and U2182 (N_2182,N_1816,N_1952);
nand U2183 (N_2183,N_1935,N_1945);
nor U2184 (N_2184,N_1989,N_1831);
nor U2185 (N_2185,N_1984,N_1828);
nor U2186 (N_2186,N_1800,N_1981);
nor U2187 (N_2187,N_1878,N_1920);
or U2188 (N_2188,N_1870,N_1990);
and U2189 (N_2189,N_1914,N_1949);
or U2190 (N_2190,N_1902,N_1839);
nor U2191 (N_2191,N_1944,N_1955);
nand U2192 (N_2192,N_1979,N_1881);
nor U2193 (N_2193,N_1895,N_1932);
nand U2194 (N_2194,N_1891,N_1861);
nand U2195 (N_2195,N_1818,N_1826);
nor U2196 (N_2196,N_1880,N_1944);
xor U2197 (N_2197,N_1815,N_1848);
or U2198 (N_2198,N_1811,N_1945);
and U2199 (N_2199,N_1996,N_1921);
nand U2200 (N_2200,N_2166,N_2195);
or U2201 (N_2201,N_2051,N_2174);
nand U2202 (N_2202,N_2160,N_2128);
nand U2203 (N_2203,N_2086,N_2062);
or U2204 (N_2204,N_2104,N_2190);
or U2205 (N_2205,N_2061,N_2025);
xnor U2206 (N_2206,N_2198,N_2108);
nand U2207 (N_2207,N_2076,N_2168);
xnor U2208 (N_2208,N_2175,N_2002);
and U2209 (N_2209,N_2043,N_2155);
xor U2210 (N_2210,N_2112,N_2094);
or U2211 (N_2211,N_2079,N_2069);
and U2212 (N_2212,N_2030,N_2129);
xor U2213 (N_2213,N_2167,N_2189);
or U2214 (N_2214,N_2145,N_2115);
nand U2215 (N_2215,N_2153,N_2091);
nand U2216 (N_2216,N_2044,N_2009);
or U2217 (N_2217,N_2151,N_2125);
and U2218 (N_2218,N_2032,N_2133);
and U2219 (N_2219,N_2197,N_2154);
or U2220 (N_2220,N_2029,N_2144);
or U2221 (N_2221,N_2005,N_2057);
nor U2222 (N_2222,N_2063,N_2089);
and U2223 (N_2223,N_2078,N_2090);
or U2224 (N_2224,N_2182,N_2018);
and U2225 (N_2225,N_2105,N_2085);
nand U2226 (N_2226,N_2040,N_2184);
or U2227 (N_2227,N_2081,N_2056);
and U2228 (N_2228,N_2045,N_2121);
nor U2229 (N_2229,N_2047,N_2074);
and U2230 (N_2230,N_2180,N_2116);
nand U2231 (N_2231,N_2146,N_2077);
nand U2232 (N_2232,N_2082,N_2120);
nor U2233 (N_2233,N_2194,N_2021);
nor U2234 (N_2234,N_2013,N_2124);
xor U2235 (N_2235,N_2165,N_2114);
or U2236 (N_2236,N_2031,N_2024);
xnor U2237 (N_2237,N_2000,N_2141);
and U2238 (N_2238,N_2126,N_2117);
xor U2239 (N_2239,N_2033,N_2035);
or U2240 (N_2240,N_2132,N_2148);
nand U2241 (N_2241,N_2158,N_2064);
xor U2242 (N_2242,N_2176,N_2007);
xor U2243 (N_2243,N_2138,N_2008);
and U2244 (N_2244,N_2017,N_2097);
and U2245 (N_2245,N_2075,N_2173);
and U2246 (N_2246,N_2011,N_2123);
nand U2247 (N_2247,N_2119,N_2196);
or U2248 (N_2248,N_2058,N_2172);
and U2249 (N_2249,N_2059,N_2037);
and U2250 (N_2250,N_2068,N_2093);
or U2251 (N_2251,N_2080,N_2046);
and U2252 (N_2252,N_2187,N_2052);
xor U2253 (N_2253,N_2053,N_2071);
nand U2254 (N_2254,N_2065,N_2183);
and U2255 (N_2255,N_2050,N_2060);
and U2256 (N_2256,N_2098,N_2113);
xor U2257 (N_2257,N_2101,N_2072);
nand U2258 (N_2258,N_2073,N_2162);
nand U2259 (N_2259,N_2041,N_2088);
and U2260 (N_2260,N_2022,N_2039);
or U2261 (N_2261,N_2163,N_2066);
or U2262 (N_2262,N_2042,N_2134);
and U2263 (N_2263,N_2193,N_2135);
nor U2264 (N_2264,N_2014,N_2122);
nor U2265 (N_2265,N_2107,N_2103);
xnor U2266 (N_2266,N_2136,N_2012);
and U2267 (N_2267,N_2001,N_2164);
or U2268 (N_2268,N_2054,N_2087);
xnor U2269 (N_2269,N_2055,N_2131);
xor U2270 (N_2270,N_2178,N_2192);
and U2271 (N_2271,N_2161,N_2156);
nand U2272 (N_2272,N_2004,N_2099);
nor U2273 (N_2273,N_2179,N_2102);
and U2274 (N_2274,N_2048,N_2177);
nand U2275 (N_2275,N_2109,N_2152);
xor U2276 (N_2276,N_2095,N_2027);
nand U2277 (N_2277,N_2150,N_2169);
or U2278 (N_2278,N_2100,N_2159);
and U2279 (N_2279,N_2067,N_2015);
nand U2280 (N_2280,N_2096,N_2147);
nand U2281 (N_2281,N_2016,N_2111);
nor U2282 (N_2282,N_2139,N_2185);
and U2283 (N_2283,N_2191,N_2110);
and U2284 (N_2284,N_2020,N_2049);
or U2285 (N_2285,N_2023,N_2130);
and U2286 (N_2286,N_2010,N_2026);
xor U2287 (N_2287,N_2170,N_2019);
and U2288 (N_2288,N_2083,N_2149);
xor U2289 (N_2289,N_2118,N_2106);
nor U2290 (N_2290,N_2028,N_2181);
or U2291 (N_2291,N_2186,N_2084);
or U2292 (N_2292,N_2157,N_2142);
or U2293 (N_2293,N_2140,N_2171);
or U2294 (N_2294,N_2092,N_2036);
xnor U2295 (N_2295,N_2143,N_2003);
nor U2296 (N_2296,N_2137,N_2006);
or U2297 (N_2297,N_2038,N_2199);
or U2298 (N_2298,N_2127,N_2070);
nand U2299 (N_2299,N_2034,N_2188);
and U2300 (N_2300,N_2073,N_2021);
or U2301 (N_2301,N_2005,N_2069);
xnor U2302 (N_2302,N_2082,N_2137);
and U2303 (N_2303,N_2100,N_2042);
or U2304 (N_2304,N_2119,N_2128);
and U2305 (N_2305,N_2192,N_2090);
xnor U2306 (N_2306,N_2108,N_2004);
or U2307 (N_2307,N_2038,N_2048);
nor U2308 (N_2308,N_2159,N_2188);
or U2309 (N_2309,N_2138,N_2096);
nor U2310 (N_2310,N_2116,N_2006);
nand U2311 (N_2311,N_2137,N_2129);
or U2312 (N_2312,N_2069,N_2001);
xnor U2313 (N_2313,N_2165,N_2175);
or U2314 (N_2314,N_2098,N_2022);
or U2315 (N_2315,N_2066,N_2015);
or U2316 (N_2316,N_2199,N_2148);
or U2317 (N_2317,N_2074,N_2058);
nand U2318 (N_2318,N_2086,N_2199);
or U2319 (N_2319,N_2062,N_2156);
or U2320 (N_2320,N_2128,N_2010);
xnor U2321 (N_2321,N_2194,N_2060);
or U2322 (N_2322,N_2012,N_2180);
and U2323 (N_2323,N_2179,N_2123);
nor U2324 (N_2324,N_2045,N_2032);
xnor U2325 (N_2325,N_2009,N_2029);
and U2326 (N_2326,N_2139,N_2069);
and U2327 (N_2327,N_2088,N_2104);
or U2328 (N_2328,N_2077,N_2141);
and U2329 (N_2329,N_2147,N_2056);
xnor U2330 (N_2330,N_2069,N_2004);
or U2331 (N_2331,N_2181,N_2195);
nor U2332 (N_2332,N_2071,N_2042);
or U2333 (N_2333,N_2020,N_2050);
nand U2334 (N_2334,N_2143,N_2046);
and U2335 (N_2335,N_2130,N_2101);
nand U2336 (N_2336,N_2102,N_2169);
nand U2337 (N_2337,N_2046,N_2075);
nor U2338 (N_2338,N_2112,N_2071);
and U2339 (N_2339,N_2177,N_2001);
xor U2340 (N_2340,N_2110,N_2096);
xnor U2341 (N_2341,N_2147,N_2079);
nand U2342 (N_2342,N_2005,N_2101);
or U2343 (N_2343,N_2136,N_2072);
or U2344 (N_2344,N_2196,N_2003);
and U2345 (N_2345,N_2184,N_2117);
or U2346 (N_2346,N_2130,N_2155);
nor U2347 (N_2347,N_2172,N_2127);
or U2348 (N_2348,N_2199,N_2010);
xor U2349 (N_2349,N_2161,N_2107);
and U2350 (N_2350,N_2111,N_2015);
xor U2351 (N_2351,N_2113,N_2172);
nand U2352 (N_2352,N_2165,N_2071);
nand U2353 (N_2353,N_2108,N_2164);
nand U2354 (N_2354,N_2064,N_2122);
xor U2355 (N_2355,N_2176,N_2161);
nand U2356 (N_2356,N_2188,N_2193);
and U2357 (N_2357,N_2143,N_2101);
nand U2358 (N_2358,N_2060,N_2006);
and U2359 (N_2359,N_2084,N_2065);
xnor U2360 (N_2360,N_2169,N_2056);
and U2361 (N_2361,N_2128,N_2058);
nand U2362 (N_2362,N_2060,N_2092);
or U2363 (N_2363,N_2188,N_2010);
nand U2364 (N_2364,N_2099,N_2058);
xor U2365 (N_2365,N_2077,N_2032);
nand U2366 (N_2366,N_2100,N_2133);
or U2367 (N_2367,N_2152,N_2139);
and U2368 (N_2368,N_2121,N_2063);
or U2369 (N_2369,N_2149,N_2067);
nor U2370 (N_2370,N_2056,N_2040);
nand U2371 (N_2371,N_2063,N_2031);
xor U2372 (N_2372,N_2105,N_2086);
and U2373 (N_2373,N_2020,N_2085);
nand U2374 (N_2374,N_2155,N_2023);
xor U2375 (N_2375,N_2110,N_2091);
nor U2376 (N_2376,N_2129,N_2051);
and U2377 (N_2377,N_2098,N_2195);
nand U2378 (N_2378,N_2123,N_2111);
nor U2379 (N_2379,N_2176,N_2169);
nand U2380 (N_2380,N_2088,N_2121);
and U2381 (N_2381,N_2112,N_2017);
and U2382 (N_2382,N_2064,N_2073);
xor U2383 (N_2383,N_2024,N_2101);
xnor U2384 (N_2384,N_2031,N_2119);
nand U2385 (N_2385,N_2061,N_2139);
nand U2386 (N_2386,N_2126,N_2181);
nand U2387 (N_2387,N_2101,N_2033);
nor U2388 (N_2388,N_2081,N_2136);
xor U2389 (N_2389,N_2152,N_2141);
nor U2390 (N_2390,N_2019,N_2103);
and U2391 (N_2391,N_2081,N_2167);
xnor U2392 (N_2392,N_2001,N_2052);
and U2393 (N_2393,N_2138,N_2165);
or U2394 (N_2394,N_2107,N_2143);
xnor U2395 (N_2395,N_2090,N_2057);
xor U2396 (N_2396,N_2018,N_2025);
nor U2397 (N_2397,N_2006,N_2134);
xnor U2398 (N_2398,N_2064,N_2183);
nand U2399 (N_2399,N_2056,N_2117);
nor U2400 (N_2400,N_2394,N_2309);
nor U2401 (N_2401,N_2390,N_2310);
xor U2402 (N_2402,N_2325,N_2367);
nand U2403 (N_2403,N_2202,N_2270);
nor U2404 (N_2404,N_2350,N_2303);
xnor U2405 (N_2405,N_2340,N_2339);
xor U2406 (N_2406,N_2263,N_2330);
xor U2407 (N_2407,N_2268,N_2200);
nand U2408 (N_2408,N_2292,N_2341);
or U2409 (N_2409,N_2369,N_2229);
nand U2410 (N_2410,N_2354,N_2274);
nand U2411 (N_2411,N_2223,N_2289);
xnor U2412 (N_2412,N_2294,N_2320);
nand U2413 (N_2413,N_2252,N_2284);
nand U2414 (N_2414,N_2346,N_2238);
and U2415 (N_2415,N_2269,N_2352);
and U2416 (N_2416,N_2312,N_2226);
or U2417 (N_2417,N_2286,N_2281);
or U2418 (N_2418,N_2391,N_2398);
or U2419 (N_2419,N_2323,N_2243);
nor U2420 (N_2420,N_2258,N_2218);
and U2421 (N_2421,N_2212,N_2392);
nor U2422 (N_2422,N_2311,N_2383);
or U2423 (N_2423,N_2228,N_2373);
or U2424 (N_2424,N_2201,N_2355);
xor U2425 (N_2425,N_2318,N_2375);
nor U2426 (N_2426,N_2211,N_2272);
nor U2427 (N_2427,N_2280,N_2271);
or U2428 (N_2428,N_2363,N_2384);
and U2429 (N_2429,N_2347,N_2360);
nor U2430 (N_2430,N_2255,N_2351);
xnor U2431 (N_2431,N_2216,N_2248);
nand U2432 (N_2432,N_2316,N_2277);
nand U2433 (N_2433,N_2356,N_2285);
nand U2434 (N_2434,N_2365,N_2338);
nand U2435 (N_2435,N_2334,N_2247);
xor U2436 (N_2436,N_2397,N_2307);
xnor U2437 (N_2437,N_2332,N_2329);
or U2438 (N_2438,N_2293,N_2237);
nand U2439 (N_2439,N_2287,N_2209);
xor U2440 (N_2440,N_2396,N_2336);
nor U2441 (N_2441,N_2388,N_2317);
or U2442 (N_2442,N_2227,N_2377);
xor U2443 (N_2443,N_2386,N_2379);
or U2444 (N_2444,N_2273,N_2308);
nor U2445 (N_2445,N_2245,N_2244);
nand U2446 (N_2446,N_2264,N_2306);
xnor U2447 (N_2447,N_2222,N_2239);
nor U2448 (N_2448,N_2385,N_2328);
or U2449 (N_2449,N_2275,N_2297);
xnor U2450 (N_2450,N_2298,N_2235);
xnor U2451 (N_2451,N_2305,N_2358);
or U2452 (N_2452,N_2300,N_2389);
nor U2453 (N_2453,N_2242,N_2378);
or U2454 (N_2454,N_2261,N_2319);
nor U2455 (N_2455,N_2322,N_2232);
xnor U2456 (N_2456,N_2224,N_2205);
xor U2457 (N_2457,N_2314,N_2236);
xor U2458 (N_2458,N_2208,N_2324);
xor U2459 (N_2459,N_2246,N_2331);
or U2460 (N_2460,N_2374,N_2395);
and U2461 (N_2461,N_2370,N_2299);
nor U2462 (N_2462,N_2254,N_2234);
nor U2463 (N_2463,N_2206,N_2204);
nand U2464 (N_2464,N_2219,N_2344);
xnor U2465 (N_2465,N_2262,N_2296);
nor U2466 (N_2466,N_2362,N_2326);
or U2467 (N_2467,N_2315,N_2295);
xnor U2468 (N_2468,N_2221,N_2371);
and U2469 (N_2469,N_2203,N_2220);
xor U2470 (N_2470,N_2333,N_2380);
or U2471 (N_2471,N_2256,N_2345);
nor U2472 (N_2472,N_2327,N_2357);
nand U2473 (N_2473,N_2349,N_2278);
and U2474 (N_2474,N_2387,N_2207);
and U2475 (N_2475,N_2257,N_2260);
xor U2476 (N_2476,N_2214,N_2215);
and U2477 (N_2477,N_2361,N_2279);
nor U2478 (N_2478,N_2267,N_2399);
or U2479 (N_2479,N_2233,N_2240);
nand U2480 (N_2480,N_2359,N_2366);
and U2481 (N_2481,N_2230,N_2290);
or U2482 (N_2482,N_2376,N_2335);
xor U2483 (N_2483,N_2353,N_2259);
nor U2484 (N_2484,N_2381,N_2253);
or U2485 (N_2485,N_2217,N_2321);
nor U2486 (N_2486,N_2291,N_2342);
nand U2487 (N_2487,N_2231,N_2393);
and U2488 (N_2488,N_2313,N_2251);
xnor U2489 (N_2489,N_2250,N_2265);
nand U2490 (N_2490,N_2266,N_2301);
nand U2491 (N_2491,N_2276,N_2210);
and U2492 (N_2492,N_2337,N_2288);
nand U2493 (N_2493,N_2225,N_2304);
xor U2494 (N_2494,N_2364,N_2213);
and U2495 (N_2495,N_2249,N_2343);
nand U2496 (N_2496,N_2302,N_2382);
nor U2497 (N_2497,N_2348,N_2282);
xnor U2498 (N_2498,N_2372,N_2283);
xnor U2499 (N_2499,N_2368,N_2241);
nand U2500 (N_2500,N_2358,N_2275);
or U2501 (N_2501,N_2255,N_2239);
nand U2502 (N_2502,N_2220,N_2295);
nor U2503 (N_2503,N_2359,N_2345);
xor U2504 (N_2504,N_2352,N_2275);
nor U2505 (N_2505,N_2305,N_2324);
or U2506 (N_2506,N_2350,N_2397);
and U2507 (N_2507,N_2363,N_2313);
nor U2508 (N_2508,N_2251,N_2377);
nand U2509 (N_2509,N_2255,N_2265);
or U2510 (N_2510,N_2246,N_2322);
nand U2511 (N_2511,N_2297,N_2353);
or U2512 (N_2512,N_2365,N_2226);
xor U2513 (N_2513,N_2378,N_2368);
or U2514 (N_2514,N_2318,N_2342);
and U2515 (N_2515,N_2310,N_2345);
nor U2516 (N_2516,N_2280,N_2208);
nand U2517 (N_2517,N_2348,N_2212);
xor U2518 (N_2518,N_2208,N_2219);
or U2519 (N_2519,N_2229,N_2228);
xnor U2520 (N_2520,N_2247,N_2305);
nor U2521 (N_2521,N_2225,N_2335);
nor U2522 (N_2522,N_2261,N_2241);
nor U2523 (N_2523,N_2269,N_2281);
nand U2524 (N_2524,N_2305,N_2303);
nor U2525 (N_2525,N_2285,N_2265);
and U2526 (N_2526,N_2242,N_2247);
or U2527 (N_2527,N_2351,N_2219);
or U2528 (N_2528,N_2398,N_2245);
nand U2529 (N_2529,N_2297,N_2339);
and U2530 (N_2530,N_2255,N_2262);
nor U2531 (N_2531,N_2245,N_2370);
nand U2532 (N_2532,N_2300,N_2256);
and U2533 (N_2533,N_2371,N_2329);
xnor U2534 (N_2534,N_2262,N_2364);
and U2535 (N_2535,N_2324,N_2252);
xor U2536 (N_2536,N_2246,N_2391);
nand U2537 (N_2537,N_2358,N_2265);
nand U2538 (N_2538,N_2300,N_2387);
nor U2539 (N_2539,N_2215,N_2206);
nand U2540 (N_2540,N_2223,N_2310);
nand U2541 (N_2541,N_2361,N_2284);
and U2542 (N_2542,N_2294,N_2342);
xor U2543 (N_2543,N_2215,N_2288);
and U2544 (N_2544,N_2209,N_2233);
or U2545 (N_2545,N_2328,N_2370);
or U2546 (N_2546,N_2325,N_2265);
nand U2547 (N_2547,N_2330,N_2333);
xnor U2548 (N_2548,N_2315,N_2338);
and U2549 (N_2549,N_2333,N_2320);
nand U2550 (N_2550,N_2212,N_2370);
or U2551 (N_2551,N_2241,N_2328);
xor U2552 (N_2552,N_2209,N_2322);
nor U2553 (N_2553,N_2389,N_2321);
and U2554 (N_2554,N_2339,N_2272);
and U2555 (N_2555,N_2309,N_2258);
nand U2556 (N_2556,N_2338,N_2357);
or U2557 (N_2557,N_2370,N_2263);
or U2558 (N_2558,N_2349,N_2252);
nand U2559 (N_2559,N_2338,N_2256);
nor U2560 (N_2560,N_2219,N_2215);
and U2561 (N_2561,N_2286,N_2337);
or U2562 (N_2562,N_2205,N_2272);
nor U2563 (N_2563,N_2390,N_2284);
nor U2564 (N_2564,N_2266,N_2275);
xnor U2565 (N_2565,N_2386,N_2282);
xor U2566 (N_2566,N_2289,N_2357);
or U2567 (N_2567,N_2229,N_2368);
or U2568 (N_2568,N_2380,N_2288);
nor U2569 (N_2569,N_2374,N_2220);
nor U2570 (N_2570,N_2212,N_2272);
and U2571 (N_2571,N_2241,N_2284);
or U2572 (N_2572,N_2224,N_2260);
nor U2573 (N_2573,N_2399,N_2296);
nor U2574 (N_2574,N_2293,N_2233);
nand U2575 (N_2575,N_2235,N_2241);
nand U2576 (N_2576,N_2336,N_2372);
nand U2577 (N_2577,N_2313,N_2286);
and U2578 (N_2578,N_2378,N_2317);
xnor U2579 (N_2579,N_2236,N_2233);
and U2580 (N_2580,N_2349,N_2391);
and U2581 (N_2581,N_2232,N_2243);
xnor U2582 (N_2582,N_2297,N_2342);
and U2583 (N_2583,N_2224,N_2303);
nand U2584 (N_2584,N_2265,N_2260);
xor U2585 (N_2585,N_2240,N_2284);
nand U2586 (N_2586,N_2223,N_2202);
nand U2587 (N_2587,N_2334,N_2276);
and U2588 (N_2588,N_2272,N_2354);
or U2589 (N_2589,N_2242,N_2356);
or U2590 (N_2590,N_2284,N_2358);
nor U2591 (N_2591,N_2279,N_2332);
xnor U2592 (N_2592,N_2303,N_2321);
xnor U2593 (N_2593,N_2383,N_2367);
or U2594 (N_2594,N_2266,N_2353);
or U2595 (N_2595,N_2311,N_2356);
and U2596 (N_2596,N_2299,N_2319);
nand U2597 (N_2597,N_2227,N_2386);
nor U2598 (N_2598,N_2269,N_2349);
nand U2599 (N_2599,N_2330,N_2368);
nor U2600 (N_2600,N_2429,N_2436);
or U2601 (N_2601,N_2533,N_2494);
nor U2602 (N_2602,N_2537,N_2517);
xor U2603 (N_2603,N_2557,N_2415);
or U2604 (N_2604,N_2541,N_2456);
nor U2605 (N_2605,N_2575,N_2571);
or U2606 (N_2606,N_2562,N_2523);
xnor U2607 (N_2607,N_2572,N_2465);
or U2608 (N_2608,N_2510,N_2447);
nor U2609 (N_2609,N_2591,N_2538);
or U2610 (N_2610,N_2569,N_2402);
or U2611 (N_2611,N_2525,N_2430);
nand U2612 (N_2612,N_2583,N_2567);
nand U2613 (N_2613,N_2428,N_2514);
and U2614 (N_2614,N_2473,N_2549);
xnor U2615 (N_2615,N_2527,N_2558);
nor U2616 (N_2616,N_2524,N_2544);
nand U2617 (N_2617,N_2552,N_2573);
nor U2618 (N_2618,N_2487,N_2400);
nand U2619 (N_2619,N_2422,N_2542);
or U2620 (N_2620,N_2505,N_2516);
nor U2621 (N_2621,N_2464,N_2521);
nand U2622 (N_2622,N_2498,N_2564);
nand U2623 (N_2623,N_2410,N_2589);
or U2624 (N_2624,N_2471,N_2502);
nand U2625 (N_2625,N_2519,N_2529);
nand U2626 (N_2626,N_2545,N_2508);
nand U2627 (N_2627,N_2509,N_2488);
or U2628 (N_2628,N_2461,N_2448);
and U2629 (N_2629,N_2458,N_2452);
and U2630 (N_2630,N_2401,N_2576);
xnor U2631 (N_2631,N_2595,N_2520);
nand U2632 (N_2632,N_2423,N_2584);
nand U2633 (N_2633,N_2561,N_2474);
nand U2634 (N_2634,N_2582,N_2518);
and U2635 (N_2635,N_2421,N_2592);
and U2636 (N_2636,N_2563,N_2426);
and U2637 (N_2637,N_2486,N_2424);
and U2638 (N_2638,N_2570,N_2543);
nor U2639 (N_2639,N_2556,N_2450);
or U2640 (N_2640,N_2483,N_2462);
xnor U2641 (N_2641,N_2500,N_2443);
nor U2642 (N_2642,N_2417,N_2440);
nor U2643 (N_2643,N_2586,N_2504);
xor U2644 (N_2644,N_2412,N_2414);
nor U2645 (N_2645,N_2548,N_2416);
nor U2646 (N_2646,N_2501,N_2490);
nand U2647 (N_2647,N_2511,N_2475);
nor U2648 (N_2648,N_2580,N_2434);
nand U2649 (N_2649,N_2431,N_2405);
nand U2650 (N_2650,N_2407,N_2420);
or U2651 (N_2651,N_2531,N_2437);
nor U2652 (N_2652,N_2418,N_2492);
nand U2653 (N_2653,N_2596,N_2528);
nand U2654 (N_2654,N_2587,N_2491);
or U2655 (N_2655,N_2459,N_2585);
nand U2656 (N_2656,N_2535,N_2594);
nor U2657 (N_2657,N_2435,N_2427);
or U2658 (N_2658,N_2481,N_2451);
nor U2659 (N_2659,N_2534,N_2578);
nand U2660 (N_2660,N_2539,N_2574);
nand U2661 (N_2661,N_2593,N_2477);
nor U2662 (N_2662,N_2526,N_2468);
or U2663 (N_2663,N_2455,N_2588);
xnor U2664 (N_2664,N_2536,N_2597);
nor U2665 (N_2665,N_2467,N_2512);
or U2666 (N_2666,N_2559,N_2479);
or U2667 (N_2667,N_2485,N_2555);
and U2668 (N_2668,N_2463,N_2425);
xor U2669 (N_2669,N_2449,N_2470);
nor U2670 (N_2670,N_2466,N_2581);
nor U2671 (N_2671,N_2506,N_2547);
nor U2672 (N_2672,N_2441,N_2579);
nor U2673 (N_2673,N_2553,N_2546);
and U2674 (N_2674,N_2411,N_2499);
or U2675 (N_2675,N_2550,N_2496);
nor U2676 (N_2676,N_2476,N_2522);
and U2677 (N_2677,N_2442,N_2454);
nand U2678 (N_2678,N_2484,N_2445);
or U2679 (N_2679,N_2403,N_2540);
nor U2680 (N_2680,N_2554,N_2446);
nor U2681 (N_2681,N_2408,N_2513);
or U2682 (N_2682,N_2404,N_2413);
xnor U2683 (N_2683,N_2453,N_2472);
and U2684 (N_2684,N_2590,N_2460);
xor U2685 (N_2685,N_2469,N_2530);
nor U2686 (N_2686,N_2503,N_2568);
or U2687 (N_2687,N_2507,N_2439);
or U2688 (N_2688,N_2532,N_2478);
xnor U2689 (N_2689,N_2497,N_2433);
and U2690 (N_2690,N_2457,N_2566);
or U2691 (N_2691,N_2599,N_2565);
nand U2692 (N_2692,N_2438,N_2493);
and U2693 (N_2693,N_2495,N_2598);
and U2694 (N_2694,N_2515,N_2419);
nand U2695 (N_2695,N_2432,N_2489);
xnor U2696 (N_2696,N_2444,N_2577);
xor U2697 (N_2697,N_2480,N_2551);
nand U2698 (N_2698,N_2409,N_2482);
nor U2699 (N_2699,N_2406,N_2560);
or U2700 (N_2700,N_2570,N_2512);
nand U2701 (N_2701,N_2421,N_2490);
or U2702 (N_2702,N_2542,N_2553);
xor U2703 (N_2703,N_2515,N_2403);
nor U2704 (N_2704,N_2539,N_2426);
or U2705 (N_2705,N_2554,N_2400);
nand U2706 (N_2706,N_2569,N_2553);
or U2707 (N_2707,N_2568,N_2536);
nand U2708 (N_2708,N_2482,N_2425);
and U2709 (N_2709,N_2537,N_2556);
xor U2710 (N_2710,N_2506,N_2593);
and U2711 (N_2711,N_2473,N_2467);
and U2712 (N_2712,N_2522,N_2513);
xor U2713 (N_2713,N_2528,N_2513);
or U2714 (N_2714,N_2425,N_2587);
nand U2715 (N_2715,N_2568,N_2446);
or U2716 (N_2716,N_2414,N_2430);
nor U2717 (N_2717,N_2446,N_2459);
nor U2718 (N_2718,N_2438,N_2495);
or U2719 (N_2719,N_2528,N_2471);
and U2720 (N_2720,N_2413,N_2541);
nor U2721 (N_2721,N_2599,N_2441);
or U2722 (N_2722,N_2564,N_2567);
nand U2723 (N_2723,N_2512,N_2559);
nor U2724 (N_2724,N_2458,N_2422);
or U2725 (N_2725,N_2541,N_2468);
xor U2726 (N_2726,N_2530,N_2436);
nand U2727 (N_2727,N_2446,N_2519);
xnor U2728 (N_2728,N_2576,N_2540);
nor U2729 (N_2729,N_2400,N_2419);
xor U2730 (N_2730,N_2587,N_2570);
nand U2731 (N_2731,N_2585,N_2417);
nor U2732 (N_2732,N_2591,N_2405);
xnor U2733 (N_2733,N_2493,N_2504);
xor U2734 (N_2734,N_2562,N_2544);
xor U2735 (N_2735,N_2481,N_2441);
xnor U2736 (N_2736,N_2437,N_2489);
nor U2737 (N_2737,N_2583,N_2536);
xnor U2738 (N_2738,N_2517,N_2555);
xnor U2739 (N_2739,N_2570,N_2439);
and U2740 (N_2740,N_2520,N_2489);
xor U2741 (N_2741,N_2521,N_2555);
nor U2742 (N_2742,N_2449,N_2576);
and U2743 (N_2743,N_2565,N_2430);
and U2744 (N_2744,N_2464,N_2448);
nand U2745 (N_2745,N_2558,N_2569);
nor U2746 (N_2746,N_2526,N_2469);
and U2747 (N_2747,N_2544,N_2512);
and U2748 (N_2748,N_2464,N_2598);
and U2749 (N_2749,N_2545,N_2450);
nand U2750 (N_2750,N_2525,N_2436);
and U2751 (N_2751,N_2558,N_2409);
or U2752 (N_2752,N_2527,N_2579);
xor U2753 (N_2753,N_2533,N_2596);
nand U2754 (N_2754,N_2407,N_2408);
xnor U2755 (N_2755,N_2587,N_2486);
or U2756 (N_2756,N_2438,N_2401);
nor U2757 (N_2757,N_2525,N_2553);
nand U2758 (N_2758,N_2482,N_2550);
nand U2759 (N_2759,N_2429,N_2516);
and U2760 (N_2760,N_2570,N_2552);
and U2761 (N_2761,N_2443,N_2546);
and U2762 (N_2762,N_2557,N_2450);
nand U2763 (N_2763,N_2575,N_2424);
and U2764 (N_2764,N_2524,N_2590);
and U2765 (N_2765,N_2440,N_2549);
xnor U2766 (N_2766,N_2599,N_2449);
nor U2767 (N_2767,N_2572,N_2437);
nor U2768 (N_2768,N_2492,N_2564);
or U2769 (N_2769,N_2565,N_2438);
nor U2770 (N_2770,N_2468,N_2465);
xor U2771 (N_2771,N_2453,N_2540);
nor U2772 (N_2772,N_2443,N_2424);
or U2773 (N_2773,N_2497,N_2535);
nand U2774 (N_2774,N_2571,N_2471);
or U2775 (N_2775,N_2572,N_2489);
or U2776 (N_2776,N_2521,N_2434);
nor U2777 (N_2777,N_2475,N_2471);
xor U2778 (N_2778,N_2484,N_2498);
nand U2779 (N_2779,N_2462,N_2402);
nand U2780 (N_2780,N_2585,N_2496);
nand U2781 (N_2781,N_2565,N_2592);
or U2782 (N_2782,N_2569,N_2408);
or U2783 (N_2783,N_2532,N_2589);
xnor U2784 (N_2784,N_2563,N_2412);
and U2785 (N_2785,N_2453,N_2455);
nor U2786 (N_2786,N_2401,N_2449);
and U2787 (N_2787,N_2420,N_2546);
nand U2788 (N_2788,N_2528,N_2544);
xor U2789 (N_2789,N_2442,N_2586);
or U2790 (N_2790,N_2438,N_2507);
or U2791 (N_2791,N_2497,N_2530);
and U2792 (N_2792,N_2451,N_2411);
and U2793 (N_2793,N_2465,N_2452);
nand U2794 (N_2794,N_2425,N_2461);
nor U2795 (N_2795,N_2589,N_2466);
xnor U2796 (N_2796,N_2417,N_2403);
nand U2797 (N_2797,N_2429,N_2487);
nand U2798 (N_2798,N_2550,N_2522);
nor U2799 (N_2799,N_2430,N_2453);
nand U2800 (N_2800,N_2687,N_2698);
nand U2801 (N_2801,N_2702,N_2738);
and U2802 (N_2802,N_2724,N_2737);
or U2803 (N_2803,N_2636,N_2790);
nand U2804 (N_2804,N_2797,N_2762);
nand U2805 (N_2805,N_2719,N_2717);
or U2806 (N_2806,N_2784,N_2773);
and U2807 (N_2807,N_2639,N_2642);
or U2808 (N_2808,N_2750,N_2619);
or U2809 (N_2809,N_2769,N_2714);
nand U2810 (N_2810,N_2761,N_2666);
and U2811 (N_2811,N_2691,N_2779);
xor U2812 (N_2812,N_2701,N_2785);
and U2813 (N_2813,N_2766,N_2681);
or U2814 (N_2814,N_2771,N_2754);
and U2815 (N_2815,N_2699,N_2692);
nand U2816 (N_2816,N_2782,N_2614);
or U2817 (N_2817,N_2621,N_2679);
nand U2818 (N_2818,N_2652,N_2690);
xor U2819 (N_2819,N_2677,N_2630);
nor U2820 (N_2820,N_2758,N_2631);
or U2821 (N_2821,N_2693,N_2694);
nand U2822 (N_2822,N_2615,N_2608);
nand U2823 (N_2823,N_2676,N_2674);
nand U2824 (N_2824,N_2658,N_2747);
or U2825 (N_2825,N_2603,N_2613);
xor U2826 (N_2826,N_2728,N_2726);
and U2827 (N_2827,N_2796,N_2755);
nor U2828 (N_2828,N_2672,N_2640);
and U2829 (N_2829,N_2633,N_2680);
nand U2830 (N_2830,N_2638,N_2629);
nand U2831 (N_2831,N_2705,N_2723);
or U2832 (N_2832,N_2742,N_2753);
nor U2833 (N_2833,N_2739,N_2684);
xor U2834 (N_2834,N_2734,N_2641);
xnor U2835 (N_2835,N_2767,N_2781);
nor U2836 (N_2836,N_2668,N_2743);
and U2837 (N_2837,N_2645,N_2703);
nand U2838 (N_2838,N_2776,N_2665);
xnor U2839 (N_2839,N_2664,N_2775);
or U2840 (N_2840,N_2626,N_2602);
nand U2841 (N_2841,N_2685,N_2605);
nor U2842 (N_2842,N_2735,N_2765);
xor U2843 (N_2843,N_2760,N_2682);
or U2844 (N_2844,N_2659,N_2733);
nor U2845 (N_2845,N_2601,N_2740);
nand U2846 (N_2846,N_2662,N_2770);
or U2847 (N_2847,N_2721,N_2774);
nand U2848 (N_2848,N_2625,N_2610);
nand U2849 (N_2849,N_2763,N_2695);
nand U2850 (N_2850,N_2706,N_2612);
nand U2851 (N_2851,N_2731,N_2669);
or U2852 (N_2852,N_2741,N_2634);
and U2853 (N_2853,N_2711,N_2748);
and U2854 (N_2854,N_2757,N_2647);
nand U2855 (N_2855,N_2736,N_2718);
nand U2856 (N_2856,N_2607,N_2795);
or U2857 (N_2857,N_2772,N_2678);
nor U2858 (N_2858,N_2788,N_2725);
and U2859 (N_2859,N_2646,N_2604);
xor U2860 (N_2860,N_2793,N_2632);
nand U2861 (N_2861,N_2786,N_2732);
and U2862 (N_2862,N_2622,N_2611);
or U2863 (N_2863,N_2712,N_2704);
nand U2864 (N_2864,N_2789,N_2657);
or U2865 (N_2865,N_2609,N_2783);
nor U2866 (N_2866,N_2799,N_2722);
xor U2867 (N_2867,N_2643,N_2756);
and U2868 (N_2868,N_2606,N_2720);
xnor U2869 (N_2869,N_2600,N_2655);
nand U2870 (N_2870,N_2661,N_2745);
or U2871 (N_2871,N_2656,N_2710);
nand U2872 (N_2872,N_2649,N_2637);
nand U2873 (N_2873,N_2617,N_2648);
nor U2874 (N_2874,N_2667,N_2751);
xor U2875 (N_2875,N_2675,N_2709);
xor U2876 (N_2876,N_2729,N_2764);
nor U2877 (N_2877,N_2791,N_2628);
and U2878 (N_2878,N_2616,N_2794);
and U2879 (N_2879,N_2651,N_2623);
nand U2880 (N_2880,N_2696,N_2798);
xnor U2881 (N_2881,N_2749,N_2780);
nor U2882 (N_2882,N_2620,N_2683);
or U2883 (N_2883,N_2730,N_2746);
nand U2884 (N_2884,N_2644,N_2624);
and U2885 (N_2885,N_2654,N_2778);
nor U2886 (N_2886,N_2635,N_2689);
xor U2887 (N_2887,N_2686,N_2663);
and U2888 (N_2888,N_2708,N_2697);
nand U2889 (N_2889,N_2752,N_2768);
and U2890 (N_2890,N_2700,N_2792);
and U2891 (N_2891,N_2713,N_2777);
or U2892 (N_2892,N_2707,N_2671);
xnor U2893 (N_2893,N_2759,N_2653);
nor U2894 (N_2894,N_2744,N_2618);
or U2895 (N_2895,N_2727,N_2715);
or U2896 (N_2896,N_2650,N_2670);
and U2897 (N_2897,N_2673,N_2716);
nor U2898 (N_2898,N_2688,N_2627);
nor U2899 (N_2899,N_2787,N_2660);
nand U2900 (N_2900,N_2720,N_2746);
nor U2901 (N_2901,N_2799,N_2771);
nor U2902 (N_2902,N_2753,N_2731);
nand U2903 (N_2903,N_2602,N_2778);
and U2904 (N_2904,N_2766,N_2628);
xnor U2905 (N_2905,N_2770,N_2717);
and U2906 (N_2906,N_2646,N_2750);
and U2907 (N_2907,N_2620,N_2682);
or U2908 (N_2908,N_2794,N_2776);
xnor U2909 (N_2909,N_2727,N_2679);
nand U2910 (N_2910,N_2602,N_2677);
nand U2911 (N_2911,N_2629,N_2678);
and U2912 (N_2912,N_2626,N_2662);
and U2913 (N_2913,N_2798,N_2786);
or U2914 (N_2914,N_2614,N_2754);
nand U2915 (N_2915,N_2670,N_2783);
and U2916 (N_2916,N_2659,N_2654);
xnor U2917 (N_2917,N_2793,N_2716);
xnor U2918 (N_2918,N_2675,N_2627);
nand U2919 (N_2919,N_2691,N_2678);
nor U2920 (N_2920,N_2756,N_2744);
nand U2921 (N_2921,N_2639,N_2777);
and U2922 (N_2922,N_2622,N_2732);
nand U2923 (N_2923,N_2779,N_2753);
nor U2924 (N_2924,N_2644,N_2623);
nor U2925 (N_2925,N_2600,N_2695);
or U2926 (N_2926,N_2711,N_2799);
or U2927 (N_2927,N_2672,N_2705);
nand U2928 (N_2928,N_2738,N_2648);
nor U2929 (N_2929,N_2799,N_2682);
nand U2930 (N_2930,N_2794,N_2618);
nand U2931 (N_2931,N_2752,N_2702);
or U2932 (N_2932,N_2680,N_2671);
or U2933 (N_2933,N_2664,N_2722);
xor U2934 (N_2934,N_2742,N_2760);
xnor U2935 (N_2935,N_2702,N_2709);
and U2936 (N_2936,N_2678,N_2706);
nand U2937 (N_2937,N_2777,N_2780);
and U2938 (N_2938,N_2731,N_2796);
nand U2939 (N_2939,N_2619,N_2675);
xnor U2940 (N_2940,N_2755,N_2623);
and U2941 (N_2941,N_2607,N_2606);
or U2942 (N_2942,N_2721,N_2751);
or U2943 (N_2943,N_2666,N_2608);
nand U2944 (N_2944,N_2752,N_2732);
nor U2945 (N_2945,N_2605,N_2759);
nor U2946 (N_2946,N_2776,N_2671);
xnor U2947 (N_2947,N_2670,N_2736);
xor U2948 (N_2948,N_2615,N_2628);
or U2949 (N_2949,N_2767,N_2779);
xnor U2950 (N_2950,N_2706,N_2679);
xor U2951 (N_2951,N_2691,N_2704);
xnor U2952 (N_2952,N_2756,N_2629);
nor U2953 (N_2953,N_2697,N_2636);
and U2954 (N_2954,N_2709,N_2794);
nor U2955 (N_2955,N_2654,N_2725);
nor U2956 (N_2956,N_2604,N_2721);
nand U2957 (N_2957,N_2601,N_2671);
and U2958 (N_2958,N_2760,N_2671);
nand U2959 (N_2959,N_2791,N_2773);
nand U2960 (N_2960,N_2720,N_2738);
nor U2961 (N_2961,N_2602,N_2768);
nor U2962 (N_2962,N_2771,N_2770);
xor U2963 (N_2963,N_2778,N_2749);
and U2964 (N_2964,N_2656,N_2780);
xnor U2965 (N_2965,N_2767,N_2741);
nand U2966 (N_2966,N_2630,N_2627);
or U2967 (N_2967,N_2632,N_2785);
nor U2968 (N_2968,N_2696,N_2719);
xor U2969 (N_2969,N_2701,N_2673);
nand U2970 (N_2970,N_2763,N_2732);
nor U2971 (N_2971,N_2742,N_2786);
xor U2972 (N_2972,N_2787,N_2749);
nor U2973 (N_2973,N_2607,N_2654);
nand U2974 (N_2974,N_2700,N_2791);
nor U2975 (N_2975,N_2624,N_2680);
nand U2976 (N_2976,N_2624,N_2616);
nor U2977 (N_2977,N_2722,N_2651);
nor U2978 (N_2978,N_2653,N_2627);
or U2979 (N_2979,N_2609,N_2626);
nand U2980 (N_2980,N_2727,N_2637);
nand U2981 (N_2981,N_2710,N_2644);
xor U2982 (N_2982,N_2730,N_2631);
xor U2983 (N_2983,N_2652,N_2645);
xnor U2984 (N_2984,N_2763,N_2793);
and U2985 (N_2985,N_2756,N_2747);
xor U2986 (N_2986,N_2705,N_2775);
nor U2987 (N_2987,N_2760,N_2647);
xnor U2988 (N_2988,N_2742,N_2765);
or U2989 (N_2989,N_2772,N_2713);
or U2990 (N_2990,N_2631,N_2609);
xor U2991 (N_2991,N_2676,N_2728);
nand U2992 (N_2992,N_2781,N_2716);
nor U2993 (N_2993,N_2646,N_2695);
nor U2994 (N_2994,N_2610,N_2784);
and U2995 (N_2995,N_2636,N_2696);
nand U2996 (N_2996,N_2665,N_2761);
or U2997 (N_2997,N_2715,N_2713);
xor U2998 (N_2998,N_2754,N_2767);
or U2999 (N_2999,N_2671,N_2752);
or UO_0 (O_0,N_2994,N_2845);
xnor UO_1 (O_1,N_2958,N_2875);
and UO_2 (O_2,N_2962,N_2915);
xnor UO_3 (O_3,N_2841,N_2967);
nand UO_4 (O_4,N_2897,N_2810);
xor UO_5 (O_5,N_2891,N_2895);
or UO_6 (O_6,N_2951,N_2830);
or UO_7 (O_7,N_2862,N_2870);
xor UO_8 (O_8,N_2995,N_2846);
nor UO_9 (O_9,N_2826,N_2977);
nand UO_10 (O_10,N_2914,N_2939);
and UO_11 (O_11,N_2964,N_2824);
nor UO_12 (O_12,N_2868,N_2910);
and UO_13 (O_13,N_2924,N_2865);
nor UO_14 (O_14,N_2950,N_2877);
nand UO_15 (O_15,N_2942,N_2815);
or UO_16 (O_16,N_2975,N_2816);
and UO_17 (O_17,N_2954,N_2884);
nand UO_18 (O_18,N_2963,N_2850);
and UO_19 (O_19,N_2907,N_2869);
nor UO_20 (O_20,N_2825,N_2874);
or UO_21 (O_21,N_2828,N_2844);
and UO_22 (O_22,N_2834,N_2819);
or UO_23 (O_23,N_2934,N_2996);
nand UO_24 (O_24,N_2970,N_2808);
or UO_25 (O_25,N_2945,N_2998);
xor UO_26 (O_26,N_2925,N_2827);
nor UO_27 (O_27,N_2873,N_2888);
and UO_28 (O_28,N_2823,N_2820);
or UO_29 (O_29,N_2978,N_2922);
xor UO_30 (O_30,N_2836,N_2804);
xnor UO_31 (O_31,N_2903,N_2800);
nor UO_32 (O_32,N_2885,N_2920);
and UO_33 (O_33,N_2984,N_2807);
nand UO_34 (O_34,N_2878,N_2851);
or UO_35 (O_35,N_2979,N_2968);
xnor UO_36 (O_36,N_2981,N_2902);
and UO_37 (O_37,N_2938,N_2918);
or UO_38 (O_38,N_2840,N_2940);
or UO_39 (O_39,N_2943,N_2831);
nand UO_40 (O_40,N_2953,N_2930);
nor UO_41 (O_41,N_2947,N_2848);
or UO_42 (O_42,N_2933,N_2919);
nand UO_43 (O_43,N_2833,N_2906);
or UO_44 (O_44,N_2813,N_2913);
nor UO_45 (O_45,N_2852,N_2936);
and UO_46 (O_46,N_2961,N_2932);
or UO_47 (O_47,N_2960,N_2842);
nand UO_48 (O_48,N_2946,N_2849);
and UO_49 (O_49,N_2832,N_2837);
and UO_50 (O_50,N_2853,N_2973);
and UO_51 (O_51,N_2992,N_2811);
or UO_52 (O_52,N_2887,N_2916);
xnor UO_53 (O_53,N_2969,N_2863);
and UO_54 (O_54,N_2821,N_2904);
nand UO_55 (O_55,N_2883,N_2856);
and UO_56 (O_56,N_2941,N_2948);
xor UO_57 (O_57,N_2864,N_2923);
nor UO_58 (O_58,N_2829,N_2989);
nand UO_59 (O_59,N_2892,N_2876);
nor UO_60 (O_60,N_2917,N_2806);
and UO_61 (O_61,N_2928,N_2986);
nand UO_62 (O_62,N_2817,N_2982);
and UO_63 (O_63,N_2944,N_2872);
xnor UO_64 (O_64,N_2926,N_2909);
nor UO_65 (O_65,N_2857,N_2854);
or UO_66 (O_66,N_2937,N_2931);
and UO_67 (O_67,N_2974,N_2991);
nor UO_68 (O_68,N_2838,N_2809);
or UO_69 (O_69,N_2812,N_2858);
or UO_70 (O_70,N_2900,N_2980);
or UO_71 (O_71,N_2955,N_2965);
xnor UO_72 (O_72,N_2921,N_2957);
and UO_73 (O_73,N_2966,N_2929);
and UO_74 (O_74,N_2999,N_2855);
and UO_75 (O_75,N_2990,N_2949);
nand UO_76 (O_76,N_2976,N_2893);
nor UO_77 (O_77,N_2843,N_2866);
or UO_78 (O_78,N_2898,N_2890);
nor UO_79 (O_79,N_2882,N_2988);
nand UO_80 (O_80,N_2905,N_2801);
xnor UO_81 (O_81,N_2959,N_2879);
or UO_82 (O_82,N_2952,N_2839);
xnor UO_83 (O_83,N_2859,N_2886);
xor UO_84 (O_84,N_2985,N_2894);
and UO_85 (O_85,N_2871,N_2803);
xnor UO_86 (O_86,N_2867,N_2880);
xor UO_87 (O_87,N_2896,N_2901);
and UO_88 (O_88,N_2908,N_2805);
or UO_89 (O_89,N_2818,N_2912);
xnor UO_90 (O_90,N_2972,N_2814);
xnor UO_91 (O_91,N_2935,N_2860);
xor UO_92 (O_92,N_2889,N_2802);
nand UO_93 (O_93,N_2956,N_2911);
xor UO_94 (O_94,N_2993,N_2997);
or UO_95 (O_95,N_2881,N_2861);
and UO_96 (O_96,N_2847,N_2835);
nor UO_97 (O_97,N_2971,N_2983);
xor UO_98 (O_98,N_2822,N_2927);
nor UO_99 (O_99,N_2987,N_2899);
xnor UO_100 (O_100,N_2836,N_2805);
and UO_101 (O_101,N_2879,N_2907);
nand UO_102 (O_102,N_2984,N_2863);
or UO_103 (O_103,N_2831,N_2810);
or UO_104 (O_104,N_2957,N_2845);
nor UO_105 (O_105,N_2875,N_2943);
and UO_106 (O_106,N_2854,N_2894);
or UO_107 (O_107,N_2911,N_2870);
and UO_108 (O_108,N_2887,N_2865);
or UO_109 (O_109,N_2845,N_2930);
xor UO_110 (O_110,N_2885,N_2930);
xor UO_111 (O_111,N_2868,N_2934);
and UO_112 (O_112,N_2884,N_2832);
or UO_113 (O_113,N_2902,N_2827);
nand UO_114 (O_114,N_2997,N_2925);
and UO_115 (O_115,N_2845,N_2879);
or UO_116 (O_116,N_2988,N_2809);
or UO_117 (O_117,N_2941,N_2986);
or UO_118 (O_118,N_2926,N_2809);
and UO_119 (O_119,N_2895,N_2899);
or UO_120 (O_120,N_2870,N_2968);
nand UO_121 (O_121,N_2957,N_2998);
and UO_122 (O_122,N_2836,N_2968);
nand UO_123 (O_123,N_2960,N_2835);
or UO_124 (O_124,N_2876,N_2973);
or UO_125 (O_125,N_2850,N_2925);
and UO_126 (O_126,N_2810,N_2989);
nand UO_127 (O_127,N_2920,N_2865);
and UO_128 (O_128,N_2848,N_2879);
xor UO_129 (O_129,N_2977,N_2834);
and UO_130 (O_130,N_2824,N_2872);
and UO_131 (O_131,N_2883,N_2882);
or UO_132 (O_132,N_2950,N_2857);
and UO_133 (O_133,N_2986,N_2897);
or UO_134 (O_134,N_2803,N_2808);
and UO_135 (O_135,N_2847,N_2808);
nand UO_136 (O_136,N_2993,N_2883);
nor UO_137 (O_137,N_2920,N_2968);
nand UO_138 (O_138,N_2980,N_2992);
and UO_139 (O_139,N_2960,N_2834);
xor UO_140 (O_140,N_2855,N_2941);
or UO_141 (O_141,N_2877,N_2868);
nand UO_142 (O_142,N_2812,N_2801);
xnor UO_143 (O_143,N_2900,N_2896);
xor UO_144 (O_144,N_2935,N_2821);
or UO_145 (O_145,N_2872,N_2947);
xnor UO_146 (O_146,N_2927,N_2863);
nand UO_147 (O_147,N_2853,N_2934);
xor UO_148 (O_148,N_2821,N_2846);
and UO_149 (O_149,N_2817,N_2865);
or UO_150 (O_150,N_2978,N_2892);
nor UO_151 (O_151,N_2999,N_2973);
and UO_152 (O_152,N_2873,N_2927);
and UO_153 (O_153,N_2814,N_2935);
or UO_154 (O_154,N_2901,N_2815);
xnor UO_155 (O_155,N_2823,N_2905);
xor UO_156 (O_156,N_2920,N_2906);
nand UO_157 (O_157,N_2945,N_2810);
nor UO_158 (O_158,N_2933,N_2977);
nor UO_159 (O_159,N_2874,N_2815);
and UO_160 (O_160,N_2987,N_2970);
and UO_161 (O_161,N_2876,N_2912);
and UO_162 (O_162,N_2918,N_2946);
or UO_163 (O_163,N_2948,N_2830);
or UO_164 (O_164,N_2880,N_2907);
nand UO_165 (O_165,N_2865,N_2906);
or UO_166 (O_166,N_2979,N_2810);
nor UO_167 (O_167,N_2820,N_2993);
nand UO_168 (O_168,N_2921,N_2886);
xnor UO_169 (O_169,N_2894,N_2963);
and UO_170 (O_170,N_2972,N_2950);
and UO_171 (O_171,N_2923,N_2908);
or UO_172 (O_172,N_2854,N_2870);
or UO_173 (O_173,N_2963,N_2975);
nor UO_174 (O_174,N_2887,N_2816);
nand UO_175 (O_175,N_2811,N_2948);
and UO_176 (O_176,N_2928,N_2857);
and UO_177 (O_177,N_2869,N_2936);
nand UO_178 (O_178,N_2842,N_2874);
nor UO_179 (O_179,N_2861,N_2924);
nor UO_180 (O_180,N_2993,N_2877);
and UO_181 (O_181,N_2867,N_2814);
and UO_182 (O_182,N_2810,N_2876);
nand UO_183 (O_183,N_2988,N_2910);
and UO_184 (O_184,N_2840,N_2824);
nor UO_185 (O_185,N_2982,N_2894);
or UO_186 (O_186,N_2802,N_2887);
nand UO_187 (O_187,N_2852,N_2857);
and UO_188 (O_188,N_2831,N_2804);
and UO_189 (O_189,N_2856,N_2970);
or UO_190 (O_190,N_2991,N_2845);
nand UO_191 (O_191,N_2989,N_2841);
and UO_192 (O_192,N_2933,N_2962);
nand UO_193 (O_193,N_2850,N_2830);
and UO_194 (O_194,N_2839,N_2802);
xnor UO_195 (O_195,N_2869,N_2903);
nand UO_196 (O_196,N_2885,N_2816);
nor UO_197 (O_197,N_2882,N_2841);
nand UO_198 (O_198,N_2945,N_2857);
xor UO_199 (O_199,N_2905,N_2835);
or UO_200 (O_200,N_2861,N_2899);
or UO_201 (O_201,N_2879,N_2826);
or UO_202 (O_202,N_2992,N_2841);
nand UO_203 (O_203,N_2809,N_2997);
nor UO_204 (O_204,N_2860,N_2861);
and UO_205 (O_205,N_2965,N_2911);
and UO_206 (O_206,N_2895,N_2988);
or UO_207 (O_207,N_2838,N_2912);
nor UO_208 (O_208,N_2868,N_2979);
or UO_209 (O_209,N_2852,N_2886);
nand UO_210 (O_210,N_2942,N_2911);
nor UO_211 (O_211,N_2974,N_2813);
nor UO_212 (O_212,N_2989,N_2992);
nor UO_213 (O_213,N_2867,N_2912);
nor UO_214 (O_214,N_2914,N_2889);
and UO_215 (O_215,N_2820,N_2960);
nand UO_216 (O_216,N_2886,N_2913);
nand UO_217 (O_217,N_2932,N_2817);
nand UO_218 (O_218,N_2919,N_2872);
nand UO_219 (O_219,N_2952,N_2979);
nand UO_220 (O_220,N_2959,N_2955);
and UO_221 (O_221,N_2871,N_2846);
xor UO_222 (O_222,N_2981,N_2875);
xnor UO_223 (O_223,N_2835,N_2969);
and UO_224 (O_224,N_2954,N_2808);
xor UO_225 (O_225,N_2922,N_2825);
or UO_226 (O_226,N_2908,N_2994);
nor UO_227 (O_227,N_2963,N_2943);
xor UO_228 (O_228,N_2811,N_2878);
and UO_229 (O_229,N_2901,N_2957);
nor UO_230 (O_230,N_2853,N_2843);
and UO_231 (O_231,N_2858,N_2815);
or UO_232 (O_232,N_2956,N_2907);
nand UO_233 (O_233,N_2894,N_2893);
xor UO_234 (O_234,N_2994,N_2915);
and UO_235 (O_235,N_2939,N_2978);
nand UO_236 (O_236,N_2952,N_2944);
nor UO_237 (O_237,N_2812,N_2943);
nor UO_238 (O_238,N_2901,N_2979);
or UO_239 (O_239,N_2830,N_2972);
nand UO_240 (O_240,N_2939,N_2830);
nand UO_241 (O_241,N_2934,N_2846);
or UO_242 (O_242,N_2991,N_2966);
nor UO_243 (O_243,N_2970,N_2979);
or UO_244 (O_244,N_2822,N_2978);
nand UO_245 (O_245,N_2926,N_2911);
or UO_246 (O_246,N_2849,N_2835);
nand UO_247 (O_247,N_2914,N_2800);
xnor UO_248 (O_248,N_2859,N_2915);
xnor UO_249 (O_249,N_2975,N_2937);
and UO_250 (O_250,N_2801,N_2960);
and UO_251 (O_251,N_2925,N_2924);
or UO_252 (O_252,N_2928,N_2850);
nor UO_253 (O_253,N_2861,N_2874);
xnor UO_254 (O_254,N_2841,N_2892);
or UO_255 (O_255,N_2876,N_2891);
nor UO_256 (O_256,N_2968,N_2975);
nor UO_257 (O_257,N_2907,N_2813);
or UO_258 (O_258,N_2948,N_2893);
and UO_259 (O_259,N_2895,N_2966);
or UO_260 (O_260,N_2984,N_2917);
and UO_261 (O_261,N_2807,N_2800);
and UO_262 (O_262,N_2845,N_2864);
xnor UO_263 (O_263,N_2884,N_2859);
nand UO_264 (O_264,N_2817,N_2928);
nand UO_265 (O_265,N_2851,N_2805);
nor UO_266 (O_266,N_2823,N_2822);
nand UO_267 (O_267,N_2890,N_2905);
and UO_268 (O_268,N_2991,N_2828);
xor UO_269 (O_269,N_2978,N_2908);
nand UO_270 (O_270,N_2868,N_2924);
or UO_271 (O_271,N_2963,N_2988);
and UO_272 (O_272,N_2881,N_2949);
xnor UO_273 (O_273,N_2929,N_2940);
or UO_274 (O_274,N_2867,N_2958);
nor UO_275 (O_275,N_2931,N_2829);
nor UO_276 (O_276,N_2861,N_2930);
and UO_277 (O_277,N_2887,N_2983);
and UO_278 (O_278,N_2935,N_2873);
xor UO_279 (O_279,N_2864,N_2801);
nor UO_280 (O_280,N_2876,N_2803);
and UO_281 (O_281,N_2918,N_2928);
nand UO_282 (O_282,N_2892,N_2860);
xor UO_283 (O_283,N_2812,N_2892);
xnor UO_284 (O_284,N_2950,N_2934);
xnor UO_285 (O_285,N_2948,N_2997);
or UO_286 (O_286,N_2883,N_2946);
and UO_287 (O_287,N_2815,N_2882);
nor UO_288 (O_288,N_2877,N_2964);
or UO_289 (O_289,N_2972,N_2911);
nor UO_290 (O_290,N_2891,N_2945);
nor UO_291 (O_291,N_2862,N_2897);
xor UO_292 (O_292,N_2963,N_2876);
nor UO_293 (O_293,N_2819,N_2902);
xor UO_294 (O_294,N_2926,N_2831);
or UO_295 (O_295,N_2876,N_2864);
or UO_296 (O_296,N_2945,N_2958);
or UO_297 (O_297,N_2888,N_2843);
xor UO_298 (O_298,N_2800,N_2892);
and UO_299 (O_299,N_2813,N_2938);
xnor UO_300 (O_300,N_2999,N_2902);
nor UO_301 (O_301,N_2801,N_2882);
xor UO_302 (O_302,N_2904,N_2824);
nand UO_303 (O_303,N_2939,N_2840);
nand UO_304 (O_304,N_2821,N_2815);
xor UO_305 (O_305,N_2981,N_2939);
and UO_306 (O_306,N_2897,N_2865);
and UO_307 (O_307,N_2908,N_2980);
nor UO_308 (O_308,N_2817,N_2831);
and UO_309 (O_309,N_2985,N_2912);
xnor UO_310 (O_310,N_2891,N_2946);
nand UO_311 (O_311,N_2911,N_2800);
xor UO_312 (O_312,N_2841,N_2840);
or UO_313 (O_313,N_2945,N_2892);
nor UO_314 (O_314,N_2993,N_2858);
xor UO_315 (O_315,N_2939,N_2949);
nor UO_316 (O_316,N_2949,N_2807);
and UO_317 (O_317,N_2842,N_2827);
nor UO_318 (O_318,N_2865,N_2826);
nor UO_319 (O_319,N_2922,N_2812);
nand UO_320 (O_320,N_2877,N_2891);
and UO_321 (O_321,N_2998,N_2986);
xor UO_322 (O_322,N_2846,N_2884);
nor UO_323 (O_323,N_2953,N_2850);
and UO_324 (O_324,N_2909,N_2900);
nand UO_325 (O_325,N_2831,N_2954);
nor UO_326 (O_326,N_2955,N_2913);
or UO_327 (O_327,N_2928,N_2815);
nor UO_328 (O_328,N_2967,N_2919);
nor UO_329 (O_329,N_2999,N_2992);
or UO_330 (O_330,N_2818,N_2825);
and UO_331 (O_331,N_2907,N_2818);
nand UO_332 (O_332,N_2848,N_2831);
and UO_333 (O_333,N_2978,N_2868);
nand UO_334 (O_334,N_2920,N_2880);
xor UO_335 (O_335,N_2826,N_2877);
and UO_336 (O_336,N_2855,N_2862);
and UO_337 (O_337,N_2827,N_2831);
nand UO_338 (O_338,N_2966,N_2812);
nand UO_339 (O_339,N_2983,N_2822);
xor UO_340 (O_340,N_2953,N_2874);
nor UO_341 (O_341,N_2867,N_2830);
xnor UO_342 (O_342,N_2936,N_2835);
xnor UO_343 (O_343,N_2920,N_2963);
nor UO_344 (O_344,N_2811,N_2860);
or UO_345 (O_345,N_2913,N_2928);
and UO_346 (O_346,N_2865,N_2820);
nand UO_347 (O_347,N_2870,N_2882);
or UO_348 (O_348,N_2949,N_2923);
nand UO_349 (O_349,N_2974,N_2832);
nor UO_350 (O_350,N_2815,N_2862);
or UO_351 (O_351,N_2820,N_2822);
or UO_352 (O_352,N_2953,N_2875);
nand UO_353 (O_353,N_2905,N_2846);
nor UO_354 (O_354,N_2864,N_2835);
nor UO_355 (O_355,N_2967,N_2864);
nor UO_356 (O_356,N_2905,N_2925);
and UO_357 (O_357,N_2970,N_2996);
nor UO_358 (O_358,N_2944,N_2970);
nor UO_359 (O_359,N_2819,N_2899);
and UO_360 (O_360,N_2858,N_2864);
xor UO_361 (O_361,N_2830,N_2831);
xor UO_362 (O_362,N_2994,N_2858);
and UO_363 (O_363,N_2901,N_2975);
nand UO_364 (O_364,N_2921,N_2999);
and UO_365 (O_365,N_2962,N_2830);
and UO_366 (O_366,N_2954,N_2966);
or UO_367 (O_367,N_2914,N_2853);
or UO_368 (O_368,N_2820,N_2958);
or UO_369 (O_369,N_2957,N_2842);
nor UO_370 (O_370,N_2809,N_2807);
or UO_371 (O_371,N_2828,N_2903);
nor UO_372 (O_372,N_2931,N_2950);
nor UO_373 (O_373,N_2926,N_2883);
xnor UO_374 (O_374,N_2999,N_2977);
nand UO_375 (O_375,N_2892,N_2809);
nand UO_376 (O_376,N_2843,N_2814);
xnor UO_377 (O_377,N_2894,N_2859);
and UO_378 (O_378,N_2890,N_2869);
xor UO_379 (O_379,N_2837,N_2803);
and UO_380 (O_380,N_2871,N_2839);
or UO_381 (O_381,N_2952,N_2809);
or UO_382 (O_382,N_2848,N_2921);
xor UO_383 (O_383,N_2890,N_2891);
nor UO_384 (O_384,N_2926,N_2813);
xor UO_385 (O_385,N_2918,N_2844);
xor UO_386 (O_386,N_2974,N_2984);
or UO_387 (O_387,N_2906,N_2889);
nand UO_388 (O_388,N_2925,N_2921);
nor UO_389 (O_389,N_2969,N_2821);
nor UO_390 (O_390,N_2867,N_2837);
nand UO_391 (O_391,N_2933,N_2801);
nand UO_392 (O_392,N_2889,N_2921);
or UO_393 (O_393,N_2902,N_2871);
or UO_394 (O_394,N_2959,N_2915);
or UO_395 (O_395,N_2816,N_2927);
or UO_396 (O_396,N_2803,N_2991);
or UO_397 (O_397,N_2868,N_2961);
or UO_398 (O_398,N_2879,N_2888);
nand UO_399 (O_399,N_2979,N_2981);
and UO_400 (O_400,N_2874,N_2812);
and UO_401 (O_401,N_2984,N_2940);
xnor UO_402 (O_402,N_2910,N_2926);
or UO_403 (O_403,N_2908,N_2888);
and UO_404 (O_404,N_2905,N_2959);
and UO_405 (O_405,N_2871,N_2924);
nor UO_406 (O_406,N_2971,N_2961);
and UO_407 (O_407,N_2844,N_2943);
or UO_408 (O_408,N_2855,N_2910);
or UO_409 (O_409,N_2866,N_2990);
or UO_410 (O_410,N_2954,N_2969);
nand UO_411 (O_411,N_2852,N_2889);
or UO_412 (O_412,N_2888,N_2878);
nand UO_413 (O_413,N_2992,N_2915);
or UO_414 (O_414,N_2879,N_2916);
and UO_415 (O_415,N_2868,N_2822);
or UO_416 (O_416,N_2838,N_2908);
xnor UO_417 (O_417,N_2853,N_2881);
nor UO_418 (O_418,N_2863,N_2814);
xnor UO_419 (O_419,N_2903,N_2819);
nand UO_420 (O_420,N_2904,N_2975);
and UO_421 (O_421,N_2933,N_2972);
xnor UO_422 (O_422,N_2869,N_2889);
nor UO_423 (O_423,N_2936,N_2886);
or UO_424 (O_424,N_2914,N_2979);
and UO_425 (O_425,N_2932,N_2848);
nor UO_426 (O_426,N_2836,N_2924);
and UO_427 (O_427,N_2948,N_2892);
xor UO_428 (O_428,N_2867,N_2882);
or UO_429 (O_429,N_2892,N_2923);
nor UO_430 (O_430,N_2895,N_2856);
and UO_431 (O_431,N_2917,N_2961);
nand UO_432 (O_432,N_2921,N_2894);
xnor UO_433 (O_433,N_2812,N_2945);
or UO_434 (O_434,N_2898,N_2924);
nor UO_435 (O_435,N_2848,N_2880);
nand UO_436 (O_436,N_2996,N_2874);
nor UO_437 (O_437,N_2979,N_2938);
xor UO_438 (O_438,N_2898,N_2910);
nor UO_439 (O_439,N_2860,N_2965);
and UO_440 (O_440,N_2852,N_2986);
nor UO_441 (O_441,N_2959,N_2916);
nand UO_442 (O_442,N_2812,N_2908);
nand UO_443 (O_443,N_2907,N_2923);
and UO_444 (O_444,N_2959,N_2807);
nor UO_445 (O_445,N_2942,N_2848);
and UO_446 (O_446,N_2900,N_2926);
nor UO_447 (O_447,N_2818,N_2893);
or UO_448 (O_448,N_2899,N_2818);
or UO_449 (O_449,N_2924,N_2845);
and UO_450 (O_450,N_2956,N_2961);
and UO_451 (O_451,N_2988,N_2972);
or UO_452 (O_452,N_2810,N_2956);
or UO_453 (O_453,N_2993,N_2843);
or UO_454 (O_454,N_2973,N_2953);
xnor UO_455 (O_455,N_2951,N_2923);
nand UO_456 (O_456,N_2996,N_2929);
and UO_457 (O_457,N_2803,N_2954);
xor UO_458 (O_458,N_2924,N_2844);
and UO_459 (O_459,N_2999,N_2978);
xnor UO_460 (O_460,N_2979,N_2860);
or UO_461 (O_461,N_2947,N_2908);
xor UO_462 (O_462,N_2980,N_2948);
or UO_463 (O_463,N_2986,N_2830);
nand UO_464 (O_464,N_2861,N_2940);
nand UO_465 (O_465,N_2889,N_2848);
nand UO_466 (O_466,N_2900,N_2947);
nand UO_467 (O_467,N_2987,N_2998);
xor UO_468 (O_468,N_2940,N_2954);
or UO_469 (O_469,N_2818,N_2836);
nor UO_470 (O_470,N_2968,N_2973);
xor UO_471 (O_471,N_2866,N_2996);
or UO_472 (O_472,N_2959,N_2921);
nand UO_473 (O_473,N_2821,N_2920);
nor UO_474 (O_474,N_2871,N_2919);
or UO_475 (O_475,N_2829,N_2978);
nand UO_476 (O_476,N_2815,N_2905);
nand UO_477 (O_477,N_2885,N_2884);
or UO_478 (O_478,N_2914,N_2927);
or UO_479 (O_479,N_2878,N_2910);
and UO_480 (O_480,N_2958,N_2949);
xor UO_481 (O_481,N_2959,N_2848);
nor UO_482 (O_482,N_2953,N_2984);
and UO_483 (O_483,N_2939,N_2842);
or UO_484 (O_484,N_2975,N_2995);
nand UO_485 (O_485,N_2943,N_2822);
nor UO_486 (O_486,N_2942,N_2931);
or UO_487 (O_487,N_2976,N_2897);
and UO_488 (O_488,N_2811,N_2854);
or UO_489 (O_489,N_2870,N_2804);
xor UO_490 (O_490,N_2937,N_2950);
nand UO_491 (O_491,N_2919,N_2962);
or UO_492 (O_492,N_2998,N_2920);
and UO_493 (O_493,N_2902,N_2941);
nor UO_494 (O_494,N_2923,N_2885);
nor UO_495 (O_495,N_2875,N_2959);
nand UO_496 (O_496,N_2971,N_2830);
and UO_497 (O_497,N_2876,N_2977);
nor UO_498 (O_498,N_2853,N_2947);
nand UO_499 (O_499,N_2955,N_2998);
endmodule