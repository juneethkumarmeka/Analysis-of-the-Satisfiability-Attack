module basic_1500_15000_2000_5_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1394,In_523);
nor U1 (N_1,In_830,In_1120);
nand U2 (N_2,In_551,In_1305);
nor U3 (N_3,In_235,In_1159);
or U4 (N_4,In_1295,In_1026);
nand U5 (N_5,In_349,In_1409);
or U6 (N_6,In_1298,In_64);
or U7 (N_7,In_1271,In_49);
or U8 (N_8,In_1307,In_1452);
or U9 (N_9,In_531,In_607);
nor U10 (N_10,In_1486,In_368);
nand U11 (N_11,In_1015,In_1468);
nand U12 (N_12,In_1333,In_653);
nor U13 (N_13,In_1377,In_930);
or U14 (N_14,In_1442,In_205);
nor U15 (N_15,In_44,In_1337);
and U16 (N_16,In_1275,In_701);
or U17 (N_17,In_1050,In_1174);
xor U18 (N_18,In_1283,In_877);
nand U19 (N_19,In_1098,In_1138);
nand U20 (N_20,In_908,In_1172);
nor U21 (N_21,In_645,In_103);
or U22 (N_22,In_1383,In_1386);
nand U23 (N_23,In_479,In_1144);
nor U24 (N_24,In_646,In_613);
nand U25 (N_25,In_612,In_1041);
nor U26 (N_26,In_730,In_710);
nor U27 (N_27,In_1462,In_27);
nor U28 (N_28,In_36,In_1148);
nand U29 (N_29,In_324,In_1330);
nor U30 (N_30,In_703,In_804);
nor U31 (N_31,In_131,In_942);
or U32 (N_32,In_670,In_808);
and U33 (N_33,In_1170,In_1140);
and U34 (N_34,In_977,In_746);
or U35 (N_35,In_11,In_1167);
and U36 (N_36,In_1200,In_1475);
and U37 (N_37,In_845,In_232);
nor U38 (N_38,In_1469,In_1079);
and U39 (N_39,In_1425,In_571);
nand U40 (N_40,In_775,In_1178);
nand U41 (N_41,In_582,In_937);
nand U42 (N_42,In_337,In_1341);
and U43 (N_43,In_1395,In_776);
nand U44 (N_44,In_1109,In_1433);
nor U45 (N_45,In_268,In_798);
and U46 (N_46,In_456,In_1422);
and U47 (N_47,In_1491,In_1097);
and U48 (N_48,In_1334,In_1368);
nand U49 (N_49,In_358,In_505);
or U50 (N_50,In_108,In_853);
and U51 (N_51,In_375,In_150);
nand U52 (N_52,In_81,In_549);
nor U53 (N_53,In_533,In_1460);
nor U54 (N_54,In_524,In_940);
nand U55 (N_55,In_1241,In_144);
nand U56 (N_56,In_239,In_511);
nor U57 (N_57,In_951,In_660);
nand U58 (N_58,In_469,In_943);
and U59 (N_59,In_1185,In_674);
nor U60 (N_60,In_1029,In_1443);
nor U61 (N_61,In_248,In_734);
or U62 (N_62,In_139,In_679);
nand U63 (N_63,In_1093,In_802);
and U64 (N_64,In_818,In_957);
nand U65 (N_65,In_480,In_859);
nand U66 (N_66,In_443,In_729);
and U67 (N_67,In_1106,In_870);
or U68 (N_68,In_1251,In_764);
nor U69 (N_69,In_1127,In_526);
nand U70 (N_70,In_771,In_514);
nor U71 (N_71,In_611,In_1081);
nor U72 (N_72,In_733,In_477);
nand U73 (N_73,In_720,In_792);
or U74 (N_74,In_796,In_185);
and U75 (N_75,In_873,In_793);
or U76 (N_76,In_998,In_462);
nand U77 (N_77,In_140,In_962);
and U78 (N_78,In_1182,In_1338);
or U79 (N_79,In_201,In_1036);
nand U80 (N_80,In_418,In_899);
or U81 (N_81,In_953,In_69);
and U82 (N_82,In_852,In_364);
nor U83 (N_83,In_1480,In_334);
and U84 (N_84,In_237,In_1256);
or U85 (N_85,In_1009,In_106);
and U86 (N_86,In_767,In_979);
xnor U87 (N_87,In_992,In_636);
or U88 (N_88,In_1155,In_1217);
nand U89 (N_89,In_465,In_675);
nand U90 (N_90,In_1125,In_1309);
nand U91 (N_91,In_532,In_1115);
or U92 (N_92,In_227,In_601);
nand U93 (N_93,In_109,In_445);
and U94 (N_94,In_838,In_823);
and U95 (N_95,In_616,In_790);
nor U96 (N_96,In_1487,In_286);
or U97 (N_97,In_331,In_102);
nor U98 (N_98,In_693,In_651);
nand U99 (N_99,In_593,In_1080);
nand U100 (N_100,In_217,In_883);
nand U101 (N_101,In_1410,In_23);
nand U102 (N_102,In_671,In_279);
nand U103 (N_103,In_595,In_1435);
nand U104 (N_104,In_906,In_322);
and U105 (N_105,In_271,In_1160);
xor U106 (N_106,In_391,In_748);
nand U107 (N_107,In_856,In_762);
nand U108 (N_108,In_1089,In_639);
nor U109 (N_109,In_918,In_936);
and U110 (N_110,In_1419,In_633);
or U111 (N_111,In_1088,In_78);
and U112 (N_112,In_863,In_233);
or U113 (N_113,In_1180,In_211);
nor U114 (N_114,In_1324,In_986);
nor U115 (N_115,In_656,In_1484);
nor U116 (N_116,In_1303,In_712);
or U117 (N_117,In_1450,In_252);
or U118 (N_118,In_1370,In_118);
or U119 (N_119,In_344,In_661);
nor U120 (N_120,In_470,In_801);
and U121 (N_121,In_777,In_1357);
or U122 (N_122,In_26,In_1471);
or U123 (N_123,In_40,In_190);
or U124 (N_124,In_981,In_1454);
and U125 (N_125,In_839,In_1280);
nor U126 (N_126,In_789,In_1215);
nor U127 (N_127,In_1226,In_259);
and U128 (N_128,In_946,In_1427);
nor U129 (N_129,In_373,In_1342);
nor U130 (N_130,In_1008,In_1047);
nand U131 (N_131,In_1406,In_837);
and U132 (N_132,In_99,In_978);
nor U133 (N_133,In_708,In_345);
nor U134 (N_134,In_1229,In_902);
and U135 (N_135,In_740,In_410);
and U136 (N_136,In_1028,In_1465);
or U137 (N_137,In_199,In_359);
or U138 (N_138,In_141,In_396);
or U139 (N_139,In_468,In_1428);
xor U140 (N_140,In_824,In_1329);
nand U141 (N_141,In_604,In_791);
and U142 (N_142,In_1183,In_642);
or U143 (N_143,In_1448,In_403);
or U144 (N_144,In_128,In_433);
or U145 (N_145,In_1085,In_483);
or U146 (N_146,In_952,In_785);
nor U147 (N_147,In_541,In_984);
nand U148 (N_148,In_1068,In_1104);
or U149 (N_149,In_246,In_615);
or U150 (N_150,In_1240,In_1322);
or U151 (N_151,In_736,In_1002);
nand U152 (N_152,In_963,In_274);
and U153 (N_153,In_262,In_12);
nor U154 (N_154,In_1071,In_457);
and U155 (N_155,In_1224,In_95);
and U156 (N_156,In_200,In_494);
and U157 (N_157,In_581,In_861);
nand U158 (N_158,In_917,In_731);
and U159 (N_159,In_1248,In_735);
and U160 (N_160,In_1114,In_301);
and U161 (N_161,In_451,In_423);
nand U162 (N_162,In_369,In_754);
or U163 (N_163,In_875,In_1472);
or U164 (N_164,In_104,In_473);
or U165 (N_165,In_1063,In_1137);
and U166 (N_166,In_181,In_1020);
and U167 (N_167,In_386,In_1139);
nand U168 (N_168,In_1122,In_496);
nor U169 (N_169,In_980,In_1268);
and U170 (N_170,In_1389,In_1306);
and U171 (N_171,In_1398,In_220);
and U172 (N_172,In_959,In_114);
or U173 (N_173,In_53,In_849);
nand U174 (N_174,In_1392,In_968);
or U175 (N_175,In_699,In_1413);
or U176 (N_176,In_1128,In_1317);
xor U177 (N_177,In_1175,In_1353);
or U178 (N_178,In_74,In_1470);
or U179 (N_179,In_698,In_1243);
or U180 (N_180,In_744,In_732);
and U181 (N_181,In_967,In_1107);
or U182 (N_182,In_41,In_1213);
xor U183 (N_183,In_93,In_618);
nor U184 (N_184,In_289,In_475);
nand U185 (N_185,In_1231,In_1230);
xor U186 (N_186,In_1262,In_1250);
nor U187 (N_187,In_22,In_1003);
nand U188 (N_188,In_1034,In_1042);
nor U189 (N_189,In_1117,In_1287);
and U190 (N_190,In_58,In_159);
nand U191 (N_191,In_174,In_1077);
and U192 (N_192,In_1135,In_910);
or U193 (N_193,In_1221,In_915);
and U194 (N_194,In_809,In_122);
nor U195 (N_195,In_449,In_33);
or U196 (N_196,In_1380,In_637);
and U197 (N_197,In_1432,In_1136);
nor U198 (N_198,In_1105,In_1446);
or U199 (N_199,In_1012,In_1388);
nand U200 (N_200,In_164,In_1142);
nor U201 (N_201,In_76,In_506);
and U202 (N_202,In_1190,In_586);
and U203 (N_203,In_24,In_1367);
and U204 (N_204,In_307,In_1005);
or U205 (N_205,In_464,In_606);
xor U206 (N_206,In_1430,In_1132);
or U207 (N_207,In_146,In_1426);
and U208 (N_208,In_562,In_319);
or U209 (N_209,In_620,In_195);
or U210 (N_210,In_1103,In_6);
xnor U211 (N_211,In_1345,In_800);
xnor U212 (N_212,In_380,In_113);
and U213 (N_213,In_871,In_1455);
or U214 (N_214,In_1112,In_715);
or U215 (N_215,In_488,In_434);
and U216 (N_216,In_395,In_415);
nor U217 (N_217,In_151,In_71);
nor U218 (N_218,In_544,In_857);
and U219 (N_219,In_152,In_1116);
nand U220 (N_220,In_356,In_1164);
nor U221 (N_221,In_343,In_1326);
or U222 (N_222,In_276,In_657);
and U223 (N_223,In_961,In_354);
nand U224 (N_224,In_121,In_133);
nor U225 (N_225,In_405,In_508);
nor U226 (N_226,In_567,In_588);
and U227 (N_227,In_497,In_895);
and U228 (N_228,In_757,In_326);
or U229 (N_229,In_1019,In_1208);
nand U230 (N_230,In_148,In_1412);
and U231 (N_231,In_230,In_817);
nor U232 (N_232,In_719,In_342);
or U233 (N_233,In_1263,In_1315);
nand U234 (N_234,In_360,In_59);
nor U235 (N_235,In_982,In_1343);
nand U236 (N_236,In_896,In_1288);
nand U237 (N_237,In_1385,In_367);
or U238 (N_238,In_388,In_716);
and U239 (N_239,In_86,In_564);
and U240 (N_240,In_1211,In_1024);
nand U241 (N_241,In_202,In_786);
nor U242 (N_242,In_363,In_515);
nor U243 (N_243,In_1133,In_62);
nor U244 (N_244,In_1485,In_452);
nand U245 (N_245,In_944,In_1049);
nand U246 (N_246,In_1356,In_408);
nor U247 (N_247,In_854,In_739);
xnor U248 (N_248,In_640,In_440);
nand U249 (N_249,In_382,In_561);
or U250 (N_250,In_1014,In_858);
xnor U251 (N_251,In_577,In_1044);
and U252 (N_252,In_466,In_450);
or U253 (N_253,In_1234,In_323);
or U254 (N_254,In_621,In_1111);
nand U255 (N_255,In_273,In_1362);
or U256 (N_256,In_594,In_1048);
nor U257 (N_257,In_80,In_1463);
xnor U258 (N_258,In_713,In_1282);
nand U259 (N_259,In_1101,In_149);
or U260 (N_260,In_1483,In_1130);
or U261 (N_261,In_659,In_467);
or U262 (N_262,In_662,In_865);
or U263 (N_263,In_568,In_1269);
and U264 (N_264,In_1102,In_283);
nand U265 (N_265,In_21,In_893);
or U266 (N_266,In_717,In_655);
nand U267 (N_267,In_528,In_376);
nor U268 (N_268,In_724,In_1156);
or U269 (N_269,In_35,In_843);
nand U270 (N_270,In_836,In_1233);
or U271 (N_271,In_647,In_1411);
xnor U272 (N_272,In_350,In_1267);
and U273 (N_273,In_339,In_797);
and U274 (N_274,In_1196,In_387);
nor U275 (N_275,In_117,In_318);
nand U276 (N_276,In_1018,In_658);
or U277 (N_277,In_503,In_691);
or U278 (N_278,In_1118,In_512);
nor U279 (N_279,In_129,In_1065);
and U280 (N_280,In_1149,In_1261);
nor U281 (N_281,In_1163,In_427);
nand U282 (N_282,In_897,In_154);
and U283 (N_283,In_79,In_0);
nand U284 (N_284,In_1286,In_600);
nor U285 (N_285,In_258,In_370);
nand U286 (N_286,In_576,In_1265);
or U287 (N_287,In_28,In_1021);
nor U288 (N_288,In_48,In_654);
and U289 (N_289,In_155,In_628);
nand U290 (N_290,In_965,In_472);
and U291 (N_291,In_1437,In_787);
and U292 (N_292,In_242,In_598);
nand U293 (N_293,In_107,In_1498);
nand U294 (N_294,In_50,In_1266);
nor U295 (N_295,In_1058,In_756);
and U296 (N_296,In_543,In_684);
nand U297 (N_297,In_1055,In_1339);
nand U298 (N_298,In_1399,In_1083);
and U299 (N_299,In_377,In_194);
nor U300 (N_300,In_752,In_964);
nor U301 (N_301,In_428,In_309);
nor U302 (N_302,In_224,In_1219);
or U303 (N_303,In_285,In_461);
nor U304 (N_304,In_687,In_442);
or U305 (N_305,In_741,In_711);
nor U306 (N_306,In_1173,In_1314);
or U307 (N_307,In_1284,In_247);
and U308 (N_308,In_814,In_495);
or U309 (N_309,In_384,In_579);
nor U310 (N_310,In_142,In_643);
nand U311 (N_311,In_138,In_1320);
nand U312 (N_312,In_177,In_850);
or U313 (N_313,In_414,In_1264);
xnor U314 (N_314,In_975,In_192);
and U315 (N_315,In_1131,In_298);
and U316 (N_316,In_1096,In_933);
nand U317 (N_317,In_288,In_1497);
or U318 (N_318,In_277,In_73);
nor U319 (N_319,In_1276,In_1436);
or U320 (N_320,In_905,In_463);
or U321 (N_321,In_348,In_291);
or U322 (N_322,In_1204,In_7);
xnor U323 (N_323,In_137,In_250);
nor U324 (N_324,In_207,In_603);
and U325 (N_325,In_1328,In_1161);
nor U326 (N_326,In_888,In_1247);
and U327 (N_327,In_419,In_1272);
nor U328 (N_328,In_1242,In_750);
nor U329 (N_329,In_763,In_904);
and U330 (N_330,In_105,In_821);
nor U331 (N_331,In_1331,In_1216);
nand U332 (N_332,In_448,In_572);
and U333 (N_333,In_1023,In_1360);
nor U334 (N_334,In_778,In_610);
or U335 (N_335,In_1281,In_822);
or U336 (N_336,In_983,In_196);
nor U337 (N_337,In_884,In_1344);
and U338 (N_338,In_312,In_504);
nand U339 (N_339,In_1205,In_846);
or U340 (N_340,In_726,In_1207);
or U341 (N_341,In_1073,In_678);
xor U342 (N_342,In_898,In_238);
and U343 (N_343,In_120,In_1400);
nand U344 (N_344,In_632,In_446);
nand U345 (N_345,In_799,In_614);
nor U346 (N_346,In_257,In_1121);
nand U347 (N_347,In_1255,In_556);
and U348 (N_348,In_1078,In_587);
nor U349 (N_349,In_243,In_1499);
nand U350 (N_350,In_4,In_1223);
nor U351 (N_351,In_1358,In_265);
and U352 (N_352,In_295,In_75);
nand U353 (N_353,In_136,In_999);
and U354 (N_354,In_1010,In_160);
nand U355 (N_355,In_275,In_1304);
nor U356 (N_356,In_1473,In_245);
nand U357 (N_357,In_1209,In_1391);
and U358 (N_358,In_517,In_1332);
nand U359 (N_359,In_125,In_92);
nand U360 (N_360,In_1253,In_1212);
and U361 (N_361,In_333,In_1067);
and U362 (N_362,In_759,In_438);
nand U363 (N_363,In_650,In_540);
or U364 (N_364,In_695,In_539);
nand U365 (N_365,In_168,In_1060);
xor U366 (N_366,In_825,In_519);
nand U367 (N_367,In_599,In_989);
and U368 (N_368,In_412,In_1007);
nand U369 (N_369,In_320,In_170);
or U370 (N_370,In_87,In_1274);
and U371 (N_371,In_29,In_175);
and U372 (N_372,In_886,In_841);
and U373 (N_373,In_700,In_1053);
nand U374 (N_374,In_1092,In_832);
nand U375 (N_375,In_1278,In_145);
nor U376 (N_376,In_811,In_530);
or U377 (N_377,In_1404,In_1218);
and U378 (N_378,In_1293,In_157);
or U379 (N_379,In_45,In_686);
nand U380 (N_380,In_1405,In_676);
and U381 (N_381,In_197,In_974);
nand U382 (N_382,In_1277,In_537);
nor U383 (N_383,In_969,In_641);
nand U384 (N_384,In_429,In_566);
nand U385 (N_385,In_1237,In_683);
and U386 (N_386,In_72,In_218);
nor U387 (N_387,In_135,In_482);
and U388 (N_388,In_987,In_198);
and U389 (N_389,In_810,In_100);
or U390 (N_390,In_1194,In_958);
and U391 (N_391,In_1227,In_18);
or U392 (N_392,In_216,In_1000);
or U393 (N_393,In_203,In_165);
and U394 (N_394,In_1294,In_110);
or U395 (N_395,In_1246,In_492);
nor U396 (N_396,In_1171,In_1254);
and U397 (N_397,In_82,In_204);
and U398 (N_398,In_553,In_714);
nor U399 (N_399,In_903,In_546);
or U400 (N_400,In_425,In_707);
or U401 (N_401,In_592,In_1192);
or U402 (N_402,In_591,In_635);
and U403 (N_403,In_630,In_251);
or U404 (N_404,In_560,In_879);
nand U405 (N_405,In_311,In_555);
nand U406 (N_406,In_609,In_14);
nor U407 (N_407,In_956,In_1099);
or U408 (N_408,In_1441,In_631);
and U409 (N_409,In_1033,In_945);
nand U410 (N_410,In_939,In_955);
or U411 (N_411,In_383,In_1378);
nor U412 (N_412,In_314,In_327);
and U413 (N_413,In_1193,In_876);
nand U414 (N_414,In_1206,In_42);
nand U415 (N_415,In_124,In_1381);
and U416 (N_416,In_536,In_772);
and U417 (N_417,In_278,In_1372);
nand U418 (N_418,In_302,In_420);
or U419 (N_419,In_747,In_214);
or U420 (N_420,In_1292,In_436);
nor U421 (N_421,In_1091,In_61);
xor U422 (N_422,In_111,In_439);
nand U423 (N_423,In_971,In_266);
or U424 (N_424,In_890,In_63);
nand U425 (N_425,In_749,In_626);
nand U426 (N_426,In_848,In_923);
nand U427 (N_427,In_1051,In_17);
or U428 (N_428,In_255,In_704);
or U429 (N_429,In_885,In_527);
nor U430 (N_430,In_1084,In_55);
nor U431 (N_431,In_835,In_1474);
and U432 (N_432,In_290,In_229);
nor U433 (N_433,In_1363,In_1424);
and U434 (N_434,In_1408,In_455);
or U435 (N_435,In_1318,In_894);
or U436 (N_436,In_1260,In_413);
and U437 (N_437,In_116,In_1201);
and U438 (N_438,In_281,In_892);
nand U439 (N_439,In_1082,In_795);
and U440 (N_440,In_1075,In_437);
nand U441 (N_441,In_928,In_163);
nand U442 (N_442,In_453,In_263);
nor U443 (N_443,In_550,In_935);
and U444 (N_444,In_585,In_417);
and U445 (N_445,In_37,In_673);
or U446 (N_446,In_206,In_1232);
nand U447 (N_447,In_187,In_1346);
xnor U448 (N_448,In_1371,In_347);
nand U449 (N_449,In_887,In_1016);
or U450 (N_450,In_548,In_1416);
or U451 (N_451,In_559,In_1393);
or U452 (N_452,In_1364,In_1312);
and U453 (N_453,In_855,In_573);
and U454 (N_454,In_1369,In_1032);
and U455 (N_455,In_287,In_816);
and U456 (N_456,In_1466,In_38);
or U457 (N_457,In_689,In_834);
nand U458 (N_458,In_1129,In_751);
or U459 (N_459,In_1108,In_1057);
nor U460 (N_460,In_435,In_507);
nand U461 (N_461,In_409,In_328);
and U462 (N_462,In_794,In_1496);
or U463 (N_463,In_1488,In_976);
and U464 (N_464,In_1239,In_1095);
and U465 (N_465,In_991,In_694);
and U466 (N_466,In_490,In_126);
nor U467 (N_467,In_1062,In_529);
or U468 (N_468,In_305,In_666);
nand U469 (N_469,In_1202,In_1297);
nand U470 (N_470,In_1373,In_1382);
nand U471 (N_471,In_30,In_426);
or U472 (N_472,In_166,In_912);
nor U473 (N_473,In_1188,In_803);
nand U474 (N_474,In_520,In_1176);
xnor U475 (N_475,In_1451,In_1147);
nor U476 (N_476,In_167,In_94);
xor U477 (N_477,In_329,In_2);
nand U478 (N_478,In_677,In_680);
nand U479 (N_479,In_421,In_19);
nor U480 (N_480,In_1258,In_1059);
nor U481 (N_481,In_1152,In_1257);
or U482 (N_482,In_231,In_1401);
nor U483 (N_483,In_134,In_1197);
xnor U484 (N_484,In_20,In_925);
nor U485 (N_485,In_5,In_1335);
or U486 (N_486,In_1126,In_1056);
or U487 (N_487,In_213,In_171);
nand U488 (N_488,In_574,In_221);
and U489 (N_489,In_374,In_422);
nor U490 (N_490,In_538,In_702);
nand U491 (N_491,In_1245,In_1157);
or U492 (N_492,In_1222,In_1198);
nand U493 (N_493,In_299,In_847);
and U494 (N_494,In_706,In_869);
or U495 (N_495,In_597,In_390);
nand U496 (N_496,In_510,In_162);
and U497 (N_497,In_254,In_584);
nand U498 (N_498,In_590,In_919);
or U499 (N_499,In_1415,In_1110);
or U500 (N_500,In_1165,In_489);
or U501 (N_501,In_340,In_223);
and U502 (N_502,In_634,In_67);
nor U503 (N_503,In_1225,In_525);
nand U504 (N_504,In_1403,In_357);
or U505 (N_505,In_995,In_1072);
nor U506 (N_506,In_1375,In_296);
and U507 (N_507,In_179,In_1429);
nor U508 (N_508,In_430,In_578);
nor U509 (N_509,In_270,In_569);
nor U510 (N_510,In_1220,In_742);
nor U511 (N_511,In_1030,In_234);
nor U512 (N_512,In_253,In_297);
nor U513 (N_513,In_781,In_1352);
and U514 (N_514,In_608,In_460);
nor U515 (N_515,In_70,In_1479);
nand U516 (N_516,In_827,In_696);
nor U517 (N_517,In_1327,In_638);
and U518 (N_518,In_685,In_1445);
and U519 (N_519,In_361,In_1431);
or U520 (N_520,In_481,In_225);
or U521 (N_521,In_303,In_156);
nor U522 (N_522,In_176,In_1249);
or U523 (N_523,In_173,In_371);
nor U524 (N_524,In_335,In_881);
nor U525 (N_525,In_833,In_306);
or U526 (N_526,In_1407,In_407);
nand U527 (N_527,In_161,In_222);
nor U528 (N_528,In_901,In_1402);
and U529 (N_529,In_619,In_697);
nor U530 (N_530,In_1476,In_459);
and U531 (N_531,In_1374,In_1038);
or U532 (N_532,In_65,In_669);
nand U533 (N_533,In_1444,In_954);
or U534 (N_534,In_1195,In_997);
and U535 (N_535,In_513,In_668);
and U536 (N_536,In_563,In_1296);
and U537 (N_537,In_1124,In_509);
nand U538 (N_538,In_1291,In_191);
xnor U539 (N_539,In_927,In_378);
and U540 (N_540,In_900,In_317);
nor U541 (N_541,In_143,In_189);
nand U542 (N_542,In_1066,In_602);
nand U543 (N_543,In_1177,In_1094);
nand U544 (N_544,In_914,In_77);
or U545 (N_545,In_1414,In_1039);
nor U546 (N_546,In_31,In_493);
or U547 (N_547,In_690,In_90);
or U548 (N_548,In_589,In_1158);
nand U549 (N_549,In_663,In_441);
nand U550 (N_550,In_966,In_1325);
and U551 (N_551,In_769,In_1273);
and U552 (N_552,In_219,In_1025);
nor U553 (N_553,In_624,In_178);
and U554 (N_554,In_891,In_547);
or U555 (N_555,In_313,In_623);
nand U556 (N_556,In_1181,In_1361);
and U557 (N_557,In_728,In_761);
and U558 (N_558,In_8,In_753);
or U559 (N_559,In_1031,In_1489);
and U560 (N_560,In_1313,In_321);
nand U561 (N_561,In_1397,In_664);
and U562 (N_562,In_1365,In_476);
xor U563 (N_563,In_1141,In_580);
nor U564 (N_564,In_209,In_1153);
and U565 (N_565,In_498,In_487);
or U566 (N_566,In_1453,In_127);
xnor U567 (N_567,In_1347,In_874);
nor U568 (N_568,In_1,In_46);
and U569 (N_569,In_264,In_432);
xnor U570 (N_570,In_362,In_1308);
and U571 (N_571,In_336,In_779);
and U572 (N_572,In_644,In_1123);
nor U573 (N_573,In_332,In_575);
and U574 (N_574,In_501,In_931);
or U575 (N_575,In_183,In_1458);
nor U576 (N_576,In_880,In_499);
and U577 (N_577,In_1351,In_629);
nand U578 (N_578,In_1100,In_866);
or U579 (N_579,In_381,In_878);
and U580 (N_580,In_921,In_596);
nand U581 (N_581,In_788,In_929);
and U582 (N_582,In_554,In_826);
and U583 (N_583,In_721,In_970);
nor U584 (N_584,In_416,In_985);
or U585 (N_585,In_471,In_502);
xnor U586 (N_586,In_1006,In_397);
nor U587 (N_587,In_1064,In_988);
and U588 (N_588,In_1259,In_552);
and U589 (N_589,In_938,In_365);
nor U590 (N_590,In_119,In_123);
or U591 (N_591,In_478,In_272);
nor U592 (N_592,In_300,In_1087);
nand U593 (N_593,In_1418,In_1438);
or U594 (N_594,In_782,In_458);
and U595 (N_595,In_130,In_147);
nand U596 (N_596,In_1186,In_1235);
nand U597 (N_597,In_1070,In_972);
nor U598 (N_598,In_557,In_84);
or U599 (N_599,In_484,In_1310);
or U600 (N_600,In_960,In_98);
nor U601 (N_601,In_115,In_1001);
nand U602 (N_602,In_1168,In_310);
and U603 (N_603,In_1495,In_911);
and U604 (N_604,In_924,In_705);
nor U605 (N_605,In_284,In_1045);
or U606 (N_606,In_316,In_112);
xor U607 (N_607,In_184,In_1439);
nand U608 (N_608,In_1022,In_1423);
nor U609 (N_609,In_1054,In_212);
nand U610 (N_610,In_16,In_1494);
nand U611 (N_611,In_1214,In_424);
or U612 (N_612,In_132,In_52);
nor U613 (N_613,In_1166,In_916);
nor U614 (N_614,In_54,In_725);
or U615 (N_615,In_1421,In_920);
nand U616 (N_616,In_649,In_862);
xnor U617 (N_617,In_583,In_1493);
nor U618 (N_618,In_864,In_868);
nor U619 (N_619,In_215,In_709);
nand U620 (N_620,In_228,In_1300);
or U621 (N_621,In_907,In_934);
xnor U622 (N_622,In_169,In_89);
and U623 (N_623,In_353,In_261);
xor U624 (N_624,In_1013,In_1390);
or U625 (N_625,In_622,In_394);
nand U626 (N_626,In_34,In_393);
and U627 (N_627,In_269,In_43);
nand U628 (N_628,In_1354,In_68);
nand U629 (N_629,In_188,In_1457);
and U630 (N_630,In_948,In_851);
and U631 (N_631,In_535,In_570);
and U632 (N_632,In_282,In_1299);
or U633 (N_633,In_341,In_97);
and U634 (N_634,In_1043,In_518);
or U635 (N_635,In_60,In_1046);
nor U636 (N_636,In_1323,In_153);
nor U637 (N_637,In_860,In_1076);
nand U638 (N_638,In_780,In_994);
and U639 (N_639,In_820,In_1228);
xor U640 (N_640,In_627,In_1464);
and U641 (N_641,In_1449,In_1290);
or U642 (N_642,In_831,In_88);
or U643 (N_643,In_973,In_766);
or U644 (N_644,In_1420,In_346);
nor U645 (N_645,In_249,In_351);
or U646 (N_646,In_47,In_1359);
nand U647 (N_647,In_39,In_1199);
or U648 (N_648,In_682,In_10);
nand U649 (N_649,In_745,In_996);
nor U650 (N_650,In_401,In_913);
and U651 (N_651,In_180,In_1011);
nand U652 (N_652,In_1113,In_1069);
nand U653 (N_653,In_1191,In_806);
nor U654 (N_654,In_882,In_829);
nand U655 (N_655,In_193,In_1461);
nor U656 (N_656,In_770,In_947);
and U657 (N_657,In_1210,In_1244);
or U658 (N_658,In_565,In_1179);
nand U659 (N_659,In_1184,In_1311);
nand U660 (N_660,In_372,In_236);
nand U661 (N_661,In_304,In_840);
or U662 (N_662,In_760,In_1143);
or U663 (N_663,In_815,In_605);
and U664 (N_664,In_737,In_56);
nand U665 (N_665,In_226,In_404);
nor U666 (N_666,In_867,In_1145);
and U667 (N_667,In_1396,In_765);
and U668 (N_668,In_722,In_819);
nand U669 (N_669,In_454,In_1492);
or U670 (N_670,In_922,In_1162);
nor U671 (N_671,In_813,In_1187);
and U672 (N_672,In_210,In_308);
nor U673 (N_673,In_280,In_941);
or U674 (N_674,In_1379,In_1252);
nand U675 (N_675,In_241,In_727);
and U676 (N_676,In_1417,In_718);
or U677 (N_677,In_1040,In_1302);
and U678 (N_678,In_1376,In_1440);
nand U679 (N_679,In_665,In_516);
xor U680 (N_680,In_256,In_889);
or U681 (N_681,In_625,In_244);
nor U682 (N_682,In_805,In_293);
and U683 (N_683,In_842,In_534);
nor U684 (N_684,In_1336,In_431);
nand U685 (N_685,In_406,In_1482);
nand U686 (N_686,In_91,In_366);
or U687 (N_687,In_1017,In_1316);
nor U688 (N_688,In_1467,In_1348);
or U689 (N_689,In_338,In_32);
or U690 (N_690,In_400,In_1134);
nor U691 (N_691,In_688,In_1090);
nor U692 (N_692,In_773,In_1349);
nor U693 (N_693,In_325,In_1189);
xor U694 (N_694,In_993,In_1037);
nor U695 (N_695,In_96,In_1366);
and U696 (N_696,In_743,In_292);
or U697 (N_697,In_25,In_267);
nand U698 (N_698,In_932,In_444);
nor U699 (N_699,In_783,In_1319);
and U700 (N_700,In_1289,In_389);
nand U701 (N_701,In_1434,In_558);
or U702 (N_702,In_158,In_1301);
nand U703 (N_703,In_85,In_83);
nand U704 (N_704,In_392,In_774);
nand U705 (N_705,In_1119,In_186);
nor U706 (N_706,In_1035,In_15);
or U707 (N_707,In_758,In_1074);
or U708 (N_708,In_385,In_807);
nand U709 (N_709,In_13,In_1150);
and U710 (N_710,In_1052,In_1285);
and U711 (N_711,In_909,In_1477);
and U712 (N_712,In_1490,In_1340);
nor U713 (N_713,In_755,In_1387);
xor U714 (N_714,In_3,In_542);
and U715 (N_715,In_692,In_1321);
or U716 (N_716,In_398,In_828);
nand U717 (N_717,In_240,In_990);
and U718 (N_718,In_447,In_1086);
and U719 (N_719,In_379,In_784);
nand U720 (N_720,In_738,In_355);
xor U721 (N_721,In_1270,In_617);
and U722 (N_722,In_399,In_667);
or U723 (N_723,In_1154,In_1027);
and U724 (N_724,In_1236,In_723);
or U725 (N_725,In_768,In_315);
and U726 (N_726,In_1384,In_294);
and U727 (N_727,In_522,In_101);
nor U728 (N_728,In_500,In_330);
nor U729 (N_729,In_486,In_1350);
nand U730 (N_730,In_9,In_648);
or U731 (N_731,In_1355,In_172);
nand U732 (N_732,In_1169,In_491);
nor U733 (N_733,In_1456,In_485);
nand U734 (N_734,In_652,In_260);
and U735 (N_735,In_1151,In_57);
nor U736 (N_736,In_352,In_208);
nor U737 (N_737,In_1447,In_402);
nand U738 (N_738,In_545,In_1146);
and U739 (N_739,In_51,In_1279);
nand U740 (N_740,In_1203,In_1238);
or U741 (N_741,In_1481,In_474);
and U742 (N_742,In_926,In_182);
nand U743 (N_743,In_521,In_1459);
nand U744 (N_744,In_844,In_812);
nand U745 (N_745,In_1478,In_1004);
nand U746 (N_746,In_949,In_872);
nor U747 (N_747,In_1061,In_681);
and U748 (N_748,In_672,In_66);
nand U749 (N_749,In_950,In_411);
nand U750 (N_750,In_99,In_341);
nand U751 (N_751,In_960,In_1309);
nand U752 (N_752,In_556,In_1113);
nand U753 (N_753,In_478,In_771);
or U754 (N_754,In_992,In_1394);
or U755 (N_755,In_512,In_1111);
nor U756 (N_756,In_922,In_563);
or U757 (N_757,In_1172,In_584);
nand U758 (N_758,In_1281,In_1323);
nor U759 (N_759,In_680,In_331);
nor U760 (N_760,In_800,In_780);
or U761 (N_761,In_435,In_1056);
nand U762 (N_762,In_77,In_1294);
nor U763 (N_763,In_1229,In_536);
nand U764 (N_764,In_1314,In_363);
or U765 (N_765,In_1069,In_1349);
nor U766 (N_766,In_210,In_755);
nand U767 (N_767,In_1232,In_1060);
and U768 (N_768,In_341,In_1289);
nor U769 (N_769,In_833,In_561);
nand U770 (N_770,In_1352,In_262);
and U771 (N_771,In_1392,In_825);
and U772 (N_772,In_806,In_983);
nor U773 (N_773,In_1154,In_457);
nand U774 (N_774,In_645,In_87);
nor U775 (N_775,In_1493,In_539);
or U776 (N_776,In_1328,In_412);
nor U777 (N_777,In_323,In_1144);
nor U778 (N_778,In_1394,In_233);
nand U779 (N_779,In_916,In_1423);
nand U780 (N_780,In_1129,In_760);
or U781 (N_781,In_1498,In_724);
nand U782 (N_782,In_1294,In_125);
nor U783 (N_783,In_12,In_696);
nor U784 (N_784,In_205,In_746);
nor U785 (N_785,In_155,In_705);
or U786 (N_786,In_681,In_10);
nand U787 (N_787,In_731,In_1310);
nand U788 (N_788,In_247,In_670);
nor U789 (N_789,In_978,In_742);
or U790 (N_790,In_156,In_179);
nand U791 (N_791,In_643,In_912);
nand U792 (N_792,In_593,In_1208);
nor U793 (N_793,In_499,In_1128);
nor U794 (N_794,In_1440,In_1038);
nand U795 (N_795,In_266,In_1468);
and U796 (N_796,In_798,In_1498);
nor U797 (N_797,In_760,In_260);
or U798 (N_798,In_343,In_698);
nor U799 (N_799,In_760,In_973);
and U800 (N_800,In_313,In_473);
and U801 (N_801,In_911,In_687);
xnor U802 (N_802,In_1340,In_80);
nor U803 (N_803,In_1414,In_385);
nor U804 (N_804,In_681,In_1234);
nand U805 (N_805,In_1009,In_111);
nor U806 (N_806,In_186,In_953);
and U807 (N_807,In_1422,In_1488);
and U808 (N_808,In_116,In_1087);
or U809 (N_809,In_1052,In_553);
and U810 (N_810,In_312,In_304);
nor U811 (N_811,In_1159,In_312);
and U812 (N_812,In_950,In_926);
or U813 (N_813,In_1075,In_1160);
nand U814 (N_814,In_399,In_502);
nor U815 (N_815,In_361,In_215);
nand U816 (N_816,In_1487,In_1044);
nor U817 (N_817,In_343,In_20);
or U818 (N_818,In_115,In_738);
or U819 (N_819,In_1013,In_993);
and U820 (N_820,In_1477,In_393);
xnor U821 (N_821,In_1404,In_1124);
nor U822 (N_822,In_1361,In_1478);
xor U823 (N_823,In_1017,In_130);
nand U824 (N_824,In_113,In_975);
or U825 (N_825,In_521,In_774);
nand U826 (N_826,In_1259,In_1316);
nand U827 (N_827,In_617,In_1028);
nor U828 (N_828,In_8,In_413);
or U829 (N_829,In_317,In_1258);
or U830 (N_830,In_302,In_1251);
xnor U831 (N_831,In_1117,In_284);
nand U832 (N_832,In_629,In_714);
and U833 (N_833,In_1116,In_489);
nand U834 (N_834,In_526,In_1435);
nor U835 (N_835,In_615,In_676);
xnor U836 (N_836,In_290,In_383);
nor U837 (N_837,In_702,In_1082);
or U838 (N_838,In_840,In_204);
nand U839 (N_839,In_935,In_297);
and U840 (N_840,In_20,In_1364);
xor U841 (N_841,In_1036,In_622);
nand U842 (N_842,In_361,In_325);
nor U843 (N_843,In_1430,In_464);
and U844 (N_844,In_912,In_630);
and U845 (N_845,In_313,In_582);
nand U846 (N_846,In_123,In_1474);
nand U847 (N_847,In_473,In_1128);
or U848 (N_848,In_4,In_753);
nor U849 (N_849,In_1406,In_232);
nor U850 (N_850,In_311,In_650);
nor U851 (N_851,In_1012,In_821);
and U852 (N_852,In_1011,In_748);
nor U853 (N_853,In_1306,In_859);
or U854 (N_854,In_959,In_809);
or U855 (N_855,In_852,In_782);
nand U856 (N_856,In_953,In_1164);
or U857 (N_857,In_237,In_830);
or U858 (N_858,In_17,In_1462);
and U859 (N_859,In_275,In_473);
or U860 (N_860,In_802,In_63);
nand U861 (N_861,In_782,In_370);
nor U862 (N_862,In_404,In_383);
nor U863 (N_863,In_582,In_534);
nand U864 (N_864,In_259,In_310);
nand U865 (N_865,In_86,In_663);
or U866 (N_866,In_152,In_601);
and U867 (N_867,In_937,In_1173);
nor U868 (N_868,In_334,In_44);
nand U869 (N_869,In_982,In_1231);
xor U870 (N_870,In_272,In_1442);
nand U871 (N_871,In_73,In_1038);
and U872 (N_872,In_435,In_1479);
nand U873 (N_873,In_1355,In_592);
nand U874 (N_874,In_1350,In_931);
and U875 (N_875,In_383,In_761);
and U876 (N_876,In_1138,In_1214);
and U877 (N_877,In_1348,In_909);
nor U878 (N_878,In_175,In_83);
nor U879 (N_879,In_415,In_507);
or U880 (N_880,In_661,In_674);
and U881 (N_881,In_1350,In_1253);
nand U882 (N_882,In_726,In_1052);
nand U883 (N_883,In_494,In_1450);
nor U884 (N_884,In_363,In_1343);
nor U885 (N_885,In_713,In_234);
nand U886 (N_886,In_280,In_551);
and U887 (N_887,In_1210,In_1344);
or U888 (N_888,In_734,In_623);
nor U889 (N_889,In_827,In_632);
nor U890 (N_890,In_811,In_1171);
nand U891 (N_891,In_1039,In_734);
nand U892 (N_892,In_949,In_1111);
or U893 (N_893,In_1074,In_564);
nand U894 (N_894,In_361,In_297);
or U895 (N_895,In_369,In_820);
nor U896 (N_896,In_417,In_882);
nor U897 (N_897,In_1461,In_1236);
and U898 (N_898,In_166,In_607);
nand U899 (N_899,In_765,In_380);
nand U900 (N_900,In_435,In_1375);
nor U901 (N_901,In_540,In_1362);
xor U902 (N_902,In_1223,In_1059);
and U903 (N_903,In_748,In_460);
and U904 (N_904,In_1414,In_1377);
or U905 (N_905,In_1228,In_1005);
nand U906 (N_906,In_704,In_702);
nor U907 (N_907,In_1179,In_967);
or U908 (N_908,In_1449,In_1443);
or U909 (N_909,In_1429,In_413);
or U910 (N_910,In_1007,In_1499);
and U911 (N_911,In_251,In_1319);
nand U912 (N_912,In_866,In_1132);
nand U913 (N_913,In_858,In_335);
and U914 (N_914,In_670,In_172);
or U915 (N_915,In_1037,In_885);
nand U916 (N_916,In_178,In_317);
nor U917 (N_917,In_1099,In_183);
xor U918 (N_918,In_1415,In_315);
or U919 (N_919,In_1244,In_1441);
or U920 (N_920,In_1438,In_190);
nor U921 (N_921,In_156,In_671);
or U922 (N_922,In_89,In_1472);
or U923 (N_923,In_349,In_442);
and U924 (N_924,In_260,In_858);
or U925 (N_925,In_798,In_64);
or U926 (N_926,In_288,In_837);
nand U927 (N_927,In_1350,In_855);
nor U928 (N_928,In_423,In_1213);
nor U929 (N_929,In_892,In_997);
or U930 (N_930,In_26,In_1283);
nand U931 (N_931,In_1451,In_159);
and U932 (N_932,In_266,In_1070);
and U933 (N_933,In_213,In_1058);
and U934 (N_934,In_314,In_638);
and U935 (N_935,In_1071,In_1385);
or U936 (N_936,In_220,In_329);
and U937 (N_937,In_665,In_175);
nand U938 (N_938,In_1317,In_1382);
and U939 (N_939,In_897,In_1370);
and U940 (N_940,In_1433,In_225);
xor U941 (N_941,In_918,In_290);
or U942 (N_942,In_388,In_374);
xnor U943 (N_943,In_755,In_1409);
nor U944 (N_944,In_1026,In_182);
or U945 (N_945,In_451,In_908);
and U946 (N_946,In_172,In_1048);
nor U947 (N_947,In_66,In_876);
nand U948 (N_948,In_39,In_323);
nand U949 (N_949,In_1407,In_622);
or U950 (N_950,In_494,In_1128);
and U951 (N_951,In_500,In_259);
and U952 (N_952,In_1300,In_32);
and U953 (N_953,In_868,In_1284);
nor U954 (N_954,In_825,In_915);
and U955 (N_955,In_973,In_520);
or U956 (N_956,In_170,In_1309);
or U957 (N_957,In_1240,In_1462);
and U958 (N_958,In_1078,In_908);
nor U959 (N_959,In_210,In_780);
nor U960 (N_960,In_76,In_990);
and U961 (N_961,In_379,In_168);
nand U962 (N_962,In_1360,In_1461);
and U963 (N_963,In_1454,In_493);
nand U964 (N_964,In_386,In_926);
or U965 (N_965,In_347,In_1386);
nand U966 (N_966,In_79,In_330);
or U967 (N_967,In_316,In_937);
and U968 (N_968,In_716,In_333);
nor U969 (N_969,In_641,In_70);
nand U970 (N_970,In_207,In_457);
nand U971 (N_971,In_1355,In_1412);
nor U972 (N_972,In_699,In_982);
nor U973 (N_973,In_544,In_461);
nor U974 (N_974,In_85,In_1095);
nand U975 (N_975,In_1267,In_484);
nor U976 (N_976,In_171,In_908);
and U977 (N_977,In_274,In_228);
nand U978 (N_978,In_129,In_147);
nor U979 (N_979,In_409,In_1149);
nor U980 (N_980,In_1061,In_1100);
nor U981 (N_981,In_868,In_155);
nor U982 (N_982,In_1197,In_1028);
or U983 (N_983,In_1007,In_76);
and U984 (N_984,In_877,In_1222);
nand U985 (N_985,In_912,In_793);
nand U986 (N_986,In_954,In_345);
nand U987 (N_987,In_172,In_190);
nor U988 (N_988,In_909,In_388);
and U989 (N_989,In_1072,In_917);
or U990 (N_990,In_295,In_634);
or U991 (N_991,In_1245,In_1197);
and U992 (N_992,In_534,In_39);
and U993 (N_993,In_320,In_255);
or U994 (N_994,In_784,In_391);
nand U995 (N_995,In_570,In_1294);
nand U996 (N_996,In_1272,In_902);
and U997 (N_997,In_1096,In_502);
xnor U998 (N_998,In_794,In_1180);
xnor U999 (N_999,In_1276,In_927);
nor U1000 (N_1000,In_971,In_612);
and U1001 (N_1001,In_473,In_1029);
or U1002 (N_1002,In_1219,In_1189);
nand U1003 (N_1003,In_1452,In_716);
or U1004 (N_1004,In_1314,In_327);
nor U1005 (N_1005,In_1284,In_53);
or U1006 (N_1006,In_260,In_67);
nor U1007 (N_1007,In_1192,In_1445);
and U1008 (N_1008,In_1291,In_979);
nor U1009 (N_1009,In_1172,In_534);
and U1010 (N_1010,In_489,In_898);
and U1011 (N_1011,In_1019,In_503);
and U1012 (N_1012,In_809,In_155);
and U1013 (N_1013,In_278,In_1405);
nor U1014 (N_1014,In_140,In_1270);
and U1015 (N_1015,In_1355,In_755);
or U1016 (N_1016,In_191,In_1);
or U1017 (N_1017,In_757,In_651);
nor U1018 (N_1018,In_949,In_1168);
nor U1019 (N_1019,In_746,In_867);
and U1020 (N_1020,In_522,In_5);
and U1021 (N_1021,In_501,In_137);
nor U1022 (N_1022,In_208,In_465);
and U1023 (N_1023,In_1428,In_1091);
and U1024 (N_1024,In_396,In_1074);
nor U1025 (N_1025,In_315,In_125);
and U1026 (N_1026,In_28,In_1358);
nand U1027 (N_1027,In_1305,In_1473);
nor U1028 (N_1028,In_635,In_437);
nor U1029 (N_1029,In_95,In_1232);
or U1030 (N_1030,In_1219,In_673);
and U1031 (N_1031,In_644,In_759);
nor U1032 (N_1032,In_269,In_814);
nand U1033 (N_1033,In_932,In_164);
nor U1034 (N_1034,In_954,In_786);
and U1035 (N_1035,In_657,In_1163);
nor U1036 (N_1036,In_428,In_315);
nor U1037 (N_1037,In_510,In_1207);
or U1038 (N_1038,In_769,In_465);
nand U1039 (N_1039,In_1438,In_1434);
nand U1040 (N_1040,In_752,In_448);
or U1041 (N_1041,In_983,In_1263);
and U1042 (N_1042,In_169,In_537);
nand U1043 (N_1043,In_1177,In_80);
nor U1044 (N_1044,In_341,In_669);
or U1045 (N_1045,In_1097,In_305);
nand U1046 (N_1046,In_1408,In_1060);
and U1047 (N_1047,In_1293,In_771);
and U1048 (N_1048,In_585,In_1157);
or U1049 (N_1049,In_341,In_950);
nor U1050 (N_1050,In_135,In_1045);
nor U1051 (N_1051,In_145,In_903);
nor U1052 (N_1052,In_712,In_876);
or U1053 (N_1053,In_770,In_801);
xnor U1054 (N_1054,In_301,In_34);
nor U1055 (N_1055,In_899,In_779);
nor U1056 (N_1056,In_1419,In_683);
or U1057 (N_1057,In_380,In_727);
nand U1058 (N_1058,In_277,In_154);
or U1059 (N_1059,In_1424,In_593);
or U1060 (N_1060,In_438,In_88);
nand U1061 (N_1061,In_686,In_973);
nand U1062 (N_1062,In_236,In_448);
nor U1063 (N_1063,In_397,In_1238);
nor U1064 (N_1064,In_423,In_1163);
xor U1065 (N_1065,In_780,In_1362);
or U1066 (N_1066,In_621,In_1147);
and U1067 (N_1067,In_458,In_767);
nor U1068 (N_1068,In_745,In_738);
xor U1069 (N_1069,In_997,In_1258);
xnor U1070 (N_1070,In_699,In_1005);
nand U1071 (N_1071,In_360,In_1279);
and U1072 (N_1072,In_1044,In_376);
or U1073 (N_1073,In_858,In_298);
nor U1074 (N_1074,In_1410,In_697);
and U1075 (N_1075,In_1248,In_871);
nand U1076 (N_1076,In_1152,In_995);
nand U1077 (N_1077,In_1260,In_1287);
or U1078 (N_1078,In_1257,In_350);
nand U1079 (N_1079,In_1467,In_1337);
or U1080 (N_1080,In_970,In_46);
and U1081 (N_1081,In_638,In_45);
and U1082 (N_1082,In_1194,In_1054);
nand U1083 (N_1083,In_733,In_1156);
and U1084 (N_1084,In_1447,In_349);
and U1085 (N_1085,In_1273,In_408);
nor U1086 (N_1086,In_1248,In_1419);
and U1087 (N_1087,In_397,In_485);
nand U1088 (N_1088,In_214,In_1358);
and U1089 (N_1089,In_548,In_4);
or U1090 (N_1090,In_316,In_1200);
nand U1091 (N_1091,In_489,In_5);
nand U1092 (N_1092,In_235,In_1058);
or U1093 (N_1093,In_1108,In_192);
nor U1094 (N_1094,In_37,In_1124);
nand U1095 (N_1095,In_531,In_1217);
or U1096 (N_1096,In_834,In_504);
or U1097 (N_1097,In_1362,In_913);
xor U1098 (N_1098,In_885,In_1340);
nor U1099 (N_1099,In_755,In_668);
and U1100 (N_1100,In_516,In_1316);
xnor U1101 (N_1101,In_321,In_37);
and U1102 (N_1102,In_197,In_1414);
and U1103 (N_1103,In_748,In_1135);
xor U1104 (N_1104,In_1418,In_1202);
or U1105 (N_1105,In_1479,In_839);
nand U1106 (N_1106,In_659,In_1204);
nand U1107 (N_1107,In_818,In_670);
xnor U1108 (N_1108,In_1284,In_592);
or U1109 (N_1109,In_28,In_1195);
or U1110 (N_1110,In_538,In_1075);
or U1111 (N_1111,In_721,In_1128);
and U1112 (N_1112,In_481,In_883);
or U1113 (N_1113,In_1157,In_1336);
and U1114 (N_1114,In_659,In_396);
and U1115 (N_1115,In_1,In_702);
nor U1116 (N_1116,In_1035,In_261);
and U1117 (N_1117,In_621,In_216);
or U1118 (N_1118,In_1198,In_73);
or U1119 (N_1119,In_1051,In_1312);
nand U1120 (N_1120,In_585,In_1093);
nand U1121 (N_1121,In_1477,In_991);
and U1122 (N_1122,In_849,In_96);
and U1123 (N_1123,In_423,In_1285);
nor U1124 (N_1124,In_1458,In_1009);
nor U1125 (N_1125,In_775,In_910);
nand U1126 (N_1126,In_496,In_1028);
nor U1127 (N_1127,In_1408,In_550);
and U1128 (N_1128,In_244,In_619);
nand U1129 (N_1129,In_819,In_701);
and U1130 (N_1130,In_124,In_257);
or U1131 (N_1131,In_1234,In_1427);
and U1132 (N_1132,In_939,In_88);
and U1133 (N_1133,In_1483,In_1087);
xnor U1134 (N_1134,In_757,In_971);
nor U1135 (N_1135,In_537,In_123);
or U1136 (N_1136,In_273,In_840);
nand U1137 (N_1137,In_466,In_985);
nor U1138 (N_1138,In_36,In_469);
or U1139 (N_1139,In_35,In_1286);
nand U1140 (N_1140,In_893,In_412);
nand U1141 (N_1141,In_507,In_513);
nor U1142 (N_1142,In_1401,In_97);
and U1143 (N_1143,In_360,In_407);
nor U1144 (N_1144,In_105,In_887);
or U1145 (N_1145,In_458,In_594);
nor U1146 (N_1146,In_579,In_1382);
and U1147 (N_1147,In_1067,In_955);
nor U1148 (N_1148,In_766,In_893);
and U1149 (N_1149,In_302,In_798);
or U1150 (N_1150,In_150,In_874);
and U1151 (N_1151,In_590,In_199);
nor U1152 (N_1152,In_1467,In_1183);
nor U1153 (N_1153,In_897,In_1101);
or U1154 (N_1154,In_266,In_614);
or U1155 (N_1155,In_141,In_1109);
nand U1156 (N_1156,In_916,In_360);
nand U1157 (N_1157,In_814,In_763);
nand U1158 (N_1158,In_1175,In_319);
nor U1159 (N_1159,In_131,In_311);
nand U1160 (N_1160,In_219,In_639);
nand U1161 (N_1161,In_1258,In_950);
nor U1162 (N_1162,In_393,In_243);
and U1163 (N_1163,In_597,In_85);
and U1164 (N_1164,In_69,In_1352);
and U1165 (N_1165,In_239,In_1267);
nand U1166 (N_1166,In_704,In_740);
or U1167 (N_1167,In_548,In_845);
nor U1168 (N_1168,In_927,In_553);
nand U1169 (N_1169,In_273,In_159);
nand U1170 (N_1170,In_240,In_1317);
and U1171 (N_1171,In_673,In_311);
or U1172 (N_1172,In_839,In_317);
nand U1173 (N_1173,In_1416,In_686);
nor U1174 (N_1174,In_614,In_326);
nand U1175 (N_1175,In_916,In_800);
nand U1176 (N_1176,In_1,In_797);
and U1177 (N_1177,In_1048,In_1220);
nor U1178 (N_1178,In_1323,In_552);
nor U1179 (N_1179,In_1073,In_989);
xnor U1180 (N_1180,In_1000,In_855);
and U1181 (N_1181,In_109,In_771);
and U1182 (N_1182,In_218,In_1068);
or U1183 (N_1183,In_245,In_1034);
and U1184 (N_1184,In_1115,In_1334);
nor U1185 (N_1185,In_1109,In_580);
and U1186 (N_1186,In_632,In_1141);
and U1187 (N_1187,In_98,In_1149);
nor U1188 (N_1188,In_407,In_1111);
xnor U1189 (N_1189,In_468,In_848);
nor U1190 (N_1190,In_1387,In_534);
and U1191 (N_1191,In_694,In_388);
and U1192 (N_1192,In_1282,In_974);
nand U1193 (N_1193,In_674,In_523);
nand U1194 (N_1194,In_791,In_729);
nand U1195 (N_1195,In_1481,In_678);
or U1196 (N_1196,In_517,In_198);
nand U1197 (N_1197,In_1374,In_767);
nand U1198 (N_1198,In_1161,In_768);
and U1199 (N_1199,In_1358,In_1411);
nand U1200 (N_1200,In_1272,In_1050);
nor U1201 (N_1201,In_1051,In_694);
and U1202 (N_1202,In_158,In_577);
nand U1203 (N_1203,In_840,In_1012);
nand U1204 (N_1204,In_1116,In_1098);
and U1205 (N_1205,In_1351,In_31);
and U1206 (N_1206,In_529,In_932);
nor U1207 (N_1207,In_736,In_1479);
nor U1208 (N_1208,In_219,In_754);
nand U1209 (N_1209,In_1272,In_717);
and U1210 (N_1210,In_1489,In_1467);
nor U1211 (N_1211,In_811,In_884);
or U1212 (N_1212,In_862,In_1195);
or U1213 (N_1213,In_813,In_722);
nand U1214 (N_1214,In_941,In_158);
nor U1215 (N_1215,In_290,In_264);
nand U1216 (N_1216,In_1279,In_1401);
and U1217 (N_1217,In_1091,In_1419);
nor U1218 (N_1218,In_1027,In_93);
and U1219 (N_1219,In_944,In_520);
nor U1220 (N_1220,In_155,In_1434);
nor U1221 (N_1221,In_498,In_1217);
nand U1222 (N_1222,In_1410,In_332);
nor U1223 (N_1223,In_31,In_891);
and U1224 (N_1224,In_591,In_334);
and U1225 (N_1225,In_1231,In_1474);
nor U1226 (N_1226,In_406,In_1345);
nor U1227 (N_1227,In_386,In_680);
nand U1228 (N_1228,In_1290,In_731);
and U1229 (N_1229,In_1387,In_1309);
and U1230 (N_1230,In_1464,In_944);
nor U1231 (N_1231,In_787,In_338);
nand U1232 (N_1232,In_485,In_332);
or U1233 (N_1233,In_1424,In_368);
nor U1234 (N_1234,In_1084,In_750);
or U1235 (N_1235,In_970,In_405);
or U1236 (N_1236,In_208,In_317);
and U1237 (N_1237,In_558,In_571);
nor U1238 (N_1238,In_711,In_334);
or U1239 (N_1239,In_9,In_1345);
nor U1240 (N_1240,In_799,In_304);
or U1241 (N_1241,In_1397,In_157);
nor U1242 (N_1242,In_489,In_1055);
and U1243 (N_1243,In_1269,In_1066);
or U1244 (N_1244,In_306,In_1193);
nand U1245 (N_1245,In_968,In_674);
nor U1246 (N_1246,In_1195,In_1021);
nor U1247 (N_1247,In_312,In_102);
nand U1248 (N_1248,In_1419,In_1388);
nor U1249 (N_1249,In_309,In_741);
and U1250 (N_1250,In_523,In_600);
and U1251 (N_1251,In_879,In_780);
or U1252 (N_1252,In_878,In_1156);
and U1253 (N_1253,In_162,In_1264);
and U1254 (N_1254,In_369,In_1198);
nor U1255 (N_1255,In_1218,In_617);
nand U1256 (N_1256,In_55,In_741);
nor U1257 (N_1257,In_1491,In_1037);
or U1258 (N_1258,In_1415,In_979);
nor U1259 (N_1259,In_192,In_1211);
and U1260 (N_1260,In_1293,In_1280);
nor U1261 (N_1261,In_1436,In_922);
or U1262 (N_1262,In_430,In_170);
and U1263 (N_1263,In_412,In_920);
or U1264 (N_1264,In_1376,In_784);
xnor U1265 (N_1265,In_693,In_1093);
nor U1266 (N_1266,In_592,In_526);
nand U1267 (N_1267,In_95,In_312);
or U1268 (N_1268,In_470,In_15);
or U1269 (N_1269,In_1023,In_829);
or U1270 (N_1270,In_1201,In_1468);
nand U1271 (N_1271,In_1391,In_681);
nor U1272 (N_1272,In_610,In_725);
nor U1273 (N_1273,In_1456,In_313);
and U1274 (N_1274,In_423,In_1276);
or U1275 (N_1275,In_1384,In_751);
nor U1276 (N_1276,In_486,In_1202);
nand U1277 (N_1277,In_458,In_1110);
nand U1278 (N_1278,In_1425,In_101);
nor U1279 (N_1279,In_711,In_229);
nand U1280 (N_1280,In_594,In_1066);
and U1281 (N_1281,In_1375,In_728);
nor U1282 (N_1282,In_710,In_997);
or U1283 (N_1283,In_371,In_765);
and U1284 (N_1284,In_478,In_676);
or U1285 (N_1285,In_517,In_316);
nand U1286 (N_1286,In_1290,In_112);
and U1287 (N_1287,In_694,In_518);
nor U1288 (N_1288,In_266,In_229);
and U1289 (N_1289,In_69,In_1160);
and U1290 (N_1290,In_423,In_318);
nor U1291 (N_1291,In_840,In_804);
nand U1292 (N_1292,In_969,In_1432);
or U1293 (N_1293,In_655,In_947);
or U1294 (N_1294,In_1081,In_203);
nor U1295 (N_1295,In_418,In_166);
or U1296 (N_1296,In_581,In_244);
or U1297 (N_1297,In_1130,In_731);
nor U1298 (N_1298,In_1085,In_832);
or U1299 (N_1299,In_976,In_677);
and U1300 (N_1300,In_1084,In_680);
or U1301 (N_1301,In_876,In_953);
and U1302 (N_1302,In_450,In_1448);
and U1303 (N_1303,In_1123,In_446);
or U1304 (N_1304,In_1478,In_596);
or U1305 (N_1305,In_1288,In_233);
nand U1306 (N_1306,In_1029,In_1235);
and U1307 (N_1307,In_1038,In_1003);
and U1308 (N_1308,In_1151,In_662);
or U1309 (N_1309,In_374,In_574);
nor U1310 (N_1310,In_793,In_1206);
nand U1311 (N_1311,In_1395,In_768);
nand U1312 (N_1312,In_950,In_939);
or U1313 (N_1313,In_1298,In_71);
and U1314 (N_1314,In_373,In_671);
nand U1315 (N_1315,In_886,In_790);
nand U1316 (N_1316,In_240,In_885);
and U1317 (N_1317,In_709,In_232);
nand U1318 (N_1318,In_227,In_148);
and U1319 (N_1319,In_382,In_10);
nand U1320 (N_1320,In_1260,In_662);
nand U1321 (N_1321,In_732,In_462);
nand U1322 (N_1322,In_1461,In_1124);
and U1323 (N_1323,In_1390,In_689);
and U1324 (N_1324,In_494,In_1489);
nor U1325 (N_1325,In_1021,In_1486);
or U1326 (N_1326,In_1436,In_1469);
and U1327 (N_1327,In_280,In_1377);
nor U1328 (N_1328,In_367,In_1092);
or U1329 (N_1329,In_1235,In_1042);
nor U1330 (N_1330,In_1082,In_436);
nor U1331 (N_1331,In_40,In_1412);
nand U1332 (N_1332,In_862,In_39);
xor U1333 (N_1333,In_774,In_770);
nor U1334 (N_1334,In_1104,In_1163);
or U1335 (N_1335,In_1459,In_626);
and U1336 (N_1336,In_745,In_1188);
or U1337 (N_1337,In_458,In_579);
or U1338 (N_1338,In_271,In_1476);
nand U1339 (N_1339,In_979,In_401);
xor U1340 (N_1340,In_3,In_1332);
and U1341 (N_1341,In_65,In_942);
and U1342 (N_1342,In_1452,In_1023);
nor U1343 (N_1343,In_505,In_1027);
or U1344 (N_1344,In_207,In_286);
nand U1345 (N_1345,In_586,In_1100);
and U1346 (N_1346,In_1377,In_476);
and U1347 (N_1347,In_239,In_104);
nor U1348 (N_1348,In_1004,In_1273);
nor U1349 (N_1349,In_737,In_462);
nand U1350 (N_1350,In_729,In_270);
or U1351 (N_1351,In_1444,In_1315);
and U1352 (N_1352,In_796,In_568);
nand U1353 (N_1353,In_1100,In_878);
nand U1354 (N_1354,In_144,In_1312);
nand U1355 (N_1355,In_1137,In_169);
nor U1356 (N_1356,In_667,In_1354);
nor U1357 (N_1357,In_550,In_843);
and U1358 (N_1358,In_75,In_784);
nand U1359 (N_1359,In_26,In_502);
nand U1360 (N_1360,In_428,In_35);
or U1361 (N_1361,In_361,In_48);
nand U1362 (N_1362,In_701,In_1304);
or U1363 (N_1363,In_518,In_902);
nand U1364 (N_1364,In_1469,In_218);
nor U1365 (N_1365,In_985,In_1255);
or U1366 (N_1366,In_152,In_1171);
and U1367 (N_1367,In_436,In_775);
nor U1368 (N_1368,In_158,In_510);
or U1369 (N_1369,In_1312,In_973);
nor U1370 (N_1370,In_692,In_73);
nor U1371 (N_1371,In_1300,In_452);
or U1372 (N_1372,In_288,In_494);
nor U1373 (N_1373,In_271,In_742);
and U1374 (N_1374,In_1348,In_457);
or U1375 (N_1375,In_764,In_863);
or U1376 (N_1376,In_1112,In_459);
and U1377 (N_1377,In_1370,In_423);
nor U1378 (N_1378,In_1258,In_434);
and U1379 (N_1379,In_659,In_787);
nand U1380 (N_1380,In_464,In_28);
nand U1381 (N_1381,In_193,In_1347);
and U1382 (N_1382,In_1001,In_1360);
nand U1383 (N_1383,In_1060,In_748);
and U1384 (N_1384,In_1408,In_242);
or U1385 (N_1385,In_456,In_1412);
nor U1386 (N_1386,In_1112,In_1021);
nor U1387 (N_1387,In_1162,In_1202);
nand U1388 (N_1388,In_890,In_605);
and U1389 (N_1389,In_334,In_1498);
or U1390 (N_1390,In_119,In_824);
or U1391 (N_1391,In_722,In_450);
and U1392 (N_1392,In_1065,In_333);
nand U1393 (N_1393,In_50,In_461);
and U1394 (N_1394,In_508,In_27);
and U1395 (N_1395,In_513,In_329);
or U1396 (N_1396,In_530,In_1176);
or U1397 (N_1397,In_555,In_1224);
nand U1398 (N_1398,In_576,In_358);
nor U1399 (N_1399,In_1334,In_1285);
nor U1400 (N_1400,In_767,In_56);
and U1401 (N_1401,In_830,In_1065);
and U1402 (N_1402,In_1437,In_616);
and U1403 (N_1403,In_1227,In_1331);
nor U1404 (N_1404,In_428,In_1375);
nand U1405 (N_1405,In_766,In_629);
or U1406 (N_1406,In_1168,In_224);
nand U1407 (N_1407,In_724,In_287);
or U1408 (N_1408,In_182,In_675);
or U1409 (N_1409,In_1342,In_295);
nand U1410 (N_1410,In_1106,In_726);
nor U1411 (N_1411,In_343,In_519);
or U1412 (N_1412,In_1365,In_657);
or U1413 (N_1413,In_140,In_493);
and U1414 (N_1414,In_706,In_117);
xor U1415 (N_1415,In_1496,In_369);
nand U1416 (N_1416,In_37,In_1242);
nand U1417 (N_1417,In_1090,In_317);
nand U1418 (N_1418,In_286,In_780);
nand U1419 (N_1419,In_221,In_428);
nand U1420 (N_1420,In_522,In_7);
nand U1421 (N_1421,In_369,In_149);
nand U1422 (N_1422,In_753,In_1414);
nand U1423 (N_1423,In_295,In_674);
or U1424 (N_1424,In_1371,In_660);
nand U1425 (N_1425,In_492,In_910);
or U1426 (N_1426,In_149,In_56);
nand U1427 (N_1427,In_1445,In_257);
nor U1428 (N_1428,In_838,In_1307);
and U1429 (N_1429,In_796,In_319);
and U1430 (N_1430,In_335,In_547);
nand U1431 (N_1431,In_531,In_1027);
nand U1432 (N_1432,In_437,In_1192);
nand U1433 (N_1433,In_933,In_682);
or U1434 (N_1434,In_1069,In_1363);
and U1435 (N_1435,In_9,In_957);
and U1436 (N_1436,In_1206,In_542);
or U1437 (N_1437,In_839,In_826);
or U1438 (N_1438,In_1375,In_590);
and U1439 (N_1439,In_1247,In_1362);
or U1440 (N_1440,In_1428,In_143);
or U1441 (N_1441,In_376,In_919);
nand U1442 (N_1442,In_392,In_166);
nor U1443 (N_1443,In_601,In_515);
nand U1444 (N_1444,In_756,In_541);
nor U1445 (N_1445,In_839,In_454);
nand U1446 (N_1446,In_360,In_718);
and U1447 (N_1447,In_1329,In_405);
nor U1448 (N_1448,In_13,In_825);
nand U1449 (N_1449,In_346,In_774);
nand U1450 (N_1450,In_999,In_275);
or U1451 (N_1451,In_688,In_40);
nor U1452 (N_1452,In_1038,In_660);
xnor U1453 (N_1453,In_219,In_146);
and U1454 (N_1454,In_500,In_930);
and U1455 (N_1455,In_150,In_1025);
nand U1456 (N_1456,In_212,In_922);
and U1457 (N_1457,In_1346,In_595);
or U1458 (N_1458,In_92,In_1343);
nor U1459 (N_1459,In_1100,In_421);
nand U1460 (N_1460,In_649,In_395);
and U1461 (N_1461,In_526,In_594);
or U1462 (N_1462,In_429,In_695);
or U1463 (N_1463,In_1075,In_364);
or U1464 (N_1464,In_470,In_1262);
or U1465 (N_1465,In_622,In_963);
nand U1466 (N_1466,In_1155,In_805);
and U1467 (N_1467,In_741,In_481);
or U1468 (N_1468,In_798,In_1461);
and U1469 (N_1469,In_884,In_1476);
and U1470 (N_1470,In_878,In_42);
and U1471 (N_1471,In_768,In_198);
nand U1472 (N_1472,In_1160,In_298);
or U1473 (N_1473,In_261,In_865);
nor U1474 (N_1474,In_1308,In_950);
nand U1475 (N_1475,In_1318,In_1226);
xnor U1476 (N_1476,In_304,In_893);
xor U1477 (N_1477,In_1102,In_1410);
nor U1478 (N_1478,In_1274,In_625);
nand U1479 (N_1479,In_1126,In_681);
nand U1480 (N_1480,In_797,In_343);
nand U1481 (N_1481,In_346,In_1135);
and U1482 (N_1482,In_241,In_901);
or U1483 (N_1483,In_1187,In_1080);
and U1484 (N_1484,In_154,In_101);
nor U1485 (N_1485,In_731,In_666);
nor U1486 (N_1486,In_555,In_569);
nor U1487 (N_1487,In_1250,In_735);
nand U1488 (N_1488,In_690,In_206);
and U1489 (N_1489,In_1072,In_250);
and U1490 (N_1490,In_1125,In_1196);
nand U1491 (N_1491,In_852,In_1397);
and U1492 (N_1492,In_275,In_1202);
or U1493 (N_1493,In_31,In_958);
or U1494 (N_1494,In_771,In_346);
nand U1495 (N_1495,In_703,In_594);
and U1496 (N_1496,In_713,In_1167);
nor U1497 (N_1497,In_839,In_93);
and U1498 (N_1498,In_1149,In_366);
or U1499 (N_1499,In_950,In_438);
xor U1500 (N_1500,In_1427,In_1073);
or U1501 (N_1501,In_367,In_1083);
or U1502 (N_1502,In_1460,In_26);
or U1503 (N_1503,In_945,In_692);
nor U1504 (N_1504,In_1423,In_897);
nand U1505 (N_1505,In_545,In_721);
nand U1506 (N_1506,In_299,In_802);
or U1507 (N_1507,In_142,In_1114);
and U1508 (N_1508,In_89,In_1070);
nand U1509 (N_1509,In_642,In_100);
nand U1510 (N_1510,In_1137,In_859);
nor U1511 (N_1511,In_449,In_948);
and U1512 (N_1512,In_902,In_346);
nand U1513 (N_1513,In_1105,In_1085);
nor U1514 (N_1514,In_1045,In_912);
or U1515 (N_1515,In_266,In_973);
and U1516 (N_1516,In_831,In_1400);
or U1517 (N_1517,In_454,In_253);
nand U1518 (N_1518,In_502,In_679);
nand U1519 (N_1519,In_175,In_1082);
or U1520 (N_1520,In_738,In_467);
nand U1521 (N_1521,In_798,In_947);
or U1522 (N_1522,In_1321,In_722);
nand U1523 (N_1523,In_846,In_809);
nor U1524 (N_1524,In_1339,In_758);
and U1525 (N_1525,In_1103,In_1012);
and U1526 (N_1526,In_1372,In_919);
or U1527 (N_1527,In_725,In_763);
or U1528 (N_1528,In_267,In_860);
nand U1529 (N_1529,In_482,In_919);
nor U1530 (N_1530,In_1366,In_1338);
or U1531 (N_1531,In_630,In_509);
or U1532 (N_1532,In_535,In_1379);
nand U1533 (N_1533,In_293,In_510);
nand U1534 (N_1534,In_366,In_1036);
and U1535 (N_1535,In_248,In_504);
and U1536 (N_1536,In_1160,In_644);
or U1537 (N_1537,In_474,In_703);
and U1538 (N_1538,In_1103,In_1411);
nand U1539 (N_1539,In_198,In_755);
or U1540 (N_1540,In_1337,In_572);
or U1541 (N_1541,In_314,In_910);
and U1542 (N_1542,In_1414,In_346);
or U1543 (N_1543,In_216,In_669);
nor U1544 (N_1544,In_738,In_515);
nand U1545 (N_1545,In_1090,In_1000);
nor U1546 (N_1546,In_1099,In_630);
nand U1547 (N_1547,In_726,In_87);
nor U1548 (N_1548,In_1210,In_227);
or U1549 (N_1549,In_309,In_383);
and U1550 (N_1550,In_926,In_884);
nand U1551 (N_1551,In_800,In_967);
nand U1552 (N_1552,In_1250,In_1384);
and U1553 (N_1553,In_1458,In_613);
and U1554 (N_1554,In_1366,In_385);
nor U1555 (N_1555,In_653,In_1470);
and U1556 (N_1556,In_1104,In_643);
nand U1557 (N_1557,In_448,In_547);
or U1558 (N_1558,In_336,In_545);
and U1559 (N_1559,In_379,In_1460);
nand U1560 (N_1560,In_50,In_456);
nand U1561 (N_1561,In_1018,In_746);
nor U1562 (N_1562,In_1179,In_624);
or U1563 (N_1563,In_1460,In_1425);
and U1564 (N_1564,In_1296,In_1381);
and U1565 (N_1565,In_568,In_1109);
nor U1566 (N_1566,In_361,In_1348);
or U1567 (N_1567,In_1208,In_31);
nand U1568 (N_1568,In_623,In_610);
and U1569 (N_1569,In_1061,In_164);
nand U1570 (N_1570,In_1062,In_560);
nor U1571 (N_1571,In_694,In_184);
nand U1572 (N_1572,In_413,In_982);
xor U1573 (N_1573,In_1186,In_848);
nand U1574 (N_1574,In_113,In_30);
nand U1575 (N_1575,In_286,In_439);
nand U1576 (N_1576,In_1121,In_1162);
nand U1577 (N_1577,In_95,In_678);
or U1578 (N_1578,In_1178,In_1193);
nand U1579 (N_1579,In_1118,In_1129);
or U1580 (N_1580,In_1456,In_464);
and U1581 (N_1581,In_1043,In_857);
and U1582 (N_1582,In_408,In_1318);
and U1583 (N_1583,In_75,In_673);
xnor U1584 (N_1584,In_1394,In_1072);
nor U1585 (N_1585,In_650,In_319);
or U1586 (N_1586,In_1316,In_960);
nor U1587 (N_1587,In_190,In_722);
and U1588 (N_1588,In_1307,In_637);
nand U1589 (N_1589,In_316,In_1243);
or U1590 (N_1590,In_692,In_527);
nand U1591 (N_1591,In_790,In_437);
and U1592 (N_1592,In_638,In_1003);
nor U1593 (N_1593,In_308,In_382);
or U1594 (N_1594,In_1414,In_1310);
and U1595 (N_1595,In_1293,In_1247);
nand U1596 (N_1596,In_1020,In_541);
nand U1597 (N_1597,In_238,In_163);
nor U1598 (N_1598,In_280,In_705);
or U1599 (N_1599,In_1182,In_630);
xnor U1600 (N_1600,In_1142,In_157);
nand U1601 (N_1601,In_1085,In_440);
nand U1602 (N_1602,In_291,In_530);
or U1603 (N_1603,In_605,In_641);
nor U1604 (N_1604,In_712,In_358);
or U1605 (N_1605,In_621,In_491);
nor U1606 (N_1606,In_410,In_860);
nor U1607 (N_1607,In_1449,In_922);
nand U1608 (N_1608,In_917,In_110);
nand U1609 (N_1609,In_359,In_252);
nand U1610 (N_1610,In_1116,In_874);
and U1611 (N_1611,In_1459,In_5);
nand U1612 (N_1612,In_41,In_781);
or U1613 (N_1613,In_559,In_516);
and U1614 (N_1614,In_773,In_1255);
and U1615 (N_1615,In_175,In_1490);
or U1616 (N_1616,In_346,In_1461);
xnor U1617 (N_1617,In_1089,In_149);
nand U1618 (N_1618,In_1088,In_1126);
xnor U1619 (N_1619,In_1247,In_1183);
nor U1620 (N_1620,In_625,In_1487);
nand U1621 (N_1621,In_1166,In_988);
nor U1622 (N_1622,In_983,In_260);
nor U1623 (N_1623,In_1080,In_1436);
nand U1624 (N_1624,In_1465,In_825);
or U1625 (N_1625,In_231,In_837);
nand U1626 (N_1626,In_103,In_1103);
nor U1627 (N_1627,In_819,In_249);
or U1628 (N_1628,In_1349,In_50);
nor U1629 (N_1629,In_113,In_164);
or U1630 (N_1630,In_1382,In_1252);
and U1631 (N_1631,In_18,In_733);
or U1632 (N_1632,In_156,In_703);
nor U1633 (N_1633,In_93,In_599);
or U1634 (N_1634,In_554,In_553);
and U1635 (N_1635,In_694,In_726);
nand U1636 (N_1636,In_185,In_70);
nand U1637 (N_1637,In_1392,In_338);
nand U1638 (N_1638,In_1265,In_1156);
nand U1639 (N_1639,In_1427,In_321);
and U1640 (N_1640,In_453,In_305);
or U1641 (N_1641,In_1169,In_734);
nand U1642 (N_1642,In_955,In_144);
and U1643 (N_1643,In_901,In_919);
and U1644 (N_1644,In_682,In_263);
nor U1645 (N_1645,In_283,In_1261);
nor U1646 (N_1646,In_1456,In_1059);
nand U1647 (N_1647,In_875,In_351);
nor U1648 (N_1648,In_827,In_30);
or U1649 (N_1649,In_528,In_1499);
nor U1650 (N_1650,In_1341,In_1129);
and U1651 (N_1651,In_683,In_1383);
or U1652 (N_1652,In_1369,In_143);
xor U1653 (N_1653,In_362,In_953);
or U1654 (N_1654,In_549,In_1273);
or U1655 (N_1655,In_273,In_198);
or U1656 (N_1656,In_412,In_945);
and U1657 (N_1657,In_931,In_830);
nor U1658 (N_1658,In_832,In_1375);
or U1659 (N_1659,In_895,In_535);
nand U1660 (N_1660,In_199,In_9);
nor U1661 (N_1661,In_1200,In_71);
nor U1662 (N_1662,In_715,In_757);
and U1663 (N_1663,In_730,In_1495);
nand U1664 (N_1664,In_138,In_381);
or U1665 (N_1665,In_1000,In_170);
and U1666 (N_1666,In_474,In_831);
nor U1667 (N_1667,In_290,In_1453);
nand U1668 (N_1668,In_422,In_788);
or U1669 (N_1669,In_324,In_162);
nand U1670 (N_1670,In_490,In_1428);
and U1671 (N_1671,In_235,In_466);
nand U1672 (N_1672,In_74,In_1406);
or U1673 (N_1673,In_1207,In_1124);
nor U1674 (N_1674,In_568,In_520);
or U1675 (N_1675,In_141,In_1075);
and U1676 (N_1676,In_558,In_1426);
or U1677 (N_1677,In_862,In_610);
nor U1678 (N_1678,In_1076,In_751);
nand U1679 (N_1679,In_251,In_913);
or U1680 (N_1680,In_879,In_553);
or U1681 (N_1681,In_1427,In_115);
nand U1682 (N_1682,In_147,In_1291);
nor U1683 (N_1683,In_68,In_298);
nor U1684 (N_1684,In_611,In_4);
nand U1685 (N_1685,In_517,In_1);
or U1686 (N_1686,In_138,In_5);
nor U1687 (N_1687,In_1496,In_1102);
nand U1688 (N_1688,In_239,In_992);
nand U1689 (N_1689,In_943,In_1003);
nand U1690 (N_1690,In_1090,In_674);
nor U1691 (N_1691,In_1241,In_227);
nand U1692 (N_1692,In_97,In_1433);
nand U1693 (N_1693,In_603,In_240);
nand U1694 (N_1694,In_1298,In_477);
nand U1695 (N_1695,In_877,In_93);
or U1696 (N_1696,In_1113,In_600);
xor U1697 (N_1697,In_166,In_924);
nand U1698 (N_1698,In_100,In_1194);
nor U1699 (N_1699,In_315,In_320);
and U1700 (N_1700,In_1084,In_1404);
nor U1701 (N_1701,In_823,In_1349);
nand U1702 (N_1702,In_1439,In_131);
and U1703 (N_1703,In_158,In_792);
or U1704 (N_1704,In_1034,In_306);
nand U1705 (N_1705,In_948,In_1024);
xnor U1706 (N_1706,In_856,In_1286);
and U1707 (N_1707,In_1158,In_1388);
and U1708 (N_1708,In_1486,In_127);
and U1709 (N_1709,In_409,In_1174);
nor U1710 (N_1710,In_344,In_430);
and U1711 (N_1711,In_258,In_1423);
nor U1712 (N_1712,In_252,In_1173);
nand U1713 (N_1713,In_44,In_1198);
nand U1714 (N_1714,In_558,In_1025);
nand U1715 (N_1715,In_1474,In_379);
nand U1716 (N_1716,In_490,In_144);
xor U1717 (N_1717,In_1008,In_284);
nand U1718 (N_1718,In_1054,In_2);
or U1719 (N_1719,In_901,In_640);
and U1720 (N_1720,In_1269,In_1195);
nor U1721 (N_1721,In_1290,In_921);
or U1722 (N_1722,In_1342,In_1061);
nand U1723 (N_1723,In_784,In_1006);
or U1724 (N_1724,In_548,In_362);
nand U1725 (N_1725,In_314,In_1202);
and U1726 (N_1726,In_1375,In_18);
or U1727 (N_1727,In_194,In_1280);
nand U1728 (N_1728,In_317,In_354);
or U1729 (N_1729,In_564,In_197);
or U1730 (N_1730,In_826,In_211);
or U1731 (N_1731,In_260,In_677);
or U1732 (N_1732,In_46,In_549);
nand U1733 (N_1733,In_762,In_749);
and U1734 (N_1734,In_1325,In_115);
nand U1735 (N_1735,In_414,In_1002);
nand U1736 (N_1736,In_1241,In_1336);
nand U1737 (N_1737,In_473,In_1233);
nor U1738 (N_1738,In_1088,In_1273);
nor U1739 (N_1739,In_823,In_1162);
or U1740 (N_1740,In_491,In_12);
nand U1741 (N_1741,In_746,In_1170);
nor U1742 (N_1742,In_1473,In_1015);
nand U1743 (N_1743,In_332,In_710);
nand U1744 (N_1744,In_568,In_1100);
nor U1745 (N_1745,In_1234,In_930);
and U1746 (N_1746,In_485,In_1025);
nor U1747 (N_1747,In_1076,In_756);
nand U1748 (N_1748,In_323,In_318);
nor U1749 (N_1749,In_856,In_887);
nor U1750 (N_1750,In_102,In_1090);
or U1751 (N_1751,In_1492,In_628);
nor U1752 (N_1752,In_464,In_1187);
nor U1753 (N_1753,In_1033,In_52);
and U1754 (N_1754,In_105,In_457);
nor U1755 (N_1755,In_136,In_1150);
and U1756 (N_1756,In_1474,In_220);
nor U1757 (N_1757,In_108,In_993);
or U1758 (N_1758,In_370,In_1353);
or U1759 (N_1759,In_94,In_581);
nor U1760 (N_1760,In_1083,In_887);
nand U1761 (N_1761,In_644,In_1104);
nor U1762 (N_1762,In_955,In_1484);
nor U1763 (N_1763,In_1297,In_831);
nor U1764 (N_1764,In_931,In_461);
or U1765 (N_1765,In_261,In_395);
or U1766 (N_1766,In_475,In_909);
nor U1767 (N_1767,In_638,In_547);
and U1768 (N_1768,In_1396,In_92);
nand U1769 (N_1769,In_441,In_983);
or U1770 (N_1770,In_606,In_441);
and U1771 (N_1771,In_547,In_257);
and U1772 (N_1772,In_499,In_609);
and U1773 (N_1773,In_1250,In_782);
xnor U1774 (N_1774,In_1137,In_1207);
and U1775 (N_1775,In_784,In_972);
xor U1776 (N_1776,In_261,In_576);
or U1777 (N_1777,In_1114,In_1446);
and U1778 (N_1778,In_989,In_60);
or U1779 (N_1779,In_1376,In_1311);
nor U1780 (N_1780,In_265,In_1431);
or U1781 (N_1781,In_794,In_1025);
or U1782 (N_1782,In_420,In_791);
or U1783 (N_1783,In_1321,In_965);
and U1784 (N_1784,In_418,In_91);
and U1785 (N_1785,In_1306,In_552);
nand U1786 (N_1786,In_546,In_1475);
or U1787 (N_1787,In_1176,In_1094);
or U1788 (N_1788,In_434,In_256);
nor U1789 (N_1789,In_672,In_895);
and U1790 (N_1790,In_367,In_225);
and U1791 (N_1791,In_187,In_758);
and U1792 (N_1792,In_163,In_309);
or U1793 (N_1793,In_975,In_327);
and U1794 (N_1794,In_467,In_1011);
nand U1795 (N_1795,In_1370,In_1006);
or U1796 (N_1796,In_78,In_1188);
nand U1797 (N_1797,In_1459,In_412);
nor U1798 (N_1798,In_1305,In_1130);
nor U1799 (N_1799,In_402,In_533);
nand U1800 (N_1800,In_254,In_1032);
and U1801 (N_1801,In_1160,In_386);
nand U1802 (N_1802,In_286,In_119);
and U1803 (N_1803,In_1353,In_313);
nand U1804 (N_1804,In_1289,In_1152);
or U1805 (N_1805,In_140,In_1341);
nor U1806 (N_1806,In_1152,In_72);
or U1807 (N_1807,In_913,In_626);
nor U1808 (N_1808,In_44,In_773);
and U1809 (N_1809,In_616,In_1475);
xnor U1810 (N_1810,In_981,In_5);
nor U1811 (N_1811,In_1246,In_115);
nor U1812 (N_1812,In_168,In_629);
nand U1813 (N_1813,In_275,In_284);
and U1814 (N_1814,In_246,In_427);
or U1815 (N_1815,In_960,In_923);
or U1816 (N_1816,In_1295,In_521);
and U1817 (N_1817,In_785,In_521);
or U1818 (N_1818,In_837,In_82);
nand U1819 (N_1819,In_233,In_1354);
or U1820 (N_1820,In_1397,In_855);
or U1821 (N_1821,In_11,In_1425);
and U1822 (N_1822,In_230,In_775);
nor U1823 (N_1823,In_1251,In_1389);
and U1824 (N_1824,In_347,In_595);
and U1825 (N_1825,In_129,In_922);
nand U1826 (N_1826,In_187,In_97);
nand U1827 (N_1827,In_976,In_1040);
and U1828 (N_1828,In_1369,In_642);
nor U1829 (N_1829,In_1179,In_514);
nor U1830 (N_1830,In_447,In_385);
nand U1831 (N_1831,In_965,In_792);
and U1832 (N_1832,In_319,In_663);
nor U1833 (N_1833,In_1237,In_430);
nor U1834 (N_1834,In_792,In_1071);
and U1835 (N_1835,In_435,In_1010);
xor U1836 (N_1836,In_248,In_786);
nor U1837 (N_1837,In_650,In_231);
and U1838 (N_1838,In_1224,In_106);
nand U1839 (N_1839,In_203,In_1360);
or U1840 (N_1840,In_457,In_771);
nand U1841 (N_1841,In_606,In_1400);
nand U1842 (N_1842,In_15,In_881);
nor U1843 (N_1843,In_690,In_624);
or U1844 (N_1844,In_421,In_1139);
and U1845 (N_1845,In_323,In_41);
nand U1846 (N_1846,In_887,In_437);
or U1847 (N_1847,In_459,In_525);
and U1848 (N_1848,In_805,In_229);
or U1849 (N_1849,In_1438,In_776);
or U1850 (N_1850,In_1396,In_564);
nor U1851 (N_1851,In_1454,In_556);
nor U1852 (N_1852,In_755,In_1445);
nand U1853 (N_1853,In_872,In_1046);
nor U1854 (N_1854,In_651,In_1077);
nor U1855 (N_1855,In_629,In_900);
and U1856 (N_1856,In_1263,In_1118);
or U1857 (N_1857,In_1481,In_1378);
and U1858 (N_1858,In_147,In_1357);
and U1859 (N_1859,In_1188,In_1091);
nor U1860 (N_1860,In_547,In_969);
nand U1861 (N_1861,In_446,In_373);
nand U1862 (N_1862,In_986,In_381);
nor U1863 (N_1863,In_869,In_619);
nand U1864 (N_1864,In_936,In_455);
nor U1865 (N_1865,In_334,In_379);
nand U1866 (N_1866,In_107,In_1395);
nor U1867 (N_1867,In_1183,In_1491);
and U1868 (N_1868,In_917,In_170);
and U1869 (N_1869,In_1034,In_699);
nand U1870 (N_1870,In_105,In_350);
nor U1871 (N_1871,In_927,In_1228);
and U1872 (N_1872,In_464,In_195);
nor U1873 (N_1873,In_177,In_638);
nand U1874 (N_1874,In_1422,In_294);
and U1875 (N_1875,In_122,In_1405);
nand U1876 (N_1876,In_625,In_3);
xor U1877 (N_1877,In_1427,In_259);
nand U1878 (N_1878,In_268,In_588);
nor U1879 (N_1879,In_1402,In_1191);
nor U1880 (N_1880,In_1090,In_1320);
nand U1881 (N_1881,In_407,In_736);
or U1882 (N_1882,In_839,In_1247);
or U1883 (N_1883,In_1487,In_773);
or U1884 (N_1884,In_725,In_1064);
or U1885 (N_1885,In_890,In_1432);
and U1886 (N_1886,In_611,In_1032);
nand U1887 (N_1887,In_661,In_271);
or U1888 (N_1888,In_1470,In_888);
nor U1889 (N_1889,In_23,In_194);
and U1890 (N_1890,In_204,In_1084);
nand U1891 (N_1891,In_1182,In_1122);
xnor U1892 (N_1892,In_1388,In_1329);
and U1893 (N_1893,In_1121,In_306);
or U1894 (N_1894,In_1386,In_1210);
nor U1895 (N_1895,In_174,In_393);
nor U1896 (N_1896,In_1247,In_758);
or U1897 (N_1897,In_771,In_813);
nand U1898 (N_1898,In_896,In_1406);
and U1899 (N_1899,In_783,In_1002);
nand U1900 (N_1900,In_104,In_1179);
nand U1901 (N_1901,In_362,In_732);
nand U1902 (N_1902,In_673,In_419);
and U1903 (N_1903,In_583,In_33);
nand U1904 (N_1904,In_1015,In_625);
and U1905 (N_1905,In_989,In_1431);
xnor U1906 (N_1906,In_1159,In_1428);
nand U1907 (N_1907,In_1147,In_714);
or U1908 (N_1908,In_1012,In_485);
nor U1909 (N_1909,In_1006,In_44);
or U1910 (N_1910,In_783,In_1301);
and U1911 (N_1911,In_726,In_1022);
and U1912 (N_1912,In_660,In_236);
and U1913 (N_1913,In_811,In_1458);
and U1914 (N_1914,In_987,In_230);
nor U1915 (N_1915,In_623,In_699);
or U1916 (N_1916,In_1365,In_1206);
nor U1917 (N_1917,In_1413,In_1205);
nor U1918 (N_1918,In_1361,In_299);
nor U1919 (N_1919,In_883,In_320);
nand U1920 (N_1920,In_1250,In_859);
or U1921 (N_1921,In_266,In_888);
nand U1922 (N_1922,In_976,In_883);
and U1923 (N_1923,In_863,In_394);
and U1924 (N_1924,In_590,In_419);
and U1925 (N_1925,In_458,In_1193);
or U1926 (N_1926,In_1288,In_1362);
or U1927 (N_1927,In_971,In_1220);
or U1928 (N_1928,In_249,In_3);
or U1929 (N_1929,In_39,In_82);
and U1930 (N_1930,In_802,In_1214);
and U1931 (N_1931,In_630,In_456);
nor U1932 (N_1932,In_1404,In_775);
nor U1933 (N_1933,In_804,In_897);
and U1934 (N_1934,In_342,In_64);
and U1935 (N_1935,In_514,In_882);
nor U1936 (N_1936,In_1433,In_406);
or U1937 (N_1937,In_1025,In_1148);
nor U1938 (N_1938,In_351,In_1045);
nor U1939 (N_1939,In_287,In_1319);
and U1940 (N_1940,In_53,In_961);
nand U1941 (N_1941,In_79,In_1006);
nor U1942 (N_1942,In_1165,In_1425);
nand U1943 (N_1943,In_1172,In_598);
nand U1944 (N_1944,In_283,In_1382);
nand U1945 (N_1945,In_172,In_1210);
nand U1946 (N_1946,In_1458,In_889);
nand U1947 (N_1947,In_987,In_707);
nor U1948 (N_1948,In_1158,In_1035);
nor U1949 (N_1949,In_705,In_304);
nor U1950 (N_1950,In_1047,In_325);
nand U1951 (N_1951,In_1174,In_702);
xor U1952 (N_1952,In_68,In_1158);
nor U1953 (N_1953,In_1156,In_288);
nor U1954 (N_1954,In_461,In_1337);
or U1955 (N_1955,In_831,In_693);
nand U1956 (N_1956,In_840,In_215);
nand U1957 (N_1957,In_1168,In_258);
nand U1958 (N_1958,In_622,In_902);
or U1959 (N_1959,In_718,In_195);
or U1960 (N_1960,In_60,In_133);
or U1961 (N_1961,In_985,In_98);
and U1962 (N_1962,In_464,In_796);
nor U1963 (N_1963,In_506,In_294);
nand U1964 (N_1964,In_1110,In_691);
or U1965 (N_1965,In_288,In_1121);
nor U1966 (N_1966,In_908,In_291);
and U1967 (N_1967,In_877,In_427);
xnor U1968 (N_1968,In_998,In_1369);
nand U1969 (N_1969,In_1483,In_612);
nand U1970 (N_1970,In_1248,In_842);
nor U1971 (N_1971,In_373,In_246);
nand U1972 (N_1972,In_567,In_1253);
or U1973 (N_1973,In_39,In_1124);
or U1974 (N_1974,In_388,In_1262);
or U1975 (N_1975,In_477,In_1110);
nand U1976 (N_1976,In_445,In_1101);
and U1977 (N_1977,In_279,In_1399);
nand U1978 (N_1978,In_126,In_1017);
nand U1979 (N_1979,In_171,In_1319);
nor U1980 (N_1980,In_1015,In_1341);
and U1981 (N_1981,In_1207,In_1231);
nor U1982 (N_1982,In_950,In_870);
and U1983 (N_1983,In_333,In_947);
and U1984 (N_1984,In_1040,In_231);
and U1985 (N_1985,In_1129,In_579);
or U1986 (N_1986,In_597,In_31);
nand U1987 (N_1987,In_80,In_117);
nor U1988 (N_1988,In_1482,In_324);
nand U1989 (N_1989,In_1087,In_164);
or U1990 (N_1990,In_120,In_1004);
nand U1991 (N_1991,In_1216,In_690);
nor U1992 (N_1992,In_1123,In_1121);
nor U1993 (N_1993,In_167,In_615);
nor U1994 (N_1994,In_554,In_1190);
or U1995 (N_1995,In_385,In_1383);
nor U1996 (N_1996,In_985,In_1026);
nand U1997 (N_1997,In_845,In_165);
and U1998 (N_1998,In_24,In_151);
nand U1999 (N_1999,In_428,In_695);
nand U2000 (N_2000,In_1068,In_939);
and U2001 (N_2001,In_289,In_647);
or U2002 (N_2002,In_29,In_196);
nand U2003 (N_2003,In_131,In_689);
nand U2004 (N_2004,In_577,In_76);
or U2005 (N_2005,In_1256,In_506);
and U2006 (N_2006,In_245,In_149);
and U2007 (N_2007,In_613,In_810);
nand U2008 (N_2008,In_1191,In_281);
and U2009 (N_2009,In_60,In_1386);
nand U2010 (N_2010,In_391,In_297);
or U2011 (N_2011,In_297,In_87);
or U2012 (N_2012,In_848,In_1388);
or U2013 (N_2013,In_1429,In_142);
and U2014 (N_2014,In_51,In_677);
nor U2015 (N_2015,In_1013,In_347);
nand U2016 (N_2016,In_1497,In_826);
and U2017 (N_2017,In_543,In_1239);
nand U2018 (N_2018,In_260,In_1349);
nand U2019 (N_2019,In_477,In_1255);
or U2020 (N_2020,In_1365,In_133);
and U2021 (N_2021,In_890,In_939);
and U2022 (N_2022,In_229,In_262);
or U2023 (N_2023,In_287,In_806);
or U2024 (N_2024,In_1448,In_401);
or U2025 (N_2025,In_914,In_1318);
nor U2026 (N_2026,In_223,In_740);
and U2027 (N_2027,In_1359,In_461);
nor U2028 (N_2028,In_917,In_1244);
nand U2029 (N_2029,In_602,In_231);
and U2030 (N_2030,In_1143,In_300);
xnor U2031 (N_2031,In_1068,In_1351);
xor U2032 (N_2032,In_859,In_1185);
nor U2033 (N_2033,In_1003,In_764);
xor U2034 (N_2034,In_134,In_669);
and U2035 (N_2035,In_606,In_533);
or U2036 (N_2036,In_371,In_1079);
nand U2037 (N_2037,In_560,In_39);
or U2038 (N_2038,In_1005,In_1211);
nor U2039 (N_2039,In_401,In_477);
nand U2040 (N_2040,In_21,In_951);
nor U2041 (N_2041,In_532,In_317);
nand U2042 (N_2042,In_254,In_701);
and U2043 (N_2043,In_773,In_1169);
and U2044 (N_2044,In_1394,In_1015);
nor U2045 (N_2045,In_850,In_27);
nor U2046 (N_2046,In_798,In_1199);
and U2047 (N_2047,In_267,In_1320);
nor U2048 (N_2048,In_39,In_806);
or U2049 (N_2049,In_506,In_1307);
nor U2050 (N_2050,In_1461,In_141);
or U2051 (N_2051,In_971,In_1309);
nor U2052 (N_2052,In_408,In_1327);
and U2053 (N_2053,In_1321,In_664);
xnor U2054 (N_2054,In_312,In_1235);
nor U2055 (N_2055,In_1093,In_1101);
or U2056 (N_2056,In_653,In_1201);
nor U2057 (N_2057,In_1473,In_1220);
nor U2058 (N_2058,In_752,In_1330);
nor U2059 (N_2059,In_732,In_1407);
nor U2060 (N_2060,In_928,In_1140);
and U2061 (N_2061,In_1371,In_1266);
or U2062 (N_2062,In_729,In_845);
nand U2063 (N_2063,In_157,In_933);
nand U2064 (N_2064,In_715,In_1429);
or U2065 (N_2065,In_723,In_344);
and U2066 (N_2066,In_69,In_1201);
and U2067 (N_2067,In_740,In_124);
and U2068 (N_2068,In_1156,In_421);
and U2069 (N_2069,In_1442,In_992);
nor U2070 (N_2070,In_1059,In_915);
nor U2071 (N_2071,In_596,In_229);
nand U2072 (N_2072,In_1030,In_762);
nand U2073 (N_2073,In_779,In_1356);
nand U2074 (N_2074,In_642,In_596);
nand U2075 (N_2075,In_821,In_1119);
nand U2076 (N_2076,In_950,In_1362);
or U2077 (N_2077,In_383,In_1163);
nand U2078 (N_2078,In_382,In_142);
and U2079 (N_2079,In_946,In_1426);
nor U2080 (N_2080,In_189,In_1198);
nor U2081 (N_2081,In_184,In_739);
and U2082 (N_2082,In_245,In_1367);
nand U2083 (N_2083,In_405,In_1433);
nand U2084 (N_2084,In_404,In_446);
and U2085 (N_2085,In_1128,In_841);
and U2086 (N_2086,In_569,In_57);
and U2087 (N_2087,In_957,In_886);
nor U2088 (N_2088,In_199,In_197);
nor U2089 (N_2089,In_1280,In_764);
or U2090 (N_2090,In_509,In_1261);
nand U2091 (N_2091,In_344,In_673);
nand U2092 (N_2092,In_1484,In_397);
nor U2093 (N_2093,In_561,In_1152);
nor U2094 (N_2094,In_275,In_447);
and U2095 (N_2095,In_695,In_1070);
and U2096 (N_2096,In_585,In_339);
or U2097 (N_2097,In_638,In_15);
nor U2098 (N_2098,In_842,In_834);
nor U2099 (N_2099,In_1494,In_783);
nand U2100 (N_2100,In_559,In_924);
nor U2101 (N_2101,In_662,In_702);
or U2102 (N_2102,In_888,In_46);
nor U2103 (N_2103,In_739,In_1466);
or U2104 (N_2104,In_1148,In_1376);
nand U2105 (N_2105,In_566,In_482);
or U2106 (N_2106,In_560,In_54);
or U2107 (N_2107,In_681,In_611);
nand U2108 (N_2108,In_1105,In_1132);
nand U2109 (N_2109,In_1456,In_1179);
xnor U2110 (N_2110,In_773,In_122);
or U2111 (N_2111,In_1363,In_418);
nor U2112 (N_2112,In_258,In_923);
and U2113 (N_2113,In_89,In_1307);
nor U2114 (N_2114,In_541,In_1192);
nand U2115 (N_2115,In_862,In_1490);
or U2116 (N_2116,In_498,In_1409);
nor U2117 (N_2117,In_831,In_1368);
nand U2118 (N_2118,In_1342,In_367);
nor U2119 (N_2119,In_1281,In_1400);
nand U2120 (N_2120,In_1242,In_258);
or U2121 (N_2121,In_771,In_1396);
xnor U2122 (N_2122,In_1153,In_61);
or U2123 (N_2123,In_410,In_563);
and U2124 (N_2124,In_665,In_683);
nand U2125 (N_2125,In_1032,In_245);
nor U2126 (N_2126,In_350,In_540);
and U2127 (N_2127,In_786,In_450);
nor U2128 (N_2128,In_1131,In_1014);
nor U2129 (N_2129,In_383,In_40);
and U2130 (N_2130,In_0,In_990);
nor U2131 (N_2131,In_154,In_1254);
and U2132 (N_2132,In_1032,In_1290);
or U2133 (N_2133,In_574,In_78);
and U2134 (N_2134,In_470,In_1166);
nand U2135 (N_2135,In_1462,In_667);
nor U2136 (N_2136,In_1425,In_1341);
and U2137 (N_2137,In_1173,In_1458);
or U2138 (N_2138,In_1410,In_945);
or U2139 (N_2139,In_70,In_1373);
nand U2140 (N_2140,In_823,In_1145);
nand U2141 (N_2141,In_1421,In_128);
nand U2142 (N_2142,In_947,In_172);
and U2143 (N_2143,In_118,In_1241);
nor U2144 (N_2144,In_684,In_370);
nand U2145 (N_2145,In_129,In_1082);
and U2146 (N_2146,In_423,In_894);
nor U2147 (N_2147,In_752,In_1383);
nand U2148 (N_2148,In_834,In_569);
and U2149 (N_2149,In_1377,In_848);
and U2150 (N_2150,In_242,In_854);
nand U2151 (N_2151,In_1449,In_1206);
or U2152 (N_2152,In_509,In_23);
nor U2153 (N_2153,In_951,In_602);
and U2154 (N_2154,In_928,In_1476);
and U2155 (N_2155,In_932,In_1419);
or U2156 (N_2156,In_79,In_258);
nand U2157 (N_2157,In_1094,In_90);
and U2158 (N_2158,In_808,In_178);
nand U2159 (N_2159,In_480,In_184);
or U2160 (N_2160,In_1164,In_388);
nand U2161 (N_2161,In_1375,In_1180);
and U2162 (N_2162,In_56,In_849);
or U2163 (N_2163,In_787,In_1242);
nand U2164 (N_2164,In_593,In_471);
nor U2165 (N_2165,In_1298,In_1291);
or U2166 (N_2166,In_1068,In_1105);
nor U2167 (N_2167,In_1318,In_30);
or U2168 (N_2168,In_113,In_1101);
or U2169 (N_2169,In_932,In_1444);
nand U2170 (N_2170,In_1038,In_92);
or U2171 (N_2171,In_863,In_607);
nor U2172 (N_2172,In_1342,In_725);
or U2173 (N_2173,In_685,In_22);
nor U2174 (N_2174,In_159,In_370);
or U2175 (N_2175,In_984,In_1285);
or U2176 (N_2176,In_245,In_1214);
nand U2177 (N_2177,In_1142,In_35);
nand U2178 (N_2178,In_679,In_345);
nand U2179 (N_2179,In_676,In_627);
nand U2180 (N_2180,In_407,In_379);
nand U2181 (N_2181,In_20,In_1304);
and U2182 (N_2182,In_1030,In_1394);
xor U2183 (N_2183,In_366,In_681);
nor U2184 (N_2184,In_1234,In_439);
or U2185 (N_2185,In_1353,In_389);
nor U2186 (N_2186,In_675,In_155);
or U2187 (N_2187,In_510,In_1046);
or U2188 (N_2188,In_984,In_1421);
nor U2189 (N_2189,In_1354,In_1329);
and U2190 (N_2190,In_898,In_1354);
nand U2191 (N_2191,In_53,In_806);
nand U2192 (N_2192,In_1402,In_358);
and U2193 (N_2193,In_555,In_647);
or U2194 (N_2194,In_370,In_1472);
and U2195 (N_2195,In_555,In_914);
nand U2196 (N_2196,In_793,In_1306);
or U2197 (N_2197,In_444,In_345);
nand U2198 (N_2198,In_477,In_1353);
or U2199 (N_2199,In_174,In_1293);
nand U2200 (N_2200,In_802,In_952);
and U2201 (N_2201,In_1025,In_88);
nor U2202 (N_2202,In_1162,In_1408);
or U2203 (N_2203,In_134,In_970);
nor U2204 (N_2204,In_716,In_27);
and U2205 (N_2205,In_1051,In_515);
xor U2206 (N_2206,In_597,In_740);
and U2207 (N_2207,In_1293,In_485);
nand U2208 (N_2208,In_507,In_659);
and U2209 (N_2209,In_551,In_232);
nor U2210 (N_2210,In_409,In_885);
or U2211 (N_2211,In_1278,In_1315);
xor U2212 (N_2212,In_994,In_1171);
nand U2213 (N_2213,In_1381,In_291);
nand U2214 (N_2214,In_823,In_1365);
and U2215 (N_2215,In_448,In_469);
and U2216 (N_2216,In_515,In_574);
nand U2217 (N_2217,In_1061,In_370);
nand U2218 (N_2218,In_373,In_1130);
and U2219 (N_2219,In_383,In_161);
and U2220 (N_2220,In_1336,In_912);
nand U2221 (N_2221,In_371,In_1482);
or U2222 (N_2222,In_913,In_56);
and U2223 (N_2223,In_1405,In_1495);
nand U2224 (N_2224,In_143,In_2);
nor U2225 (N_2225,In_900,In_923);
or U2226 (N_2226,In_275,In_1489);
and U2227 (N_2227,In_22,In_1315);
and U2228 (N_2228,In_179,In_747);
nor U2229 (N_2229,In_1294,In_1425);
nand U2230 (N_2230,In_1347,In_135);
and U2231 (N_2231,In_727,In_99);
and U2232 (N_2232,In_1480,In_1008);
or U2233 (N_2233,In_239,In_741);
or U2234 (N_2234,In_84,In_681);
nor U2235 (N_2235,In_1012,In_295);
nor U2236 (N_2236,In_752,In_971);
nor U2237 (N_2237,In_982,In_406);
and U2238 (N_2238,In_899,In_290);
nor U2239 (N_2239,In_856,In_1405);
or U2240 (N_2240,In_1496,In_457);
nand U2241 (N_2241,In_634,In_64);
nand U2242 (N_2242,In_956,In_1146);
nor U2243 (N_2243,In_584,In_1286);
and U2244 (N_2244,In_440,In_683);
nor U2245 (N_2245,In_903,In_60);
nor U2246 (N_2246,In_1073,In_1200);
nand U2247 (N_2247,In_696,In_481);
nand U2248 (N_2248,In_395,In_669);
nand U2249 (N_2249,In_1373,In_333);
nor U2250 (N_2250,In_710,In_627);
and U2251 (N_2251,In_857,In_612);
and U2252 (N_2252,In_577,In_465);
and U2253 (N_2253,In_1149,In_1186);
nand U2254 (N_2254,In_618,In_312);
nand U2255 (N_2255,In_586,In_745);
or U2256 (N_2256,In_867,In_194);
nand U2257 (N_2257,In_1224,In_411);
nand U2258 (N_2258,In_1233,In_1250);
or U2259 (N_2259,In_338,In_1057);
or U2260 (N_2260,In_778,In_331);
nand U2261 (N_2261,In_595,In_1466);
or U2262 (N_2262,In_605,In_590);
nand U2263 (N_2263,In_1166,In_57);
and U2264 (N_2264,In_364,In_1282);
nand U2265 (N_2265,In_742,In_497);
nand U2266 (N_2266,In_1219,In_1134);
nand U2267 (N_2267,In_909,In_1419);
nor U2268 (N_2268,In_1278,In_465);
or U2269 (N_2269,In_1144,In_278);
nor U2270 (N_2270,In_909,In_1330);
nor U2271 (N_2271,In_1348,In_1362);
or U2272 (N_2272,In_138,In_584);
nor U2273 (N_2273,In_631,In_439);
xnor U2274 (N_2274,In_1394,In_222);
and U2275 (N_2275,In_1105,In_1095);
and U2276 (N_2276,In_26,In_1365);
xor U2277 (N_2277,In_691,In_144);
nand U2278 (N_2278,In_1022,In_569);
nor U2279 (N_2279,In_254,In_460);
xor U2280 (N_2280,In_1070,In_340);
nor U2281 (N_2281,In_1109,In_1000);
nand U2282 (N_2282,In_891,In_273);
or U2283 (N_2283,In_565,In_1204);
nand U2284 (N_2284,In_1433,In_607);
nor U2285 (N_2285,In_1156,In_616);
nand U2286 (N_2286,In_1072,In_932);
nor U2287 (N_2287,In_206,In_922);
and U2288 (N_2288,In_428,In_917);
nand U2289 (N_2289,In_656,In_850);
and U2290 (N_2290,In_53,In_399);
nand U2291 (N_2291,In_211,In_1462);
nand U2292 (N_2292,In_1070,In_331);
and U2293 (N_2293,In_443,In_23);
nor U2294 (N_2294,In_1285,In_462);
nand U2295 (N_2295,In_37,In_1394);
or U2296 (N_2296,In_893,In_632);
or U2297 (N_2297,In_1471,In_661);
nor U2298 (N_2298,In_951,In_1326);
and U2299 (N_2299,In_385,In_1081);
nand U2300 (N_2300,In_727,In_966);
and U2301 (N_2301,In_230,In_300);
and U2302 (N_2302,In_481,In_1499);
or U2303 (N_2303,In_1267,In_205);
and U2304 (N_2304,In_409,In_1025);
or U2305 (N_2305,In_642,In_675);
and U2306 (N_2306,In_531,In_995);
nor U2307 (N_2307,In_1349,In_289);
and U2308 (N_2308,In_990,In_384);
nor U2309 (N_2309,In_149,In_1419);
and U2310 (N_2310,In_993,In_911);
and U2311 (N_2311,In_248,In_1118);
and U2312 (N_2312,In_25,In_1355);
nor U2313 (N_2313,In_537,In_1008);
nor U2314 (N_2314,In_386,In_1197);
or U2315 (N_2315,In_387,In_1123);
nor U2316 (N_2316,In_1096,In_526);
and U2317 (N_2317,In_580,In_662);
nor U2318 (N_2318,In_1416,In_579);
or U2319 (N_2319,In_33,In_1221);
and U2320 (N_2320,In_153,In_748);
or U2321 (N_2321,In_1326,In_1164);
and U2322 (N_2322,In_109,In_166);
or U2323 (N_2323,In_310,In_1152);
and U2324 (N_2324,In_180,In_1070);
or U2325 (N_2325,In_1390,In_1356);
nand U2326 (N_2326,In_1293,In_754);
nand U2327 (N_2327,In_350,In_311);
nand U2328 (N_2328,In_974,In_224);
or U2329 (N_2329,In_1221,In_1005);
and U2330 (N_2330,In_863,In_375);
or U2331 (N_2331,In_106,In_644);
nor U2332 (N_2332,In_178,In_473);
xor U2333 (N_2333,In_1439,In_127);
nor U2334 (N_2334,In_463,In_1224);
nand U2335 (N_2335,In_58,In_1203);
and U2336 (N_2336,In_156,In_562);
and U2337 (N_2337,In_857,In_199);
nor U2338 (N_2338,In_1111,In_985);
or U2339 (N_2339,In_14,In_268);
and U2340 (N_2340,In_285,In_178);
nor U2341 (N_2341,In_1257,In_847);
nor U2342 (N_2342,In_508,In_164);
nand U2343 (N_2343,In_319,In_396);
or U2344 (N_2344,In_410,In_1093);
nand U2345 (N_2345,In_752,In_866);
and U2346 (N_2346,In_1356,In_553);
nor U2347 (N_2347,In_1499,In_513);
or U2348 (N_2348,In_682,In_1393);
nor U2349 (N_2349,In_820,In_616);
and U2350 (N_2350,In_717,In_332);
or U2351 (N_2351,In_412,In_186);
or U2352 (N_2352,In_424,In_1397);
nand U2353 (N_2353,In_575,In_170);
nor U2354 (N_2354,In_385,In_969);
nor U2355 (N_2355,In_1121,In_1396);
and U2356 (N_2356,In_619,In_1314);
or U2357 (N_2357,In_1077,In_1112);
xnor U2358 (N_2358,In_1389,In_1395);
or U2359 (N_2359,In_743,In_1193);
or U2360 (N_2360,In_1012,In_1470);
and U2361 (N_2361,In_1003,In_529);
nor U2362 (N_2362,In_389,In_1124);
and U2363 (N_2363,In_982,In_1073);
nor U2364 (N_2364,In_386,In_186);
nor U2365 (N_2365,In_6,In_514);
nand U2366 (N_2366,In_1380,In_116);
nor U2367 (N_2367,In_152,In_125);
nor U2368 (N_2368,In_1023,In_210);
and U2369 (N_2369,In_1257,In_726);
or U2370 (N_2370,In_996,In_29);
nand U2371 (N_2371,In_51,In_767);
or U2372 (N_2372,In_26,In_1182);
nand U2373 (N_2373,In_1405,In_808);
or U2374 (N_2374,In_1174,In_1201);
or U2375 (N_2375,In_1181,In_1321);
nand U2376 (N_2376,In_1143,In_673);
nand U2377 (N_2377,In_551,In_97);
nor U2378 (N_2378,In_218,In_648);
and U2379 (N_2379,In_1430,In_1107);
xnor U2380 (N_2380,In_1003,In_518);
or U2381 (N_2381,In_918,In_910);
and U2382 (N_2382,In_516,In_569);
or U2383 (N_2383,In_1495,In_207);
and U2384 (N_2384,In_682,In_1178);
nand U2385 (N_2385,In_103,In_446);
or U2386 (N_2386,In_1214,In_901);
or U2387 (N_2387,In_886,In_645);
nor U2388 (N_2388,In_206,In_804);
and U2389 (N_2389,In_1370,In_315);
nor U2390 (N_2390,In_589,In_272);
and U2391 (N_2391,In_351,In_1138);
or U2392 (N_2392,In_1272,In_473);
or U2393 (N_2393,In_1092,In_1054);
and U2394 (N_2394,In_352,In_938);
or U2395 (N_2395,In_1364,In_830);
nor U2396 (N_2396,In_1352,In_708);
nor U2397 (N_2397,In_1268,In_86);
and U2398 (N_2398,In_790,In_548);
and U2399 (N_2399,In_72,In_1302);
and U2400 (N_2400,In_1292,In_890);
nor U2401 (N_2401,In_1113,In_978);
or U2402 (N_2402,In_201,In_472);
and U2403 (N_2403,In_1346,In_982);
nand U2404 (N_2404,In_783,In_1063);
nand U2405 (N_2405,In_930,In_1062);
nor U2406 (N_2406,In_113,In_1185);
and U2407 (N_2407,In_1059,In_255);
nand U2408 (N_2408,In_1209,In_590);
nor U2409 (N_2409,In_1232,In_658);
or U2410 (N_2410,In_1338,In_1077);
nor U2411 (N_2411,In_1399,In_1058);
or U2412 (N_2412,In_1356,In_14);
nand U2413 (N_2413,In_1357,In_406);
and U2414 (N_2414,In_1361,In_1463);
nand U2415 (N_2415,In_1473,In_1045);
or U2416 (N_2416,In_1451,In_340);
or U2417 (N_2417,In_470,In_865);
nand U2418 (N_2418,In_519,In_1231);
or U2419 (N_2419,In_1170,In_1438);
nor U2420 (N_2420,In_1186,In_1384);
or U2421 (N_2421,In_627,In_594);
or U2422 (N_2422,In_545,In_919);
and U2423 (N_2423,In_1156,In_386);
nor U2424 (N_2424,In_170,In_763);
nand U2425 (N_2425,In_822,In_867);
and U2426 (N_2426,In_33,In_98);
nor U2427 (N_2427,In_721,In_1081);
and U2428 (N_2428,In_614,In_1473);
nand U2429 (N_2429,In_957,In_728);
or U2430 (N_2430,In_241,In_605);
or U2431 (N_2431,In_783,In_407);
nor U2432 (N_2432,In_57,In_1273);
nand U2433 (N_2433,In_1464,In_559);
and U2434 (N_2434,In_180,In_993);
nand U2435 (N_2435,In_823,In_505);
nand U2436 (N_2436,In_1362,In_123);
and U2437 (N_2437,In_411,In_224);
nor U2438 (N_2438,In_42,In_482);
nor U2439 (N_2439,In_818,In_549);
nand U2440 (N_2440,In_1459,In_340);
nand U2441 (N_2441,In_435,In_968);
or U2442 (N_2442,In_111,In_1275);
nor U2443 (N_2443,In_97,In_138);
nor U2444 (N_2444,In_78,In_23);
nor U2445 (N_2445,In_659,In_1130);
nor U2446 (N_2446,In_706,In_815);
nor U2447 (N_2447,In_721,In_548);
nand U2448 (N_2448,In_570,In_656);
nor U2449 (N_2449,In_1425,In_293);
nor U2450 (N_2450,In_1131,In_1002);
or U2451 (N_2451,In_1123,In_1486);
nor U2452 (N_2452,In_1301,In_1087);
or U2453 (N_2453,In_625,In_814);
nor U2454 (N_2454,In_557,In_1205);
and U2455 (N_2455,In_374,In_932);
nor U2456 (N_2456,In_1223,In_1185);
xor U2457 (N_2457,In_1186,In_650);
or U2458 (N_2458,In_154,In_1306);
nand U2459 (N_2459,In_990,In_641);
nor U2460 (N_2460,In_1024,In_174);
nand U2461 (N_2461,In_1472,In_369);
nor U2462 (N_2462,In_1235,In_894);
or U2463 (N_2463,In_1233,In_1318);
and U2464 (N_2464,In_955,In_80);
or U2465 (N_2465,In_1113,In_26);
nor U2466 (N_2466,In_1309,In_688);
nand U2467 (N_2467,In_1014,In_1415);
and U2468 (N_2468,In_724,In_996);
nor U2469 (N_2469,In_1077,In_982);
and U2470 (N_2470,In_431,In_448);
or U2471 (N_2471,In_35,In_675);
and U2472 (N_2472,In_1068,In_1182);
xnor U2473 (N_2473,In_1220,In_354);
or U2474 (N_2474,In_997,In_1081);
or U2475 (N_2475,In_741,In_391);
xnor U2476 (N_2476,In_1155,In_415);
nand U2477 (N_2477,In_647,In_363);
or U2478 (N_2478,In_1394,In_123);
nand U2479 (N_2479,In_1230,In_722);
nand U2480 (N_2480,In_564,In_125);
nor U2481 (N_2481,In_347,In_1499);
or U2482 (N_2482,In_1179,In_746);
and U2483 (N_2483,In_1358,In_4);
nand U2484 (N_2484,In_1212,In_873);
nor U2485 (N_2485,In_1092,In_168);
or U2486 (N_2486,In_503,In_934);
and U2487 (N_2487,In_237,In_422);
or U2488 (N_2488,In_1442,In_474);
and U2489 (N_2489,In_7,In_659);
nand U2490 (N_2490,In_618,In_622);
and U2491 (N_2491,In_323,In_89);
and U2492 (N_2492,In_983,In_145);
nor U2493 (N_2493,In_583,In_252);
nor U2494 (N_2494,In_1002,In_674);
nor U2495 (N_2495,In_1492,In_1089);
nor U2496 (N_2496,In_1239,In_663);
and U2497 (N_2497,In_973,In_1022);
or U2498 (N_2498,In_528,In_181);
nand U2499 (N_2499,In_190,In_600);
nand U2500 (N_2500,In_476,In_1276);
nand U2501 (N_2501,In_1340,In_498);
or U2502 (N_2502,In_1413,In_173);
nand U2503 (N_2503,In_1463,In_1003);
or U2504 (N_2504,In_1497,In_152);
or U2505 (N_2505,In_403,In_585);
and U2506 (N_2506,In_1014,In_393);
and U2507 (N_2507,In_1148,In_1305);
nand U2508 (N_2508,In_1288,In_1446);
and U2509 (N_2509,In_485,In_78);
xor U2510 (N_2510,In_768,In_281);
nand U2511 (N_2511,In_423,In_599);
or U2512 (N_2512,In_876,In_1252);
xnor U2513 (N_2513,In_469,In_51);
nand U2514 (N_2514,In_57,In_269);
nand U2515 (N_2515,In_54,In_240);
or U2516 (N_2516,In_931,In_1128);
nand U2517 (N_2517,In_399,In_966);
nor U2518 (N_2518,In_1066,In_856);
nor U2519 (N_2519,In_981,In_1081);
and U2520 (N_2520,In_678,In_1492);
nand U2521 (N_2521,In_1467,In_623);
nand U2522 (N_2522,In_483,In_275);
nand U2523 (N_2523,In_463,In_1173);
or U2524 (N_2524,In_731,In_445);
and U2525 (N_2525,In_932,In_602);
and U2526 (N_2526,In_1148,In_1004);
nor U2527 (N_2527,In_1448,In_507);
nor U2528 (N_2528,In_1247,In_377);
or U2529 (N_2529,In_856,In_781);
and U2530 (N_2530,In_1413,In_967);
nand U2531 (N_2531,In_1496,In_815);
nand U2532 (N_2532,In_891,In_467);
and U2533 (N_2533,In_446,In_77);
and U2534 (N_2534,In_466,In_350);
and U2535 (N_2535,In_1365,In_1210);
nand U2536 (N_2536,In_1324,In_387);
nand U2537 (N_2537,In_542,In_17);
and U2538 (N_2538,In_1028,In_44);
nand U2539 (N_2539,In_1381,In_1222);
or U2540 (N_2540,In_1370,In_1363);
nand U2541 (N_2541,In_473,In_755);
and U2542 (N_2542,In_814,In_258);
nor U2543 (N_2543,In_371,In_455);
nor U2544 (N_2544,In_1011,In_140);
and U2545 (N_2545,In_188,In_775);
and U2546 (N_2546,In_849,In_1154);
or U2547 (N_2547,In_174,In_743);
nor U2548 (N_2548,In_996,In_423);
or U2549 (N_2549,In_1289,In_793);
nand U2550 (N_2550,In_123,In_1495);
nor U2551 (N_2551,In_1311,In_244);
and U2552 (N_2552,In_1097,In_738);
and U2553 (N_2553,In_1418,In_200);
or U2554 (N_2554,In_916,In_94);
and U2555 (N_2555,In_844,In_1174);
nor U2556 (N_2556,In_242,In_270);
nor U2557 (N_2557,In_9,In_470);
nor U2558 (N_2558,In_268,In_1327);
nand U2559 (N_2559,In_1301,In_686);
xnor U2560 (N_2560,In_497,In_890);
nand U2561 (N_2561,In_267,In_127);
and U2562 (N_2562,In_1370,In_1405);
nor U2563 (N_2563,In_912,In_354);
and U2564 (N_2564,In_653,In_1332);
nor U2565 (N_2565,In_143,In_530);
nor U2566 (N_2566,In_908,In_1193);
nand U2567 (N_2567,In_1461,In_1081);
nand U2568 (N_2568,In_299,In_459);
nand U2569 (N_2569,In_652,In_1373);
nand U2570 (N_2570,In_686,In_1216);
or U2571 (N_2571,In_813,In_1028);
and U2572 (N_2572,In_857,In_738);
nand U2573 (N_2573,In_662,In_1427);
and U2574 (N_2574,In_1043,In_592);
nor U2575 (N_2575,In_46,In_840);
and U2576 (N_2576,In_1074,In_819);
or U2577 (N_2577,In_578,In_630);
or U2578 (N_2578,In_1358,In_227);
and U2579 (N_2579,In_139,In_178);
nor U2580 (N_2580,In_1205,In_842);
and U2581 (N_2581,In_245,In_476);
or U2582 (N_2582,In_568,In_419);
nand U2583 (N_2583,In_724,In_565);
nand U2584 (N_2584,In_1058,In_725);
nor U2585 (N_2585,In_160,In_757);
nand U2586 (N_2586,In_157,In_1427);
and U2587 (N_2587,In_221,In_967);
nand U2588 (N_2588,In_1033,In_120);
nor U2589 (N_2589,In_1237,In_40);
and U2590 (N_2590,In_754,In_518);
and U2591 (N_2591,In_1019,In_332);
and U2592 (N_2592,In_483,In_1145);
nand U2593 (N_2593,In_293,In_617);
nor U2594 (N_2594,In_1326,In_985);
nand U2595 (N_2595,In_1354,In_586);
and U2596 (N_2596,In_652,In_258);
nand U2597 (N_2597,In_1223,In_872);
xor U2598 (N_2598,In_1101,In_83);
or U2599 (N_2599,In_1067,In_1089);
or U2600 (N_2600,In_1031,In_589);
or U2601 (N_2601,In_1235,In_472);
and U2602 (N_2602,In_1292,In_837);
or U2603 (N_2603,In_1093,In_199);
and U2604 (N_2604,In_466,In_443);
xor U2605 (N_2605,In_192,In_457);
nand U2606 (N_2606,In_971,In_1348);
or U2607 (N_2607,In_1464,In_272);
nor U2608 (N_2608,In_584,In_1046);
or U2609 (N_2609,In_629,In_1201);
nor U2610 (N_2610,In_1430,In_1179);
or U2611 (N_2611,In_673,In_43);
or U2612 (N_2612,In_630,In_706);
or U2613 (N_2613,In_337,In_689);
nor U2614 (N_2614,In_744,In_1260);
nand U2615 (N_2615,In_953,In_562);
nand U2616 (N_2616,In_1182,In_297);
or U2617 (N_2617,In_1,In_378);
or U2618 (N_2618,In_1324,In_1092);
nor U2619 (N_2619,In_884,In_783);
nor U2620 (N_2620,In_1307,In_161);
or U2621 (N_2621,In_654,In_1000);
nand U2622 (N_2622,In_557,In_333);
or U2623 (N_2623,In_1379,In_1063);
nor U2624 (N_2624,In_768,In_1412);
or U2625 (N_2625,In_1377,In_1207);
nand U2626 (N_2626,In_1240,In_488);
nand U2627 (N_2627,In_617,In_250);
and U2628 (N_2628,In_1058,In_818);
nor U2629 (N_2629,In_1297,In_765);
nor U2630 (N_2630,In_935,In_445);
nor U2631 (N_2631,In_812,In_163);
nor U2632 (N_2632,In_57,In_1011);
nor U2633 (N_2633,In_695,In_268);
nand U2634 (N_2634,In_487,In_9);
or U2635 (N_2635,In_1248,In_445);
nand U2636 (N_2636,In_607,In_139);
and U2637 (N_2637,In_670,In_1098);
and U2638 (N_2638,In_568,In_1056);
and U2639 (N_2639,In_774,In_899);
nor U2640 (N_2640,In_851,In_746);
or U2641 (N_2641,In_341,In_450);
nor U2642 (N_2642,In_980,In_1376);
and U2643 (N_2643,In_405,In_884);
nor U2644 (N_2644,In_999,In_1298);
or U2645 (N_2645,In_619,In_342);
or U2646 (N_2646,In_1014,In_819);
or U2647 (N_2647,In_26,In_1323);
nand U2648 (N_2648,In_420,In_671);
nand U2649 (N_2649,In_806,In_133);
nor U2650 (N_2650,In_410,In_708);
or U2651 (N_2651,In_195,In_1386);
nand U2652 (N_2652,In_1189,In_1101);
or U2653 (N_2653,In_488,In_15);
nor U2654 (N_2654,In_415,In_1047);
nor U2655 (N_2655,In_1370,In_842);
nor U2656 (N_2656,In_1426,In_399);
nor U2657 (N_2657,In_856,In_158);
and U2658 (N_2658,In_340,In_242);
and U2659 (N_2659,In_914,In_95);
nand U2660 (N_2660,In_439,In_319);
or U2661 (N_2661,In_243,In_701);
or U2662 (N_2662,In_1096,In_580);
nand U2663 (N_2663,In_921,In_151);
or U2664 (N_2664,In_1065,In_1279);
nor U2665 (N_2665,In_31,In_210);
and U2666 (N_2666,In_646,In_18);
or U2667 (N_2667,In_1293,In_515);
nor U2668 (N_2668,In_1051,In_675);
nand U2669 (N_2669,In_425,In_102);
nand U2670 (N_2670,In_638,In_1007);
nor U2671 (N_2671,In_600,In_568);
nand U2672 (N_2672,In_1292,In_1371);
or U2673 (N_2673,In_1104,In_392);
and U2674 (N_2674,In_1084,In_264);
and U2675 (N_2675,In_407,In_1105);
or U2676 (N_2676,In_144,In_1480);
nand U2677 (N_2677,In_488,In_1496);
nand U2678 (N_2678,In_790,In_953);
and U2679 (N_2679,In_721,In_1002);
nor U2680 (N_2680,In_17,In_352);
nor U2681 (N_2681,In_327,In_263);
nor U2682 (N_2682,In_859,In_662);
nor U2683 (N_2683,In_1187,In_1115);
or U2684 (N_2684,In_1331,In_738);
nor U2685 (N_2685,In_1323,In_264);
nand U2686 (N_2686,In_347,In_320);
nand U2687 (N_2687,In_47,In_1118);
nor U2688 (N_2688,In_1230,In_689);
nor U2689 (N_2689,In_706,In_1261);
nand U2690 (N_2690,In_169,In_939);
nor U2691 (N_2691,In_884,In_337);
nor U2692 (N_2692,In_644,In_35);
or U2693 (N_2693,In_541,In_761);
xnor U2694 (N_2694,In_1387,In_391);
and U2695 (N_2695,In_1437,In_583);
nor U2696 (N_2696,In_528,In_1056);
and U2697 (N_2697,In_318,In_397);
or U2698 (N_2698,In_263,In_1136);
or U2699 (N_2699,In_872,In_127);
or U2700 (N_2700,In_146,In_1076);
and U2701 (N_2701,In_608,In_980);
nor U2702 (N_2702,In_1034,In_257);
nor U2703 (N_2703,In_214,In_1254);
and U2704 (N_2704,In_778,In_1353);
nand U2705 (N_2705,In_1379,In_467);
xor U2706 (N_2706,In_799,In_873);
or U2707 (N_2707,In_8,In_1328);
and U2708 (N_2708,In_671,In_1190);
nor U2709 (N_2709,In_382,In_708);
nor U2710 (N_2710,In_790,In_866);
and U2711 (N_2711,In_530,In_1278);
or U2712 (N_2712,In_802,In_1459);
and U2713 (N_2713,In_368,In_656);
and U2714 (N_2714,In_1071,In_1302);
nor U2715 (N_2715,In_1103,In_296);
nand U2716 (N_2716,In_984,In_1055);
nor U2717 (N_2717,In_137,In_1263);
and U2718 (N_2718,In_238,In_217);
nor U2719 (N_2719,In_367,In_249);
and U2720 (N_2720,In_811,In_1325);
nor U2721 (N_2721,In_304,In_1464);
and U2722 (N_2722,In_574,In_1217);
or U2723 (N_2723,In_320,In_634);
xor U2724 (N_2724,In_71,In_1162);
or U2725 (N_2725,In_236,In_291);
nor U2726 (N_2726,In_1134,In_435);
and U2727 (N_2727,In_107,In_457);
or U2728 (N_2728,In_1324,In_145);
and U2729 (N_2729,In_662,In_1324);
or U2730 (N_2730,In_768,In_289);
and U2731 (N_2731,In_219,In_480);
or U2732 (N_2732,In_770,In_1488);
nor U2733 (N_2733,In_1144,In_248);
and U2734 (N_2734,In_1182,In_45);
nor U2735 (N_2735,In_216,In_823);
nor U2736 (N_2736,In_682,In_616);
or U2737 (N_2737,In_861,In_972);
or U2738 (N_2738,In_1226,In_246);
or U2739 (N_2739,In_506,In_552);
or U2740 (N_2740,In_1272,In_470);
nor U2741 (N_2741,In_332,In_874);
nor U2742 (N_2742,In_136,In_1268);
nor U2743 (N_2743,In_243,In_914);
nor U2744 (N_2744,In_264,In_957);
or U2745 (N_2745,In_937,In_544);
or U2746 (N_2746,In_582,In_1419);
nand U2747 (N_2747,In_333,In_752);
nor U2748 (N_2748,In_1460,In_1032);
and U2749 (N_2749,In_679,In_834);
or U2750 (N_2750,In_1039,In_233);
nor U2751 (N_2751,In_1104,In_150);
or U2752 (N_2752,In_137,In_1166);
nand U2753 (N_2753,In_233,In_351);
nor U2754 (N_2754,In_1269,In_514);
nand U2755 (N_2755,In_795,In_172);
or U2756 (N_2756,In_393,In_1252);
or U2757 (N_2757,In_653,In_519);
xnor U2758 (N_2758,In_798,In_342);
and U2759 (N_2759,In_1206,In_72);
nor U2760 (N_2760,In_225,In_643);
and U2761 (N_2761,In_209,In_71);
nor U2762 (N_2762,In_796,In_899);
or U2763 (N_2763,In_56,In_1398);
nor U2764 (N_2764,In_652,In_1441);
and U2765 (N_2765,In_1371,In_378);
or U2766 (N_2766,In_1189,In_1274);
or U2767 (N_2767,In_549,In_365);
nor U2768 (N_2768,In_1453,In_1343);
and U2769 (N_2769,In_768,In_1068);
nand U2770 (N_2770,In_12,In_988);
nor U2771 (N_2771,In_1037,In_649);
or U2772 (N_2772,In_106,In_865);
nand U2773 (N_2773,In_47,In_470);
nor U2774 (N_2774,In_503,In_711);
nor U2775 (N_2775,In_1043,In_447);
xnor U2776 (N_2776,In_274,In_1240);
nor U2777 (N_2777,In_1490,In_572);
or U2778 (N_2778,In_1261,In_1103);
or U2779 (N_2779,In_370,In_1304);
nor U2780 (N_2780,In_103,In_1300);
and U2781 (N_2781,In_251,In_278);
xnor U2782 (N_2782,In_1325,In_844);
or U2783 (N_2783,In_440,In_90);
nor U2784 (N_2784,In_1103,In_1405);
and U2785 (N_2785,In_1350,In_748);
or U2786 (N_2786,In_1357,In_1200);
nand U2787 (N_2787,In_410,In_712);
and U2788 (N_2788,In_1337,In_689);
nand U2789 (N_2789,In_926,In_355);
or U2790 (N_2790,In_899,In_628);
and U2791 (N_2791,In_63,In_196);
and U2792 (N_2792,In_1076,In_1242);
nor U2793 (N_2793,In_1290,In_320);
or U2794 (N_2794,In_111,In_723);
nor U2795 (N_2795,In_1237,In_47);
and U2796 (N_2796,In_1463,In_1187);
nand U2797 (N_2797,In_1266,In_854);
or U2798 (N_2798,In_983,In_666);
nand U2799 (N_2799,In_282,In_1317);
and U2800 (N_2800,In_1446,In_230);
and U2801 (N_2801,In_355,In_1014);
nand U2802 (N_2802,In_1436,In_871);
nor U2803 (N_2803,In_74,In_928);
nand U2804 (N_2804,In_1409,In_673);
and U2805 (N_2805,In_1048,In_124);
nand U2806 (N_2806,In_1145,In_1452);
nor U2807 (N_2807,In_1249,In_649);
and U2808 (N_2808,In_376,In_1108);
or U2809 (N_2809,In_1211,In_109);
nand U2810 (N_2810,In_113,In_1158);
nand U2811 (N_2811,In_446,In_1047);
nor U2812 (N_2812,In_219,In_497);
nand U2813 (N_2813,In_1051,In_659);
or U2814 (N_2814,In_371,In_1498);
and U2815 (N_2815,In_610,In_382);
or U2816 (N_2816,In_645,In_207);
and U2817 (N_2817,In_649,In_1274);
nor U2818 (N_2818,In_1231,In_287);
nor U2819 (N_2819,In_1005,In_1071);
and U2820 (N_2820,In_1384,In_1330);
or U2821 (N_2821,In_68,In_252);
nand U2822 (N_2822,In_745,In_254);
or U2823 (N_2823,In_1088,In_1139);
and U2824 (N_2824,In_26,In_134);
nor U2825 (N_2825,In_611,In_1232);
nor U2826 (N_2826,In_1493,In_643);
and U2827 (N_2827,In_954,In_729);
and U2828 (N_2828,In_1153,In_1423);
or U2829 (N_2829,In_320,In_240);
and U2830 (N_2830,In_1321,In_540);
nor U2831 (N_2831,In_775,In_423);
or U2832 (N_2832,In_83,In_1291);
and U2833 (N_2833,In_686,In_930);
nor U2834 (N_2834,In_1395,In_1133);
and U2835 (N_2835,In_392,In_1303);
or U2836 (N_2836,In_719,In_1307);
nand U2837 (N_2837,In_1473,In_97);
or U2838 (N_2838,In_1380,In_741);
or U2839 (N_2839,In_7,In_464);
nand U2840 (N_2840,In_577,In_1293);
nor U2841 (N_2841,In_578,In_998);
and U2842 (N_2842,In_188,In_324);
nor U2843 (N_2843,In_752,In_188);
and U2844 (N_2844,In_685,In_420);
nor U2845 (N_2845,In_1469,In_1495);
nand U2846 (N_2846,In_749,In_298);
nor U2847 (N_2847,In_1155,In_173);
nor U2848 (N_2848,In_329,In_464);
and U2849 (N_2849,In_888,In_1498);
or U2850 (N_2850,In_357,In_1268);
or U2851 (N_2851,In_1154,In_754);
nand U2852 (N_2852,In_835,In_577);
nand U2853 (N_2853,In_187,In_291);
or U2854 (N_2854,In_588,In_928);
nor U2855 (N_2855,In_632,In_24);
nand U2856 (N_2856,In_911,In_427);
or U2857 (N_2857,In_257,In_816);
nand U2858 (N_2858,In_492,In_1401);
nand U2859 (N_2859,In_573,In_65);
and U2860 (N_2860,In_1346,In_1274);
nor U2861 (N_2861,In_1009,In_1131);
nor U2862 (N_2862,In_42,In_439);
and U2863 (N_2863,In_767,In_148);
nand U2864 (N_2864,In_1415,In_1382);
and U2865 (N_2865,In_645,In_1420);
or U2866 (N_2866,In_1290,In_835);
or U2867 (N_2867,In_695,In_86);
and U2868 (N_2868,In_1235,In_1436);
nand U2869 (N_2869,In_1458,In_1477);
nand U2870 (N_2870,In_13,In_1019);
or U2871 (N_2871,In_1454,In_538);
nand U2872 (N_2872,In_785,In_845);
nor U2873 (N_2873,In_741,In_330);
nand U2874 (N_2874,In_343,In_771);
or U2875 (N_2875,In_1101,In_672);
nand U2876 (N_2876,In_616,In_256);
and U2877 (N_2877,In_1308,In_1483);
nand U2878 (N_2878,In_448,In_83);
or U2879 (N_2879,In_367,In_477);
nor U2880 (N_2880,In_998,In_66);
or U2881 (N_2881,In_376,In_909);
nand U2882 (N_2882,In_46,In_192);
nand U2883 (N_2883,In_100,In_880);
and U2884 (N_2884,In_1125,In_576);
or U2885 (N_2885,In_1198,In_613);
nor U2886 (N_2886,In_851,In_1325);
nor U2887 (N_2887,In_1201,In_1309);
nand U2888 (N_2888,In_716,In_490);
or U2889 (N_2889,In_924,In_1071);
or U2890 (N_2890,In_770,In_342);
nand U2891 (N_2891,In_1201,In_40);
nand U2892 (N_2892,In_222,In_1441);
nor U2893 (N_2893,In_15,In_1450);
nand U2894 (N_2894,In_422,In_1093);
and U2895 (N_2895,In_584,In_544);
and U2896 (N_2896,In_310,In_1095);
nor U2897 (N_2897,In_1245,In_17);
and U2898 (N_2898,In_1142,In_1314);
nor U2899 (N_2899,In_549,In_966);
or U2900 (N_2900,In_1077,In_338);
and U2901 (N_2901,In_935,In_1297);
or U2902 (N_2902,In_334,In_1143);
or U2903 (N_2903,In_1335,In_422);
or U2904 (N_2904,In_971,In_1100);
nor U2905 (N_2905,In_518,In_343);
or U2906 (N_2906,In_193,In_1268);
and U2907 (N_2907,In_1478,In_1318);
nand U2908 (N_2908,In_1127,In_1498);
nor U2909 (N_2909,In_777,In_1484);
or U2910 (N_2910,In_1369,In_1304);
nand U2911 (N_2911,In_725,In_103);
nand U2912 (N_2912,In_1035,In_748);
or U2913 (N_2913,In_525,In_790);
and U2914 (N_2914,In_385,In_965);
or U2915 (N_2915,In_217,In_442);
nand U2916 (N_2916,In_153,In_262);
or U2917 (N_2917,In_656,In_765);
or U2918 (N_2918,In_1192,In_618);
or U2919 (N_2919,In_1019,In_1170);
nand U2920 (N_2920,In_855,In_241);
nor U2921 (N_2921,In_994,In_401);
nand U2922 (N_2922,In_1099,In_991);
nand U2923 (N_2923,In_1087,In_526);
or U2924 (N_2924,In_97,In_31);
or U2925 (N_2925,In_458,In_486);
or U2926 (N_2926,In_839,In_344);
and U2927 (N_2927,In_883,In_348);
and U2928 (N_2928,In_796,In_393);
nand U2929 (N_2929,In_1097,In_270);
nor U2930 (N_2930,In_1039,In_121);
nand U2931 (N_2931,In_1285,In_1379);
and U2932 (N_2932,In_110,In_545);
nand U2933 (N_2933,In_479,In_61);
or U2934 (N_2934,In_1248,In_226);
or U2935 (N_2935,In_358,In_79);
nand U2936 (N_2936,In_1370,In_683);
and U2937 (N_2937,In_582,In_185);
or U2938 (N_2938,In_1127,In_639);
nand U2939 (N_2939,In_266,In_49);
nand U2940 (N_2940,In_208,In_1000);
nor U2941 (N_2941,In_1366,In_1241);
or U2942 (N_2942,In_731,In_1357);
nand U2943 (N_2943,In_715,In_689);
nand U2944 (N_2944,In_518,In_1274);
nor U2945 (N_2945,In_1157,In_731);
or U2946 (N_2946,In_899,In_871);
and U2947 (N_2947,In_722,In_279);
or U2948 (N_2948,In_1083,In_332);
or U2949 (N_2949,In_564,In_9);
and U2950 (N_2950,In_1237,In_1428);
or U2951 (N_2951,In_182,In_584);
nor U2952 (N_2952,In_184,In_1217);
or U2953 (N_2953,In_1300,In_248);
or U2954 (N_2954,In_1197,In_560);
or U2955 (N_2955,In_681,In_115);
nand U2956 (N_2956,In_756,In_1031);
nand U2957 (N_2957,In_1411,In_1399);
and U2958 (N_2958,In_128,In_1319);
nor U2959 (N_2959,In_775,In_407);
nand U2960 (N_2960,In_1041,In_87);
or U2961 (N_2961,In_859,In_938);
nor U2962 (N_2962,In_1360,In_1289);
nand U2963 (N_2963,In_143,In_861);
or U2964 (N_2964,In_295,In_511);
nand U2965 (N_2965,In_433,In_394);
or U2966 (N_2966,In_774,In_332);
and U2967 (N_2967,In_1154,In_653);
nand U2968 (N_2968,In_799,In_1349);
and U2969 (N_2969,In_353,In_420);
or U2970 (N_2970,In_1353,In_495);
nand U2971 (N_2971,In_97,In_3);
nand U2972 (N_2972,In_484,In_969);
or U2973 (N_2973,In_986,In_131);
or U2974 (N_2974,In_164,In_1393);
nor U2975 (N_2975,In_158,In_1354);
nand U2976 (N_2976,In_243,In_924);
or U2977 (N_2977,In_1008,In_650);
or U2978 (N_2978,In_489,In_617);
or U2979 (N_2979,In_358,In_750);
nor U2980 (N_2980,In_769,In_519);
nand U2981 (N_2981,In_507,In_193);
nor U2982 (N_2982,In_758,In_547);
nand U2983 (N_2983,In_294,In_422);
nor U2984 (N_2984,In_846,In_1435);
nor U2985 (N_2985,In_488,In_1095);
and U2986 (N_2986,In_828,In_196);
and U2987 (N_2987,In_1386,In_1056);
nor U2988 (N_2988,In_1143,In_177);
nand U2989 (N_2989,In_582,In_767);
nor U2990 (N_2990,In_385,In_1090);
nand U2991 (N_2991,In_280,In_272);
nand U2992 (N_2992,In_580,In_1105);
nor U2993 (N_2993,In_1101,In_1307);
or U2994 (N_2994,In_628,In_693);
or U2995 (N_2995,In_1129,In_844);
nor U2996 (N_2996,In_129,In_749);
nor U2997 (N_2997,In_566,In_369);
nor U2998 (N_2998,In_175,In_743);
or U2999 (N_2999,In_1090,In_1089);
and U3000 (N_3000,N_375,N_567);
and U3001 (N_3001,N_913,N_197);
nand U3002 (N_3002,N_1134,N_235);
nand U3003 (N_3003,N_276,N_1100);
nand U3004 (N_3004,N_2912,N_1892);
and U3005 (N_3005,N_2466,N_412);
nand U3006 (N_3006,N_2120,N_194);
and U3007 (N_3007,N_1769,N_2858);
nand U3008 (N_3008,N_2831,N_2659);
nor U3009 (N_3009,N_42,N_1060);
nand U3010 (N_3010,N_2539,N_1259);
or U3011 (N_3011,N_1506,N_1280);
nor U3012 (N_3012,N_746,N_2010);
nor U3013 (N_3013,N_144,N_2583);
nand U3014 (N_3014,N_1193,N_358);
nor U3015 (N_3015,N_2594,N_2615);
nand U3016 (N_3016,N_894,N_1065);
or U3017 (N_3017,N_390,N_1514);
and U3018 (N_3018,N_2427,N_2037);
nand U3019 (N_3019,N_613,N_1614);
and U3020 (N_3020,N_1716,N_2392);
and U3021 (N_3021,N_2048,N_2782);
or U3022 (N_3022,N_1090,N_2051);
nand U3023 (N_3023,N_139,N_1706);
or U3024 (N_3024,N_2582,N_2820);
and U3025 (N_3025,N_494,N_99);
or U3026 (N_3026,N_2043,N_406);
nor U3027 (N_3027,N_1057,N_2564);
nor U3028 (N_3028,N_2029,N_1351);
nand U3029 (N_3029,N_1550,N_767);
or U3030 (N_3030,N_1670,N_754);
or U3031 (N_3031,N_1684,N_1927);
nand U3032 (N_3032,N_695,N_665);
nand U3033 (N_3033,N_410,N_2959);
nand U3034 (N_3034,N_1136,N_2910);
or U3035 (N_3035,N_2137,N_507);
xor U3036 (N_3036,N_2590,N_979);
and U3037 (N_3037,N_2900,N_813);
and U3038 (N_3038,N_681,N_2380);
nand U3039 (N_3039,N_2842,N_648);
nand U3040 (N_3040,N_2686,N_72);
or U3041 (N_3041,N_938,N_409);
nor U3042 (N_3042,N_1099,N_1638);
and U3043 (N_3043,N_503,N_163);
nand U3044 (N_3044,N_1559,N_36);
or U3045 (N_3045,N_511,N_1226);
nor U3046 (N_3046,N_525,N_1500);
nand U3047 (N_3047,N_1821,N_467);
or U3048 (N_3048,N_1202,N_1128);
nand U3049 (N_3049,N_1875,N_2335);
and U3050 (N_3050,N_690,N_1776);
nor U3051 (N_3051,N_1019,N_745);
nand U3052 (N_3052,N_330,N_2053);
nand U3053 (N_3053,N_1110,N_1388);
nor U3054 (N_3054,N_1436,N_1497);
xor U3055 (N_3055,N_1204,N_2290);
nand U3056 (N_3056,N_620,N_642);
nor U3057 (N_3057,N_167,N_291);
nor U3058 (N_3058,N_2089,N_2836);
nor U3059 (N_3059,N_1268,N_2189);
and U3060 (N_3060,N_580,N_1391);
nand U3061 (N_3061,N_699,N_1669);
nor U3062 (N_3062,N_2862,N_600);
nand U3063 (N_3063,N_856,N_2094);
nor U3064 (N_3064,N_1303,N_2517);
or U3065 (N_3065,N_2390,N_1722);
and U3066 (N_3066,N_1718,N_416);
nor U3067 (N_3067,N_1146,N_257);
and U3068 (N_3068,N_1984,N_211);
nor U3069 (N_3069,N_1794,N_1362);
nand U3070 (N_3070,N_2738,N_2944);
or U3071 (N_3071,N_2976,N_2062);
and U3072 (N_3072,N_840,N_1400);
or U3073 (N_3073,N_2462,N_2047);
xnor U3074 (N_3074,N_1572,N_1066);
or U3075 (N_3075,N_817,N_1829);
and U3076 (N_3076,N_164,N_2835);
nand U3077 (N_3077,N_2244,N_2515);
nor U3078 (N_3078,N_2599,N_1975);
or U3079 (N_3079,N_446,N_1331);
or U3080 (N_3080,N_433,N_214);
and U3081 (N_3081,N_2557,N_1624);
nand U3082 (N_3082,N_1929,N_2343);
and U3083 (N_3083,N_1819,N_1895);
xnor U3084 (N_3084,N_646,N_1055);
nor U3085 (N_3085,N_1820,N_2199);
or U3086 (N_3086,N_2591,N_2793);
nor U3087 (N_3087,N_1884,N_308);
or U3088 (N_3088,N_2018,N_807);
nand U3089 (N_3089,N_2485,N_2394);
and U3090 (N_3090,N_1507,N_1796);
nor U3091 (N_3091,N_2409,N_2629);
nand U3092 (N_3092,N_2084,N_2324);
nor U3093 (N_3093,N_1373,N_921);
and U3094 (N_3094,N_307,N_700);
or U3095 (N_3095,N_1471,N_2059);
nor U3096 (N_3096,N_778,N_1833);
and U3097 (N_3097,N_2116,N_659);
or U3098 (N_3098,N_2844,N_1904);
nand U3099 (N_3099,N_2351,N_2241);
nor U3100 (N_3100,N_2925,N_2428);
and U3101 (N_3101,N_289,N_1224);
and U3102 (N_3102,N_1167,N_2724);
nand U3103 (N_3103,N_657,N_1304);
nand U3104 (N_3104,N_2797,N_268);
nand U3105 (N_3105,N_2649,N_2839);
and U3106 (N_3106,N_254,N_533);
and U3107 (N_3107,N_2832,N_1971);
nand U3108 (N_3108,N_985,N_1192);
and U3109 (N_3109,N_1586,N_1120);
nor U3110 (N_3110,N_2891,N_1994);
or U3111 (N_3111,N_1360,N_246);
or U3112 (N_3112,N_2531,N_1551);
and U3113 (N_3113,N_1420,N_1006);
and U3114 (N_3114,N_1095,N_1288);
and U3115 (N_3115,N_942,N_2677);
nand U3116 (N_3116,N_2500,N_2093);
xnor U3117 (N_3117,N_1751,N_2081);
nand U3118 (N_3118,N_39,N_1594);
or U3119 (N_3119,N_2936,N_73);
and U3120 (N_3120,N_2830,N_1246);
nand U3121 (N_3121,N_1313,N_46);
nand U3122 (N_3122,N_1069,N_143);
nor U3123 (N_3123,N_2345,N_2363);
or U3124 (N_3124,N_1163,N_1284);
nor U3125 (N_3125,N_93,N_316);
nand U3126 (N_3126,N_2402,N_462);
nor U3127 (N_3127,N_270,N_1449);
nor U3128 (N_3128,N_2665,N_48);
nor U3129 (N_3129,N_1775,N_1107);
nor U3130 (N_3130,N_1656,N_1073);
and U3131 (N_3131,N_1000,N_2581);
and U3132 (N_3132,N_174,N_373);
nor U3133 (N_3133,N_1882,N_2651);
nand U3134 (N_3134,N_293,N_355);
nor U3135 (N_3135,N_2707,N_21);
xnor U3136 (N_3136,N_44,N_88);
nand U3137 (N_3137,N_1426,N_715);
and U3138 (N_3138,N_165,N_1860);
and U3139 (N_3139,N_571,N_1615);
or U3140 (N_3140,N_1340,N_2109);
and U3141 (N_3141,N_388,N_2433);
and U3142 (N_3142,N_1952,N_2494);
or U3143 (N_3143,N_2681,N_1538);
nor U3144 (N_3144,N_1503,N_509);
nand U3145 (N_3145,N_1423,N_2332);
and U3146 (N_3146,N_106,N_2745);
nand U3147 (N_3147,N_2328,N_1770);
and U3148 (N_3148,N_1205,N_801);
nor U3149 (N_3149,N_2076,N_2796);
nand U3150 (N_3150,N_1189,N_2320);
and U3151 (N_3151,N_28,N_798);
nor U3152 (N_3152,N_2854,N_184);
nand U3153 (N_3153,N_1879,N_429);
nor U3154 (N_3154,N_1413,N_2156);
nand U3155 (N_3155,N_2237,N_1077);
nand U3156 (N_3156,N_1747,N_2027);
or U3157 (N_3157,N_2104,N_666);
nor U3158 (N_3158,N_1477,N_2175);
nand U3159 (N_3159,N_1002,N_1935);
nand U3160 (N_3160,N_1864,N_2180);
nand U3161 (N_3161,N_1618,N_245);
nand U3162 (N_3162,N_1940,N_2764);
xnor U3163 (N_3163,N_1050,N_1393);
xnor U3164 (N_3164,N_2661,N_1665);
nor U3165 (N_3165,N_1767,N_1789);
and U3166 (N_3166,N_2833,N_160);
and U3167 (N_3167,N_545,N_1611);
or U3168 (N_3168,N_1143,N_1384);
and U3169 (N_3169,N_2049,N_336);
nor U3170 (N_3170,N_2323,N_1662);
and U3171 (N_3171,N_1451,N_1790);
or U3172 (N_3172,N_842,N_115);
nand U3173 (N_3173,N_304,N_2269);
nor U3174 (N_3174,N_628,N_634);
and U3175 (N_3175,N_679,N_2715);
or U3176 (N_3176,N_103,N_2040);
or U3177 (N_3177,N_2553,N_2792);
xnor U3178 (N_3178,N_1680,N_937);
nand U3179 (N_3179,N_1554,N_2355);
nor U3180 (N_3180,N_258,N_1173);
nand U3181 (N_3181,N_2003,N_1628);
and U3182 (N_3182,N_712,N_1759);
and U3183 (N_3183,N_1292,N_2578);
and U3184 (N_3184,N_2924,N_70);
nor U3185 (N_3185,N_2790,N_122);
nor U3186 (N_3186,N_3,N_841);
and U3187 (N_3187,N_569,N_1082);
and U3188 (N_3188,N_598,N_2304);
and U3189 (N_3189,N_247,N_2456);
nor U3190 (N_3190,N_2684,N_2032);
nand U3191 (N_3191,N_1710,N_2756);
nand U3192 (N_3192,N_2901,N_279);
nand U3193 (N_3193,N_2859,N_2044);
or U3194 (N_3194,N_2486,N_346);
or U3195 (N_3195,N_1894,N_2713);
or U3196 (N_3196,N_1035,N_251);
and U3197 (N_3197,N_2683,N_1936);
nand U3198 (N_3198,N_2856,N_2788);
or U3199 (N_3199,N_1934,N_344);
nand U3200 (N_3200,N_2077,N_2876);
nand U3201 (N_3201,N_1792,N_846);
nand U3202 (N_3202,N_1979,N_547);
nor U3203 (N_3203,N_2277,N_1238);
or U3204 (N_3204,N_458,N_1933);
nand U3205 (N_3205,N_2149,N_2103);
nand U3206 (N_3206,N_783,N_2384);
nand U3207 (N_3207,N_2215,N_2245);
or U3208 (N_3208,N_2100,N_1116);
and U3209 (N_3209,N_74,N_87);
or U3210 (N_3210,N_908,N_652);
or U3211 (N_3211,N_845,N_2798);
nor U3212 (N_3212,N_2947,N_2650);
xor U3213 (N_3213,N_422,N_812);
or U3214 (N_3214,N_608,N_1653);
nor U3215 (N_3215,N_799,N_1956);
or U3216 (N_3216,N_1697,N_2732);
and U3217 (N_3217,N_2755,N_1237);
and U3218 (N_3218,N_2408,N_2775);
nor U3219 (N_3219,N_1299,N_1330);
or U3220 (N_3220,N_1909,N_1972);
xor U3221 (N_3221,N_1197,N_2701);
nor U3222 (N_3222,N_1880,N_590);
or U3223 (N_3223,N_321,N_546);
or U3224 (N_3224,N_2075,N_2412);
and U3225 (N_3225,N_519,N_2501);
or U3226 (N_3226,N_1369,N_2586);
or U3227 (N_3227,N_2102,N_177);
nor U3228 (N_3228,N_1954,N_1080);
nor U3229 (N_3229,N_1920,N_454);
or U3230 (N_3230,N_1513,N_1402);
and U3231 (N_3231,N_890,N_1166);
nor U3232 (N_3232,N_773,N_743);
nand U3233 (N_3233,N_2902,N_1948);
nor U3234 (N_3234,N_925,N_116);
nand U3235 (N_3235,N_1876,N_2791);
nor U3236 (N_3236,N_2297,N_98);
and U3237 (N_3237,N_2635,N_185);
or U3238 (N_3238,N_2827,N_1406);
nand U3239 (N_3239,N_870,N_461);
nor U3240 (N_3240,N_1648,N_1172);
nand U3241 (N_3241,N_915,N_1034);
xor U3242 (N_3242,N_914,N_2685);
nand U3243 (N_3243,N_1587,N_52);
and U3244 (N_3244,N_238,N_770);
nand U3245 (N_3245,N_1481,N_717);
nand U3246 (N_3246,N_1443,N_2054);
and U3247 (N_3247,N_1982,N_2817);
and U3248 (N_3248,N_1553,N_53);
nand U3249 (N_3249,N_627,N_784);
or U3250 (N_3250,N_1315,N_1639);
nor U3251 (N_3251,N_1977,N_1112);
and U3252 (N_3252,N_1563,N_1612);
nand U3253 (N_3253,N_671,N_1516);
or U3254 (N_3254,N_2082,N_2369);
or U3255 (N_3255,N_1686,N_777);
or U3256 (N_3256,N_809,N_1270);
or U3257 (N_3257,N_2640,N_2203);
or U3258 (N_3258,N_2927,N_718);
nand U3259 (N_3259,N_1811,N_2331);
or U3260 (N_3260,N_1125,N_1962);
nand U3261 (N_3261,N_852,N_2783);
or U3262 (N_3262,N_1574,N_234);
nor U3263 (N_3263,N_472,N_2449);
nand U3264 (N_3264,N_2789,N_630);
nor U3265 (N_3265,N_788,N_1029);
and U3266 (N_3266,N_105,N_867);
and U3267 (N_3267,N_2816,N_107);
or U3268 (N_3268,N_1001,N_1139);
or U3269 (N_3269,N_2413,N_266);
nor U3270 (N_3270,N_1741,N_1054);
nor U3271 (N_3271,N_1729,N_2751);
or U3272 (N_3272,N_101,N_2155);
or U3273 (N_3273,N_1140,N_2522);
nand U3274 (N_3274,N_1549,N_68);
or U3275 (N_3275,N_1106,N_274);
nor U3276 (N_3276,N_1676,N_797);
and U3277 (N_3277,N_1872,N_1926);
or U3278 (N_3278,N_916,N_1673);
nor U3279 (N_3279,N_384,N_2425);
and U3280 (N_3280,N_574,N_486);
and U3281 (N_3281,N_2562,N_360);
nand U3282 (N_3282,N_2346,N_67);
or U3283 (N_3283,N_2802,N_1316);
and U3284 (N_3284,N_2857,N_231);
nand U3285 (N_3285,N_997,N_1901);
nor U3286 (N_3286,N_2024,N_2339);
nand U3287 (N_3287,N_1319,N_1523);
nor U3288 (N_3288,N_918,N_2248);
or U3289 (N_3289,N_1242,N_265);
xnor U3290 (N_3290,N_1508,N_2917);
nand U3291 (N_3291,N_435,N_742);
and U3292 (N_3292,N_248,N_1185);
nor U3293 (N_3293,N_831,N_2334);
nand U3294 (N_3294,N_2502,N_1309);
xor U3295 (N_3295,N_2992,N_1218);
or U3296 (N_3296,N_528,N_1414);
or U3297 (N_3297,N_1448,N_1087);
and U3298 (N_3298,N_1221,N_1543);
or U3299 (N_3299,N_2918,N_586);
or U3300 (N_3300,N_804,N_2747);
or U3301 (N_3301,N_2490,N_527);
nand U3302 (N_3302,N_477,N_2946);
or U3303 (N_3303,N_935,N_973);
and U3304 (N_3304,N_2092,N_1326);
or U3305 (N_3305,N_2060,N_720);
and U3306 (N_3306,N_1296,N_2679);
and U3307 (N_3307,N_860,N_959);
or U3308 (N_3308,N_2892,N_1736);
nand U3309 (N_3309,N_32,N_2209);
xnor U3310 (N_3310,N_676,N_84);
and U3311 (N_3311,N_2916,N_611);
xor U3312 (N_3312,N_549,N_1142);
nand U3313 (N_3313,N_1924,N_685);
and U3314 (N_3314,N_379,N_1943);
and U3315 (N_3315,N_1137,N_1078);
nand U3316 (N_3316,N_2023,N_529);
nor U3317 (N_3317,N_168,N_1417);
and U3318 (N_3318,N_1757,N_992);
and U3319 (N_3319,N_880,N_1668);
nand U3320 (N_3320,N_2487,N_1993);
and U3321 (N_3321,N_1306,N_148);
or U3322 (N_3322,N_2556,N_1126);
and U3323 (N_3323,N_2544,N_761);
nand U3324 (N_3324,N_1438,N_1051);
xnor U3325 (N_3325,N_1492,N_1235);
or U3326 (N_3326,N_1210,N_2829);
nand U3327 (N_3327,N_1375,N_2080);
nor U3328 (N_3328,N_172,N_697);
nor U3329 (N_3329,N_426,N_626);
nor U3330 (N_3330,N_255,N_1717);
or U3331 (N_3331,N_2949,N_2309);
nand U3332 (N_3332,N_2693,N_2377);
and U3333 (N_3333,N_2682,N_305);
or U3334 (N_3334,N_885,N_1004);
and U3335 (N_3335,N_162,N_1632);
nand U3336 (N_3336,N_201,N_591);
and U3337 (N_3337,N_1188,N_110);
nor U3338 (N_3338,N_1873,N_2688);
or U3339 (N_3339,N_242,N_2541);
nand U3340 (N_3340,N_1597,N_2253);
or U3341 (N_3341,N_1496,N_460);
or U3342 (N_3342,N_1441,N_2008);
or U3343 (N_3343,N_1247,N_2400);
and U3344 (N_3344,N_541,N_2875);
and U3345 (N_3345,N_2288,N_1236);
nand U3346 (N_3346,N_662,N_1970);
and U3347 (N_3347,N_114,N_170);
nand U3348 (N_3348,N_2496,N_2937);
nor U3349 (N_3349,N_601,N_998);
or U3350 (N_3350,N_275,N_1740);
nand U3351 (N_3351,N_296,N_1658);
and U3352 (N_3352,N_2663,N_1661);
or U3353 (N_3353,N_965,N_1735);
nand U3354 (N_3354,N_847,N_1130);
and U3355 (N_3355,N_1501,N_647);
or U3356 (N_3356,N_2056,N_1701);
nand U3357 (N_3357,N_609,N_2318);
or U3358 (N_3358,N_1083,N_815);
or U3359 (N_3359,N_1260,N_1990);
nor U3360 (N_3360,N_2317,N_644);
nor U3361 (N_3361,N_558,N_2198);
nor U3362 (N_3362,N_2904,N_2670);
and U3363 (N_3363,N_1267,N_2143);
or U3364 (N_3364,N_1510,N_1081);
nand U3365 (N_3365,N_883,N_1325);
and U3366 (N_3366,N_877,N_2554);
nand U3367 (N_3367,N_1617,N_1682);
or U3368 (N_3368,N_1424,N_1067);
nor U3369 (N_3369,N_2152,N_2628);
and U3370 (N_3370,N_1076,N_1435);
nor U3371 (N_3371,N_1533,N_1967);
and U3372 (N_3372,N_2687,N_1942);
nor U3373 (N_3373,N_2115,N_1817);
nor U3374 (N_3374,N_1337,N_2885);
or U3375 (N_3375,N_1455,N_300);
and U3376 (N_3376,N_1634,N_2860);
and U3377 (N_3377,N_902,N_2888);
or U3378 (N_3378,N_2382,N_2015);
and U3379 (N_3379,N_2610,N_599);
and U3380 (N_3380,N_443,N_1502);
or U3381 (N_3381,N_2162,N_1630);
nor U3382 (N_3382,N_1953,N_1743);
and U3383 (N_3383,N_1902,N_2471);
and U3384 (N_3384,N_1842,N_1932);
or U3385 (N_3385,N_1119,N_343);
nand U3386 (N_3386,N_2654,N_2480);
nand U3387 (N_3387,N_1432,N_181);
or U3388 (N_3388,N_928,N_1801);
nand U3389 (N_3389,N_1613,N_578);
nor U3390 (N_3390,N_2243,N_361);
nand U3391 (N_3391,N_1225,N_1871);
nor U3392 (N_3392,N_418,N_362);
xor U3393 (N_3393,N_733,N_1036);
nand U3394 (N_3394,N_943,N_1281);
or U3395 (N_3395,N_2216,N_889);
nor U3396 (N_3396,N_872,N_563);
or U3397 (N_3397,N_1969,N_749);
nor U3398 (N_3398,N_672,N_1203);
and U3399 (N_3399,N_1763,N_351);
nand U3400 (N_3400,N_1261,N_2527);
nor U3401 (N_3401,N_193,N_2705);
and U3402 (N_3402,N_1294,N_2647);
or U3403 (N_3403,N_1305,N_993);
nand U3404 (N_3404,N_982,N_1409);
or U3405 (N_3405,N_2621,N_1385);
nor U3406 (N_3406,N_1158,N_573);
xor U3407 (N_3407,N_2126,N_2587);
or U3408 (N_3408,N_2899,N_724);
and U3409 (N_3409,N_497,N_961);
nor U3410 (N_3410,N_1071,N_983);
nand U3411 (N_3411,N_399,N_331);
nand U3412 (N_3412,N_635,N_2020);
nand U3413 (N_3413,N_2930,N_121);
and U3414 (N_3414,N_2994,N_2370);
nand U3415 (N_3415,N_977,N_714);
or U3416 (N_3416,N_1122,N_2302);
nor U3417 (N_3417,N_2604,N_405);
or U3418 (N_3418,N_789,N_1715);
or U3419 (N_3419,N_178,N_111);
or U3420 (N_3420,N_385,N_638);
and U3421 (N_3421,N_2287,N_1249);
and U3422 (N_3422,N_15,N_1773);
and U3423 (N_3423,N_2064,N_2219);
and U3424 (N_3424,N_808,N_508);
and U3425 (N_3425,N_2823,N_1037);
or U3426 (N_3426,N_484,N_1764);
xor U3427 (N_3427,N_2593,N_865);
nand U3428 (N_3428,N_470,N_2671);
or U3429 (N_3429,N_1703,N_221);
and U3430 (N_3430,N_2736,N_22);
nand U3431 (N_3431,N_2251,N_2372);
or U3432 (N_3432,N_1998,N_1946);
nor U3433 (N_3433,N_1487,N_2799);
nand U3434 (N_3434,N_2499,N_868);
xor U3435 (N_3435,N_1643,N_2450);
nand U3436 (N_3436,N_2913,N_2634);
and U3437 (N_3437,N_1031,N_971);
and U3438 (N_3438,N_1485,N_2837);
or U3439 (N_3439,N_1804,N_886);
nand U3440 (N_3440,N_1870,N_1347);
nor U3441 (N_3441,N_2118,N_1694);
nor U3442 (N_3442,N_619,N_2250);
nor U3443 (N_3443,N_1986,N_2626);
and U3444 (N_3444,N_1580,N_515);
and U3445 (N_3445,N_1704,N_1457);
nand U3446 (N_3446,N_2616,N_2222);
or U3447 (N_3447,N_2519,N_2815);
nand U3448 (N_3448,N_2753,N_329);
nand U3449 (N_3449,N_2470,N_2666);
or U3450 (N_3450,N_423,N_2000);
or U3451 (N_3451,N_2579,N_1453);
and U3452 (N_3452,N_866,N_2723);
or U3453 (N_3453,N_1368,N_2220);
nor U3454 (N_3454,N_1928,N_2617);
nor U3455 (N_3455,N_2153,N_2795);
nor U3456 (N_3456,N_2619,N_427);
and U3457 (N_3457,N_2236,N_597);
and U3458 (N_3458,N_543,N_1484);
or U3459 (N_3459,N_1540,N_755);
nor U3460 (N_3460,N_625,N_1672);
nor U3461 (N_3461,N_1328,N_2877);
or U3462 (N_3462,N_1620,N_1381);
or U3463 (N_3463,N_2555,N_1849);
nor U3464 (N_3464,N_118,N_244);
nor U3465 (N_3465,N_2415,N_2125);
nor U3466 (N_3466,N_2239,N_1068);
or U3467 (N_3467,N_763,N_157);
or U3468 (N_3468,N_1963,N_2371);
or U3469 (N_3469,N_436,N_2605);
nor U3470 (N_3470,N_1227,N_1271);
and U3471 (N_3471,N_893,N_1696);
nor U3472 (N_3472,N_2945,N_2627);
and U3473 (N_3473,N_834,N_1269);
nand U3474 (N_3474,N_2463,N_2459);
nand U3475 (N_3475,N_91,N_2672);
nand U3476 (N_3476,N_2855,N_1355);
and U3477 (N_3477,N_1008,N_1760);
or U3478 (N_3478,N_595,N_2066);
or U3479 (N_3479,N_1725,N_2375);
nor U3480 (N_3480,N_2508,N_158);
and U3481 (N_3481,N_2041,N_1059);
nand U3482 (N_3482,N_2431,N_2187);
nand U3483 (N_3483,N_1631,N_2689);
nor U3484 (N_3484,N_2235,N_1096);
and U3485 (N_3485,N_58,N_1797);
or U3486 (N_3486,N_502,N_780);
and U3487 (N_3487,N_1843,N_323);
or U3488 (N_3488,N_779,N_1458);
or U3489 (N_3489,N_1622,N_135);
nand U3490 (N_3490,N_2366,N_1626);
nor U3491 (N_3491,N_756,N_878);
nor U3492 (N_3492,N_830,N_2221);
and U3493 (N_3493,N_2974,N_250);
nor U3494 (N_3494,N_2819,N_1522);
nand U3495 (N_3495,N_1010,N_2070);
and U3496 (N_3496,N_2543,N_1765);
nor U3497 (N_3497,N_318,N_2646);
or U3498 (N_3498,N_577,N_758);
nor U3499 (N_3499,N_54,N_707);
nand U3500 (N_3500,N_879,N_861);
and U3501 (N_3501,N_2883,N_1798);
or U3502 (N_3502,N_2442,N_2388);
and U3503 (N_3503,N_2252,N_1475);
and U3504 (N_3504,N_2356,N_1846);
and U3505 (N_3505,N_2866,N_1132);
or U3506 (N_3506,N_33,N_1179);
nor U3507 (N_3507,N_1361,N_90);
nor U3508 (N_3508,N_1250,N_1957);
nand U3509 (N_3509,N_881,N_1756);
xor U3510 (N_3510,N_520,N_565);
nand U3511 (N_3511,N_2188,N_1900);
nand U3512 (N_3512,N_217,N_636);
or U3513 (N_3513,N_438,N_1907);
and U3514 (N_3514,N_2914,N_104);
nand U3515 (N_3515,N_1577,N_19);
or U3516 (N_3516,N_516,N_2184);
and U3517 (N_3517,N_1589,N_750);
nor U3518 (N_3518,N_1687,N_2690);
nor U3519 (N_3519,N_1024,N_480);
and U3520 (N_3520,N_1016,N_735);
and U3521 (N_3521,N_2869,N_1645);
nor U3522 (N_3522,N_2240,N_694);
or U3523 (N_3523,N_748,N_873);
nand U3524 (N_3524,N_2454,N_2204);
or U3525 (N_3525,N_588,N_2349);
and U3526 (N_3526,N_730,N_774);
or U3527 (N_3527,N_1652,N_267);
nand U3528 (N_3528,N_703,N_2987);
nor U3529 (N_3529,N_1575,N_451);
nand U3530 (N_3530,N_71,N_1198);
nor U3531 (N_3531,N_825,N_1230);
nor U3532 (N_3532,N_414,N_2341);
nand U3533 (N_3533,N_999,N_532);
nand U3534 (N_3534,N_2563,N_59);
or U3535 (N_3535,N_76,N_2733);
nor U3536 (N_3536,N_2295,N_1366);
and U3537 (N_3537,N_2192,N_692);
or U3538 (N_3538,N_218,N_1463);
nand U3539 (N_3539,N_1646,N_1468);
or U3540 (N_3540,N_469,N_1411);
nor U3541 (N_3541,N_1675,N_1434);
nand U3542 (N_3542,N_1590,N_1840);
or U3543 (N_3543,N_131,N_955);
nand U3544 (N_3544,N_391,N_1182);
nand U3545 (N_3545,N_795,N_156);
nor U3546 (N_3546,N_2880,N_1495);
nor U3547 (N_3547,N_814,N_448);
nor U3548 (N_3548,N_668,N_1195);
nor U3549 (N_3549,N_2893,N_513);
nand U3550 (N_3550,N_2028,N_1691);
nor U3551 (N_3551,N_1965,N_63);
or U3552 (N_3552,N_906,N_612);
and U3553 (N_3553,N_113,N_327);
and U3554 (N_3554,N_1573,N_622);
xor U3555 (N_3555,N_2061,N_1987);
or U3556 (N_3556,N_2310,N_1108);
nor U3557 (N_3557,N_2329,N_1779);
nand U3558 (N_3558,N_2348,N_1308);
nand U3559 (N_3559,N_2213,N_1109);
xnor U3560 (N_3560,N_1585,N_2737);
nor U3561 (N_3561,N_2483,N_2529);
nand U3562 (N_3562,N_1466,N_615);
and U3563 (N_3563,N_1431,N_2140);
and U3564 (N_3564,N_952,N_161);
and U3565 (N_3565,N_2603,N_196);
nor U3566 (N_3566,N_382,N_2352);
nand U3567 (N_3567,N_411,N_1584);
nor U3568 (N_3568,N_1421,N_1750);
and U3569 (N_3569,N_2809,N_1307);
and U3570 (N_3570,N_149,N_2865);
nor U3571 (N_3571,N_372,N_978);
or U3572 (N_3572,N_1088,N_1983);
nor U3573 (N_3573,N_688,N_510);
and U3574 (N_3574,N_536,N_781);
nor U3575 (N_3575,N_2656,N_2598);
nor U3576 (N_3576,N_26,N_2403);
or U3577 (N_3577,N_1372,N_2364);
and U3578 (N_3578,N_492,N_2492);
and U3579 (N_3579,N_1053,N_933);
nand U3580 (N_3580,N_934,N_987);
nor U3581 (N_3581,N_18,N_1908);
or U3582 (N_3582,N_1898,N_2217);
nor U3583 (N_3583,N_97,N_731);
or U3584 (N_3584,N_2573,N_2105);
and U3585 (N_3585,N_1150,N_23);
and U3586 (N_3586,N_1647,N_352);
and U3587 (N_3587,N_2620,N_920);
nor U3588 (N_3588,N_1815,N_2322);
and U3589 (N_3589,N_2521,N_805);
or U3590 (N_3590,N_760,N_1058);
nor U3591 (N_3591,N_1123,N_848);
nor U3592 (N_3592,N_728,N_576);
nand U3593 (N_3593,N_696,N_556);
nor U3594 (N_3594,N_986,N_281);
and U3595 (N_3595,N_1548,N_2678);
nor U3596 (N_3596,N_2358,N_2472);
nor U3597 (N_3597,N_109,N_1228);
and U3598 (N_3598,N_1245,N_2291);
nor U3599 (N_3599,N_1118,N_1278);
or U3600 (N_3600,N_1659,N_936);
or U3601 (N_3601,N_286,N_1407);
nand U3602 (N_3602,N_2004,N_2196);
nand U3603 (N_3603,N_2354,N_1015);
nor U3604 (N_3604,N_1440,N_2478);
nand U3605 (N_3605,N_2709,N_1854);
nor U3606 (N_3606,N_1038,N_2031);
nor U3607 (N_3607,N_1713,N_2419);
or U3608 (N_3608,N_1552,N_557);
or U3609 (N_3609,N_2307,N_2313);
nor U3610 (N_3610,N_2638,N_2067);
nand U3611 (N_3611,N_526,N_1277);
nand U3612 (N_3612,N_4,N_2814);
nand U3613 (N_3613,N_452,N_1127);
and U3614 (N_3614,N_2767,N_2446);
nand U3615 (N_3615,N_280,N_1350);
and U3616 (N_3616,N_1209,N_1408);
or U3617 (N_3617,N_1297,N_292);
and U3618 (N_3618,N_1364,N_176);
and U3619 (N_3619,N_1859,N_332);
and U3620 (N_3620,N_2482,N_849);
or U3621 (N_3621,N_1022,N_561);
and U3622 (N_3622,N_2197,N_2759);
or U3623 (N_3623,N_1469,N_2457);
nand U3624 (N_3624,N_2151,N_593);
nand U3625 (N_3625,N_1064,N_2845);
and U3626 (N_3626,N_1806,N_869);
xor U3627 (N_3627,N_2697,N_1483);
or U3628 (N_3628,N_517,N_485);
or U3629 (N_3629,N_1746,N_378);
nor U3630 (N_3630,N_2337,N_1598);
or U3631 (N_3631,N_403,N_1791);
nand U3632 (N_3632,N_1737,N_1921);
and U3633 (N_3633,N_1222,N_1201);
nor U3634 (N_3634,N_1101,N_1795);
nor U3635 (N_3635,N_1711,N_277);
or U3636 (N_3636,N_2975,N_2387);
or U3637 (N_3637,N_2712,N_1155);
and U3638 (N_3638,N_775,N_912);
and U3639 (N_3639,N_1520,N_2418);
nand U3640 (N_3640,N_970,N_737);
nand U3641 (N_3641,N_1482,N_1752);
xor U3642 (N_3642,N_2136,N_2757);
nor U3643 (N_3643,N_958,N_192);
or U3644 (N_3644,N_1416,N_2662);
nand U3645 (N_3645,N_2969,N_704);
or U3646 (N_3646,N_2357,N_9);
nor U3647 (N_3647,N_2567,N_2803);
nor U3648 (N_3648,N_273,N_2021);
nor U3649 (N_3649,N_1356,N_618);
and U3650 (N_3650,N_325,N_345);
nor U3651 (N_3651,N_1149,N_1442);
or U3652 (N_3652,N_1607,N_2652);
xnor U3653 (N_3653,N_2943,N_2536);
nor U3654 (N_3654,N_2623,N_1883);
and U3655 (N_3655,N_402,N_2130);
xnor U3656 (N_3656,N_1886,N_2810);
nor U3657 (N_3657,N_2022,N_2141);
and U3658 (N_3658,N_450,N_2849);
or U3659 (N_3659,N_1814,N_2227);
and U3660 (N_3660,N_2750,N_392);
or U3661 (N_3661,N_14,N_2129);
nor U3662 (N_3662,N_1478,N_820);
nor U3663 (N_3663,N_2447,N_2559);
and U3664 (N_3664,N_2410,N_2973);
nor U3665 (N_3665,N_133,N_2171);
nand U3666 (N_3666,N_1605,N_2898);
and U3667 (N_3667,N_2964,N_187);
or U3668 (N_3668,N_371,N_1214);
or U3669 (N_3669,N_1302,N_1847);
and U3670 (N_3670,N_2811,N_2399);
nand U3671 (N_3671,N_2207,N_47);
or U3672 (N_3672,N_2850,N_339);
and U3673 (N_3673,N_288,N_261);
and U3674 (N_3674,N_832,N_1855);
nand U3675 (N_3675,N_2231,N_2545);
and U3676 (N_3676,N_794,N_1145);
nor U3677 (N_3677,N_1459,N_669);
nor U3678 (N_3678,N_2005,N_874);
and U3679 (N_3679,N_534,N_2282);
nand U3680 (N_3680,N_357,N_2326);
nor U3681 (N_3681,N_2762,N_2595);
or U3682 (N_3682,N_2978,N_1234);
nor U3683 (N_3683,N_988,N_698);
and U3684 (N_3684,N_186,N_637);
nand U3685 (N_3685,N_2921,N_1637);
or U3686 (N_3686,N_691,N_1263);
and U3687 (N_3687,N_2401,N_1196);
or U3688 (N_3688,N_776,N_991);
xor U3689 (N_3689,N_2391,N_1988);
nor U3690 (N_3690,N_1745,N_40);
nand U3691 (N_3691,N_1519,N_1175);
nand U3692 (N_3692,N_1856,N_2406);
nor U3693 (N_3693,N_1276,N_400);
and U3694 (N_3694,N_278,N_2624);
nand U3695 (N_3695,N_1845,N_2396);
nand U3696 (N_3696,N_2259,N_705);
and U3697 (N_3697,N_2905,N_367);
nand U3698 (N_3698,N_844,N_440);
nor U3699 (N_3699,N_2660,N_445);
or U3700 (N_3700,N_1063,N_1535);
nor U3701 (N_3701,N_1256,N_891);
nand U3702 (N_3702,N_2655,N_501);
nand U3703 (N_3703,N_806,N_673);
and U3704 (N_3704,N_322,N_2825);
nor U3705 (N_3705,N_1300,N_2692);
nor U3706 (N_3706,N_1489,N_2769);
or U3707 (N_3707,N_1283,N_2706);
nand U3708 (N_3708,N_826,N_1723);
nor U3709 (N_3709,N_2451,N_159);
and U3710 (N_3710,N_65,N_119);
and U3711 (N_3711,N_828,N_2948);
or U3712 (N_3712,N_1959,N_2142);
nand U3713 (N_3713,N_1344,N_2760);
or U3714 (N_3714,N_2330,N_2731);
nand U3715 (N_3715,N_2389,N_898);
or U3716 (N_3716,N_2042,N_479);
or U3717 (N_3717,N_537,N_2800);
nand U3718 (N_3718,N_2607,N_559);
and U3719 (N_3719,N_2928,N_2719);
nor U3720 (N_3720,N_2532,N_141);
nor U3721 (N_3721,N_2383,N_1262);
nand U3722 (N_3722,N_736,N_1616);
or U3723 (N_3723,N_51,N_2643);
nor U3724 (N_3724,N_2397,N_1699);
and U3725 (N_3725,N_1509,N_324);
and U3726 (N_3726,N_2727,N_2333);
nor U3727 (N_3727,N_2982,N_1721);
nand U3728 (N_3728,N_1917,N_1265);
or U3729 (N_3729,N_1766,N_498);
nand U3730 (N_3730,N_839,N_1040);
or U3731 (N_3731,N_1838,N_199);
nand U3732 (N_3732,N_1810,N_582);
nor U3733 (N_3733,N_2560,N_837);
and U3734 (N_3734,N_1666,N_604);
nand U3735 (N_3735,N_2489,N_2163);
nand U3736 (N_3736,N_83,N_478);
nor U3737 (N_3737,N_1786,N_1822);
nand U3738 (N_3738,N_2098,N_1651);
and U3739 (N_3739,N_96,N_643);
or U3740 (N_3740,N_1905,N_729);
nand U3741 (N_3741,N_722,N_2744);
nand U3742 (N_3742,N_2897,N_786);
xnor U3743 (N_3743,N_1515,N_2101);
xor U3744 (N_3744,N_132,N_2518);
nor U3745 (N_3745,N_1363,N_539);
and U3746 (N_3746,N_2718,N_772);
or U3747 (N_3747,N_1911,N_1094);
or U3748 (N_3748,N_1635,N_56);
and U3749 (N_3749,N_301,N_233);
nor U3750 (N_3750,N_2512,N_1529);
xor U3751 (N_3751,N_2950,N_762);
nand U3752 (N_3752,N_1153,N_2618);
or U3753 (N_3753,N_1461,N_1322);
nor U3754 (N_3754,N_1357,N_5);
nor U3755 (N_3755,N_397,N_1141);
and U3756 (N_3756,N_2881,N_313);
nor U3757 (N_3757,N_2983,N_328);
nor U3758 (N_3758,N_1396,N_2147);
or U3759 (N_3759,N_2768,N_2589);
or U3760 (N_3760,N_2090,N_2477);
nor U3761 (N_3761,N_364,N_2068);
and U3762 (N_3762,N_606,N_592);
nor U3763 (N_3763,N_726,N_1863);
nand U3764 (N_3764,N_540,N_1376);
or U3765 (N_3765,N_1097,N_223);
or U3766 (N_3766,N_1,N_1018);
and U3767 (N_3767,N_2131,N_2113);
nand U3768 (N_3768,N_2218,N_1966);
or U3769 (N_3769,N_1976,N_1784);
nand U3770 (N_3770,N_686,N_1091);
and U3771 (N_3771,N_1973,N_2214);
nand U3772 (N_3772,N_850,N_2404);
nor U3773 (N_3773,N_560,N_1705);
or U3774 (N_3774,N_1074,N_2514);
nand U3775 (N_3775,N_1947,N_2429);
or U3776 (N_3776,N_1190,N_960);
nand U3777 (N_3777,N_1181,N_95);
or U3778 (N_3778,N_995,N_1916);
or U3779 (N_3779,N_2440,N_205);
or U3780 (N_3780,N_1671,N_2378);
nor U3781 (N_3781,N_932,N_1642);
nand U3782 (N_3782,N_2099,N_1380);
or U3783 (N_3783,N_851,N_2046);
and U3784 (N_3784,N_64,N_354);
nand U3785 (N_3785,N_2294,N_2985);
nand U3786 (N_3786,N_1348,N_1619);
and U3787 (N_3787,N_2896,N_2255);
nor U3788 (N_3788,N_1610,N_1320);
or U3789 (N_3789,N_811,N_1217);
and U3790 (N_3790,N_1674,N_425);
or U3791 (N_3791,N_239,N_941);
nor U3792 (N_3792,N_295,N_948);
and U3793 (N_3793,N_2909,N_1663);
nand U3794 (N_3794,N_1578,N_1239);
nor U3795 (N_3795,N_2017,N_1279);
nand U3796 (N_3796,N_2193,N_1404);
nor U3797 (N_3797,N_1318,N_182);
nor U3798 (N_3798,N_1156,N_1005);
or U3799 (N_3799,N_2725,N_2903);
and U3800 (N_3800,N_2523,N_2954);
nor U3801 (N_3801,N_903,N_61);
or U3802 (N_3802,N_2121,N_1582);
nor U3803 (N_3803,N_123,N_1922);
and U3804 (N_3804,N_1079,N_1061);
or U3805 (N_3805,N_711,N_670);
or U3806 (N_3806,N_946,N_398);
nand U3807 (N_3807,N_1446,N_2752);
or U3808 (N_3808,N_2609,N_2691);
nand U3809 (N_3809,N_689,N_1683);
and U3810 (N_3810,N_1042,N_1028);
nor U3811 (N_3811,N_190,N_2931);
nand U3812 (N_3812,N_69,N_2182);
or U3813 (N_3813,N_253,N_2170);
or U3814 (N_3814,N_677,N_2016);
xor U3815 (N_3815,N_2540,N_2002);
nor U3816 (N_3816,N_1558,N_200);
nand U3817 (N_3817,N_1365,N_675);
and U3818 (N_3818,N_1874,N_1124);
nand U3819 (N_3819,N_2955,N_1208);
nor U3820 (N_3820,N_1212,N_1274);
or U3821 (N_3821,N_1241,N_864);
nand U3822 (N_3822,N_518,N_663);
nand U3823 (N_3823,N_2934,N_2749);
or U3824 (N_3824,N_904,N_2734);
and U3825 (N_3825,N_2432,N_1462);
or U3826 (N_3826,N_1913,N_535);
nand U3827 (N_3827,N_1467,N_2848);
or U3828 (N_3828,N_2458,N_1223);
nor U3829 (N_3829,N_2907,N_2952);
and U3830 (N_3830,N_2368,N_2998);
or U3831 (N_3831,N_2699,N_896);
and U3832 (N_3832,N_654,N_562);
or U3833 (N_3833,N_2439,N_2779);
xnor U3834 (N_3834,N_1877,N_1433);
nand U3835 (N_3835,N_2468,N_2286);
nand U3836 (N_3836,N_2474,N_464);
and U3837 (N_3837,N_2208,N_2386);
and U3838 (N_3838,N_1255,N_1889);
nand U3839 (N_3839,N_741,N_793);
xor U3840 (N_3840,N_2644,N_2919);
and U3841 (N_3841,N_1649,N_2119);
or U3842 (N_3842,N_1333,N_2072);
and U3843 (N_3843,N_2577,N_2871);
or U3844 (N_3844,N_1761,N_1349);
and U3845 (N_3845,N_2096,N_2704);
or U3846 (N_3846,N_1869,N_1780);
nor U3847 (N_3847,N_1564,N_996);
and U3848 (N_3848,N_2895,N_1989);
nor U3849 (N_3849,N_2966,N_2367);
nor U3850 (N_3850,N_2144,N_512);
or U3851 (N_3851,N_2641,N_431);
and U3852 (N_3852,N_2161,N_198);
or U3853 (N_3853,N_49,N_802);
nand U3854 (N_3854,N_1848,N_684);
or U3855 (N_3855,N_2036,N_1479);
nand U3856 (N_3856,N_2013,N_2476);
nand U3857 (N_3857,N_764,N_751);
or U3858 (N_3858,N_314,N_1240);
nand U3859 (N_3859,N_1601,N_145);
nand U3860 (N_3860,N_2283,N_2488);
xor U3861 (N_3861,N_2247,N_1151);
or U3862 (N_3862,N_204,N_2264);
or U3863 (N_3863,N_2703,N_125);
xnor U3864 (N_3864,N_2030,N_2258);
and U3865 (N_3865,N_1293,N_2773);
or U3866 (N_3866,N_919,N_2284);
and U3867 (N_3867,N_1650,N_153);
nor U3868 (N_3868,N_1272,N_203);
nor U3869 (N_3869,N_1830,N_413);
or U3870 (N_3870,N_1186,N_2424);
nor U3871 (N_3871,N_2807,N_463);
or U3872 (N_3872,N_2552,N_1014);
nand U3873 (N_3873,N_1923,N_1392);
and U3874 (N_3874,N_2185,N_1170);
and U3875 (N_3875,N_2327,N_734);
and U3876 (N_3876,N_752,N_2696);
nor U3877 (N_3877,N_1720,N_553);
nand U3878 (N_3878,N_387,N_1207);
nor U3879 (N_3879,N_2606,N_290);
nor U3880 (N_3880,N_495,N_945);
and U3881 (N_3881,N_1345,N_459);
and U3882 (N_3882,N_2700,N_2786);
or U3883 (N_3883,N_2069,N_655);
nor U3884 (N_3884,N_241,N_1727);
nand U3885 (N_3885,N_2645,N_2513);
nor U3886 (N_3886,N_1832,N_1390);
or U3887 (N_3887,N_2884,N_1897);
or U3888 (N_3888,N_2576,N_816);
and U3889 (N_3889,N_2279,N_2205);
xor U3890 (N_3890,N_907,N_2511);
and U3891 (N_3891,N_1336,N_262);
nand U3892 (N_3892,N_2159,N_1915);
nand U3893 (N_3893,N_876,N_2739);
nand U3894 (N_3894,N_1289,N_2780);
nand U3895 (N_3895,N_1861,N_2438);
or U3896 (N_3896,N_1690,N_1353);
nand U3897 (N_3897,N_2395,N_2537);
and U3898 (N_3898,N_1772,N_1473);
or U3899 (N_3899,N_2863,N_2172);
or U3900 (N_3900,N_1056,N_2957);
and U3901 (N_3901,N_2735,N_1374);
or U3902 (N_3902,N_1692,N_723);
or U3903 (N_3903,N_1298,N_2495);
or U3904 (N_3904,N_491,N_766);
nand U3905 (N_3905,N_1311,N_1499);
xor U3906 (N_3906,N_1282,N_1839);
and U3907 (N_3907,N_16,N_950);
or U3908 (N_3908,N_20,N_2083);
or U3909 (N_3909,N_1395,N_191);
or U3910 (N_3910,N_1334,N_79);
nor U3911 (N_3911,N_823,N_2528);
or U3912 (N_3912,N_765,N_2289);
and U3913 (N_3913,N_2498,N_1343);
nand U3914 (N_3914,N_285,N_2122);
nor U3915 (N_3915,N_1324,N_1154);
nand U3916 (N_3916,N_2808,N_1999);
nand U3917 (N_3917,N_311,N_1596);
or U3918 (N_3918,N_1144,N_206);
or U3919 (N_3919,N_1335,N_1534);
nor U3920 (N_3920,N_1231,N_810);
nor U3921 (N_3921,N_2596,N_2422);
nor U3922 (N_3922,N_150,N_829);
and U3923 (N_3923,N_2546,N_2273);
nand U3924 (N_3924,N_2942,N_368);
nand U3925 (N_3925,N_1851,N_2547);
nand U3926 (N_3926,N_1807,N_522);
nor U3927 (N_3927,N_1945,N_709);
nor U3928 (N_3928,N_1117,N_1472);
nor U3929 (N_3929,N_875,N_2664);
and U3930 (N_3930,N_2267,N_2906);
nor U3931 (N_3931,N_2063,N_2232);
or U3932 (N_3932,N_603,N_1049);
or U3933 (N_3933,N_1329,N_2325);
nand U3934 (N_3934,N_2772,N_1273);
or U3935 (N_3935,N_1958,N_1657);
nor U3936 (N_3936,N_183,N_126);
and U3937 (N_3937,N_1072,N_1169);
or U3938 (N_3938,N_1621,N_1581);
nor U3939 (N_3939,N_2506,N_1700);
and U3940 (N_3940,N_2633,N_1835);
and U3941 (N_3941,N_1464,N_989);
nand U3942 (N_3942,N_2224,N_468);
nor U3943 (N_3943,N_2107,N_1456);
nor U3944 (N_3944,N_2585,N_2164);
nor U3945 (N_3945,N_2365,N_152);
nor U3946 (N_3946,N_1824,N_1176);
nor U3947 (N_3947,N_682,N_147);
or U3948 (N_3948,N_2702,N_2026);
xor U3949 (N_3949,N_1371,N_43);
nor U3950 (N_3950,N_1625,N_10);
nand U3951 (N_3951,N_2360,N_2561);
nand U3952 (N_3952,N_2710,N_2938);
nor U3953 (N_3953,N_370,N_1338);
nor U3954 (N_3954,N_2157,N_2812);
and U3955 (N_3955,N_2565,N_2319);
or U3956 (N_3956,N_29,N_2312);
or U3957 (N_3957,N_2493,N_909);
nand U3958 (N_3958,N_2292,N_857);
nand U3959 (N_3959,N_2781,N_835);
and U3960 (N_3960,N_1160,N_2716);
nor U3961 (N_3961,N_664,N_2376);
nand U3962 (N_3962,N_1113,N_1698);
nor U3963 (N_3963,N_2443,N_102);
nor U3964 (N_3964,N_1310,N_1813);
nor U3965 (N_3965,N_2951,N_366);
nor U3966 (N_3966,N_236,N_2434);
xor U3967 (N_3967,N_1397,N_2846);
nor U3968 (N_3968,N_956,N_25);
nand U3969 (N_3969,N_1708,N_7);
and U3970 (N_3970,N_859,N_1867);
and U3971 (N_3971,N_2150,N_209);
and U3972 (N_3972,N_2971,N_2999);
nor U3973 (N_3973,N_818,N_476);
xor U3974 (N_3974,N_1178,N_381);
and U3975 (N_3975,N_81,N_1949);
and U3976 (N_3976,N_1562,N_1452);
and U3977 (N_3977,N_2714,N_249);
nand U3978 (N_3978,N_1836,N_2038);
nand U3979 (N_3979,N_2516,N_2778);
and U3980 (N_3980,N_1161,N_2138);
and U3981 (N_3981,N_2894,N_417);
nor U3982 (N_3982,N_2730,N_2338);
and U3983 (N_3983,N_623,N_2436);
nor U3984 (N_3984,N_1788,N_447);
nand U3985 (N_3985,N_1098,N_2211);
nor U3986 (N_3986,N_927,N_2503);
and U3987 (N_3987,N_2979,N_1678);
nor U3988 (N_3988,N_455,N_2746);
nor U3989 (N_3989,N_923,N_747);
xnor U3990 (N_3990,N_1753,N_136);
and U3991 (N_3991,N_1925,N_2344);
or U3992 (N_3992,N_363,N_2632);
nand U3993 (N_3993,N_1754,N_1517);
nor U3994 (N_3994,N_2230,N_538);
nand U3995 (N_3995,N_2009,N_2233);
nand U3996 (N_3996,N_1853,N_1183);
and U3997 (N_3997,N_1206,N_2270);
or U3998 (N_3998,N_1266,N_1387);
nor U3999 (N_3999,N_2717,N_838);
and U4000 (N_4000,N_134,N_2960);
and U4001 (N_4001,N_542,N_785);
nand U4002 (N_4002,N_1321,N_259);
nor U4003 (N_4003,N_1512,N_962);
xnor U4004 (N_4004,N_320,N_617);
or U4005 (N_4005,N_1732,N_1229);
or U4006 (N_4006,N_2569,N_1332);
nor U4007 (N_4007,N_24,N_1491);
nand U4008 (N_4008,N_2533,N_554);
nor U4009 (N_4009,N_1086,N_2806);
and U4010 (N_4010,N_930,N_974);
or U4011 (N_4011,N_89,N_2694);
or U4012 (N_4012,N_1399,N_1470);
nor U4013 (N_4013,N_2824,N_1812);
nand U4014 (N_4014,N_957,N_151);
or U4015 (N_4015,N_2266,N_2920);
nor U4016 (N_4016,N_1748,N_2911);
or U4017 (N_4017,N_2771,N_481);
nor U4018 (N_4018,N_1354,N_1199);
nand U4019 (N_4019,N_2787,N_702);
nor U4020 (N_4020,N_863,N_1546);
nor U4021 (N_4021,N_2202,N_2711);
nand U4022 (N_4022,N_1121,N_1465);
and U4023 (N_4023,N_1505,N_2411);
nand U4024 (N_4024,N_1695,N_2667);
and U4025 (N_4025,N_127,N_2305);
or U4026 (N_4026,N_2242,N_2874);
nand U4027 (N_4027,N_2139,N_220);
or U4028 (N_4028,N_369,N_1437);
nor U4029 (N_4029,N_2570,N_1215);
and U4030 (N_4030,N_1131,N_1903);
or U4031 (N_4031,N_1603,N_596);
or U4032 (N_4032,N_309,N_2841);
and U4033 (N_4033,N_555,N_1568);
nor U4034 (N_4034,N_900,N_1606);
nand U4035 (N_4035,N_271,N_544);
nor U4036 (N_4036,N_1525,N_790);
or U4037 (N_4037,N_2915,N_2657);
nand U4038 (N_4038,N_2300,N_2524);
or U4039 (N_4039,N_2777,N_2766);
and U4040 (N_4040,N_905,N_1346);
or U4041 (N_4041,N_2984,N_940);
or U4042 (N_4042,N_2256,N_2234);
and U4043 (N_4043,N_207,N_2648);
and U4044 (N_4044,N_2006,N_2460);
nand U4045 (N_4045,N_650,N_1738);
nand U4046 (N_4046,N_910,N_1599);
nor U4047 (N_4047,N_1045,N_2088);
nor U4048 (N_4048,N_1157,N_2584);
and U4049 (N_4049,N_421,N_701);
or U4050 (N_4050,N_2804,N_1771);
or U4051 (N_4051,N_2509,N_821);
or U4052 (N_4052,N_283,N_2276);
or U4053 (N_4053,N_1219,N_1816);
or U4054 (N_4054,N_2989,N_1419);
and U4055 (N_4055,N_2754,N_1102);
nand U4056 (N_4056,N_929,N_653);
and U4057 (N_4057,N_579,N_2538);
nor U4058 (N_4058,N_757,N_86);
nor U4059 (N_4059,N_2669,N_11);
or U4060 (N_4060,N_263,N_800);
and U4061 (N_4061,N_408,N_1537);
nor U4062 (N_4062,N_2226,N_1950);
nand U4063 (N_4063,N_287,N_1129);
and U4064 (N_4064,N_1906,N_1301);
nand U4065 (N_4065,N_488,N_2050);
nor U4066 (N_4066,N_972,N_130);
or U4067 (N_4067,N_2379,N_897);
or U4068 (N_4068,N_420,N_2124);
and U4069 (N_4069,N_1944,N_2385);
nor U4070 (N_4070,N_2592,N_2843);
and U4071 (N_4071,N_146,N_624);
nor U4072 (N_4072,N_1561,N_2953);
nor U4073 (N_4073,N_2614,N_2097);
nand U4074 (N_4074,N_2271,N_1837);
nand U4075 (N_4075,N_82,N_2882);
nor U4076 (N_4076,N_1032,N_583);
or U4077 (N_4077,N_216,N_222);
and U4078 (N_4078,N_169,N_759);
and U4079 (N_4079,N_195,N_1174);
or U4080 (N_4080,N_1978,N_2078);
or U4081 (N_4081,N_1541,N_2821);
or U4082 (N_4082,N_888,N_2851);
nor U4083 (N_4083,N_348,N_548);
nor U4084 (N_4084,N_2057,N_505);
nand U4085 (N_4085,N_1138,N_2748);
or U4086 (N_4086,N_1474,N_2822);
and U4087 (N_4087,N_2296,N_284);
or U4088 (N_4088,N_1602,N_340);
and U4089 (N_4089,N_2548,N_2794);
nor U4090 (N_4090,N_2961,N_282);
nand U4091 (N_4091,N_457,N_2445);
nand U4092 (N_4092,N_2195,N_1378);
nor U4093 (N_4093,N_2525,N_2631);
nand U4094 (N_4094,N_1052,N_1062);
and U4095 (N_4095,N_128,N_2526);
nand U4096 (N_4096,N_1774,N_2801);
or U4097 (N_4097,N_2,N_1105);
nand U4098 (N_4098,N_1152,N_94);
or U4099 (N_4099,N_80,N_1490);
nand U4100 (N_4100,N_2939,N_1739);
nand U4101 (N_4101,N_2566,N_2726);
or U4102 (N_4102,N_2321,N_1476);
or U4103 (N_4103,N_2135,N_1264);
xnor U4104 (N_4104,N_2165,N_1660);
nand U4105 (N_4105,N_2611,N_1734);
or U4106 (N_4106,N_2452,N_2014);
or U4107 (N_4107,N_954,N_112);
and U4108 (N_4108,N_1104,N_2729);
nand U4109 (N_4109,N_966,N_2868);
and U4110 (N_4110,N_607,N_2784);
and U4111 (N_4111,N_442,N_2958);
and U4112 (N_4112,N_1290,N_338);
and U4113 (N_4113,N_1571,N_610);
nand U4114 (N_4114,N_771,N_2970);
nand U4115 (N_4115,N_1555,N_1046);
nand U4116 (N_4116,N_1799,N_882);
nor U4117 (N_4117,N_531,N_782);
and U4118 (N_4118,N_969,N_1591);
nor U4119 (N_4119,N_725,N_1254);
and U4120 (N_4120,N_753,N_651);
or U4121 (N_4121,N_2110,N_744);
or U4122 (N_4122,N_482,N_1044);
nor U4123 (N_4123,N_2134,N_2941);
nor U4124 (N_4124,N_260,N_2674);
nor U4125 (N_4125,N_2194,N_2260);
or U4126 (N_4126,N_564,N_990);
nand U4127 (N_4127,N_35,N_1707);
nor U4128 (N_4128,N_2178,N_1171);
or U4129 (N_4129,N_1164,N_2275);
nor U4130 (N_4130,N_1115,N_1677);
and U4131 (N_4131,N_1009,N_213);
and U4132 (N_4132,N_2133,N_640);
and U4133 (N_4133,N_2542,N_616);
and U4134 (N_4134,N_884,N_984);
or U4135 (N_4135,N_2743,N_1358);
nor U4136 (N_4136,N_911,N_1567);
nand U4137 (N_4137,N_585,N_475);
xnor U4138 (N_4138,N_34,N_1865);
and U4139 (N_4139,N_658,N_2680);
nor U4140 (N_4140,N_2977,N_2058);
or U4141 (N_4141,N_1712,N_1339);
or U4142 (N_4142,N_2673,N_1111);
nor U4143 (N_4143,N_2878,N_302);
or U4144 (N_4144,N_1013,N_2469);
or U4145 (N_4145,N_2148,N_2473);
or U4146 (N_4146,N_490,N_1447);
or U4147 (N_4147,N_1012,N_2908);
nor U4148 (N_4148,N_2306,N_2039);
and U4149 (N_4149,N_1938,N_1724);
or U4150 (N_4150,N_2886,N_2210);
and U4151 (N_4151,N_1412,N_1679);
or U4152 (N_4152,N_2601,N_2416);
xor U4153 (N_4153,N_393,N_493);
and U4154 (N_4154,N_1592,N_1544);
or U4155 (N_4155,N_1881,N_639);
nor U4156 (N_4156,N_740,N_2229);
nand U4157 (N_4157,N_2079,N_2630);
and U4158 (N_4158,N_171,N_1486);
or U4159 (N_4159,N_1248,N_437);
nor U4160 (N_4160,N_1314,N_2272);
or U4161 (N_4161,N_2491,N_1427);
or U4162 (N_4162,N_1439,N_1685);
nor U4163 (N_4163,N_1530,N_2636);
or U4164 (N_4164,N_1033,N_2407);
and U4165 (N_4165,N_2342,N_901);
or U4166 (N_4166,N_1629,N_315);
nand U4167 (N_4167,N_2183,N_2361);
and U4168 (N_4168,N_2423,N_2872);
nor U4169 (N_4169,N_1498,N_858);
nand U4170 (N_4170,N_2132,N_2879);
or U4171 (N_4171,N_1689,N_2962);
and U4172 (N_4172,N_1818,N_2052);
or U4173 (N_4173,N_976,N_1914);
nand U4174 (N_4174,N_1726,N_1995);
or U4175 (N_4175,N_1749,N_2200);
and U4176 (N_4176,N_208,N_2011);
nor U4177 (N_4177,N_120,N_2206);
nand U4178 (N_4178,N_2166,N_1165);
or U4179 (N_4179,N_521,N_2840);
nor U4180 (N_4180,N_2012,N_566);
or U4181 (N_4181,N_1048,N_1778);
or U4182 (N_4182,N_2558,N_1623);
nor U4183 (N_4183,N_347,N_2721);
or U4184 (N_4184,N_1039,N_2838);
or U4185 (N_4185,N_1878,N_269);
or U4186 (N_4186,N_1532,N_1593);
or U4187 (N_4187,N_1518,N_1253);
and U4188 (N_4188,N_1744,N_951);
and U4189 (N_4189,N_2073,N_1595);
and U4190 (N_4190,N_1560,N_2167);
and U4191 (N_4191,N_2720,N_1352);
nand U4192 (N_4192,N_2065,N_1576);
and U4193 (N_4193,N_137,N_1783);
nand U4194 (N_4194,N_2212,N_738);
nor U4195 (N_4195,N_1893,N_299);
and U4196 (N_4196,N_2776,N_2238);
nor U4197 (N_4197,N_2191,N_2722);
and U4198 (N_4198,N_2986,N_1257);
nand U4199 (N_4199,N_215,N_389);
or U4200 (N_4200,N_2128,N_2123);
or U4201 (N_4201,N_1862,N_2956);
nand U4202 (N_4202,N_2600,N_1785);
nand U4203 (N_4203,N_1782,N_1341);
and U4204 (N_4204,N_1985,N_2085);
nand U4205 (N_4205,N_1405,N_895);
or U4206 (N_4206,N_2981,N_138);
nand U4207 (N_4207,N_924,N_2996);
nor U4208 (N_4208,N_1020,N_310);
and U4209 (N_4209,N_1415,N_1858);
or U4210 (N_4210,N_926,N_2263);
nor U4211 (N_4211,N_2114,N_37);
nor U4212 (N_4212,N_980,N_2127);
xor U4213 (N_4213,N_38,N_1890);
or U4214 (N_4214,N_1627,N_1641);
or U4215 (N_4215,N_975,N_2695);
and U4216 (N_4216,N_1521,N_202);
nor U4217 (N_4217,N_2575,N_2464);
or U4218 (N_4218,N_2708,N_2728);
nor U4219 (N_4219,N_1047,N_645);
or U4220 (N_4220,N_967,N_2932);
and U4221 (N_4221,N_1454,N_1285);
nand U4222 (N_4222,N_1025,N_854);
nand U4223 (N_4223,N_2347,N_1844);
nor U4224 (N_4224,N_1444,N_2847);
and U4225 (N_4225,N_465,N_2972);
or U4226 (N_4226,N_716,N_649);
nor U4227 (N_4227,N_1997,N_312);
and U4228 (N_4228,N_981,N_237);
nand U4229 (N_4229,N_335,N_1148);
or U4230 (N_4230,N_365,N_1557);
xor U4231 (N_4231,N_298,N_1667);
and U4232 (N_4232,N_2025,N_787);
and U4233 (N_4233,N_1401,N_2177);
and U4234 (N_4234,N_2071,N_1011);
and U4235 (N_4235,N_2465,N_2813);
xnor U4236 (N_4236,N_2353,N_584);
nor U4237 (N_4237,N_2430,N_2420);
or U4238 (N_4238,N_2535,N_2461);
nor U4239 (N_4239,N_1425,N_2426);
and U4240 (N_4240,N_1180,N_1007);
and U4241 (N_4241,N_589,N_1888);
and U4242 (N_4242,N_2448,N_1445);
or U4243 (N_4243,N_2111,N_1213);
nand U4244 (N_4244,N_333,N_594);
and U4245 (N_4245,N_605,N_1184);
nor U4246 (N_4246,N_226,N_2154);
and U4247 (N_4247,N_1147,N_2504);
or U4248 (N_4248,N_2568,N_166);
or U4249 (N_4249,N_173,N_1159);
or U4250 (N_4250,N_108,N_489);
and U4251 (N_4251,N_1693,N_129);
nor U4252 (N_4252,N_1755,N_483);
nor U4253 (N_4253,N_376,N_60);
and U4254 (N_4254,N_240,N_1800);
or U4255 (N_4255,N_2625,N_66);
nor U4256 (N_4256,N_1547,N_2758);
nand U4257 (N_4257,N_1377,N_680);
nor U4258 (N_4258,N_552,N_2158);
and U4259 (N_4259,N_1382,N_2574);
nand U4260 (N_4260,N_1762,N_419);
or U4261 (N_4261,N_449,N_2828);
nor U4262 (N_4262,N_524,N_2990);
or U4263 (N_4263,N_1805,N_1389);
nand U4264 (N_4264,N_1531,N_1808);
nand U4265 (N_4265,N_2763,N_1187);
nor U4266 (N_4266,N_374,N_1070);
nand U4267 (N_4267,N_661,N_2186);
and U4268 (N_4268,N_2278,N_2095);
nand U4269 (N_4269,N_964,N_2350);
and U4270 (N_4270,N_350,N_570);
nor U4271 (N_4271,N_2108,N_227);
nand U4272 (N_4272,N_154,N_917);
nor U4273 (N_4273,N_1323,N_1912);
or U4274 (N_4274,N_1992,N_1714);
and U4275 (N_4275,N_2315,N_2642);
nand U4276 (N_4276,N_500,N_2742);
or U4277 (N_4277,N_1730,N_2299);
nand U4278 (N_4278,N_791,N_2160);
or U4279 (N_4279,N_2045,N_303);
and U4280 (N_4280,N_1961,N_2285);
or U4281 (N_4281,N_1980,N_2007);
or U4282 (N_4282,N_2765,N_1579);
nor U4283 (N_4283,N_2940,N_1891);
or U4284 (N_4284,N_1200,N_229);
nor U4285 (N_4285,N_2298,N_706);
and U4286 (N_4286,N_2074,N_12);
or U4287 (N_4287,N_1460,N_1991);
nand U4288 (N_4288,N_2571,N_2698);
nor U4289 (N_4289,N_1488,N_822);
nand U4290 (N_4290,N_2453,N_85);
nor U4291 (N_4291,N_383,N_1394);
xor U4292 (N_4292,N_514,N_1026);
nand U4293 (N_4293,N_1608,N_629);
nand U4294 (N_4294,N_2637,N_1275);
nor U4295 (N_4295,N_453,N_575);
nor U4296 (N_4296,N_256,N_2873);
nor U4297 (N_4297,N_1493,N_264);
and U4298 (N_4298,N_2308,N_1728);
or U4299 (N_4299,N_2826,N_1823);
nand U4300 (N_4300,N_1398,N_1367);
or U4301 (N_4301,N_1092,N_1787);
and U4302 (N_4302,N_2867,N_2988);
or U4303 (N_4303,N_922,N_396);
or U4304 (N_4304,N_2668,N_1327);
nor U4305 (N_4305,N_62,N_1793);
or U4306 (N_4306,N_1043,N_2249);
and U4307 (N_4307,N_2507,N_2861);
and U4308 (N_4308,N_1640,N_471);
and U4309 (N_4309,N_2639,N_30);
or U4310 (N_4310,N_1887,N_228);
and U4311 (N_4311,N_2475,N_1526);
nand U4312 (N_4312,N_708,N_2967);
nand U4313 (N_4313,N_1556,N_827);
or U4314 (N_4314,N_768,N_1542);
or U4315 (N_4315,N_2676,N_1609);
and U4316 (N_4316,N_683,N_2261);
nand U4317 (N_4317,N_632,N_2484);
nor U4318 (N_4318,N_2106,N_1386);
or U4319 (N_4319,N_17,N_326);
xnor U4320 (N_4320,N_2223,N_621);
nand U4321 (N_4321,N_2675,N_1941);
nand U4322 (N_4322,N_572,N_1803);
nor U4323 (N_4323,N_1023,N_721);
nand U4324 (N_4324,N_2653,N_2228);
nand U4325 (N_4325,N_1359,N_1731);
xnor U4326 (N_4326,N_224,N_1511);
nor U4327 (N_4327,N_963,N_2889);
and U4328 (N_4328,N_2001,N_386);
nand U4329 (N_4329,N_1233,N_2362);
and U4330 (N_4330,N_2257,N_404);
nand U4331 (N_4331,N_2980,N_2834);
xnor U4332 (N_4332,N_2741,N_2381);
and U4333 (N_4333,N_2091,N_180);
or U4334 (N_4334,N_1831,N_2580);
nand U4335 (N_4335,N_319,N_693);
nor U4336 (N_4336,N_45,N_401);
nor U4337 (N_4337,N_2254,N_41);
and U4338 (N_4338,N_892,N_2613);
nand U4339 (N_4339,N_1636,N_1974);
nand U4340 (N_4340,N_8,N_441);
and U4341 (N_4341,N_1777,N_2890);
nand U4342 (N_4342,N_92,N_769);
nand U4343 (N_4343,N_2926,N_1937);
nor U4344 (N_4344,N_1960,N_294);
or U4345 (N_4345,N_1177,N_2455);
nand U4346 (N_4346,N_432,N_862);
and U4347 (N_4347,N_1681,N_1429);
nand U4348 (N_4348,N_2818,N_631);
xor U4349 (N_4349,N_2265,N_792);
and U4350 (N_4350,N_2444,N_2146);
and U4351 (N_4351,N_947,N_2550);
and U4352 (N_4352,N_530,N_439);
xnor U4353 (N_4353,N_674,N_117);
or U4354 (N_4354,N_1964,N_1286);
and U4355 (N_4355,N_1030,N_353);
and U4356 (N_4356,N_100,N_1244);
nand U4357 (N_4357,N_1828,N_568);
nand U4358 (N_4358,N_188,N_2201);
and U4359 (N_4359,N_2393,N_55);
nand U4360 (N_4360,N_667,N_824);
nand U4361 (N_4361,N_2280,N_1569);
nor U4362 (N_4362,N_179,N_1527);
or U4363 (N_4363,N_474,N_887);
or U4364 (N_4364,N_2441,N_1370);
and U4365 (N_4365,N_1524,N_2417);
nor U4366 (N_4366,N_1841,N_2929);
nand U4367 (N_4367,N_2597,N_57);
and U4368 (N_4368,N_1825,N_2852);
or U4369 (N_4369,N_1583,N_1027);
nor U4370 (N_4370,N_1430,N_1655);
or U4371 (N_4371,N_31,N_499);
nand U4372 (N_4372,N_1968,N_1899);
nor U4373 (N_4373,N_337,N_523);
and U4374 (N_4374,N_2035,N_994);
or U4375 (N_4375,N_614,N_2968);
and U4376 (N_4376,N_2055,N_1291);
or U4377 (N_4377,N_487,N_633);
nor U4378 (N_4378,N_550,N_189);
nor U4379 (N_4379,N_1003,N_394);
and U4380 (N_4380,N_1919,N_2405);
or U4381 (N_4381,N_2421,N_2761);
nand U4382 (N_4382,N_2963,N_1733);
and U4383 (N_4383,N_2774,N_466);
nand U4384 (N_4384,N_297,N_732);
or U4385 (N_4385,N_2414,N_225);
nor U4386 (N_4386,N_342,N_424);
or U4387 (N_4387,N_1450,N_1719);
nor U4388 (N_4388,N_1866,N_1702);
nor U4389 (N_4389,N_1211,N_1379);
and U4390 (N_4390,N_2922,N_2225);
nor U4391 (N_4391,N_1688,N_2870);
or U4392 (N_4392,N_1295,N_2481);
or U4393 (N_4393,N_1939,N_1604);
and U4394 (N_4394,N_2467,N_506);
nor U4395 (N_4395,N_1220,N_1084);
or U4396 (N_4396,N_2510,N_496);
and U4397 (N_4397,N_2505,N_2281);
or U4398 (N_4398,N_1827,N_2262);
or U4399 (N_4399,N_1536,N_2359);
nor U4400 (N_4400,N_212,N_2740);
nand U4401 (N_4401,N_678,N_2034);
nor U4402 (N_4402,N_1951,N_2887);
nor U4403 (N_4403,N_219,N_78);
or U4404 (N_4404,N_2316,N_456);
nor U4405 (N_4405,N_2437,N_853);
nand U4406 (N_4406,N_2805,N_641);
nand U4407 (N_4407,N_656,N_1781);
nor U4408 (N_4408,N_2173,N_377);
nor U4409 (N_4409,N_871,N_2190);
nor U4410 (N_4410,N_2993,N_836);
xor U4411 (N_4411,N_899,N_1981);
or U4412 (N_4412,N_1664,N_359);
and U4413 (N_4413,N_341,N_232);
nand U4414 (N_4414,N_1075,N_1243);
nor U4415 (N_4415,N_6,N_1258);
and U4416 (N_4416,N_2497,N_252);
or U4417 (N_4417,N_739,N_2168);
and U4418 (N_4418,N_2622,N_1133);
nand U4419 (N_4419,N_1768,N_1930);
nor U4420 (N_4420,N_1504,N_13);
and U4421 (N_4421,N_1480,N_819);
and U4422 (N_4422,N_2179,N_1312);
or U4423 (N_4423,N_1410,N_2658);
nand U4424 (N_4424,N_1093,N_2169);
and U4425 (N_4425,N_77,N_1885);
nor U4426 (N_4426,N_602,N_407);
or U4427 (N_4427,N_710,N_142);
nor U4428 (N_4428,N_2145,N_1114);
nand U4429 (N_4429,N_1103,N_1918);
and U4430 (N_4430,N_1317,N_2117);
xnor U4431 (N_4431,N_2530,N_380);
or U4432 (N_4432,N_551,N_2853);
nand U4433 (N_4433,N_2995,N_1251);
xnor U4434 (N_4434,N_230,N_444);
or U4435 (N_4435,N_2087,N_2612);
nor U4436 (N_4436,N_2398,N_317);
and U4437 (N_4437,N_1910,N_0);
and U4438 (N_4438,N_2311,N_1852);
nand U4439 (N_4439,N_1545,N_2997);
and U4440 (N_4440,N_1566,N_395);
nand U4441 (N_4441,N_175,N_2268);
nor U4442 (N_4442,N_719,N_2933);
nor U4443 (N_4443,N_803,N_1252);
nor U4444 (N_4444,N_1422,N_2303);
and U4445 (N_4445,N_473,N_2374);
nor U4446 (N_4446,N_660,N_1570);
nor U4447 (N_4447,N_1850,N_1216);
and U4448 (N_4448,N_2785,N_349);
nor U4449 (N_4449,N_2572,N_1654);
nand U4450 (N_4450,N_2991,N_2551);
nand U4451 (N_4451,N_334,N_953);
or U4452 (N_4452,N_2935,N_1194);
nor U4453 (N_4453,N_272,N_2534);
nor U4454 (N_4454,N_27,N_713);
and U4455 (N_4455,N_1232,N_1168);
and U4456 (N_4456,N_306,N_434);
nand U4457 (N_4457,N_1809,N_1996);
and U4458 (N_4458,N_949,N_75);
nor U4459 (N_4459,N_1383,N_1528);
or U4460 (N_4460,N_2112,N_1802);
or U4461 (N_4461,N_210,N_1191);
nand U4462 (N_4462,N_855,N_944);
and U4463 (N_4463,N_2520,N_833);
nor U4464 (N_4464,N_968,N_2181);
or U4465 (N_4465,N_1857,N_356);
or U4466 (N_4466,N_1709,N_140);
nor U4467 (N_4467,N_430,N_687);
nand U4468 (N_4468,N_727,N_2314);
nand U4469 (N_4469,N_2033,N_1834);
nor U4470 (N_4470,N_2301,N_2246);
nand U4471 (N_4471,N_1418,N_124);
nor U4472 (N_4472,N_1403,N_1342);
xor U4473 (N_4473,N_2435,N_1826);
and U4474 (N_4474,N_2923,N_155);
nand U4475 (N_4475,N_1539,N_1644);
or U4476 (N_4476,N_504,N_843);
or U4477 (N_4477,N_587,N_2864);
or U4478 (N_4478,N_1742,N_2373);
nand U4479 (N_4479,N_1931,N_2176);
or U4480 (N_4480,N_1600,N_2274);
or U4481 (N_4481,N_1758,N_1868);
nand U4482 (N_4482,N_2608,N_2174);
or U4483 (N_4483,N_1955,N_2549);
nor U4484 (N_4484,N_2602,N_796);
nand U4485 (N_4485,N_50,N_1089);
or U4486 (N_4486,N_2965,N_2588);
nor U4487 (N_4487,N_1588,N_931);
or U4488 (N_4488,N_2479,N_2770);
or U4489 (N_4489,N_2340,N_1633);
or U4490 (N_4490,N_428,N_2019);
or U4491 (N_4491,N_1896,N_1041);
or U4492 (N_4492,N_415,N_1287);
nand U4493 (N_4493,N_1021,N_1135);
nor U4494 (N_4494,N_2086,N_939);
nor U4495 (N_4495,N_1162,N_1085);
or U4496 (N_4496,N_2293,N_1565);
or U4497 (N_4497,N_1017,N_243);
nor U4498 (N_4498,N_2336,N_581);
and U4499 (N_4499,N_1428,N_1494);
nand U4500 (N_4500,N_2185,N_1544);
or U4501 (N_4501,N_772,N_505);
nand U4502 (N_4502,N_47,N_474);
xor U4503 (N_4503,N_108,N_2758);
nor U4504 (N_4504,N_683,N_1313);
xor U4505 (N_4505,N_1090,N_203);
nand U4506 (N_4506,N_556,N_812);
and U4507 (N_4507,N_1520,N_2347);
nor U4508 (N_4508,N_2588,N_1833);
nand U4509 (N_4509,N_2042,N_1451);
nor U4510 (N_4510,N_703,N_1987);
nand U4511 (N_4511,N_623,N_1716);
or U4512 (N_4512,N_1827,N_1284);
nand U4513 (N_4513,N_2301,N_936);
or U4514 (N_4514,N_1146,N_1433);
or U4515 (N_4515,N_1747,N_2163);
nor U4516 (N_4516,N_494,N_805);
nand U4517 (N_4517,N_596,N_704);
xor U4518 (N_4518,N_1586,N_2912);
nor U4519 (N_4519,N_2121,N_102);
or U4520 (N_4520,N_2941,N_1565);
or U4521 (N_4521,N_2760,N_2209);
nand U4522 (N_4522,N_2621,N_240);
nand U4523 (N_4523,N_1084,N_85);
and U4524 (N_4524,N_1868,N_2239);
or U4525 (N_4525,N_2099,N_2976);
nor U4526 (N_4526,N_2723,N_2795);
nand U4527 (N_4527,N_1151,N_1422);
and U4528 (N_4528,N_1448,N_2466);
nor U4529 (N_4529,N_2206,N_63);
or U4530 (N_4530,N_1299,N_2367);
nand U4531 (N_4531,N_1579,N_1649);
xor U4532 (N_4532,N_2818,N_512);
and U4533 (N_4533,N_702,N_2744);
and U4534 (N_4534,N_1164,N_1308);
nor U4535 (N_4535,N_1356,N_2342);
xor U4536 (N_4536,N_561,N_782);
or U4537 (N_4537,N_421,N_982);
and U4538 (N_4538,N_2200,N_479);
or U4539 (N_4539,N_2765,N_512);
or U4540 (N_4540,N_300,N_466);
nor U4541 (N_4541,N_2080,N_1288);
and U4542 (N_4542,N_2934,N_1480);
and U4543 (N_4543,N_2788,N_2366);
nor U4544 (N_4544,N_250,N_931);
or U4545 (N_4545,N_2423,N_2861);
or U4546 (N_4546,N_313,N_1003);
or U4547 (N_4547,N_1793,N_1759);
nor U4548 (N_4548,N_1949,N_938);
nor U4549 (N_4549,N_301,N_2100);
and U4550 (N_4550,N_1457,N_730);
or U4551 (N_4551,N_2505,N_2673);
or U4552 (N_4552,N_2191,N_2944);
and U4553 (N_4553,N_429,N_481);
nand U4554 (N_4554,N_1275,N_910);
and U4555 (N_4555,N_676,N_312);
nand U4556 (N_4556,N_1790,N_1369);
nand U4557 (N_4557,N_79,N_631);
and U4558 (N_4558,N_1735,N_986);
or U4559 (N_4559,N_114,N_458);
nor U4560 (N_4560,N_2170,N_115);
nor U4561 (N_4561,N_1636,N_2317);
or U4562 (N_4562,N_2899,N_1950);
and U4563 (N_4563,N_422,N_2275);
nor U4564 (N_4564,N_1051,N_969);
nand U4565 (N_4565,N_108,N_390);
and U4566 (N_4566,N_548,N_2971);
or U4567 (N_4567,N_707,N_2499);
or U4568 (N_4568,N_2154,N_2837);
or U4569 (N_4569,N_1231,N_2129);
or U4570 (N_4570,N_1083,N_129);
nand U4571 (N_4571,N_301,N_1199);
nand U4572 (N_4572,N_216,N_915);
or U4573 (N_4573,N_1582,N_1345);
and U4574 (N_4574,N_104,N_2501);
nand U4575 (N_4575,N_378,N_804);
nand U4576 (N_4576,N_2955,N_2499);
or U4577 (N_4577,N_1716,N_2444);
or U4578 (N_4578,N_1391,N_2605);
nor U4579 (N_4579,N_2893,N_1803);
xnor U4580 (N_4580,N_2623,N_2303);
or U4581 (N_4581,N_1845,N_2756);
nand U4582 (N_4582,N_1655,N_1809);
nand U4583 (N_4583,N_1855,N_175);
nor U4584 (N_4584,N_2760,N_956);
nand U4585 (N_4585,N_542,N_2721);
nor U4586 (N_4586,N_2727,N_1852);
nor U4587 (N_4587,N_599,N_2667);
and U4588 (N_4588,N_1432,N_1447);
nor U4589 (N_4589,N_1799,N_2575);
or U4590 (N_4590,N_1530,N_1381);
nand U4591 (N_4591,N_1166,N_949);
xor U4592 (N_4592,N_895,N_1199);
nand U4593 (N_4593,N_606,N_1128);
nor U4594 (N_4594,N_417,N_2044);
and U4595 (N_4595,N_2866,N_2280);
nand U4596 (N_4596,N_821,N_73);
nand U4597 (N_4597,N_2010,N_1986);
and U4598 (N_4598,N_2801,N_1520);
or U4599 (N_4599,N_845,N_1702);
nor U4600 (N_4600,N_732,N_2930);
nor U4601 (N_4601,N_2842,N_1350);
nand U4602 (N_4602,N_2227,N_602);
and U4603 (N_4603,N_54,N_657);
nor U4604 (N_4604,N_2755,N_540);
and U4605 (N_4605,N_510,N_201);
nor U4606 (N_4606,N_1984,N_2179);
or U4607 (N_4607,N_2188,N_2035);
nand U4608 (N_4608,N_1312,N_1630);
and U4609 (N_4609,N_2406,N_2710);
and U4610 (N_4610,N_1332,N_2268);
nand U4611 (N_4611,N_1684,N_802);
or U4612 (N_4612,N_1258,N_246);
nand U4613 (N_4613,N_2172,N_885);
or U4614 (N_4614,N_1541,N_1372);
nor U4615 (N_4615,N_1130,N_879);
nand U4616 (N_4616,N_2427,N_1552);
or U4617 (N_4617,N_2068,N_1408);
nor U4618 (N_4618,N_835,N_2853);
and U4619 (N_4619,N_1836,N_2707);
nand U4620 (N_4620,N_1740,N_2842);
or U4621 (N_4621,N_1204,N_2680);
nor U4622 (N_4622,N_2419,N_1506);
nor U4623 (N_4623,N_881,N_1480);
nor U4624 (N_4624,N_969,N_2720);
nand U4625 (N_4625,N_2914,N_1822);
nor U4626 (N_4626,N_479,N_636);
xor U4627 (N_4627,N_2254,N_303);
nor U4628 (N_4628,N_2652,N_1785);
nand U4629 (N_4629,N_1114,N_1944);
nand U4630 (N_4630,N_2539,N_1571);
nor U4631 (N_4631,N_902,N_1913);
or U4632 (N_4632,N_2689,N_64);
nor U4633 (N_4633,N_247,N_1637);
and U4634 (N_4634,N_461,N_246);
nand U4635 (N_4635,N_117,N_442);
nor U4636 (N_4636,N_613,N_1032);
nand U4637 (N_4637,N_2665,N_793);
nand U4638 (N_4638,N_2390,N_1427);
xnor U4639 (N_4639,N_930,N_91);
nand U4640 (N_4640,N_2167,N_2162);
nor U4641 (N_4641,N_359,N_829);
nand U4642 (N_4642,N_382,N_2635);
and U4643 (N_4643,N_420,N_2095);
and U4644 (N_4644,N_59,N_831);
or U4645 (N_4645,N_1112,N_2661);
nor U4646 (N_4646,N_1114,N_390);
nand U4647 (N_4647,N_1450,N_2377);
or U4648 (N_4648,N_2241,N_1105);
nor U4649 (N_4649,N_496,N_1156);
nand U4650 (N_4650,N_99,N_496);
or U4651 (N_4651,N_1733,N_1426);
or U4652 (N_4652,N_2373,N_2227);
or U4653 (N_4653,N_1742,N_705);
and U4654 (N_4654,N_1711,N_2947);
nor U4655 (N_4655,N_2646,N_631);
and U4656 (N_4656,N_1455,N_1318);
nor U4657 (N_4657,N_2147,N_1765);
nand U4658 (N_4658,N_2942,N_2232);
and U4659 (N_4659,N_2652,N_282);
or U4660 (N_4660,N_2498,N_811);
and U4661 (N_4661,N_2182,N_2129);
nand U4662 (N_4662,N_1080,N_156);
nand U4663 (N_4663,N_503,N_1854);
or U4664 (N_4664,N_672,N_1855);
or U4665 (N_4665,N_889,N_2243);
nand U4666 (N_4666,N_1922,N_1731);
and U4667 (N_4667,N_2107,N_497);
or U4668 (N_4668,N_752,N_1955);
nand U4669 (N_4669,N_1091,N_2225);
or U4670 (N_4670,N_1791,N_2862);
xnor U4671 (N_4671,N_770,N_1898);
and U4672 (N_4672,N_2504,N_2867);
and U4673 (N_4673,N_2492,N_2571);
or U4674 (N_4674,N_410,N_847);
nor U4675 (N_4675,N_1543,N_367);
or U4676 (N_4676,N_2427,N_736);
nand U4677 (N_4677,N_1389,N_345);
xnor U4678 (N_4678,N_1624,N_644);
nor U4679 (N_4679,N_24,N_1294);
nand U4680 (N_4680,N_2892,N_317);
or U4681 (N_4681,N_569,N_1804);
or U4682 (N_4682,N_1260,N_2260);
nand U4683 (N_4683,N_177,N_1226);
nor U4684 (N_4684,N_835,N_2336);
and U4685 (N_4685,N_567,N_169);
nor U4686 (N_4686,N_607,N_1804);
nor U4687 (N_4687,N_2985,N_614);
or U4688 (N_4688,N_1032,N_586);
and U4689 (N_4689,N_1538,N_1651);
or U4690 (N_4690,N_2668,N_2368);
nand U4691 (N_4691,N_486,N_1331);
nand U4692 (N_4692,N_1592,N_1347);
nor U4693 (N_4693,N_1478,N_2499);
nor U4694 (N_4694,N_858,N_1826);
and U4695 (N_4695,N_1303,N_1655);
or U4696 (N_4696,N_441,N_681);
nor U4697 (N_4697,N_126,N_1478);
and U4698 (N_4698,N_315,N_1596);
and U4699 (N_4699,N_2679,N_2154);
or U4700 (N_4700,N_2583,N_1165);
or U4701 (N_4701,N_1004,N_2069);
and U4702 (N_4702,N_2712,N_1920);
or U4703 (N_4703,N_1344,N_2064);
nor U4704 (N_4704,N_2794,N_2946);
and U4705 (N_4705,N_317,N_184);
or U4706 (N_4706,N_2038,N_2897);
or U4707 (N_4707,N_1512,N_1599);
nand U4708 (N_4708,N_879,N_2879);
and U4709 (N_4709,N_1163,N_1435);
and U4710 (N_4710,N_1611,N_2098);
and U4711 (N_4711,N_1047,N_1486);
nor U4712 (N_4712,N_1811,N_2757);
nor U4713 (N_4713,N_564,N_457);
nor U4714 (N_4714,N_1702,N_1682);
or U4715 (N_4715,N_44,N_1479);
or U4716 (N_4716,N_2640,N_783);
and U4717 (N_4717,N_1563,N_2466);
or U4718 (N_4718,N_1582,N_1977);
nor U4719 (N_4719,N_1469,N_734);
or U4720 (N_4720,N_842,N_1402);
or U4721 (N_4721,N_1639,N_1045);
nor U4722 (N_4722,N_255,N_794);
nor U4723 (N_4723,N_2098,N_1796);
xor U4724 (N_4724,N_1207,N_501);
and U4725 (N_4725,N_8,N_1655);
and U4726 (N_4726,N_2262,N_477);
nand U4727 (N_4727,N_1672,N_2059);
and U4728 (N_4728,N_162,N_837);
nor U4729 (N_4729,N_80,N_281);
nor U4730 (N_4730,N_1640,N_287);
nand U4731 (N_4731,N_2801,N_1617);
and U4732 (N_4732,N_1667,N_2601);
nand U4733 (N_4733,N_2217,N_585);
nor U4734 (N_4734,N_1196,N_2352);
or U4735 (N_4735,N_2457,N_2060);
and U4736 (N_4736,N_1293,N_125);
or U4737 (N_4737,N_2665,N_1511);
or U4738 (N_4738,N_761,N_68);
or U4739 (N_4739,N_2022,N_2995);
nor U4740 (N_4740,N_611,N_1257);
or U4741 (N_4741,N_1992,N_1012);
nand U4742 (N_4742,N_2824,N_918);
nor U4743 (N_4743,N_25,N_1793);
nor U4744 (N_4744,N_1211,N_1166);
or U4745 (N_4745,N_264,N_2707);
or U4746 (N_4746,N_201,N_2453);
or U4747 (N_4747,N_2592,N_555);
nor U4748 (N_4748,N_2657,N_2389);
nor U4749 (N_4749,N_1374,N_952);
nor U4750 (N_4750,N_838,N_38);
or U4751 (N_4751,N_1048,N_523);
nand U4752 (N_4752,N_778,N_312);
or U4753 (N_4753,N_140,N_715);
nor U4754 (N_4754,N_2024,N_1182);
nor U4755 (N_4755,N_1051,N_501);
nand U4756 (N_4756,N_29,N_452);
nor U4757 (N_4757,N_2486,N_769);
or U4758 (N_4758,N_972,N_546);
nor U4759 (N_4759,N_2074,N_2147);
nand U4760 (N_4760,N_2833,N_2403);
and U4761 (N_4761,N_235,N_1804);
xor U4762 (N_4762,N_836,N_1898);
nor U4763 (N_4763,N_637,N_385);
nor U4764 (N_4764,N_1203,N_2865);
and U4765 (N_4765,N_2972,N_1158);
nor U4766 (N_4766,N_149,N_2725);
nor U4767 (N_4767,N_1006,N_1784);
nand U4768 (N_4768,N_281,N_184);
and U4769 (N_4769,N_648,N_1881);
nor U4770 (N_4770,N_1922,N_2650);
nor U4771 (N_4771,N_2537,N_2458);
nand U4772 (N_4772,N_1141,N_824);
and U4773 (N_4773,N_2797,N_2410);
nor U4774 (N_4774,N_2468,N_2724);
nand U4775 (N_4775,N_1874,N_2636);
nand U4776 (N_4776,N_1305,N_562);
or U4777 (N_4777,N_1122,N_1183);
nor U4778 (N_4778,N_98,N_2086);
or U4779 (N_4779,N_501,N_680);
nand U4780 (N_4780,N_2278,N_492);
nor U4781 (N_4781,N_2099,N_496);
nand U4782 (N_4782,N_1757,N_2240);
nor U4783 (N_4783,N_640,N_658);
nor U4784 (N_4784,N_1340,N_355);
nand U4785 (N_4785,N_2347,N_1085);
nand U4786 (N_4786,N_347,N_1429);
or U4787 (N_4787,N_1048,N_1210);
or U4788 (N_4788,N_2844,N_174);
nand U4789 (N_4789,N_1972,N_2751);
or U4790 (N_4790,N_353,N_1764);
nor U4791 (N_4791,N_1709,N_295);
xor U4792 (N_4792,N_1505,N_2089);
nand U4793 (N_4793,N_2194,N_918);
and U4794 (N_4794,N_1447,N_415);
and U4795 (N_4795,N_2133,N_198);
nand U4796 (N_4796,N_2940,N_936);
nor U4797 (N_4797,N_1205,N_805);
nand U4798 (N_4798,N_1692,N_2156);
nand U4799 (N_4799,N_1508,N_1288);
or U4800 (N_4800,N_1514,N_1813);
nor U4801 (N_4801,N_202,N_2283);
nand U4802 (N_4802,N_2329,N_1771);
or U4803 (N_4803,N_1116,N_2477);
nand U4804 (N_4804,N_1883,N_2250);
nor U4805 (N_4805,N_2157,N_2299);
nand U4806 (N_4806,N_1350,N_83);
nor U4807 (N_4807,N_1690,N_2375);
nor U4808 (N_4808,N_1568,N_2675);
nor U4809 (N_4809,N_2721,N_1956);
or U4810 (N_4810,N_1440,N_1409);
nand U4811 (N_4811,N_1077,N_2341);
nand U4812 (N_4812,N_2501,N_2395);
or U4813 (N_4813,N_399,N_1363);
nand U4814 (N_4814,N_287,N_2090);
nand U4815 (N_4815,N_271,N_1395);
or U4816 (N_4816,N_846,N_1943);
or U4817 (N_4817,N_604,N_1506);
or U4818 (N_4818,N_1532,N_2207);
and U4819 (N_4819,N_400,N_1036);
nand U4820 (N_4820,N_2904,N_1136);
xor U4821 (N_4821,N_353,N_1208);
nand U4822 (N_4822,N_2774,N_1651);
nand U4823 (N_4823,N_15,N_743);
nor U4824 (N_4824,N_705,N_1297);
or U4825 (N_4825,N_2228,N_1239);
or U4826 (N_4826,N_1453,N_865);
nor U4827 (N_4827,N_578,N_533);
nor U4828 (N_4828,N_2141,N_1791);
nand U4829 (N_4829,N_2994,N_1283);
or U4830 (N_4830,N_134,N_372);
nand U4831 (N_4831,N_1453,N_2459);
or U4832 (N_4832,N_1247,N_1890);
nand U4833 (N_4833,N_2048,N_422);
nor U4834 (N_4834,N_2884,N_449);
nor U4835 (N_4835,N_1755,N_809);
nand U4836 (N_4836,N_262,N_2090);
nand U4837 (N_4837,N_2091,N_2521);
nand U4838 (N_4838,N_1733,N_1219);
and U4839 (N_4839,N_2545,N_906);
nor U4840 (N_4840,N_1638,N_551);
nand U4841 (N_4841,N_857,N_2937);
nand U4842 (N_4842,N_439,N_2391);
or U4843 (N_4843,N_656,N_369);
nand U4844 (N_4844,N_1967,N_2544);
and U4845 (N_4845,N_228,N_88);
nor U4846 (N_4846,N_37,N_408);
nand U4847 (N_4847,N_49,N_963);
or U4848 (N_4848,N_2339,N_88);
or U4849 (N_4849,N_810,N_629);
xor U4850 (N_4850,N_1555,N_2678);
nand U4851 (N_4851,N_1226,N_1528);
or U4852 (N_4852,N_92,N_668);
nand U4853 (N_4853,N_2853,N_2630);
or U4854 (N_4854,N_1561,N_246);
or U4855 (N_4855,N_462,N_1216);
xor U4856 (N_4856,N_662,N_2612);
nor U4857 (N_4857,N_2253,N_313);
and U4858 (N_4858,N_701,N_480);
nand U4859 (N_4859,N_1642,N_938);
and U4860 (N_4860,N_565,N_2778);
nand U4861 (N_4861,N_1164,N_2649);
and U4862 (N_4862,N_575,N_1406);
xor U4863 (N_4863,N_1820,N_395);
nor U4864 (N_4864,N_427,N_1902);
xnor U4865 (N_4865,N_554,N_2319);
nand U4866 (N_4866,N_1642,N_2244);
and U4867 (N_4867,N_1418,N_170);
nand U4868 (N_4868,N_910,N_904);
nor U4869 (N_4869,N_1985,N_860);
nand U4870 (N_4870,N_144,N_2977);
nor U4871 (N_4871,N_1508,N_1524);
or U4872 (N_4872,N_2405,N_630);
nand U4873 (N_4873,N_608,N_1480);
nor U4874 (N_4874,N_956,N_1097);
nor U4875 (N_4875,N_1419,N_2692);
nand U4876 (N_4876,N_1327,N_2335);
and U4877 (N_4877,N_1762,N_69);
and U4878 (N_4878,N_321,N_1975);
nand U4879 (N_4879,N_2189,N_387);
nand U4880 (N_4880,N_523,N_872);
nand U4881 (N_4881,N_2515,N_363);
nor U4882 (N_4882,N_149,N_896);
or U4883 (N_4883,N_2354,N_145);
or U4884 (N_4884,N_2064,N_798);
and U4885 (N_4885,N_1209,N_401);
and U4886 (N_4886,N_527,N_2557);
and U4887 (N_4887,N_228,N_2790);
nand U4888 (N_4888,N_2215,N_2320);
nand U4889 (N_4889,N_2668,N_49);
xor U4890 (N_4890,N_2507,N_1711);
or U4891 (N_4891,N_144,N_1118);
or U4892 (N_4892,N_2594,N_805);
nor U4893 (N_4893,N_1043,N_1362);
and U4894 (N_4894,N_238,N_1608);
nand U4895 (N_4895,N_1830,N_1867);
or U4896 (N_4896,N_1467,N_2823);
or U4897 (N_4897,N_733,N_932);
or U4898 (N_4898,N_54,N_699);
and U4899 (N_4899,N_837,N_1090);
nor U4900 (N_4900,N_1128,N_909);
nor U4901 (N_4901,N_911,N_2431);
and U4902 (N_4902,N_749,N_462);
nor U4903 (N_4903,N_2455,N_1967);
and U4904 (N_4904,N_2986,N_1007);
nor U4905 (N_4905,N_2873,N_1718);
nor U4906 (N_4906,N_1076,N_688);
nand U4907 (N_4907,N_2698,N_2870);
and U4908 (N_4908,N_1946,N_694);
nand U4909 (N_4909,N_2775,N_311);
nor U4910 (N_4910,N_1650,N_2711);
or U4911 (N_4911,N_1367,N_52);
and U4912 (N_4912,N_2585,N_1790);
and U4913 (N_4913,N_216,N_307);
or U4914 (N_4914,N_2598,N_1613);
and U4915 (N_4915,N_2752,N_2882);
nand U4916 (N_4916,N_2043,N_1103);
or U4917 (N_4917,N_2684,N_591);
and U4918 (N_4918,N_2001,N_1199);
nor U4919 (N_4919,N_2178,N_842);
nor U4920 (N_4920,N_427,N_1612);
nand U4921 (N_4921,N_1078,N_1549);
or U4922 (N_4922,N_1933,N_2201);
nand U4923 (N_4923,N_2915,N_2336);
nand U4924 (N_4924,N_1933,N_613);
nand U4925 (N_4925,N_2551,N_942);
and U4926 (N_4926,N_2565,N_31);
and U4927 (N_4927,N_2284,N_2849);
nand U4928 (N_4928,N_2129,N_2826);
or U4929 (N_4929,N_1819,N_2236);
nand U4930 (N_4930,N_1842,N_2324);
nor U4931 (N_4931,N_1228,N_853);
and U4932 (N_4932,N_1482,N_2733);
or U4933 (N_4933,N_690,N_247);
nor U4934 (N_4934,N_215,N_317);
or U4935 (N_4935,N_1052,N_206);
and U4936 (N_4936,N_996,N_1401);
or U4937 (N_4937,N_801,N_67);
and U4938 (N_4938,N_1234,N_1869);
or U4939 (N_4939,N_817,N_1265);
nor U4940 (N_4940,N_2500,N_1389);
nand U4941 (N_4941,N_2153,N_2419);
nand U4942 (N_4942,N_1146,N_65);
and U4943 (N_4943,N_1394,N_938);
nor U4944 (N_4944,N_1051,N_451);
nor U4945 (N_4945,N_1753,N_1320);
nand U4946 (N_4946,N_1216,N_2219);
nor U4947 (N_4947,N_885,N_919);
nand U4948 (N_4948,N_2632,N_2051);
nand U4949 (N_4949,N_2386,N_528);
or U4950 (N_4950,N_2912,N_2871);
and U4951 (N_4951,N_2660,N_2841);
and U4952 (N_4952,N_126,N_2443);
nor U4953 (N_4953,N_2135,N_2545);
or U4954 (N_4954,N_2378,N_152);
and U4955 (N_4955,N_2842,N_2008);
nor U4956 (N_4956,N_2618,N_2725);
and U4957 (N_4957,N_1274,N_2459);
or U4958 (N_4958,N_2819,N_936);
xnor U4959 (N_4959,N_358,N_2886);
or U4960 (N_4960,N_2857,N_820);
or U4961 (N_4961,N_997,N_2031);
nor U4962 (N_4962,N_2101,N_208);
or U4963 (N_4963,N_872,N_440);
and U4964 (N_4964,N_429,N_962);
or U4965 (N_4965,N_1432,N_1135);
nand U4966 (N_4966,N_1284,N_218);
and U4967 (N_4967,N_1878,N_716);
and U4968 (N_4968,N_754,N_2138);
or U4969 (N_4969,N_2378,N_270);
and U4970 (N_4970,N_2867,N_2330);
and U4971 (N_4971,N_541,N_1649);
nor U4972 (N_4972,N_2854,N_2667);
nand U4973 (N_4973,N_605,N_2260);
nand U4974 (N_4974,N_2400,N_1922);
or U4975 (N_4975,N_2490,N_336);
and U4976 (N_4976,N_2295,N_682);
or U4977 (N_4977,N_108,N_2812);
or U4978 (N_4978,N_741,N_722);
and U4979 (N_4979,N_2950,N_1175);
nand U4980 (N_4980,N_293,N_2382);
and U4981 (N_4981,N_2078,N_2157);
xnor U4982 (N_4982,N_1505,N_2294);
and U4983 (N_4983,N_2857,N_564);
or U4984 (N_4984,N_1622,N_2665);
and U4985 (N_4985,N_2666,N_1495);
or U4986 (N_4986,N_1792,N_2566);
nor U4987 (N_4987,N_2224,N_1632);
and U4988 (N_4988,N_1850,N_2626);
or U4989 (N_4989,N_145,N_2450);
nor U4990 (N_4990,N_673,N_571);
and U4991 (N_4991,N_279,N_1425);
and U4992 (N_4992,N_2647,N_1409);
and U4993 (N_4993,N_769,N_2344);
nor U4994 (N_4994,N_2658,N_1425);
nor U4995 (N_4995,N_209,N_1896);
nor U4996 (N_4996,N_1742,N_1516);
and U4997 (N_4997,N_139,N_102);
or U4998 (N_4998,N_910,N_2645);
nand U4999 (N_4999,N_2757,N_1484);
or U5000 (N_5000,N_545,N_1363);
nand U5001 (N_5001,N_1184,N_2692);
or U5002 (N_5002,N_1396,N_335);
nand U5003 (N_5003,N_2158,N_1795);
nand U5004 (N_5004,N_1805,N_2994);
nor U5005 (N_5005,N_565,N_2132);
nand U5006 (N_5006,N_2809,N_1653);
and U5007 (N_5007,N_2994,N_11);
nand U5008 (N_5008,N_2966,N_1473);
nand U5009 (N_5009,N_884,N_614);
and U5010 (N_5010,N_1083,N_2196);
nor U5011 (N_5011,N_1496,N_2404);
nor U5012 (N_5012,N_1920,N_543);
xor U5013 (N_5013,N_248,N_1565);
nand U5014 (N_5014,N_1406,N_685);
and U5015 (N_5015,N_1864,N_197);
nor U5016 (N_5016,N_1291,N_2431);
and U5017 (N_5017,N_1935,N_2197);
nand U5018 (N_5018,N_1057,N_655);
and U5019 (N_5019,N_2350,N_1745);
or U5020 (N_5020,N_2793,N_250);
or U5021 (N_5021,N_2704,N_2466);
and U5022 (N_5022,N_2492,N_1240);
nor U5023 (N_5023,N_645,N_1762);
and U5024 (N_5024,N_1541,N_1018);
or U5025 (N_5025,N_1359,N_1134);
and U5026 (N_5026,N_970,N_1137);
nand U5027 (N_5027,N_2548,N_1469);
nand U5028 (N_5028,N_1881,N_941);
and U5029 (N_5029,N_2550,N_754);
nor U5030 (N_5030,N_2891,N_2015);
or U5031 (N_5031,N_2383,N_2396);
xor U5032 (N_5032,N_2237,N_2691);
nand U5033 (N_5033,N_822,N_1091);
xor U5034 (N_5034,N_875,N_1774);
nor U5035 (N_5035,N_2608,N_1763);
nand U5036 (N_5036,N_351,N_2718);
nor U5037 (N_5037,N_2428,N_195);
or U5038 (N_5038,N_822,N_1566);
and U5039 (N_5039,N_1057,N_1525);
nor U5040 (N_5040,N_2955,N_2742);
nand U5041 (N_5041,N_1511,N_2962);
nand U5042 (N_5042,N_2004,N_2034);
and U5043 (N_5043,N_2692,N_1235);
nor U5044 (N_5044,N_2532,N_2706);
or U5045 (N_5045,N_1847,N_1265);
nor U5046 (N_5046,N_171,N_2181);
nand U5047 (N_5047,N_2626,N_2871);
or U5048 (N_5048,N_2171,N_808);
or U5049 (N_5049,N_540,N_69);
nor U5050 (N_5050,N_1728,N_2959);
or U5051 (N_5051,N_1405,N_1050);
nand U5052 (N_5052,N_2154,N_842);
xor U5053 (N_5053,N_2256,N_1605);
and U5054 (N_5054,N_2402,N_2093);
or U5055 (N_5055,N_1795,N_1448);
or U5056 (N_5056,N_1618,N_2506);
nand U5057 (N_5057,N_1915,N_935);
nor U5058 (N_5058,N_2274,N_2617);
nor U5059 (N_5059,N_1943,N_1117);
nor U5060 (N_5060,N_1463,N_1809);
nor U5061 (N_5061,N_2667,N_1114);
xnor U5062 (N_5062,N_471,N_1701);
or U5063 (N_5063,N_2685,N_356);
nand U5064 (N_5064,N_2968,N_1330);
or U5065 (N_5065,N_621,N_2863);
nand U5066 (N_5066,N_2127,N_1387);
and U5067 (N_5067,N_689,N_1213);
nand U5068 (N_5068,N_988,N_2549);
nand U5069 (N_5069,N_2209,N_1790);
or U5070 (N_5070,N_437,N_1139);
or U5071 (N_5071,N_683,N_640);
xnor U5072 (N_5072,N_2498,N_152);
and U5073 (N_5073,N_1960,N_2248);
or U5074 (N_5074,N_712,N_1875);
nor U5075 (N_5075,N_1508,N_1122);
nor U5076 (N_5076,N_1853,N_2911);
nor U5077 (N_5077,N_2493,N_2470);
and U5078 (N_5078,N_261,N_1150);
or U5079 (N_5079,N_1816,N_1083);
nor U5080 (N_5080,N_1753,N_1597);
and U5081 (N_5081,N_2386,N_325);
xor U5082 (N_5082,N_2409,N_222);
and U5083 (N_5083,N_1875,N_1858);
or U5084 (N_5084,N_1652,N_70);
and U5085 (N_5085,N_1169,N_335);
or U5086 (N_5086,N_777,N_1287);
nor U5087 (N_5087,N_282,N_2186);
and U5088 (N_5088,N_178,N_691);
xor U5089 (N_5089,N_1095,N_1379);
or U5090 (N_5090,N_1565,N_723);
nand U5091 (N_5091,N_1751,N_2175);
and U5092 (N_5092,N_1005,N_1864);
or U5093 (N_5093,N_553,N_2577);
or U5094 (N_5094,N_277,N_1960);
or U5095 (N_5095,N_296,N_1601);
and U5096 (N_5096,N_2345,N_373);
nand U5097 (N_5097,N_2333,N_1657);
nor U5098 (N_5098,N_336,N_1476);
and U5099 (N_5099,N_1052,N_601);
nand U5100 (N_5100,N_1052,N_2450);
nand U5101 (N_5101,N_1416,N_2990);
nand U5102 (N_5102,N_104,N_1876);
nand U5103 (N_5103,N_659,N_929);
and U5104 (N_5104,N_889,N_1837);
nor U5105 (N_5105,N_2578,N_1097);
nand U5106 (N_5106,N_1733,N_808);
nor U5107 (N_5107,N_1548,N_1970);
and U5108 (N_5108,N_1289,N_1942);
or U5109 (N_5109,N_713,N_1332);
and U5110 (N_5110,N_2325,N_5);
nand U5111 (N_5111,N_1264,N_1282);
nor U5112 (N_5112,N_899,N_2647);
and U5113 (N_5113,N_61,N_2608);
nor U5114 (N_5114,N_2040,N_2128);
or U5115 (N_5115,N_2595,N_1480);
nand U5116 (N_5116,N_2521,N_2446);
and U5117 (N_5117,N_2137,N_1042);
nand U5118 (N_5118,N_2461,N_1463);
or U5119 (N_5119,N_908,N_2389);
nand U5120 (N_5120,N_1995,N_2738);
nor U5121 (N_5121,N_1001,N_2342);
nor U5122 (N_5122,N_1894,N_2200);
nand U5123 (N_5123,N_1835,N_867);
or U5124 (N_5124,N_2686,N_349);
nand U5125 (N_5125,N_2169,N_2628);
nor U5126 (N_5126,N_1584,N_728);
nand U5127 (N_5127,N_150,N_69);
and U5128 (N_5128,N_2782,N_1322);
or U5129 (N_5129,N_2636,N_2516);
nand U5130 (N_5130,N_1040,N_2634);
or U5131 (N_5131,N_1436,N_1841);
nand U5132 (N_5132,N_602,N_2533);
and U5133 (N_5133,N_664,N_666);
and U5134 (N_5134,N_534,N_1259);
nor U5135 (N_5135,N_819,N_520);
and U5136 (N_5136,N_423,N_1179);
nand U5137 (N_5137,N_632,N_2798);
and U5138 (N_5138,N_2846,N_2321);
nor U5139 (N_5139,N_1202,N_999);
or U5140 (N_5140,N_1284,N_135);
and U5141 (N_5141,N_2371,N_2584);
xor U5142 (N_5142,N_2161,N_2431);
nand U5143 (N_5143,N_2524,N_2041);
or U5144 (N_5144,N_909,N_1847);
nor U5145 (N_5145,N_2880,N_176);
nand U5146 (N_5146,N_2155,N_618);
nor U5147 (N_5147,N_1550,N_2458);
or U5148 (N_5148,N_353,N_683);
nor U5149 (N_5149,N_2363,N_628);
nor U5150 (N_5150,N_174,N_1399);
nand U5151 (N_5151,N_945,N_383);
nand U5152 (N_5152,N_936,N_1869);
nand U5153 (N_5153,N_2351,N_75);
or U5154 (N_5154,N_9,N_2462);
and U5155 (N_5155,N_2572,N_748);
or U5156 (N_5156,N_899,N_389);
or U5157 (N_5157,N_1895,N_8);
and U5158 (N_5158,N_1614,N_1624);
nand U5159 (N_5159,N_1522,N_693);
nand U5160 (N_5160,N_280,N_2025);
or U5161 (N_5161,N_2341,N_563);
or U5162 (N_5162,N_2844,N_918);
and U5163 (N_5163,N_2202,N_2751);
nor U5164 (N_5164,N_1838,N_1632);
or U5165 (N_5165,N_1692,N_1129);
and U5166 (N_5166,N_2297,N_2623);
or U5167 (N_5167,N_719,N_1772);
nand U5168 (N_5168,N_2865,N_2746);
nand U5169 (N_5169,N_2704,N_648);
or U5170 (N_5170,N_673,N_2364);
nand U5171 (N_5171,N_2556,N_702);
and U5172 (N_5172,N_425,N_65);
or U5173 (N_5173,N_1598,N_907);
nand U5174 (N_5174,N_2653,N_30);
and U5175 (N_5175,N_463,N_2573);
nor U5176 (N_5176,N_2605,N_1381);
nor U5177 (N_5177,N_1120,N_2114);
or U5178 (N_5178,N_446,N_2507);
or U5179 (N_5179,N_2685,N_130);
or U5180 (N_5180,N_2513,N_2063);
and U5181 (N_5181,N_815,N_2316);
or U5182 (N_5182,N_115,N_1667);
or U5183 (N_5183,N_1226,N_2695);
and U5184 (N_5184,N_1449,N_67);
and U5185 (N_5185,N_584,N_90);
nand U5186 (N_5186,N_708,N_571);
nor U5187 (N_5187,N_2853,N_1717);
and U5188 (N_5188,N_1969,N_2899);
and U5189 (N_5189,N_1388,N_2746);
nor U5190 (N_5190,N_695,N_861);
or U5191 (N_5191,N_2262,N_1029);
nor U5192 (N_5192,N_900,N_2868);
and U5193 (N_5193,N_137,N_878);
nor U5194 (N_5194,N_1187,N_2390);
and U5195 (N_5195,N_1619,N_1383);
nor U5196 (N_5196,N_1685,N_2516);
and U5197 (N_5197,N_2887,N_2465);
nand U5198 (N_5198,N_1807,N_884);
nor U5199 (N_5199,N_2813,N_552);
and U5200 (N_5200,N_1605,N_295);
nand U5201 (N_5201,N_186,N_1887);
nor U5202 (N_5202,N_2575,N_1462);
and U5203 (N_5203,N_2677,N_1995);
or U5204 (N_5204,N_1399,N_2470);
nand U5205 (N_5205,N_641,N_255);
and U5206 (N_5206,N_478,N_2968);
or U5207 (N_5207,N_356,N_322);
or U5208 (N_5208,N_189,N_549);
or U5209 (N_5209,N_1185,N_1875);
or U5210 (N_5210,N_28,N_767);
nor U5211 (N_5211,N_615,N_1934);
and U5212 (N_5212,N_890,N_2509);
xnor U5213 (N_5213,N_1433,N_1919);
and U5214 (N_5214,N_1220,N_154);
or U5215 (N_5215,N_200,N_2556);
and U5216 (N_5216,N_1217,N_2214);
and U5217 (N_5217,N_2534,N_2422);
nor U5218 (N_5218,N_2403,N_738);
nor U5219 (N_5219,N_2446,N_2486);
or U5220 (N_5220,N_2296,N_2304);
and U5221 (N_5221,N_1978,N_1404);
nand U5222 (N_5222,N_2601,N_1487);
nand U5223 (N_5223,N_2019,N_2707);
nor U5224 (N_5224,N_4,N_1493);
nor U5225 (N_5225,N_2034,N_370);
and U5226 (N_5226,N_588,N_1756);
nand U5227 (N_5227,N_1616,N_187);
or U5228 (N_5228,N_915,N_2949);
xor U5229 (N_5229,N_1768,N_1968);
or U5230 (N_5230,N_226,N_1980);
or U5231 (N_5231,N_1581,N_294);
nand U5232 (N_5232,N_1290,N_1958);
and U5233 (N_5233,N_2077,N_499);
nand U5234 (N_5234,N_1477,N_2924);
nand U5235 (N_5235,N_2938,N_944);
and U5236 (N_5236,N_1306,N_1479);
and U5237 (N_5237,N_1823,N_1724);
nand U5238 (N_5238,N_1979,N_2405);
nor U5239 (N_5239,N_2392,N_1989);
nor U5240 (N_5240,N_1258,N_196);
or U5241 (N_5241,N_136,N_1185);
or U5242 (N_5242,N_776,N_396);
and U5243 (N_5243,N_389,N_1650);
nor U5244 (N_5244,N_2603,N_1721);
nand U5245 (N_5245,N_341,N_480);
and U5246 (N_5246,N_288,N_2363);
or U5247 (N_5247,N_2309,N_2439);
and U5248 (N_5248,N_945,N_611);
nor U5249 (N_5249,N_490,N_2393);
nand U5250 (N_5250,N_515,N_1073);
nand U5251 (N_5251,N_2990,N_613);
nor U5252 (N_5252,N_521,N_754);
nand U5253 (N_5253,N_1054,N_1204);
or U5254 (N_5254,N_1863,N_921);
or U5255 (N_5255,N_833,N_847);
nor U5256 (N_5256,N_1294,N_2280);
nor U5257 (N_5257,N_948,N_13);
nor U5258 (N_5258,N_1409,N_1228);
nor U5259 (N_5259,N_2603,N_512);
or U5260 (N_5260,N_1494,N_655);
and U5261 (N_5261,N_2487,N_2540);
or U5262 (N_5262,N_2961,N_2509);
nand U5263 (N_5263,N_1203,N_1554);
and U5264 (N_5264,N_1964,N_2182);
nor U5265 (N_5265,N_1043,N_2285);
nand U5266 (N_5266,N_2176,N_1155);
or U5267 (N_5267,N_2311,N_1316);
and U5268 (N_5268,N_94,N_2094);
nand U5269 (N_5269,N_2035,N_1623);
or U5270 (N_5270,N_51,N_742);
nor U5271 (N_5271,N_2633,N_1567);
nand U5272 (N_5272,N_433,N_2075);
or U5273 (N_5273,N_1731,N_391);
or U5274 (N_5274,N_2591,N_2584);
nor U5275 (N_5275,N_1805,N_2868);
and U5276 (N_5276,N_888,N_1830);
nor U5277 (N_5277,N_2254,N_2398);
nand U5278 (N_5278,N_2211,N_686);
and U5279 (N_5279,N_459,N_1177);
nand U5280 (N_5280,N_36,N_2260);
nor U5281 (N_5281,N_959,N_1392);
nand U5282 (N_5282,N_1649,N_794);
nor U5283 (N_5283,N_534,N_1910);
nor U5284 (N_5284,N_904,N_365);
nand U5285 (N_5285,N_1131,N_1419);
or U5286 (N_5286,N_1891,N_2430);
nand U5287 (N_5287,N_94,N_2766);
nand U5288 (N_5288,N_2759,N_529);
nor U5289 (N_5289,N_1104,N_2505);
or U5290 (N_5290,N_2387,N_496);
and U5291 (N_5291,N_1639,N_675);
nand U5292 (N_5292,N_1925,N_1378);
nand U5293 (N_5293,N_391,N_2466);
nor U5294 (N_5294,N_2128,N_558);
nor U5295 (N_5295,N_444,N_2256);
nor U5296 (N_5296,N_2425,N_1115);
or U5297 (N_5297,N_712,N_1926);
and U5298 (N_5298,N_1667,N_801);
nor U5299 (N_5299,N_2230,N_460);
nor U5300 (N_5300,N_1742,N_2196);
and U5301 (N_5301,N_1994,N_1048);
nand U5302 (N_5302,N_2765,N_440);
nand U5303 (N_5303,N_1198,N_1977);
and U5304 (N_5304,N_1012,N_170);
and U5305 (N_5305,N_2325,N_1196);
and U5306 (N_5306,N_1813,N_807);
or U5307 (N_5307,N_594,N_2523);
nor U5308 (N_5308,N_894,N_161);
or U5309 (N_5309,N_2955,N_37);
or U5310 (N_5310,N_50,N_2130);
or U5311 (N_5311,N_2998,N_520);
nand U5312 (N_5312,N_631,N_1871);
nor U5313 (N_5313,N_649,N_2566);
nor U5314 (N_5314,N_2442,N_1576);
nor U5315 (N_5315,N_1167,N_2420);
nor U5316 (N_5316,N_1681,N_469);
or U5317 (N_5317,N_1218,N_2450);
nor U5318 (N_5318,N_1753,N_1818);
nand U5319 (N_5319,N_1755,N_264);
or U5320 (N_5320,N_1749,N_2290);
or U5321 (N_5321,N_803,N_1683);
nand U5322 (N_5322,N_856,N_1998);
nand U5323 (N_5323,N_1994,N_2081);
or U5324 (N_5324,N_2716,N_2034);
or U5325 (N_5325,N_598,N_1741);
or U5326 (N_5326,N_2655,N_2432);
nand U5327 (N_5327,N_2537,N_1796);
or U5328 (N_5328,N_2313,N_628);
nand U5329 (N_5329,N_2838,N_378);
nor U5330 (N_5330,N_373,N_1803);
xor U5331 (N_5331,N_1388,N_1088);
and U5332 (N_5332,N_562,N_222);
and U5333 (N_5333,N_2293,N_26);
xnor U5334 (N_5334,N_14,N_334);
nand U5335 (N_5335,N_1206,N_25);
or U5336 (N_5336,N_1831,N_1959);
nor U5337 (N_5337,N_1817,N_1252);
and U5338 (N_5338,N_445,N_1070);
nand U5339 (N_5339,N_137,N_901);
nand U5340 (N_5340,N_2025,N_1074);
and U5341 (N_5341,N_493,N_2434);
nor U5342 (N_5342,N_1433,N_2557);
or U5343 (N_5343,N_1335,N_60);
or U5344 (N_5344,N_2180,N_1569);
nand U5345 (N_5345,N_1280,N_1658);
or U5346 (N_5346,N_2661,N_1925);
nand U5347 (N_5347,N_685,N_425);
nor U5348 (N_5348,N_408,N_445);
nand U5349 (N_5349,N_2733,N_1607);
or U5350 (N_5350,N_2511,N_2910);
and U5351 (N_5351,N_469,N_404);
or U5352 (N_5352,N_2396,N_1366);
and U5353 (N_5353,N_2999,N_1258);
nor U5354 (N_5354,N_1880,N_2734);
and U5355 (N_5355,N_2942,N_2424);
or U5356 (N_5356,N_2204,N_918);
nand U5357 (N_5357,N_1887,N_406);
and U5358 (N_5358,N_1516,N_2573);
nor U5359 (N_5359,N_2196,N_1698);
or U5360 (N_5360,N_2559,N_158);
nand U5361 (N_5361,N_1199,N_1270);
nand U5362 (N_5362,N_5,N_96);
nor U5363 (N_5363,N_1616,N_2809);
nand U5364 (N_5364,N_1657,N_515);
or U5365 (N_5365,N_2914,N_2007);
and U5366 (N_5366,N_567,N_1892);
nand U5367 (N_5367,N_2916,N_1403);
nor U5368 (N_5368,N_2601,N_201);
and U5369 (N_5369,N_2487,N_127);
nand U5370 (N_5370,N_580,N_529);
nand U5371 (N_5371,N_1715,N_1733);
nand U5372 (N_5372,N_1115,N_1696);
and U5373 (N_5373,N_1124,N_2505);
nand U5374 (N_5374,N_2936,N_2650);
nand U5375 (N_5375,N_1246,N_136);
xor U5376 (N_5376,N_2716,N_651);
nand U5377 (N_5377,N_1779,N_2703);
or U5378 (N_5378,N_195,N_1611);
or U5379 (N_5379,N_138,N_1816);
and U5380 (N_5380,N_785,N_2840);
xor U5381 (N_5381,N_2347,N_751);
and U5382 (N_5382,N_2422,N_2292);
nor U5383 (N_5383,N_1949,N_1459);
or U5384 (N_5384,N_154,N_321);
and U5385 (N_5385,N_308,N_730);
or U5386 (N_5386,N_380,N_1163);
nor U5387 (N_5387,N_1572,N_717);
nand U5388 (N_5388,N_1598,N_255);
xor U5389 (N_5389,N_964,N_1871);
nand U5390 (N_5390,N_1737,N_939);
nor U5391 (N_5391,N_2855,N_47);
nor U5392 (N_5392,N_334,N_1100);
or U5393 (N_5393,N_381,N_2644);
nor U5394 (N_5394,N_2929,N_2898);
or U5395 (N_5395,N_495,N_1454);
nand U5396 (N_5396,N_1855,N_2653);
and U5397 (N_5397,N_1812,N_1003);
nand U5398 (N_5398,N_2948,N_225);
or U5399 (N_5399,N_2193,N_2149);
nor U5400 (N_5400,N_525,N_1890);
or U5401 (N_5401,N_1304,N_739);
and U5402 (N_5402,N_221,N_2573);
nor U5403 (N_5403,N_2830,N_135);
and U5404 (N_5404,N_2944,N_2973);
or U5405 (N_5405,N_2162,N_2892);
and U5406 (N_5406,N_1168,N_655);
and U5407 (N_5407,N_294,N_1454);
and U5408 (N_5408,N_966,N_897);
and U5409 (N_5409,N_2389,N_673);
xor U5410 (N_5410,N_1158,N_2302);
or U5411 (N_5411,N_2724,N_1008);
and U5412 (N_5412,N_455,N_2868);
or U5413 (N_5413,N_34,N_1005);
nand U5414 (N_5414,N_1085,N_621);
nand U5415 (N_5415,N_1722,N_633);
nand U5416 (N_5416,N_586,N_238);
and U5417 (N_5417,N_2928,N_351);
and U5418 (N_5418,N_2684,N_2885);
nor U5419 (N_5419,N_741,N_1459);
or U5420 (N_5420,N_1218,N_422);
nand U5421 (N_5421,N_1855,N_1833);
nor U5422 (N_5422,N_425,N_1450);
nor U5423 (N_5423,N_1097,N_486);
or U5424 (N_5424,N_342,N_2067);
nor U5425 (N_5425,N_260,N_1033);
nand U5426 (N_5426,N_1654,N_632);
and U5427 (N_5427,N_962,N_388);
nor U5428 (N_5428,N_1006,N_2329);
xnor U5429 (N_5429,N_1812,N_320);
nor U5430 (N_5430,N_81,N_1773);
and U5431 (N_5431,N_2712,N_314);
and U5432 (N_5432,N_2856,N_1563);
nor U5433 (N_5433,N_1222,N_2555);
or U5434 (N_5434,N_1160,N_899);
nor U5435 (N_5435,N_2517,N_1547);
nor U5436 (N_5436,N_722,N_2682);
nor U5437 (N_5437,N_1774,N_2390);
or U5438 (N_5438,N_1703,N_2188);
nor U5439 (N_5439,N_2557,N_1094);
and U5440 (N_5440,N_1689,N_2796);
nand U5441 (N_5441,N_1192,N_1884);
or U5442 (N_5442,N_1692,N_1184);
and U5443 (N_5443,N_1051,N_851);
and U5444 (N_5444,N_1934,N_2329);
and U5445 (N_5445,N_1975,N_1704);
nor U5446 (N_5446,N_1033,N_1803);
and U5447 (N_5447,N_2678,N_736);
or U5448 (N_5448,N_2359,N_572);
nor U5449 (N_5449,N_545,N_1439);
and U5450 (N_5450,N_1350,N_1044);
nor U5451 (N_5451,N_28,N_1406);
and U5452 (N_5452,N_1838,N_433);
and U5453 (N_5453,N_986,N_21);
nor U5454 (N_5454,N_995,N_1814);
nand U5455 (N_5455,N_1575,N_296);
xor U5456 (N_5456,N_2455,N_2167);
or U5457 (N_5457,N_1073,N_1437);
or U5458 (N_5458,N_2209,N_1753);
nor U5459 (N_5459,N_2047,N_200);
nand U5460 (N_5460,N_1310,N_2840);
or U5461 (N_5461,N_161,N_284);
and U5462 (N_5462,N_2912,N_2376);
nor U5463 (N_5463,N_2597,N_2872);
nor U5464 (N_5464,N_1411,N_2263);
nand U5465 (N_5465,N_1578,N_493);
and U5466 (N_5466,N_189,N_797);
or U5467 (N_5467,N_778,N_2969);
or U5468 (N_5468,N_2037,N_1362);
or U5469 (N_5469,N_1056,N_1875);
and U5470 (N_5470,N_476,N_2610);
and U5471 (N_5471,N_2007,N_1136);
nand U5472 (N_5472,N_2565,N_744);
and U5473 (N_5473,N_1346,N_558);
xor U5474 (N_5474,N_1886,N_727);
and U5475 (N_5475,N_1136,N_470);
nand U5476 (N_5476,N_659,N_465);
and U5477 (N_5477,N_1793,N_1574);
nor U5478 (N_5478,N_1093,N_1235);
nor U5479 (N_5479,N_1232,N_1362);
xnor U5480 (N_5480,N_2291,N_2416);
xnor U5481 (N_5481,N_2141,N_2955);
or U5482 (N_5482,N_2658,N_2278);
nor U5483 (N_5483,N_2321,N_2260);
and U5484 (N_5484,N_1118,N_2337);
and U5485 (N_5485,N_1942,N_493);
nor U5486 (N_5486,N_2402,N_742);
or U5487 (N_5487,N_325,N_1515);
nor U5488 (N_5488,N_1216,N_2551);
nand U5489 (N_5489,N_641,N_1639);
nand U5490 (N_5490,N_430,N_1404);
or U5491 (N_5491,N_1073,N_1907);
nor U5492 (N_5492,N_1971,N_2222);
or U5493 (N_5493,N_1488,N_868);
nor U5494 (N_5494,N_1985,N_494);
or U5495 (N_5495,N_801,N_1214);
nand U5496 (N_5496,N_1656,N_2774);
xnor U5497 (N_5497,N_831,N_1215);
nor U5498 (N_5498,N_2832,N_425);
nor U5499 (N_5499,N_2185,N_2946);
and U5500 (N_5500,N_1508,N_1019);
nor U5501 (N_5501,N_1321,N_1464);
or U5502 (N_5502,N_2667,N_1754);
nor U5503 (N_5503,N_2630,N_2938);
nand U5504 (N_5504,N_1709,N_1400);
and U5505 (N_5505,N_1963,N_156);
nor U5506 (N_5506,N_2537,N_2325);
nand U5507 (N_5507,N_1498,N_2830);
nor U5508 (N_5508,N_868,N_1792);
nor U5509 (N_5509,N_2937,N_1005);
or U5510 (N_5510,N_1318,N_727);
or U5511 (N_5511,N_442,N_161);
nor U5512 (N_5512,N_2999,N_1456);
nor U5513 (N_5513,N_1525,N_96);
nand U5514 (N_5514,N_1788,N_790);
nand U5515 (N_5515,N_529,N_1914);
nand U5516 (N_5516,N_2159,N_358);
nor U5517 (N_5517,N_1089,N_864);
nand U5518 (N_5518,N_297,N_2223);
nor U5519 (N_5519,N_843,N_2200);
nand U5520 (N_5520,N_1782,N_143);
nand U5521 (N_5521,N_1093,N_644);
xor U5522 (N_5522,N_2092,N_246);
nor U5523 (N_5523,N_1745,N_2268);
nor U5524 (N_5524,N_1517,N_1609);
nand U5525 (N_5525,N_1784,N_1213);
nor U5526 (N_5526,N_1117,N_2611);
nor U5527 (N_5527,N_2267,N_2413);
or U5528 (N_5528,N_522,N_1210);
nand U5529 (N_5529,N_1328,N_2321);
xor U5530 (N_5530,N_1691,N_2244);
nor U5531 (N_5531,N_2562,N_934);
and U5532 (N_5532,N_444,N_1263);
nor U5533 (N_5533,N_2155,N_2956);
nor U5534 (N_5534,N_1267,N_1899);
nand U5535 (N_5535,N_2273,N_486);
nand U5536 (N_5536,N_1494,N_1571);
nand U5537 (N_5537,N_756,N_1345);
and U5538 (N_5538,N_1311,N_1711);
and U5539 (N_5539,N_2397,N_1862);
and U5540 (N_5540,N_2412,N_1074);
or U5541 (N_5541,N_591,N_2083);
and U5542 (N_5542,N_835,N_1549);
or U5543 (N_5543,N_2727,N_2874);
or U5544 (N_5544,N_1538,N_2093);
nor U5545 (N_5545,N_136,N_2581);
and U5546 (N_5546,N_1580,N_272);
nand U5547 (N_5547,N_1612,N_38);
nand U5548 (N_5548,N_164,N_2673);
nand U5549 (N_5549,N_584,N_877);
or U5550 (N_5550,N_1048,N_2191);
xnor U5551 (N_5551,N_2689,N_2823);
and U5552 (N_5552,N_1525,N_1337);
and U5553 (N_5553,N_2871,N_1813);
nor U5554 (N_5554,N_1670,N_203);
nand U5555 (N_5555,N_1369,N_2789);
nand U5556 (N_5556,N_2400,N_842);
nand U5557 (N_5557,N_2827,N_1800);
or U5558 (N_5558,N_154,N_2583);
nor U5559 (N_5559,N_409,N_1836);
or U5560 (N_5560,N_2551,N_1034);
nand U5561 (N_5561,N_498,N_2281);
and U5562 (N_5562,N_1101,N_2737);
or U5563 (N_5563,N_566,N_2284);
nor U5564 (N_5564,N_280,N_1497);
nor U5565 (N_5565,N_1820,N_2864);
nand U5566 (N_5566,N_2682,N_2808);
nor U5567 (N_5567,N_2569,N_1293);
nand U5568 (N_5568,N_1839,N_45);
and U5569 (N_5569,N_1562,N_1856);
and U5570 (N_5570,N_1310,N_944);
or U5571 (N_5571,N_45,N_117);
nand U5572 (N_5572,N_1227,N_2898);
nand U5573 (N_5573,N_1373,N_2522);
nor U5574 (N_5574,N_1201,N_455);
nand U5575 (N_5575,N_1880,N_2279);
or U5576 (N_5576,N_278,N_1959);
and U5577 (N_5577,N_2956,N_2918);
or U5578 (N_5578,N_862,N_663);
nor U5579 (N_5579,N_1291,N_1229);
or U5580 (N_5580,N_2743,N_1009);
and U5581 (N_5581,N_1577,N_1390);
and U5582 (N_5582,N_35,N_2301);
nand U5583 (N_5583,N_1126,N_2568);
nor U5584 (N_5584,N_1420,N_728);
or U5585 (N_5585,N_1055,N_2458);
and U5586 (N_5586,N_2027,N_2616);
nor U5587 (N_5587,N_329,N_30);
or U5588 (N_5588,N_218,N_1107);
nand U5589 (N_5589,N_1182,N_1374);
nor U5590 (N_5590,N_142,N_2252);
nand U5591 (N_5591,N_2999,N_692);
or U5592 (N_5592,N_982,N_296);
xnor U5593 (N_5593,N_1491,N_169);
or U5594 (N_5594,N_557,N_260);
or U5595 (N_5595,N_1863,N_2264);
nor U5596 (N_5596,N_923,N_180);
nor U5597 (N_5597,N_2526,N_1713);
or U5598 (N_5598,N_2532,N_2298);
and U5599 (N_5599,N_874,N_2142);
or U5600 (N_5600,N_497,N_553);
nor U5601 (N_5601,N_1369,N_778);
or U5602 (N_5602,N_386,N_478);
nand U5603 (N_5603,N_1170,N_693);
and U5604 (N_5604,N_2975,N_1993);
nor U5605 (N_5605,N_1041,N_2196);
nand U5606 (N_5606,N_2188,N_452);
or U5607 (N_5607,N_1829,N_588);
or U5608 (N_5608,N_2821,N_651);
and U5609 (N_5609,N_458,N_2593);
nor U5610 (N_5610,N_1590,N_1718);
nand U5611 (N_5611,N_429,N_2378);
nand U5612 (N_5612,N_543,N_2151);
and U5613 (N_5613,N_2080,N_2603);
or U5614 (N_5614,N_1947,N_427);
nand U5615 (N_5615,N_2918,N_1849);
or U5616 (N_5616,N_2682,N_734);
and U5617 (N_5617,N_2366,N_1289);
or U5618 (N_5618,N_2360,N_2);
nor U5619 (N_5619,N_2019,N_194);
nand U5620 (N_5620,N_2335,N_1807);
nor U5621 (N_5621,N_2493,N_1497);
nor U5622 (N_5622,N_1834,N_581);
nand U5623 (N_5623,N_2878,N_1613);
and U5624 (N_5624,N_2593,N_862);
or U5625 (N_5625,N_1335,N_1824);
nor U5626 (N_5626,N_380,N_830);
and U5627 (N_5627,N_1164,N_2030);
or U5628 (N_5628,N_2945,N_1868);
nor U5629 (N_5629,N_143,N_312);
nand U5630 (N_5630,N_1085,N_2878);
nand U5631 (N_5631,N_1134,N_448);
nand U5632 (N_5632,N_2077,N_1029);
or U5633 (N_5633,N_2165,N_1592);
or U5634 (N_5634,N_22,N_2318);
or U5635 (N_5635,N_865,N_52);
xor U5636 (N_5636,N_1555,N_2995);
and U5637 (N_5637,N_1508,N_1855);
and U5638 (N_5638,N_266,N_863);
and U5639 (N_5639,N_41,N_2195);
or U5640 (N_5640,N_2146,N_1609);
and U5641 (N_5641,N_2714,N_704);
and U5642 (N_5642,N_955,N_317);
nor U5643 (N_5643,N_2894,N_648);
nor U5644 (N_5644,N_1854,N_2015);
nor U5645 (N_5645,N_1586,N_1026);
nand U5646 (N_5646,N_802,N_390);
or U5647 (N_5647,N_1663,N_880);
and U5648 (N_5648,N_137,N_1123);
nand U5649 (N_5649,N_712,N_602);
nand U5650 (N_5650,N_2800,N_1736);
nor U5651 (N_5651,N_1712,N_760);
nor U5652 (N_5652,N_915,N_1642);
or U5653 (N_5653,N_1244,N_1874);
nor U5654 (N_5654,N_578,N_1292);
or U5655 (N_5655,N_2477,N_172);
or U5656 (N_5656,N_945,N_2579);
nor U5657 (N_5657,N_2878,N_2175);
and U5658 (N_5658,N_1610,N_2516);
or U5659 (N_5659,N_123,N_1913);
nand U5660 (N_5660,N_2228,N_1247);
and U5661 (N_5661,N_762,N_812);
nor U5662 (N_5662,N_2384,N_1995);
nand U5663 (N_5663,N_2187,N_1532);
or U5664 (N_5664,N_895,N_93);
nor U5665 (N_5665,N_2586,N_1903);
nor U5666 (N_5666,N_1800,N_2239);
xor U5667 (N_5667,N_2519,N_1443);
and U5668 (N_5668,N_1841,N_2448);
nor U5669 (N_5669,N_1235,N_110);
xor U5670 (N_5670,N_363,N_2895);
or U5671 (N_5671,N_826,N_646);
nor U5672 (N_5672,N_1388,N_1075);
or U5673 (N_5673,N_1254,N_2936);
nor U5674 (N_5674,N_1696,N_386);
or U5675 (N_5675,N_2266,N_985);
xnor U5676 (N_5676,N_1191,N_1765);
nand U5677 (N_5677,N_376,N_1647);
or U5678 (N_5678,N_1714,N_694);
or U5679 (N_5679,N_1396,N_2191);
and U5680 (N_5680,N_2825,N_2111);
nand U5681 (N_5681,N_1874,N_2054);
or U5682 (N_5682,N_556,N_1583);
and U5683 (N_5683,N_2520,N_1007);
xnor U5684 (N_5684,N_844,N_70);
or U5685 (N_5685,N_2393,N_366);
nand U5686 (N_5686,N_1615,N_2804);
and U5687 (N_5687,N_1845,N_702);
nor U5688 (N_5688,N_1488,N_2547);
nand U5689 (N_5689,N_1648,N_2040);
and U5690 (N_5690,N_2708,N_806);
xor U5691 (N_5691,N_921,N_2218);
or U5692 (N_5692,N_458,N_1206);
nand U5693 (N_5693,N_1921,N_1369);
xor U5694 (N_5694,N_2561,N_2698);
nand U5695 (N_5695,N_791,N_1000);
or U5696 (N_5696,N_926,N_2244);
and U5697 (N_5697,N_2562,N_1598);
xnor U5698 (N_5698,N_1907,N_1054);
or U5699 (N_5699,N_1245,N_1018);
nand U5700 (N_5700,N_1892,N_2782);
or U5701 (N_5701,N_1474,N_2827);
nor U5702 (N_5702,N_2202,N_1758);
and U5703 (N_5703,N_2314,N_2255);
nor U5704 (N_5704,N_1005,N_130);
nand U5705 (N_5705,N_2250,N_770);
xnor U5706 (N_5706,N_467,N_782);
nand U5707 (N_5707,N_832,N_2985);
nand U5708 (N_5708,N_1992,N_2633);
and U5709 (N_5709,N_2037,N_2665);
nor U5710 (N_5710,N_2216,N_846);
and U5711 (N_5711,N_259,N_712);
and U5712 (N_5712,N_209,N_2343);
or U5713 (N_5713,N_906,N_1675);
nor U5714 (N_5714,N_1355,N_2329);
or U5715 (N_5715,N_1112,N_958);
nor U5716 (N_5716,N_1408,N_2211);
or U5717 (N_5717,N_1264,N_1128);
nor U5718 (N_5718,N_110,N_2342);
and U5719 (N_5719,N_1133,N_177);
nand U5720 (N_5720,N_1319,N_2196);
nor U5721 (N_5721,N_1774,N_1610);
nand U5722 (N_5722,N_120,N_1018);
nand U5723 (N_5723,N_707,N_2153);
or U5724 (N_5724,N_2333,N_813);
or U5725 (N_5725,N_2643,N_1922);
and U5726 (N_5726,N_1607,N_2155);
and U5727 (N_5727,N_2715,N_172);
nand U5728 (N_5728,N_2073,N_2570);
nand U5729 (N_5729,N_1742,N_819);
and U5730 (N_5730,N_2333,N_2125);
or U5731 (N_5731,N_1240,N_1813);
nor U5732 (N_5732,N_1006,N_359);
or U5733 (N_5733,N_1596,N_1464);
or U5734 (N_5734,N_1981,N_268);
and U5735 (N_5735,N_2311,N_685);
and U5736 (N_5736,N_1759,N_2115);
nor U5737 (N_5737,N_1960,N_2174);
nand U5738 (N_5738,N_2999,N_2478);
nand U5739 (N_5739,N_941,N_1514);
or U5740 (N_5740,N_1294,N_2964);
nor U5741 (N_5741,N_2169,N_954);
nor U5742 (N_5742,N_2460,N_709);
and U5743 (N_5743,N_810,N_413);
nor U5744 (N_5744,N_551,N_2224);
or U5745 (N_5745,N_357,N_1774);
nand U5746 (N_5746,N_2788,N_146);
and U5747 (N_5747,N_1003,N_1412);
xnor U5748 (N_5748,N_886,N_801);
and U5749 (N_5749,N_2962,N_1559);
nand U5750 (N_5750,N_884,N_2321);
xor U5751 (N_5751,N_910,N_1003);
or U5752 (N_5752,N_2237,N_1899);
nand U5753 (N_5753,N_1149,N_2891);
and U5754 (N_5754,N_1508,N_1892);
nor U5755 (N_5755,N_1681,N_325);
and U5756 (N_5756,N_1621,N_1142);
nand U5757 (N_5757,N_1966,N_2113);
or U5758 (N_5758,N_2140,N_821);
nor U5759 (N_5759,N_429,N_2519);
nor U5760 (N_5760,N_2348,N_1114);
and U5761 (N_5761,N_1314,N_596);
nor U5762 (N_5762,N_1931,N_1140);
or U5763 (N_5763,N_680,N_2605);
nand U5764 (N_5764,N_1811,N_2642);
nor U5765 (N_5765,N_1703,N_575);
or U5766 (N_5766,N_2886,N_1264);
nor U5767 (N_5767,N_135,N_417);
nand U5768 (N_5768,N_2745,N_601);
and U5769 (N_5769,N_1835,N_2896);
nor U5770 (N_5770,N_899,N_403);
nor U5771 (N_5771,N_1522,N_462);
nand U5772 (N_5772,N_680,N_912);
and U5773 (N_5773,N_558,N_2617);
or U5774 (N_5774,N_1066,N_1189);
nand U5775 (N_5775,N_2804,N_2385);
and U5776 (N_5776,N_1028,N_622);
or U5777 (N_5777,N_1257,N_307);
nand U5778 (N_5778,N_1331,N_795);
and U5779 (N_5779,N_2577,N_2351);
nand U5780 (N_5780,N_1792,N_562);
nor U5781 (N_5781,N_2563,N_2192);
and U5782 (N_5782,N_2095,N_1171);
or U5783 (N_5783,N_2632,N_1269);
or U5784 (N_5784,N_1518,N_1458);
and U5785 (N_5785,N_2633,N_985);
nand U5786 (N_5786,N_390,N_2641);
or U5787 (N_5787,N_1972,N_2351);
or U5788 (N_5788,N_2772,N_1888);
and U5789 (N_5789,N_2430,N_1822);
or U5790 (N_5790,N_316,N_2236);
or U5791 (N_5791,N_1227,N_193);
nand U5792 (N_5792,N_1819,N_360);
nand U5793 (N_5793,N_1724,N_1644);
nand U5794 (N_5794,N_2003,N_689);
nor U5795 (N_5795,N_940,N_2986);
or U5796 (N_5796,N_564,N_1268);
and U5797 (N_5797,N_1782,N_2276);
xor U5798 (N_5798,N_243,N_1033);
or U5799 (N_5799,N_1575,N_68);
and U5800 (N_5800,N_2990,N_366);
or U5801 (N_5801,N_394,N_1834);
nand U5802 (N_5802,N_2152,N_979);
nand U5803 (N_5803,N_134,N_10);
nor U5804 (N_5804,N_2188,N_1363);
and U5805 (N_5805,N_517,N_1827);
nand U5806 (N_5806,N_892,N_1930);
and U5807 (N_5807,N_1201,N_622);
nor U5808 (N_5808,N_143,N_2575);
and U5809 (N_5809,N_2658,N_425);
nor U5810 (N_5810,N_1582,N_2911);
nor U5811 (N_5811,N_965,N_769);
nor U5812 (N_5812,N_36,N_1965);
nand U5813 (N_5813,N_2663,N_1644);
nor U5814 (N_5814,N_2755,N_2187);
nor U5815 (N_5815,N_93,N_2495);
or U5816 (N_5816,N_2334,N_2828);
xor U5817 (N_5817,N_2294,N_2081);
or U5818 (N_5818,N_2219,N_1907);
and U5819 (N_5819,N_1734,N_2024);
nand U5820 (N_5820,N_925,N_2374);
and U5821 (N_5821,N_1105,N_140);
nor U5822 (N_5822,N_1092,N_1173);
and U5823 (N_5823,N_600,N_2601);
nor U5824 (N_5824,N_341,N_551);
or U5825 (N_5825,N_2925,N_2888);
nor U5826 (N_5826,N_624,N_914);
and U5827 (N_5827,N_1689,N_1475);
nor U5828 (N_5828,N_40,N_362);
and U5829 (N_5829,N_1685,N_1712);
and U5830 (N_5830,N_1971,N_600);
nor U5831 (N_5831,N_2470,N_1373);
nor U5832 (N_5832,N_2343,N_1155);
and U5833 (N_5833,N_924,N_654);
nor U5834 (N_5834,N_2644,N_1550);
and U5835 (N_5835,N_2186,N_2561);
or U5836 (N_5836,N_292,N_713);
xnor U5837 (N_5837,N_1128,N_555);
and U5838 (N_5838,N_1361,N_890);
nor U5839 (N_5839,N_1477,N_1482);
nor U5840 (N_5840,N_2763,N_2120);
or U5841 (N_5841,N_1477,N_543);
and U5842 (N_5842,N_547,N_1626);
and U5843 (N_5843,N_584,N_1501);
and U5844 (N_5844,N_192,N_1320);
nand U5845 (N_5845,N_421,N_1936);
nor U5846 (N_5846,N_818,N_1949);
and U5847 (N_5847,N_1113,N_2855);
nand U5848 (N_5848,N_477,N_770);
or U5849 (N_5849,N_2490,N_2534);
nor U5850 (N_5850,N_1559,N_114);
and U5851 (N_5851,N_1365,N_308);
nor U5852 (N_5852,N_697,N_2601);
nand U5853 (N_5853,N_2995,N_2948);
and U5854 (N_5854,N_2812,N_1086);
nor U5855 (N_5855,N_66,N_2555);
or U5856 (N_5856,N_1537,N_1294);
or U5857 (N_5857,N_2762,N_2992);
nand U5858 (N_5858,N_2227,N_2732);
nand U5859 (N_5859,N_616,N_1221);
nand U5860 (N_5860,N_2077,N_1132);
nand U5861 (N_5861,N_2403,N_1187);
and U5862 (N_5862,N_318,N_1864);
nor U5863 (N_5863,N_1681,N_837);
and U5864 (N_5864,N_2082,N_641);
or U5865 (N_5865,N_2659,N_2719);
nand U5866 (N_5866,N_376,N_362);
and U5867 (N_5867,N_183,N_741);
nand U5868 (N_5868,N_2104,N_2987);
nor U5869 (N_5869,N_980,N_1232);
nor U5870 (N_5870,N_1837,N_2645);
and U5871 (N_5871,N_1437,N_1200);
and U5872 (N_5872,N_1816,N_165);
nor U5873 (N_5873,N_906,N_450);
nor U5874 (N_5874,N_675,N_1943);
nor U5875 (N_5875,N_1260,N_1340);
or U5876 (N_5876,N_805,N_465);
nor U5877 (N_5877,N_2439,N_617);
nand U5878 (N_5878,N_2960,N_100);
and U5879 (N_5879,N_579,N_2294);
nand U5880 (N_5880,N_2332,N_2831);
or U5881 (N_5881,N_1207,N_1352);
nand U5882 (N_5882,N_673,N_2426);
and U5883 (N_5883,N_2766,N_954);
nor U5884 (N_5884,N_2034,N_2679);
or U5885 (N_5885,N_1849,N_804);
nand U5886 (N_5886,N_431,N_638);
nand U5887 (N_5887,N_2408,N_2027);
nor U5888 (N_5888,N_680,N_2381);
nor U5889 (N_5889,N_2082,N_2683);
nand U5890 (N_5890,N_2510,N_2793);
or U5891 (N_5891,N_525,N_853);
and U5892 (N_5892,N_2286,N_1313);
and U5893 (N_5893,N_2688,N_1390);
nand U5894 (N_5894,N_284,N_371);
and U5895 (N_5895,N_2147,N_1526);
or U5896 (N_5896,N_2594,N_2988);
xnor U5897 (N_5897,N_2320,N_1412);
or U5898 (N_5898,N_972,N_1056);
and U5899 (N_5899,N_1023,N_511);
or U5900 (N_5900,N_2959,N_937);
and U5901 (N_5901,N_1058,N_2614);
and U5902 (N_5902,N_928,N_222);
nor U5903 (N_5903,N_1846,N_1637);
nand U5904 (N_5904,N_1583,N_22);
nand U5905 (N_5905,N_1184,N_1035);
and U5906 (N_5906,N_384,N_2193);
nor U5907 (N_5907,N_2709,N_527);
nor U5908 (N_5908,N_2472,N_1512);
and U5909 (N_5909,N_545,N_1810);
nand U5910 (N_5910,N_1784,N_2707);
and U5911 (N_5911,N_1988,N_1085);
and U5912 (N_5912,N_2007,N_432);
or U5913 (N_5913,N_1100,N_1581);
nor U5914 (N_5914,N_2171,N_285);
nor U5915 (N_5915,N_2836,N_1887);
nor U5916 (N_5916,N_2091,N_2320);
and U5917 (N_5917,N_2780,N_1442);
nand U5918 (N_5918,N_594,N_1440);
and U5919 (N_5919,N_2873,N_1628);
nand U5920 (N_5920,N_1684,N_2854);
or U5921 (N_5921,N_2320,N_1211);
nor U5922 (N_5922,N_2271,N_2858);
nand U5923 (N_5923,N_1633,N_824);
and U5924 (N_5924,N_1883,N_845);
nand U5925 (N_5925,N_1286,N_671);
nor U5926 (N_5926,N_2572,N_1986);
or U5927 (N_5927,N_58,N_2526);
and U5928 (N_5928,N_2466,N_2612);
and U5929 (N_5929,N_1431,N_1080);
nor U5930 (N_5930,N_386,N_2326);
and U5931 (N_5931,N_2066,N_1468);
or U5932 (N_5932,N_2744,N_1999);
and U5933 (N_5933,N_2233,N_1524);
nor U5934 (N_5934,N_745,N_2979);
nand U5935 (N_5935,N_338,N_1601);
nor U5936 (N_5936,N_1015,N_2212);
or U5937 (N_5937,N_1320,N_2060);
nand U5938 (N_5938,N_1328,N_2041);
nor U5939 (N_5939,N_875,N_1464);
and U5940 (N_5940,N_938,N_2835);
or U5941 (N_5941,N_183,N_330);
nor U5942 (N_5942,N_326,N_441);
and U5943 (N_5943,N_748,N_1582);
or U5944 (N_5944,N_1820,N_1359);
or U5945 (N_5945,N_2825,N_2814);
nand U5946 (N_5946,N_380,N_471);
xor U5947 (N_5947,N_1719,N_2935);
or U5948 (N_5948,N_232,N_1946);
and U5949 (N_5949,N_1822,N_2485);
and U5950 (N_5950,N_2680,N_943);
nand U5951 (N_5951,N_2731,N_574);
and U5952 (N_5952,N_2485,N_2605);
and U5953 (N_5953,N_1169,N_107);
nand U5954 (N_5954,N_1310,N_1097);
or U5955 (N_5955,N_146,N_2128);
nor U5956 (N_5956,N_241,N_2142);
or U5957 (N_5957,N_947,N_117);
and U5958 (N_5958,N_2843,N_2891);
or U5959 (N_5959,N_2984,N_1004);
nand U5960 (N_5960,N_2597,N_1741);
or U5961 (N_5961,N_1501,N_1098);
nor U5962 (N_5962,N_2995,N_838);
nor U5963 (N_5963,N_1773,N_2625);
nand U5964 (N_5964,N_1016,N_1786);
nand U5965 (N_5965,N_94,N_2785);
nand U5966 (N_5966,N_870,N_734);
nor U5967 (N_5967,N_1951,N_1696);
and U5968 (N_5968,N_936,N_2217);
and U5969 (N_5969,N_2436,N_2725);
or U5970 (N_5970,N_1080,N_2291);
or U5971 (N_5971,N_1371,N_1819);
and U5972 (N_5972,N_2845,N_77);
nand U5973 (N_5973,N_2910,N_2617);
nor U5974 (N_5974,N_1020,N_433);
and U5975 (N_5975,N_1285,N_2953);
or U5976 (N_5976,N_2489,N_690);
and U5977 (N_5977,N_1434,N_2908);
and U5978 (N_5978,N_515,N_2291);
nand U5979 (N_5979,N_2559,N_317);
and U5980 (N_5980,N_2624,N_438);
or U5981 (N_5981,N_1155,N_504);
and U5982 (N_5982,N_237,N_1498);
and U5983 (N_5983,N_1939,N_2793);
and U5984 (N_5984,N_2522,N_256);
nand U5985 (N_5985,N_2697,N_1519);
and U5986 (N_5986,N_544,N_411);
or U5987 (N_5987,N_122,N_1863);
and U5988 (N_5988,N_2761,N_1929);
and U5989 (N_5989,N_1110,N_311);
nor U5990 (N_5990,N_2081,N_2214);
and U5991 (N_5991,N_288,N_268);
nor U5992 (N_5992,N_1529,N_2262);
or U5993 (N_5993,N_1687,N_2452);
or U5994 (N_5994,N_231,N_1090);
nand U5995 (N_5995,N_1463,N_1460);
or U5996 (N_5996,N_420,N_2413);
xnor U5997 (N_5997,N_665,N_1960);
or U5998 (N_5998,N_2353,N_1066);
or U5999 (N_5999,N_2621,N_390);
nor U6000 (N_6000,N_3134,N_4368);
nand U6001 (N_6001,N_3792,N_3536);
and U6002 (N_6002,N_4415,N_4215);
nand U6003 (N_6003,N_3526,N_5707);
nor U6004 (N_6004,N_5211,N_3397);
nor U6005 (N_6005,N_3079,N_4107);
or U6006 (N_6006,N_5572,N_3868);
or U6007 (N_6007,N_5874,N_4818);
or U6008 (N_6008,N_3354,N_4063);
nor U6009 (N_6009,N_4367,N_5951);
nand U6010 (N_6010,N_4621,N_3326);
or U6011 (N_6011,N_4609,N_3346);
or U6012 (N_6012,N_4757,N_3214);
or U6013 (N_6013,N_5953,N_3320);
and U6014 (N_6014,N_4387,N_5623);
nor U6015 (N_6015,N_3288,N_3297);
or U6016 (N_6016,N_5223,N_4324);
or U6017 (N_6017,N_4699,N_3208);
or U6018 (N_6018,N_4200,N_3880);
or U6019 (N_6019,N_3499,N_3154);
or U6020 (N_6020,N_5231,N_4094);
nand U6021 (N_6021,N_4546,N_4954);
nor U6022 (N_6022,N_4297,N_4773);
or U6023 (N_6023,N_5626,N_3711);
nor U6024 (N_6024,N_3764,N_5757);
or U6025 (N_6025,N_5059,N_5304);
or U6026 (N_6026,N_5183,N_5361);
and U6027 (N_6027,N_3052,N_5030);
and U6028 (N_6028,N_4979,N_4947);
nor U6029 (N_6029,N_5614,N_4296);
nand U6030 (N_6030,N_3255,N_4596);
nand U6031 (N_6031,N_3666,N_4251);
nor U6032 (N_6032,N_5739,N_5063);
or U6033 (N_6033,N_5701,N_4775);
nor U6034 (N_6034,N_4008,N_4476);
nor U6035 (N_6035,N_3658,N_3284);
or U6036 (N_6036,N_5747,N_4010);
nor U6037 (N_6037,N_5932,N_5993);
or U6038 (N_6038,N_5759,N_3864);
or U6039 (N_6039,N_5831,N_5620);
or U6040 (N_6040,N_4338,N_5206);
or U6041 (N_6041,N_4208,N_5344);
nor U6042 (N_6042,N_3589,N_5649);
nor U6043 (N_6043,N_3782,N_4743);
and U6044 (N_6044,N_3547,N_3216);
nand U6045 (N_6045,N_4982,N_4407);
and U6046 (N_6046,N_3539,N_5177);
and U6047 (N_6047,N_5306,N_3631);
nor U6048 (N_6048,N_4352,N_5131);
and U6049 (N_6049,N_4740,N_5410);
nor U6050 (N_6050,N_4915,N_3862);
and U6051 (N_6051,N_4154,N_3137);
nand U6052 (N_6052,N_3998,N_3468);
and U6053 (N_6053,N_5546,N_3237);
and U6054 (N_6054,N_5413,N_5971);
nor U6055 (N_6055,N_5693,N_4265);
nor U6056 (N_6056,N_5411,N_5233);
nand U6057 (N_6057,N_4420,N_5870);
and U6058 (N_6058,N_3135,N_5862);
and U6059 (N_6059,N_4872,N_5067);
nand U6060 (N_6060,N_5170,N_5667);
and U6061 (N_6061,N_3457,N_4319);
and U6062 (N_6062,N_5172,N_3476);
or U6063 (N_6063,N_5659,N_3256);
or U6064 (N_6064,N_5889,N_5755);
and U6065 (N_6065,N_4687,N_5289);
and U6066 (N_6066,N_4584,N_3809);
or U6067 (N_6067,N_5429,N_4845);
or U6068 (N_6068,N_5612,N_4711);
and U6069 (N_6069,N_3550,N_3357);
nor U6070 (N_6070,N_3374,N_3837);
xnor U6071 (N_6071,N_5495,N_3840);
and U6072 (N_6072,N_4460,N_5291);
nor U6073 (N_6073,N_3599,N_4388);
or U6074 (N_6074,N_5330,N_3313);
nor U6075 (N_6075,N_5363,N_5408);
xor U6076 (N_6076,N_5671,N_5664);
nor U6077 (N_6077,N_3659,N_5081);
xnor U6078 (N_6078,N_5605,N_3701);
nor U6079 (N_6079,N_3181,N_4891);
nor U6080 (N_6080,N_4466,N_4177);
nor U6081 (N_6081,N_4893,N_4372);
or U6082 (N_6082,N_3147,N_4482);
nor U6083 (N_6083,N_4676,N_5343);
and U6084 (N_6084,N_5622,N_5725);
and U6085 (N_6085,N_5143,N_5758);
nand U6086 (N_6086,N_4813,N_4253);
nor U6087 (N_6087,N_3151,N_5902);
and U6088 (N_6088,N_3083,N_4206);
nor U6089 (N_6089,N_5348,N_5196);
or U6090 (N_6090,N_4897,N_3921);
nor U6091 (N_6091,N_4789,N_4874);
or U6092 (N_6092,N_4172,N_3946);
nand U6093 (N_6093,N_4179,N_3772);
or U6094 (N_6094,N_4169,N_4403);
and U6095 (N_6095,N_3300,N_4752);
nor U6096 (N_6096,N_4939,N_5458);
nor U6097 (N_6097,N_4247,N_4192);
or U6098 (N_6098,N_5591,N_3653);
and U6099 (N_6099,N_5723,N_4349);
xnor U6100 (N_6100,N_4287,N_4158);
and U6101 (N_6101,N_4330,N_4758);
or U6102 (N_6102,N_5207,N_4877);
or U6103 (N_6103,N_4607,N_5074);
nand U6104 (N_6104,N_4853,N_4722);
and U6105 (N_6105,N_3040,N_3213);
nor U6106 (N_6106,N_3872,N_3674);
nor U6107 (N_6107,N_5409,N_4073);
nand U6108 (N_6108,N_5954,N_5270);
nand U6109 (N_6109,N_4822,N_3465);
and U6110 (N_6110,N_3249,N_3591);
nor U6111 (N_6111,N_5097,N_3408);
and U6112 (N_6112,N_3218,N_4538);
nor U6113 (N_6113,N_4619,N_4375);
and U6114 (N_6114,N_5960,N_5508);
nand U6115 (N_6115,N_4274,N_4906);
nor U6116 (N_6116,N_5851,N_4197);
nor U6117 (N_6117,N_4421,N_4439);
nand U6118 (N_6118,N_5029,N_4858);
nand U6119 (N_6119,N_4737,N_4149);
nor U6120 (N_6120,N_4186,N_3736);
nand U6121 (N_6121,N_4969,N_4955);
nor U6122 (N_6122,N_4020,N_5194);
and U6123 (N_6123,N_5997,N_5673);
and U6124 (N_6124,N_4512,N_3286);
and U6125 (N_6125,N_5630,N_3673);
xor U6126 (N_6126,N_3308,N_5446);
or U6127 (N_6127,N_5921,N_3363);
and U6128 (N_6128,N_4912,N_4762);
or U6129 (N_6129,N_3239,N_4417);
nand U6130 (N_6130,N_4385,N_5080);
or U6131 (N_6131,N_4637,N_5307);
nor U6132 (N_6132,N_5009,N_4289);
nor U6133 (N_6133,N_3209,N_5093);
or U6134 (N_6134,N_3480,N_5950);
nand U6135 (N_6135,N_5527,N_4936);
nor U6136 (N_6136,N_3765,N_3716);
and U6137 (N_6137,N_4007,N_5171);
nor U6138 (N_6138,N_4677,N_5703);
and U6139 (N_6139,N_4196,N_4889);
nor U6140 (N_6140,N_4044,N_3339);
and U6141 (N_6141,N_3632,N_3474);
and U6142 (N_6142,N_4127,N_4641);
and U6143 (N_6143,N_5140,N_4927);
nor U6144 (N_6144,N_3285,N_5749);
nor U6145 (N_6145,N_3254,N_3004);
nand U6146 (N_6146,N_3000,N_5505);
nand U6147 (N_6147,N_3478,N_3777);
nand U6148 (N_6148,N_4646,N_4854);
and U6149 (N_6149,N_3062,N_3890);
nor U6150 (N_6150,N_4561,N_3867);
and U6151 (N_6151,N_3511,N_5275);
nand U6152 (N_6152,N_4507,N_3459);
and U6153 (N_6153,N_5611,N_5876);
or U6154 (N_6154,N_4956,N_5577);
nand U6155 (N_6155,N_5991,N_5435);
and U6156 (N_6156,N_5491,N_4697);
or U6157 (N_6157,N_5051,N_5199);
or U6158 (N_6158,N_4294,N_3801);
or U6159 (N_6159,N_4662,N_5264);
nor U6160 (N_6160,N_4738,N_5047);
nand U6161 (N_6161,N_3574,N_3570);
nand U6162 (N_6162,N_5226,N_5216);
nand U6163 (N_6163,N_5853,N_4214);
or U6164 (N_6164,N_4564,N_3755);
nor U6165 (N_6165,N_4363,N_4620);
nand U6166 (N_6166,N_5012,N_3085);
or U6167 (N_6167,N_5881,N_3403);
and U6168 (N_6168,N_5235,N_3595);
and U6169 (N_6169,N_3241,N_4767);
and U6170 (N_6170,N_5316,N_5002);
nand U6171 (N_6171,N_3846,N_4068);
and U6172 (N_6172,N_3875,N_3540);
nand U6173 (N_6173,N_5838,N_3234);
nand U6174 (N_6174,N_5869,N_4978);
and U6175 (N_6175,N_4601,N_3163);
and U6176 (N_6176,N_3194,N_4503);
and U6177 (N_6177,N_3498,N_5273);
nand U6178 (N_6178,N_4292,N_4097);
and U6179 (N_6179,N_5368,N_5694);
nor U6180 (N_6180,N_5990,N_5432);
nor U6181 (N_6181,N_4949,N_4944);
nand U6182 (N_6182,N_3033,N_3871);
nand U6183 (N_6183,N_5061,N_4051);
nand U6184 (N_6184,N_4361,N_4772);
nor U6185 (N_6185,N_4993,N_4760);
xor U6186 (N_6186,N_4973,N_5357);
or U6187 (N_6187,N_3857,N_3024);
and U6188 (N_6188,N_5507,N_5462);
nand U6189 (N_6189,N_5863,N_3275);
nand U6190 (N_6190,N_4136,N_5896);
nand U6191 (N_6191,N_4272,N_3829);
nand U6192 (N_6192,N_5662,N_4353);
nor U6193 (N_6193,N_3352,N_5007);
or U6194 (N_6194,N_5371,N_4376);
nor U6195 (N_6195,N_5824,N_3379);
nor U6196 (N_6196,N_4867,N_4032);
and U6197 (N_6197,N_3876,N_3433);
nand U6198 (N_6198,N_5342,N_3334);
and U6199 (N_6199,N_3202,N_4232);
and U6200 (N_6200,N_5854,N_5310);
nand U6201 (N_6201,N_4919,N_4748);
nand U6202 (N_6202,N_5384,N_5204);
nor U6203 (N_6203,N_5492,N_3703);
or U6204 (N_6204,N_3123,N_4074);
or U6205 (N_6205,N_5980,N_3825);
and U6206 (N_6206,N_4463,N_3099);
nor U6207 (N_6207,N_4280,N_3970);
and U6208 (N_6208,N_3055,N_4050);
and U6209 (N_6209,N_4565,N_5493);
or U6210 (N_6210,N_5924,N_3232);
or U6211 (N_6211,N_4670,N_5983);
nor U6212 (N_6212,N_4930,N_4120);
nand U6213 (N_6213,N_4878,N_4021);
and U6214 (N_6214,N_4497,N_4461);
nor U6215 (N_6215,N_5778,N_5276);
nor U6216 (N_6216,N_5509,N_4147);
and U6217 (N_6217,N_3979,N_5048);
nor U6218 (N_6218,N_5102,N_4494);
and U6219 (N_6219,N_4418,N_5142);
nor U6220 (N_6220,N_4259,N_3221);
or U6221 (N_6221,N_4741,N_3307);
xnor U6222 (N_6222,N_5670,N_4254);
nor U6223 (N_6223,N_4034,N_5750);
nor U6224 (N_6224,N_4309,N_3283);
nor U6225 (N_6225,N_5958,N_5549);
nand U6226 (N_6226,N_5920,N_3974);
and U6227 (N_6227,N_4731,N_4317);
and U6228 (N_6228,N_3586,N_5443);
nand U6229 (N_6229,N_3634,N_5001);
and U6230 (N_6230,N_5871,N_4709);
or U6231 (N_6231,N_5387,N_3253);
nor U6232 (N_6232,N_3037,N_4583);
and U6233 (N_6233,N_3422,N_4163);
nand U6234 (N_6234,N_3827,N_5433);
nor U6235 (N_6235,N_3210,N_4419);
nand U6236 (N_6236,N_5710,N_4873);
nand U6237 (N_6237,N_3662,N_5114);
nor U6238 (N_6238,N_3173,N_5872);
or U6239 (N_6239,N_4673,N_5374);
and U6240 (N_6240,N_5516,N_5916);
nand U6241 (N_6241,N_4467,N_4371);
or U6242 (N_6242,N_5910,N_4125);
and U6243 (N_6243,N_3661,N_3271);
nor U6244 (N_6244,N_4411,N_4382);
or U6245 (N_6245,N_5781,N_4436);
or U6246 (N_6246,N_5089,N_5552);
nand U6247 (N_6247,N_3928,N_3937);
and U6248 (N_6248,N_5841,N_3545);
nor U6249 (N_6249,N_3458,N_3467);
or U6250 (N_6250,N_3748,N_4631);
nor U6251 (N_6251,N_5607,N_5846);
nand U6252 (N_6252,N_5379,N_5883);
nor U6253 (N_6253,N_5192,N_3046);
nor U6254 (N_6254,N_5415,N_5441);
nor U6255 (N_6255,N_5221,N_3048);
nand U6256 (N_6256,N_4487,N_4183);
and U6257 (N_6257,N_5407,N_4556);
or U6258 (N_6258,N_3053,N_5215);
and U6259 (N_6259,N_5692,N_4513);
nor U6260 (N_6260,N_5726,N_5394);
or U6261 (N_6261,N_5796,N_3312);
or U6262 (N_6262,N_4984,N_3510);
nor U6263 (N_6263,N_3966,N_4935);
nor U6264 (N_6264,N_5115,N_4322);
nor U6265 (N_6265,N_4346,N_5793);
and U6266 (N_6266,N_5949,N_4462);
and U6267 (N_6267,N_3031,N_3897);
and U6268 (N_6268,N_5298,N_4043);
and U6269 (N_6269,N_4345,N_4537);
nand U6270 (N_6270,N_3371,N_3569);
or U6271 (N_6271,N_5279,N_4568);
nor U6272 (N_6272,N_4207,N_3344);
nor U6273 (N_6273,N_3236,N_5992);
nand U6274 (N_6274,N_3315,N_3084);
nor U6275 (N_6275,N_4655,N_3245);
nor U6276 (N_6276,N_5892,N_4479);
and U6277 (N_6277,N_3565,N_3649);
or U6278 (N_6278,N_3775,N_5158);
and U6279 (N_6279,N_3988,N_4140);
nand U6280 (N_6280,N_5460,N_4155);
nor U6281 (N_6281,N_4270,N_4672);
nor U6282 (N_6282,N_3532,N_4119);
xor U6283 (N_6283,N_3906,N_4255);
or U6284 (N_6284,N_3874,N_3087);
or U6285 (N_6285,N_3566,N_3918);
and U6286 (N_6286,N_3115,N_5897);
xor U6287 (N_6287,N_3412,N_3955);
and U6288 (N_6288,N_5700,N_3528);
nor U6289 (N_6289,N_5780,N_4435);
nor U6290 (N_6290,N_3567,N_3222);
nand U6291 (N_6291,N_5644,N_4887);
and U6292 (N_6292,N_5702,N_5193);
or U6293 (N_6293,N_5331,N_4967);
and U6294 (N_6294,N_5464,N_4027);
and U6295 (N_6295,N_4799,N_3069);
nand U6296 (N_6296,N_5537,N_5174);
nand U6297 (N_6297,N_5359,N_4381);
and U6298 (N_6298,N_3907,N_4794);
nor U6299 (N_6299,N_5506,N_3542);
and U6300 (N_6300,N_3272,N_5731);
nand U6301 (N_6301,N_3851,N_4733);
and U6302 (N_6302,N_3885,N_3665);
and U6303 (N_6303,N_4938,N_5720);
nor U6304 (N_6304,N_5011,N_3296);
nand U6305 (N_6305,N_3035,N_5480);
and U6306 (N_6306,N_4855,N_3858);
nor U6307 (N_6307,N_5466,N_5256);
nand U6308 (N_6308,N_4262,N_5925);
or U6309 (N_6309,N_5165,N_5149);
and U6310 (N_6310,N_3109,N_3022);
and U6311 (N_6311,N_4100,N_5116);
or U6312 (N_6312,N_5985,N_5332);
and U6313 (N_6313,N_3602,N_5467);
nand U6314 (N_6314,N_5447,N_5996);
nor U6315 (N_6315,N_3290,N_4340);
and U6316 (N_6316,N_3699,N_4905);
and U6317 (N_6317,N_5661,N_3546);
or U6318 (N_6318,N_4827,N_3789);
or U6319 (N_6319,N_4541,N_4618);
or U6320 (N_6320,N_4424,N_5209);
or U6321 (N_6321,N_5698,N_4001);
or U6322 (N_6322,N_5683,N_5355);
and U6323 (N_6323,N_5254,N_4377);
nor U6324 (N_6324,N_4527,N_5807);
nor U6325 (N_6325,N_3977,N_3964);
and U6326 (N_6326,N_5141,N_5760);
nor U6327 (N_6327,N_4425,N_3615);
and U6328 (N_6328,N_5973,N_5322);
and U6329 (N_6329,N_5785,N_3404);
and U6330 (N_6330,N_3576,N_3002);
nor U6331 (N_6331,N_3803,N_5064);
nor U6332 (N_6332,N_4765,N_3445);
nand U6333 (N_6333,N_5634,N_5351);
nand U6334 (N_6334,N_5907,N_4937);
or U6335 (N_6335,N_3961,N_5904);
and U6336 (N_6336,N_5453,N_3332);
nor U6337 (N_6337,N_4201,N_3282);
and U6338 (N_6338,N_4329,N_4633);
nor U6339 (N_6339,N_4521,N_3618);
or U6340 (N_6340,N_3075,N_4282);
and U6341 (N_6341,N_4080,N_3912);
or U6342 (N_6342,N_5220,N_3952);
or U6343 (N_6343,N_5285,N_3783);
nor U6344 (N_6344,N_3947,N_3353);
and U6345 (N_6345,N_3351,N_4408);
nor U6346 (N_6346,N_3451,N_5303);
xnor U6347 (N_6347,N_4456,N_4263);
and U6348 (N_6348,N_3122,N_3889);
or U6349 (N_6349,N_3273,N_3621);
or U6350 (N_6350,N_3780,N_5260);
and U6351 (N_6351,N_5156,N_4380);
nand U6352 (N_6352,N_5547,N_5619);
and U6353 (N_6353,N_3042,N_4724);
and U6354 (N_6354,N_5104,N_5939);
nand U6355 (N_6355,N_3915,N_5763);
or U6356 (N_6356,N_4834,N_4328);
nor U6357 (N_6357,N_5200,N_3367);
or U6358 (N_6358,N_5034,N_3520);
nor U6359 (N_6359,N_4431,N_5403);
nor U6360 (N_6360,N_3169,N_3359);
and U6361 (N_6361,N_5367,N_3270);
or U6362 (N_6362,N_3039,N_4173);
or U6363 (N_6363,N_5642,N_5989);
nand U6364 (N_6364,N_5684,N_5272);
and U6365 (N_6365,N_5471,N_4019);
nand U6366 (N_6366,N_3014,N_5548);
or U6367 (N_6367,N_5933,N_3149);
and U6368 (N_6368,N_4028,N_4812);
and U6369 (N_6369,N_3369,N_3901);
and U6370 (N_6370,N_5370,N_3905);
nor U6371 (N_6371,N_3804,N_5008);
nor U6372 (N_6372,N_4657,N_5946);
and U6373 (N_6373,N_5789,N_4493);
or U6374 (N_6374,N_5817,N_5137);
nor U6375 (N_6375,N_5998,N_3242);
and U6376 (N_6376,N_5058,N_3795);
nor U6377 (N_6377,N_3489,N_4106);
xor U6378 (N_6378,N_5682,N_5497);
xnor U6379 (N_6379,N_3318,N_4985);
nand U6380 (N_6380,N_5062,N_5345);
nor U6381 (N_6381,N_4405,N_3933);
nor U6382 (N_6382,N_3544,N_3903);
and U6383 (N_6383,N_5969,N_3852);
or U6384 (N_6384,N_5833,N_3252);
and U6385 (N_6385,N_3244,N_5487);
nor U6386 (N_6386,N_3936,N_3409);
nor U6387 (N_6387,N_5783,N_5968);
or U6388 (N_6388,N_5406,N_5286);
and U6389 (N_6389,N_3814,N_3925);
or U6390 (N_6390,N_4747,N_3693);
and U6391 (N_6391,N_3939,N_4240);
and U6392 (N_6392,N_4252,N_5995);
nor U6393 (N_6393,N_4782,N_5772);
nand U6394 (N_6394,N_3580,N_5761);
and U6395 (N_6395,N_3924,N_4830);
or U6396 (N_6396,N_3041,N_5227);
nor U6397 (N_6397,N_5918,N_5654);
xnor U6398 (N_6398,N_3365,N_3714);
xnor U6399 (N_6399,N_5557,N_5346);
and U6400 (N_6400,N_5139,N_4053);
and U6401 (N_6401,N_5650,N_3168);
or U6402 (N_6402,N_5929,N_5773);
and U6403 (N_6403,N_4734,N_5651);
nand U6404 (N_6404,N_5603,N_3093);
or U6405 (N_6405,N_3267,N_4736);
nand U6406 (N_6406,N_3056,N_5522);
nand U6407 (N_6407,N_3295,N_4404);
nor U6408 (N_6408,N_5685,N_4800);
or U6409 (N_6409,N_4248,N_5392);
xnor U6410 (N_6410,N_3461,N_5455);
nor U6411 (N_6411,N_5043,N_5257);
xnor U6412 (N_6412,N_3140,N_4608);
nor U6413 (N_6413,N_4178,N_3951);
nor U6414 (N_6414,N_5716,N_5909);
and U6415 (N_6415,N_4249,N_4884);
nand U6416 (N_6416,N_5625,N_5556);
and U6417 (N_6417,N_4667,N_5900);
nand U6418 (N_6418,N_4303,N_4597);
or U6419 (N_6419,N_4766,N_4728);
nand U6420 (N_6420,N_4904,N_3479);
nor U6421 (N_6421,N_4438,N_3057);
nand U6422 (N_6422,N_4305,N_3101);
and U6423 (N_6423,N_4116,N_3424);
and U6424 (N_6424,N_3475,N_3562);
nand U6425 (N_6425,N_4909,N_4591);
and U6426 (N_6426,N_4841,N_3640);
nor U6427 (N_6427,N_4627,N_3483);
nand U6428 (N_6428,N_4454,N_5751);
or U6429 (N_6429,N_5737,N_4486);
nor U6430 (N_6430,N_3342,N_5105);
nor U6431 (N_6431,N_4496,N_5035);
nor U6432 (N_6432,N_3654,N_4886);
nor U6433 (N_6433,N_3677,N_3347);
and U6434 (N_6434,N_3197,N_4614);
nor U6435 (N_6435,N_5888,N_3442);
or U6436 (N_6436,N_3446,N_3579);
and U6437 (N_6437,N_3926,N_5239);
or U6438 (N_6438,N_5880,N_5228);
or U6439 (N_6439,N_5593,N_3452);
xnor U6440 (N_6440,N_5978,N_3734);
xor U6441 (N_6441,N_5500,N_5248);
nor U6442 (N_6442,N_3155,N_5135);
or U6443 (N_6443,N_4185,N_3807);
nand U6444 (N_6444,N_5952,N_5959);
and U6445 (N_6445,N_5945,N_5917);
nand U6446 (N_6446,N_3380,N_4659);
nor U6447 (N_6447,N_3005,N_5770);
and U6448 (N_6448,N_5117,N_5324);
or U6449 (N_6449,N_4603,N_5476);
nor U6450 (N_6450,N_5326,N_3657);
nor U6451 (N_6451,N_3306,N_4908);
or U6452 (N_6452,N_4558,N_3798);
nand U6453 (N_6453,N_4374,N_3484);
nor U6454 (N_6454,N_5882,N_3753);
or U6455 (N_6455,N_5456,N_3130);
nand U6456 (N_6456,N_3643,N_5887);
nand U6457 (N_6457,N_3120,N_3393);
nor U6458 (N_6458,N_4784,N_5784);
or U6459 (N_6459,N_4666,N_3899);
and U6460 (N_6460,N_5567,N_3172);
nor U6461 (N_6461,N_4778,N_3684);
nand U6462 (N_6462,N_5159,N_3455);
and U6463 (N_6463,N_5736,N_3292);
or U6464 (N_6464,N_5629,N_5844);
nor U6465 (N_6465,N_5499,N_4612);
or U6466 (N_6466,N_5004,N_4151);
and U6467 (N_6467,N_4427,N_3894);
or U6468 (N_6468,N_3248,N_4536);
or U6469 (N_6469,N_3026,N_5134);
or U6470 (N_6470,N_3166,N_5901);
nor U6471 (N_6471,N_4237,N_4002);
nand U6472 (N_6472,N_5444,N_3124);
or U6473 (N_6473,N_5999,N_3324);
and U6474 (N_6474,N_4446,N_3706);
and U6475 (N_6475,N_4219,N_5461);
xnor U6476 (N_6476,N_4242,N_4756);
or U6477 (N_6477,N_5704,N_5812);
nor U6478 (N_6478,N_5022,N_3051);
nand U6479 (N_6479,N_5049,N_4847);
and U6480 (N_6480,N_3470,N_4182);
nor U6481 (N_6481,N_3750,N_3554);
nor U6482 (N_6482,N_4428,N_3487);
and U6483 (N_6483,N_3896,N_4257);
or U6484 (N_6484,N_3118,N_4518);
nand U6485 (N_6485,N_4373,N_5964);
nand U6486 (N_6486,N_4959,N_5376);
nand U6487 (N_6487,N_4866,N_4038);
nand U6488 (N_6488,N_4194,N_4708);
and U6489 (N_6489,N_5928,N_5775);
nand U6490 (N_6490,N_4300,N_4894);
and U6491 (N_6491,N_4974,N_5600);
or U6492 (N_6492,N_5715,N_5768);
nor U6493 (N_6493,N_5318,N_5616);
nor U6494 (N_6494,N_3877,N_5294);
and U6495 (N_6495,N_3349,N_4205);
or U6496 (N_6496,N_3212,N_3806);
nor U6497 (N_6497,N_5110,N_3170);
and U6498 (N_6498,N_5563,N_3260);
and U6499 (N_6499,N_5656,N_5734);
nor U6500 (N_6500,N_5075,N_3770);
or U6501 (N_6501,N_5391,N_5938);
or U6502 (N_6502,N_3594,N_4654);
or U6503 (N_6503,N_5375,N_3377);
nand U6504 (N_6504,N_3329,N_5621);
or U6505 (N_6505,N_5293,N_5558);
nor U6506 (N_6506,N_3942,N_3145);
nand U6507 (N_6507,N_3453,N_5970);
or U6508 (N_6508,N_4774,N_4869);
and U6509 (N_6509,N_5555,N_4014);
nand U6510 (N_6510,N_5108,N_5399);
and U6511 (N_6511,N_5800,N_3269);
or U6512 (N_6512,N_5186,N_3873);
nor U6513 (N_6513,N_3086,N_3454);
nand U6514 (N_6514,N_5054,N_5631);
or U6515 (N_6515,N_5085,N_3078);
or U6516 (N_6516,N_3530,N_3590);
or U6517 (N_6517,N_5389,N_5609);
nor U6518 (N_6518,N_5756,N_5697);
and U6519 (N_6519,N_5961,N_4770);
or U6520 (N_6520,N_3639,N_3321);
nor U6521 (N_6521,N_4058,N_4628);
nor U6522 (N_6522,N_5249,N_3104);
nand U6523 (N_6523,N_3695,N_3604);
nand U6524 (N_6524,N_4171,N_4269);
nand U6525 (N_6525,N_3375,N_4828);
or U6526 (N_6526,N_5336,N_3129);
and U6527 (N_6527,N_4108,N_5419);
nor U6528 (N_6528,N_4848,N_4473);
and U6529 (N_6529,N_5060,N_4084);
nand U6530 (N_6530,N_3201,N_3663);
nor U6531 (N_6531,N_3378,N_5822);
nor U6532 (N_6532,N_3385,N_3516);
nand U6533 (N_6533,N_4003,N_4464);
or U6534 (N_6534,N_5442,N_4124);
and U6535 (N_6535,N_3886,N_5280);
and U6536 (N_6536,N_5295,N_3515);
and U6537 (N_6537,N_3449,N_4732);
nor U6538 (N_6538,N_3386,N_4323);
or U6539 (N_6539,N_5224,N_3805);
or U6540 (N_6540,N_3860,N_5674);
xnor U6541 (N_6541,N_3497,N_4085);
and U6542 (N_6542,N_4811,N_4525);
or U6543 (N_6543,N_4041,N_4776);
and U6544 (N_6544,N_4204,N_4181);
or U6545 (N_6545,N_4261,N_5559);
and U6546 (N_6546,N_4998,N_3548);
nor U6547 (N_6547,N_3094,N_3609);
or U6548 (N_6548,N_3396,N_3549);
or U6549 (N_6549,N_4318,N_4604);
or U6550 (N_6550,N_3731,N_5681);
nor U6551 (N_6551,N_5095,N_4184);
and U6552 (N_6552,N_5053,N_3192);
nand U6553 (N_6553,N_3088,N_5148);
or U6554 (N_6554,N_5994,N_3729);
nand U6555 (N_6555,N_4926,N_5263);
nor U6556 (N_6556,N_5266,N_3504);
and U6557 (N_6557,N_5618,N_3940);
or U6558 (N_6558,N_4006,N_3074);
nor U6559 (N_6559,N_5107,N_4046);
nand U6560 (N_6560,N_4600,N_4567);
or U6561 (N_6561,N_3893,N_4152);
nor U6562 (N_6562,N_5913,N_5849);
nand U6563 (N_6563,N_3223,N_5122);
and U6564 (N_6564,N_5203,N_5353);
and U6565 (N_6565,N_4190,N_5601);
nor U6566 (N_6566,N_4754,N_3191);
nand U6567 (N_6567,N_3050,N_4611);
or U6568 (N_6568,N_5023,N_5101);
nand U6569 (N_6569,N_3644,N_4160);
nand U6570 (N_6570,N_4669,N_3605);
or U6571 (N_6571,N_5769,N_5111);
or U6572 (N_6572,N_5337,N_4807);
or U6573 (N_6573,N_5823,N_3368);
nor U6574 (N_6574,N_5470,N_3635);
nor U6575 (N_6575,N_4320,N_4883);
or U6576 (N_6576,N_3622,N_4311);
nand U6577 (N_6577,N_5835,N_5561);
xnor U6578 (N_6578,N_4447,N_5155);
and U6579 (N_6579,N_4833,N_3065);
nand U6580 (N_6580,N_4634,N_5205);
nand U6581 (N_6581,N_5393,N_4490);
or U6582 (N_6582,N_4806,N_5746);
nor U6583 (N_6583,N_3848,N_4831);
nand U6584 (N_6584,N_3881,N_4815);
nor U6585 (N_6585,N_4332,N_3747);
and U6586 (N_6586,N_4065,N_4012);
and U6587 (N_6587,N_3788,N_3943);
nor U6588 (N_6588,N_4095,N_3405);
nor U6589 (N_6589,N_5082,N_4999);
and U6590 (N_6590,N_4976,N_5185);
or U6591 (N_6591,N_3543,N_5312);
nor U6592 (N_6592,N_3443,N_5740);
nand U6593 (N_6593,N_5364,N_3686);
or U6594 (N_6594,N_4267,N_3148);
and U6595 (N_6595,N_5847,N_5106);
or U6596 (N_6596,N_5752,N_3398);
nand U6597 (N_6597,N_5977,N_5127);
or U6598 (N_6598,N_4144,N_5602);
or U6599 (N_6599,N_5428,N_4729);
and U6600 (N_6600,N_4577,N_5504);
or U6601 (N_6601,N_5788,N_3537);
nor U6602 (N_6602,N_4016,N_4868);
and U6603 (N_6603,N_5606,N_3277);
and U6604 (N_6604,N_3931,N_4749);
nor U6605 (N_6605,N_3717,N_3702);
or U6606 (N_6606,N_3331,N_5613);
nor U6607 (N_6607,N_5405,N_3981);
nand U6608 (N_6608,N_3738,N_4397);
xor U6609 (N_6609,N_5573,N_3356);
and U6610 (N_6610,N_5418,N_5259);
nor U6611 (N_6611,N_5839,N_3142);
nor U6612 (N_6612,N_3991,N_3514);
nor U6613 (N_6613,N_4039,N_5242);
and U6614 (N_6614,N_4118,N_5845);
nor U6615 (N_6615,N_3150,N_3709);
nor U6616 (N_6616,N_4535,N_4203);
and U6617 (N_6617,N_4643,N_3651);
nor U6618 (N_6618,N_3821,N_5582);
nand U6619 (N_6619,N_4351,N_3448);
or U6620 (N_6620,N_5277,N_4187);
nand U6621 (N_6621,N_5586,N_3020);
or U6622 (N_6622,N_5164,N_3276);
nor U6623 (N_6623,N_4335,N_5512);
nor U6624 (N_6624,N_3888,N_5840);
nor U6625 (N_6625,N_5040,N_3413);
or U6626 (N_6626,N_3841,N_4092);
nor U6627 (N_6627,N_5315,N_4768);
and U6628 (N_6628,N_4700,N_4649);
or U6629 (N_6629,N_3938,N_4651);
or U6630 (N_6630,N_5923,N_4040);
nor U6631 (N_6631,N_3650,N_3250);
nand U6632 (N_6632,N_5792,N_3364);
nor U6633 (N_6633,N_5641,N_4958);
and U6634 (N_6634,N_4434,N_4863);
nand U6635 (N_6635,N_3362,N_5617);
or U6636 (N_6636,N_5191,N_4791);
nand U6637 (N_6637,N_3898,N_4410);
nor U6638 (N_6638,N_4804,N_5590);
and U6639 (N_6639,N_5711,N_4440);
and U6640 (N_6640,N_5297,N_4679);
nor U6641 (N_6641,N_4105,N_4980);
or U6642 (N_6642,N_5153,N_3957);
or U6643 (N_6643,N_5440,N_4458);
nand U6644 (N_6644,N_3161,N_4229);
or U6645 (N_6645,N_5672,N_5321);
nor U6646 (N_6646,N_3401,N_4553);
or U6647 (N_6647,N_5754,N_3360);
nor U6648 (N_6648,N_3010,N_5915);
nand U6649 (N_6649,N_5967,N_3724);
nor U6650 (N_6650,N_3527,N_4552);
or U6651 (N_6651,N_3138,N_4429);
nand U6652 (N_6652,N_3687,N_4457);
or U6653 (N_6653,N_5282,N_5930);
or U6654 (N_6654,N_4437,N_5163);
xor U6655 (N_6655,N_4640,N_3407);
nor U6656 (N_6656,N_5718,N_4587);
and U6657 (N_6657,N_5426,N_5748);
or U6658 (N_6658,N_3557,N_4299);
nand U6659 (N_6659,N_3495,N_3429);
and U6660 (N_6660,N_3355,N_3956);
or U6661 (N_6661,N_3646,N_3279);
nor U6662 (N_6662,N_3311,N_3815);
nand U6663 (N_6663,N_5816,N_3810);
nand U6664 (N_6664,N_3568,N_3293);
or U6665 (N_6665,N_4139,N_5890);
nand U6666 (N_6666,N_4389,N_5687);
nor U6667 (N_6667,N_3506,N_5436);
nand U6668 (N_6668,N_3660,N_4011);
nor U6669 (N_6669,N_4064,N_3972);
and U6670 (N_6670,N_3119,N_3762);
nor U6671 (N_6671,N_4717,N_4268);
or U6672 (N_6672,N_5157,N_3190);
nor U6673 (N_6673,N_4307,N_3749);
or U6674 (N_6674,N_5245,N_5457);
and U6675 (N_6675,N_3337,N_4223);
and U6676 (N_6676,N_3509,N_4316);
nor U6677 (N_6677,N_3802,N_3561);
and U6678 (N_6678,N_4759,N_3923);
or U6679 (N_6679,N_5525,N_5084);
and U6680 (N_6680,N_4639,N_5396);
or U6681 (N_6681,N_5764,N_3911);
nor U6682 (N_6682,N_4630,N_4644);
nand U6683 (N_6683,N_3882,N_5802);
and U6684 (N_6684,N_5753,N_3989);
nand U6685 (N_6685,N_4792,N_4862);
nor U6686 (N_6686,N_3064,N_5146);
nand U6687 (N_6687,N_5168,N_3471);
or U6688 (N_6688,N_5927,N_5639);
nor U6689 (N_6689,N_3188,N_5129);
or U6690 (N_6690,N_3533,N_4198);
nor U6691 (N_6691,N_4570,N_3521);
or U6692 (N_6692,N_3430,N_5501);
nor U6693 (N_6693,N_3512,N_5790);
nand U6694 (N_6694,N_3564,N_5866);
and U6695 (N_6695,N_4622,N_5320);
nor U6696 (N_6696,N_3968,N_3597);
or U6697 (N_6697,N_3559,N_5037);
and U6698 (N_6698,N_5056,N_4860);
xnor U6699 (N_6699,N_3922,N_5308);
and U6700 (N_6700,N_4531,N_3419);
or U6701 (N_6701,N_5898,N_4835);
and U6702 (N_6702,N_3127,N_5706);
or U6703 (N_6703,N_3133,N_5518);
or U6704 (N_6704,N_3975,N_3727);
and U6705 (N_6705,N_5903,N_5615);
nor U6706 (N_6706,N_5598,N_3917);
nor U6707 (N_6707,N_3183,N_3301);
and U6708 (N_6708,N_5589,N_3529);
nand U6709 (N_6709,N_5984,N_4691);
or U6710 (N_6710,N_4432,N_4802);
nor U6711 (N_6711,N_5283,N_3690);
and U6712 (N_6712,N_4642,N_5451);
nand U6713 (N_6713,N_5688,N_3844);
and U6714 (N_6714,N_5865,N_3629);
nand U6715 (N_6715,N_3689,N_4101);
and U6716 (N_6716,N_5144,N_4113);
nor U6717 (N_6717,N_4968,N_3555);
or U6718 (N_6718,N_5019,N_5328);
or U6719 (N_6719,N_3323,N_3784);
or U6720 (N_6720,N_4230,N_4209);
or U6721 (N_6721,N_5229,N_4735);
and U6722 (N_6722,N_4975,N_5079);
or U6723 (N_6723,N_4083,N_3143);
and U6724 (N_6724,N_3856,N_4067);
or U6725 (N_6725,N_5905,N_5068);
or U6726 (N_6726,N_3583,N_4715);
and U6727 (N_6727,N_5267,N_4033);
or U6728 (N_6728,N_3552,N_4036);
nand U6729 (N_6729,N_5676,N_4595);
and U6730 (N_6730,N_4961,N_3679);
xnor U6731 (N_6731,N_3251,N_4394);
and U6732 (N_6732,N_5765,N_4071);
xnor U6733 (N_6733,N_5169,N_4971);
nand U6734 (N_6734,N_5502,N_4054);
nor U6735 (N_6735,N_5100,N_4864);
and U6736 (N_6736,N_3460,N_3743);
or U6737 (N_6737,N_5583,N_3016);
nand U6738 (N_6738,N_5542,N_4952);
or U6739 (N_6739,N_5732,N_4298);
or U6740 (N_6740,N_3280,N_5517);
and U6741 (N_6741,N_5689,N_5690);
or U6742 (N_6742,N_4228,N_4217);
nand U6743 (N_6743,N_5979,N_3577);
nor U6744 (N_6744,N_5861,N_3773);
nand U6745 (N_6745,N_3818,N_5624);
and U6746 (N_6746,N_5519,N_4585);
or U6747 (N_6747,N_4055,N_5535);
nand U6748 (N_6748,N_4505,N_4304);
and U6749 (N_6749,N_4180,N_4852);
and U6750 (N_6750,N_4188,N_5121);
and U6751 (N_6751,N_4285,N_3215);
nor U6752 (N_6752,N_3153,N_3694);
nand U6753 (N_6753,N_5133,N_3633);
and U6754 (N_6754,N_5333,N_4060);
or U6755 (N_6755,N_4288,N_5125);
nor U6756 (N_6756,N_3327,N_3920);
or U6757 (N_6757,N_5118,N_3097);
nand U6758 (N_6758,N_5814,N_3211);
or U6759 (N_6759,N_3441,N_3350);
nand U6760 (N_6760,N_5338,N_3853);
nor U6761 (N_6761,N_4452,N_5894);
nor U6762 (N_6762,N_5680,N_3496);
nand U6763 (N_6763,N_4256,N_5696);
nor U6764 (N_6764,N_3675,N_3287);
or U6765 (N_6765,N_5390,N_5608);
xor U6766 (N_6766,N_5825,N_4369);
and U6767 (N_6767,N_4359,N_4781);
or U6768 (N_6768,N_3322,N_5188);
and U6769 (N_6769,N_5098,N_3167);
nor U6770 (N_6770,N_4843,N_5791);
or U6771 (N_6771,N_4616,N_4495);
or U6772 (N_6772,N_5350,N_4226);
and U6773 (N_6773,N_4920,N_3704);
or U6774 (N_6774,N_3158,N_5162);
and U6775 (N_6775,N_4885,N_3017);
nor U6776 (N_6776,N_4104,N_3719);
or U6777 (N_6777,N_5092,N_3420);
nor U6778 (N_6778,N_3910,N_4589);
nor U6779 (N_6779,N_4327,N_4689);
nor U6780 (N_6780,N_3999,N_4037);
nand U6781 (N_6781,N_4343,N_5744);
or U6782 (N_6782,N_4308,N_4337);
or U6783 (N_6783,N_5550,N_3341);
or U6784 (N_6784,N_5962,N_4880);
or U6785 (N_6785,N_3757,N_3068);
nor U6786 (N_6786,N_4114,N_3012);
and U6787 (N_6787,N_4480,N_5167);
xor U6788 (N_6788,N_5027,N_3108);
nand U6789 (N_6789,N_4808,N_4686);
nor U6790 (N_6790,N_4576,N_4519);
nor U6791 (N_6791,N_3246,N_5893);
or U6792 (N_6792,N_3389,N_3800);
nand U6793 (N_6793,N_3778,N_4578);
nor U6794 (N_6794,N_4045,N_5721);
or U6795 (N_6795,N_4810,N_3152);
or U6796 (N_6796,N_4400,N_3264);
and U6797 (N_6797,N_5398,N_3447);
xnor U6798 (N_6798,N_3713,N_4238);
nand U6799 (N_6799,N_4090,N_4750);
and U6800 (N_6800,N_5820,N_5988);
and U6801 (N_6801,N_5317,N_5536);
nand U6802 (N_6802,N_3141,N_4554);
or U6803 (N_6803,N_3541,N_3878);
or U6804 (N_6804,N_5057,N_5016);
nor U6805 (N_6805,N_5587,N_5069);
nand U6806 (N_6806,N_3902,N_5184);
nor U6807 (N_6807,N_4081,N_4879);
and U6808 (N_6808,N_3596,N_3563);
nor U6809 (N_6809,N_3518,N_4581);
nand U6810 (N_6810,N_5777,N_4995);
or U6811 (N_6811,N_5873,N_3636);
or U6812 (N_6812,N_5944,N_5511);
nor U6813 (N_6813,N_5551,N_4660);
or U6814 (N_6814,N_3382,N_5339);
or U6815 (N_6815,N_3707,N_5679);
xnor U6816 (N_6816,N_3973,N_4593);
and U6817 (N_6817,N_3100,N_5369);
and U6818 (N_6818,N_4680,N_5564);
or U6819 (N_6819,N_4725,N_3227);
nor U6820 (N_6820,N_5569,N_4326);
nand U6821 (N_6821,N_3281,N_3117);
or U6822 (N_6822,N_3929,N_5031);
nor U6823 (N_6823,N_5160,N_4395);
nor U6824 (N_6824,N_3971,N_5388);
and U6825 (N_6825,N_4940,N_3682);
or U6826 (N_6826,N_4703,N_4295);
nor U6827 (N_6827,N_3047,N_5771);
nand U6828 (N_6828,N_3060,N_3531);
xnor U6829 (N_6829,N_3335,N_3466);
and U6830 (N_6830,N_5088,N_4842);
nor U6831 (N_6831,N_5378,N_3664);
xor U6832 (N_6832,N_4972,N_3195);
and U6833 (N_6833,N_3463,N_5026);
nor U6834 (N_6834,N_3077,N_4988);
nor U6835 (N_6835,N_3584,N_3426);
nor U6836 (N_6836,N_5733,N_5843);
and U6837 (N_6837,N_4509,N_5526);
and U6838 (N_6838,N_3387,N_3667);
nor U6839 (N_6839,N_4825,N_5252);
nor U6840 (N_6840,N_4590,N_4957);
nor U6841 (N_6841,N_3722,N_5404);
nor U6842 (N_6842,N_5292,N_5305);
or U6843 (N_6843,N_4362,N_3638);
nand U6844 (N_6844,N_4365,N_4315);
or U6845 (N_6845,N_4491,N_5652);
or U6846 (N_6846,N_3090,N_5848);
nor U6847 (N_6847,N_4942,N_4645);
nand U6848 (N_6848,N_3839,N_3963);
nor U6849 (N_6849,N_3786,N_4599);
and U6850 (N_6850,N_3238,N_3865);
and U6851 (N_6851,N_4851,N_3985);
and U6852 (N_6852,N_4279,N_4225);
or U6853 (N_6853,N_4164,N_4755);
nor U6854 (N_6854,N_3128,N_3601);
and U6855 (N_6855,N_3600,N_3437);
nand U6856 (N_6856,N_5152,N_4313);
or U6857 (N_6857,N_3505,N_4191);
or U6858 (N_6858,N_5472,N_4004);
nor U6859 (N_6859,N_3820,N_4721);
and U6860 (N_6860,N_3103,N_5431);
or U6861 (N_6861,N_4764,N_5385);
or U6862 (N_6862,N_4542,N_3987);
nor U6863 (N_6863,N_3186,N_4895);
and U6864 (N_6864,N_3358,N_5762);
nand U6865 (N_6865,N_5483,N_4031);
and U6866 (N_6866,N_5834,N_5647);
nor U6867 (N_6867,N_4135,N_4474);
nor U6868 (N_6868,N_5302,N_3049);
nand U6869 (N_6869,N_4816,N_3261);
nand U6870 (N_6870,N_3900,N_4370);
xnor U6871 (N_6871,N_4981,N_4443);
or U6872 (N_6872,N_4174,N_4916);
or U6873 (N_6873,N_5850,N_3691);
nand U6874 (N_6874,N_5025,N_5633);
and U6875 (N_6875,N_3444,N_4293);
nand U6876 (N_6876,N_5786,N_4121);
and U6877 (N_6877,N_4744,N_5360);
and U6878 (N_6878,N_3610,N_3996);
or U6879 (N_6879,N_5860,N_3376);
or U6880 (N_6880,N_3179,N_3178);
nor U6881 (N_6881,N_4624,N_3950);
or U6882 (N_6882,N_4798,N_4899);
and U6883 (N_6883,N_4795,N_4665);
nand U6884 (N_6884,N_4921,N_3680);
nand U6885 (N_6885,N_4682,N_5489);
xor U6886 (N_6886,N_5212,N_4122);
nor U6887 (N_6887,N_3645,N_5448);
nor U6888 (N_6888,N_4803,N_5955);
and U6889 (N_6889,N_5728,N_4498);
and U6890 (N_6890,N_4520,N_3305);
and U6891 (N_6891,N_5678,N_4523);
and U6892 (N_6892,N_3953,N_4574);
nand U6893 (N_6893,N_5219,N_5713);
and U6894 (N_6894,N_5091,N_4876);
or U6895 (N_6895,N_5271,N_5815);
nor U6896 (N_6896,N_3501,N_4024);
nand U6897 (N_6897,N_5120,N_3105);
or U6898 (N_6898,N_4451,N_3414);
or U6899 (N_6899,N_3759,N_4052);
nor U6900 (N_6900,N_3556,N_4684);
nor U6901 (N_6901,N_3908,N_3477);
nand U6902 (N_6902,N_3008,N_4896);
or U6903 (N_6903,N_4391,N_5354);
or U6904 (N_6904,N_4286,N_3114);
and U6905 (N_6905,N_5521,N_5597);
nand U6906 (N_6906,N_5965,N_4653);
nor U6907 (N_6907,N_3833,N_4836);
nor U6908 (N_6908,N_5798,N_4386);
nor U6909 (N_6909,N_3697,N_4339);
nand U6910 (N_6910,N_3785,N_5891);
nand U6911 (N_6911,N_4814,N_4922);
or U6912 (N_6912,N_5668,N_3685);
nor U6913 (N_6913,N_3410,N_3009);
nor U6914 (N_6914,N_5899,N_3366);
nand U6915 (N_6915,N_4573,N_5094);
or U6916 (N_6916,N_3157,N_5857);
nor U6917 (N_6917,N_4069,N_4588);
or U6918 (N_6918,N_4357,N_5290);
nor U6919 (N_6919,N_3744,N_4099);
nor U6920 (N_6920,N_4606,N_4945);
or U6921 (N_6921,N_4314,N_4156);
or U6922 (N_6922,N_5222,N_5202);
or U6923 (N_6923,N_5774,N_4996);
or U6924 (N_6924,N_5213,N_3613);
and U6925 (N_6925,N_5335,N_5937);
or U6926 (N_6926,N_5284,N_3472);
nand U6927 (N_6927,N_5926,N_3824);
nor U6928 (N_6928,N_5197,N_5366);
nand U6929 (N_6929,N_3578,N_4354);
nor U6930 (N_6930,N_5400,N_4777);
nand U6931 (N_6931,N_4449,N_3198);
and U6932 (N_6932,N_4469,N_3958);
and U6933 (N_6933,N_5810,N_5837);
nor U6934 (N_6934,N_3217,N_5981);
nor U6935 (N_6935,N_5529,N_4170);
or U6936 (N_6936,N_4062,N_3257);
and U6937 (N_6937,N_5931,N_5038);
nor U6938 (N_6938,N_5072,N_4159);
or U6939 (N_6939,N_4103,N_4817);
nand U6940 (N_6940,N_3302,N_3224);
or U6941 (N_6941,N_3464,N_4244);
or U6942 (N_6942,N_5208,N_3247);
or U6943 (N_6943,N_4805,N_4638);
and U6944 (N_6944,N_5986,N_4857);
and U6945 (N_6945,N_5912,N_4134);
or U6946 (N_6946,N_3855,N_5437);
nor U6947 (N_6947,N_4098,N_3481);
and U6948 (N_6948,N_4566,N_4990);
nor U6949 (N_6949,N_4026,N_5313);
xor U6950 (N_6950,N_4783,N_3967);
or U6951 (N_6951,N_3787,N_3102);
nor U6952 (N_6952,N_4623,N_5138);
nor U6953 (N_6953,N_4079,N_4278);
xnor U6954 (N_6954,N_3073,N_4128);
nor U6955 (N_6955,N_4788,N_5454);
nor U6956 (N_6956,N_5830,N_3934);
nand U6957 (N_6957,N_5528,N_4430);
nand U6958 (N_6958,N_4334,N_5859);
nand U6959 (N_6959,N_4727,N_3626);
nand U6960 (N_6960,N_3001,N_5445);
and U6961 (N_6961,N_3585,N_3265);
xnor U6962 (N_6962,N_4907,N_3023);
nand U6963 (N_6963,N_4951,N_3978);
nand U6964 (N_6964,N_4023,N_5818);
nor U6965 (N_6965,N_5198,N_5481);
nand U6966 (N_6966,N_5943,N_4222);
and U6967 (N_6967,N_3072,N_4383);
nor U6968 (N_6968,N_4526,N_3456);
and U6969 (N_6969,N_5628,N_5151);
or U6970 (N_6970,N_4233,N_5485);
and U6971 (N_6971,N_3018,N_5238);
or U6972 (N_6972,N_3811,N_4336);
and U6973 (N_6973,N_5050,N_3945);
nor U6974 (N_6974,N_5145,N_5578);
nor U6975 (N_6975,N_5090,N_4650);
or U6976 (N_6976,N_5028,N_5166);
and U6977 (N_6977,N_4824,N_5329);
nor U6978 (N_6978,N_4030,N_4953);
and U6979 (N_6979,N_5543,N_4129);
nand U6980 (N_6980,N_3177,N_5594);
or U6981 (N_6981,N_5877,N_5225);
nor U6982 (N_6982,N_5314,N_3132);
or U6983 (N_6983,N_3808,N_3428);
nand U6984 (N_6984,N_3913,N_5813);
nor U6985 (N_6985,N_3678,N_5886);
and U6986 (N_6986,N_4517,N_3091);
nand U6987 (N_6987,N_4360,N_3884);
xnor U6988 (N_6988,N_3625,N_4671);
nand U6989 (N_6989,N_3432,N_3676);
nand U6990 (N_6990,N_5402,N_4227);
nor U6991 (N_6991,N_5189,N_3333);
and U6992 (N_6992,N_5579,N_3760);
and U6993 (N_6993,N_4489,N_3949);
and U6994 (N_6994,N_5459,N_3648);
nor U6995 (N_6995,N_5729,N_4548);
nor U6996 (N_6996,N_3199,N_4161);
nor U6997 (N_6997,N_3226,N_3732);
nand U6998 (N_6998,N_5055,N_4312);
and U6999 (N_6999,N_5420,N_4468);
nor U7000 (N_7000,N_3869,N_3061);
and U7001 (N_7001,N_4696,N_3304);
or U7002 (N_7002,N_3930,N_4793);
nor U7003 (N_7003,N_5919,N_4414);
nand U7004 (N_7004,N_5911,N_5395);
nand U7005 (N_7005,N_3310,N_5588);
and U7006 (N_7006,N_4142,N_5922);
and U7007 (N_7007,N_5627,N_5013);
nor U7008 (N_7008,N_3043,N_3794);
nor U7009 (N_7009,N_5743,N_3021);
or U7010 (N_7010,N_3228,N_4392);
nand U7011 (N_7011,N_3230,N_4832);
or U7012 (N_7012,N_4522,N_5855);
and U7013 (N_7013,N_3754,N_5427);
or U7014 (N_7014,N_4850,N_4488);
and U7015 (N_7015,N_4931,N_5042);
and U7016 (N_7016,N_3309,N_5136);
nand U7017 (N_7017,N_4017,N_4688);
and U7018 (N_7018,N_4202,N_3174);
nor U7019 (N_7019,N_4720,N_4422);
or U7020 (N_7020,N_5657,N_3816);
nand U7021 (N_7021,N_5827,N_3028);
or U7022 (N_7022,N_3692,N_4613);
and U7023 (N_7023,N_4234,N_3681);
or U7024 (N_7024,N_4168,N_5767);
or U7025 (N_7025,N_4175,N_3204);
nor U7026 (N_7026,N_4291,N_4066);
nand U7027 (N_7027,N_4218,N_3652);
nand U7028 (N_7028,N_4210,N_5832);
nor U7029 (N_7029,N_5414,N_4723);
or U7030 (N_7030,N_5592,N_4846);
nand U7031 (N_7031,N_3416,N_4617);
nor U7032 (N_7032,N_4970,N_3200);
and U7033 (N_7033,N_3608,N_3647);
nor U7034 (N_7034,N_4167,N_4668);
xor U7035 (N_7035,N_4283,N_3571);
and U7036 (N_7036,N_3299,N_3058);
nor U7037 (N_7037,N_4965,N_4545);
nor U7038 (N_7038,N_4547,N_3488);
nand U7039 (N_7039,N_4785,N_4393);
nand U7040 (N_7040,N_3206,N_3756);
nand U7041 (N_7041,N_3768,N_4534);
or U7042 (N_7042,N_4492,N_4656);
and U7043 (N_7043,N_5531,N_3259);
nand U7044 (N_7044,N_4258,N_3909);
nand U7045 (N_7045,N_5401,N_5201);
or U7046 (N_7046,N_5300,N_5187);
or U7047 (N_7047,N_4692,N_4663);
nor U7048 (N_7048,N_3418,N_4212);
and U7049 (N_7049,N_5646,N_5875);
xor U7050 (N_7050,N_5538,N_4250);
and U7051 (N_7051,N_4786,N_4911);
and U7052 (N_7052,N_4061,N_5236);
and U7053 (N_7053,N_3990,N_3623);
nor U7054 (N_7054,N_3080,N_5372);
nor U7055 (N_7055,N_3131,N_3954);
xor U7056 (N_7056,N_5632,N_4964);
or U7057 (N_7057,N_3207,N_3522);
or U7058 (N_7058,N_4875,N_5581);
or U7059 (N_7059,N_5123,N_3203);
nor U7060 (N_7060,N_4078,N_5534);
nor U7061 (N_7061,N_4290,N_3159);
or U7062 (N_7062,N_5341,N_4555);
xnor U7063 (N_7063,N_5808,N_4780);
nor U7064 (N_7064,N_3317,N_5147);
or U7065 (N_7065,N_5438,N_3965);
or U7066 (N_7066,N_5571,N_5705);
or U7067 (N_7067,N_4745,N_3156);
or U7068 (N_7068,N_4941,N_4840);
or U7069 (N_7069,N_5956,N_5562);
nand U7070 (N_7070,N_4626,N_3372);
or U7071 (N_7071,N_4636,N_4838);
or U7072 (N_7072,N_5014,N_3842);
nor U7073 (N_7073,N_3728,N_5010);
nand U7074 (N_7074,N_3492,N_4384);
nor U7075 (N_7075,N_5554,N_5132);
or U7076 (N_7076,N_5804,N_4413);
nand U7077 (N_7077,N_3628,N_3126);
xnor U7078 (N_7078,N_4378,N_4000);
nor U7079 (N_7079,N_5024,N_3417);
nand U7080 (N_7080,N_5036,N_4821);
nor U7081 (N_7081,N_3581,N_3233);
and U7082 (N_7082,N_5719,N_3125);
and U7083 (N_7083,N_4563,N_5045);
nor U7084 (N_7084,N_4550,N_5234);
and U7085 (N_7085,N_3182,N_4769);
and U7086 (N_7086,N_4035,N_5987);
or U7087 (N_7087,N_4453,N_5819);
nor U7088 (N_7088,N_4132,N_4235);
nand U7089 (N_7089,N_3919,N_3067);
nand U7090 (N_7090,N_3175,N_5585);
nor U7091 (N_7091,N_3107,N_4562);
nor U7092 (N_7092,N_5421,N_3070);
or U7093 (N_7093,N_4047,N_4072);
and U7094 (N_7094,N_4109,N_5524);
and U7095 (N_7095,N_3144,N_5574);
nand U7096 (N_7096,N_4820,N_3187);
and U7097 (N_7097,N_3025,N_3538);
nand U7098 (N_7098,N_4648,N_3348);
and U7099 (N_7099,N_5161,N_3969);
nand U7100 (N_7100,N_5250,N_4903);
or U7101 (N_7101,N_3071,N_5490);
and U7102 (N_7102,N_3225,N_3482);
or U7103 (N_7103,N_5936,N_3845);
nor U7104 (N_7104,N_5423,N_4987);
nand U7105 (N_7105,N_4632,N_5868);
nand U7106 (N_7106,N_4928,N_3136);
xor U7107 (N_7107,N_4943,N_3258);
nor U7108 (N_7108,N_5003,N_5666);
nor U7109 (N_7109,N_5544,N_5109);
and U7110 (N_7110,N_4350,N_3434);
and U7111 (N_7111,N_4882,N_4719);
and U7112 (N_7112,N_3761,N_4123);
nand U7113 (N_7113,N_4918,N_4716);
nor U7114 (N_7114,N_3614,N_3112);
or U7115 (N_7115,N_5856,N_5805);
and U7116 (N_7116,N_4871,N_4829);
nand U7117 (N_7117,N_5709,N_5301);
nand U7118 (N_7118,N_5828,N_4344);
nor U7119 (N_7119,N_4712,N_4844);
nand U7120 (N_7120,N_5766,N_4902);
nor U7121 (N_7121,N_4779,N_3160);
and U7122 (N_7122,N_5274,N_5520);
nand U7123 (N_7123,N_3373,N_3162);
and U7124 (N_7124,N_4592,N_5017);
or U7125 (N_7125,N_4652,N_5867);
and U7126 (N_7126,N_4960,N_4442);
or U7127 (N_7127,N_4049,N_3081);
xor U7128 (N_7128,N_4849,N_5181);
nor U7129 (N_7129,N_4529,N_4302);
nor U7130 (N_7130,N_4790,N_4273);
or U7131 (N_7131,N_4306,N_5319);
nand U7132 (N_7132,N_4276,N_3328);
nand U7133 (N_7133,N_5327,N_3314);
or U7134 (N_7134,N_4753,N_5020);
and U7135 (N_7135,N_4143,N_5957);
nand U7136 (N_7136,N_4325,N_3935);
nand U7137 (N_7137,N_3029,N_5000);
nand U7138 (N_7138,N_4991,N_5452);
or U7139 (N_7139,N_4924,N_5083);
and U7140 (N_7140,N_5635,N_5699);
and U7141 (N_7141,N_4888,N_5439);
nor U7142 (N_7142,N_3582,N_3751);
xnor U7143 (N_7143,N_5195,N_4658);
or U7144 (N_7144,N_3603,N_3425);
xor U7145 (N_7145,N_3345,N_5660);
nor U7146 (N_7146,N_4865,N_3193);
or U7147 (N_7147,N_3883,N_4130);
and U7148 (N_7148,N_4221,N_4932);
or U7149 (N_7149,N_3045,N_5463);
or U7150 (N_7150,N_4260,N_3303);
nor U7151 (N_7151,N_3976,N_4544);
or U7152 (N_7152,N_3044,N_5218);
nand U7153 (N_7153,N_5288,N_3850);
nand U7154 (N_7154,N_5776,N_4580);
and U7155 (N_7155,N_4423,N_5381);
xnor U7156 (N_7156,N_3607,N_4356);
and U7157 (N_7157,N_5265,N_4629);
and U7158 (N_7158,N_5934,N_5065);
nand U7159 (N_7159,N_3655,N_4569);
and U7160 (N_7160,N_4082,N_5640);
or U7161 (N_7161,N_3517,N_3294);
nand U7162 (N_7162,N_3641,N_4321);
and U7163 (N_7163,N_3849,N_3705);
or U7164 (N_7164,N_4211,N_5779);
or U7165 (N_7165,N_5809,N_5494);
or U7166 (N_7166,N_3274,N_5595);
nand U7167 (N_7167,N_3758,N_4409);
or U7168 (N_7168,N_3469,N_5349);
and U7169 (N_7169,N_5103,N_3779);
nor U7170 (N_7170,N_4165,N_5523);
or U7171 (N_7171,N_3431,N_4837);
and U7172 (N_7172,N_3394,N_5325);
and U7173 (N_7173,N_4511,N_5477);
and U7174 (N_7174,N_3771,N_5545);
or U7175 (N_7175,N_4390,N_4433);
nand U7176 (N_7176,N_5914,N_4102);
nor U7177 (N_7177,N_5496,N_5648);
nand U7178 (N_7178,N_5119,N_3519);
or U7179 (N_7179,N_4508,N_4029);
nand U7180 (N_7180,N_4056,N_3551);
or U7181 (N_7181,N_5078,N_5966);
or U7182 (N_7182,N_5373,N_3436);
or U7183 (N_7183,N_5963,N_5794);
nor U7184 (N_7184,N_3730,N_4157);
or U7185 (N_7185,N_4572,N_5479);
nor U7186 (N_7186,N_5269,N_5380);
and U7187 (N_7187,N_5669,N_4977);
and U7188 (N_7188,N_4925,N_4195);
or U7189 (N_7189,N_4146,N_4861);
or U7190 (N_7190,N_3619,N_5596);
nor U7191 (N_7191,N_5128,N_5503);
nor U7192 (N_7192,N_4787,N_4022);
nor U7193 (N_7193,N_5217,N_4070);
nor U7194 (N_7194,N_4823,N_5742);
and U7195 (N_7195,N_3863,N_5604);
or U7196 (N_7196,N_5686,N_3490);
nand U7197 (N_7197,N_3507,N_3916);
nor U7198 (N_7198,N_3558,N_3098);
or U7199 (N_7199,N_5852,N_3205);
nor U7200 (N_7200,N_3343,N_4162);
or U7201 (N_7201,N_3392,N_3745);
nand U7202 (N_7202,N_4714,N_3095);
and U7203 (N_7203,N_5532,N_5515);
nor U7204 (N_7204,N_3959,N_3003);
or U7205 (N_7205,N_5124,N_5086);
nor U7206 (N_7206,N_5210,N_5636);
nand U7207 (N_7207,N_3617,N_3962);
nand U7208 (N_7208,N_4914,N_4148);
nand U7209 (N_7209,N_3637,N_3503);
or U7210 (N_7210,N_3220,N_4138);
or U7211 (N_7211,N_3319,N_5540);
or U7212 (N_7212,N_5498,N_3671);
and U7213 (N_7213,N_5066,N_3534);
or U7214 (N_7214,N_4176,N_4506);
and U7215 (N_7215,N_3388,N_3493);
or U7216 (N_7216,N_3036,N_3185);
nand U7217 (N_7217,N_3502,N_4746);
nor U7218 (N_7218,N_3831,N_3752);
nand U7219 (N_7219,N_3861,N_3733);
nor U7220 (N_7220,N_5730,N_4594);
or U7221 (N_7221,N_4881,N_4271);
and U7222 (N_7222,N_4347,N_4983);
or U7223 (N_7223,N_3994,N_5382);
or U7224 (N_7224,N_3721,N_3500);
or U7225 (N_7225,N_5230,N_5182);
or U7226 (N_7226,N_5362,N_3229);
nand U7227 (N_7227,N_3415,N_4966);
nor U7228 (N_7228,N_4236,N_4571);
or U7229 (N_7229,N_5982,N_4647);
nor U7230 (N_7230,N_3796,N_5262);
nand U7231 (N_7231,N_4948,N_4087);
nor U7232 (N_7232,N_5258,N_3473);
nor U7233 (N_7233,N_3523,N_4528);
nor U7234 (N_7234,N_5942,N_4485);
or U7235 (N_7235,N_5478,N_3847);
and U7236 (N_7236,N_3171,N_3240);
nand U7237 (N_7237,N_5180,N_4470);
or U7238 (N_7238,N_5695,N_4484);
nor U7239 (N_7239,N_4005,N_3984);
nand U7240 (N_7240,N_5566,N_5787);
and U7241 (N_7241,N_4946,N_3836);
or U7242 (N_7242,N_3381,N_4331);
nor U7243 (N_7243,N_3325,N_4730);
and U7244 (N_7244,N_4539,N_4839);
nor U7245 (N_7245,N_5039,N_3180);
nand U7246 (N_7246,N_4605,N_5560);
or U7247 (N_7247,N_3032,N_5677);
nor U7248 (N_7248,N_5070,N_3616);
or U7249 (N_7249,N_5541,N_4448);
nand U7250 (N_7250,N_4402,N_3983);
nand U7251 (N_7251,N_4761,N_3627);
or U7252 (N_7252,N_5175,N_4220);
nand U7253 (N_7253,N_5356,N_4088);
nand U7254 (N_7254,N_3866,N_4145);
nand U7255 (N_7255,N_3063,N_5032);
nand U7256 (N_7256,N_3184,N_5434);
or U7257 (N_7257,N_4426,N_3710);
or U7258 (N_7258,N_4693,N_4450);
nand U7259 (N_7259,N_3812,N_4277);
nor U7260 (N_7260,N_3834,N_5864);
nand U7261 (N_7261,N_5190,N_5475);
and U7262 (N_7262,N_5469,N_4333);
or U7263 (N_7263,N_4742,N_3439);
nor U7264 (N_7264,N_4239,N_5425);
nor U7265 (N_7265,N_3231,N_4701);
nand U7266 (N_7266,N_5797,N_5449);
nor U7267 (N_7267,N_5021,N_5803);
and U7268 (N_7268,N_5484,N_5712);
nor U7269 (N_7269,N_4913,N_5836);
or U7270 (N_7270,N_4093,N_5247);
nand U7271 (N_7271,N_4514,N_5821);
nand U7272 (N_7272,N_4444,N_3116);
nand U7273 (N_7273,N_4532,N_5570);
nor U7274 (N_7274,N_4910,N_5309);
and U7275 (N_7275,N_4992,N_5041);
and U7276 (N_7276,N_5126,N_3944);
or U7277 (N_7277,N_3980,N_4602);
and U7278 (N_7278,N_5386,N_3243);
and U7279 (N_7279,N_3611,N_4901);
nor U7280 (N_7280,N_4934,N_5976);
nor U7281 (N_7281,N_5575,N_5576);
nand U7282 (N_7282,N_3630,N_3606);
nor U7283 (N_7283,N_4801,N_5935);
nor U7284 (N_7284,N_4900,N_3941);
nand U7285 (N_7285,N_4455,N_3914);
nand U7286 (N_7286,N_4472,N_3011);
and U7287 (N_7287,N_3406,N_5941);
or U7288 (N_7288,N_5377,N_4870);
nand U7289 (N_7289,N_4009,N_5474);
or U7290 (N_7290,N_3535,N_4398);
nor U7291 (N_7291,N_3268,N_3089);
or U7292 (N_7292,N_4530,N_3038);
nand U7293 (N_7293,N_5513,N_3106);
nand U7294 (N_7294,N_4797,N_4441);
nor U7295 (N_7295,N_4342,N_5178);
and U7296 (N_7296,N_3121,N_4150);
and U7297 (N_7297,N_3669,N_4986);
xor U7298 (N_7298,N_4763,N_5422);
and U7299 (N_7299,N_5052,N_4819);
or U7300 (N_7300,N_3763,N_3986);
or U7301 (N_7301,N_5383,N_5745);
xor U7302 (N_7302,N_5358,N_3838);
nand U7303 (N_7303,N_4091,N_3330);
and U7304 (N_7304,N_5173,N_3015);
and U7305 (N_7305,N_5975,N_3402);
nand U7306 (N_7306,N_3960,N_5972);
or U7307 (N_7307,N_4923,N_4153);
and U7308 (N_7308,N_5533,N_3624);
nand U7309 (N_7309,N_5112,N_5424);
or U7310 (N_7310,N_4465,N_3383);
and U7311 (N_7311,N_5735,N_5510);
nand U7312 (N_7312,N_4412,N_4445);
nand U7313 (N_7313,N_3688,N_5643);
or U7314 (N_7314,N_5468,N_3013);
and U7315 (N_7315,N_4898,N_5430);
nand U7316 (N_7316,N_4549,N_3390);
nor U7317 (N_7317,N_4702,N_3263);
nand U7318 (N_7318,N_3723,N_3735);
and U7319 (N_7319,N_5738,N_4533);
nand U7320 (N_7320,N_4683,N_5782);
xnor U7321 (N_7321,N_3006,N_4664);
nor U7322 (N_7322,N_5416,N_4661);
and U7323 (N_7323,N_5826,N_5154);
nand U7324 (N_7324,N_5244,N_5323);
nand U7325 (N_7325,N_4582,N_5176);
nor U7326 (N_7326,N_3826,N_5727);
xor U7327 (N_7327,N_3781,N_3879);
or U7328 (N_7328,N_5658,N_4086);
or U7329 (N_7329,N_3508,N_3421);
nand U7330 (N_7330,N_4366,N_4690);
nand U7331 (N_7331,N_5675,N_4598);
or U7332 (N_7332,N_4695,N_3438);
or U7333 (N_7333,N_4963,N_4475);
nand U7334 (N_7334,N_3740,N_4025);
nor U7335 (N_7335,N_3034,N_3113);
nand U7336 (N_7336,N_4560,N_3164);
and U7337 (N_7337,N_4364,N_4989);
and U7338 (N_7338,N_4076,N_3553);
nor U7339 (N_7339,N_4707,N_5397);
or U7340 (N_7340,N_3769,N_3790);
nor U7341 (N_7341,N_4859,N_4189);
nand U7342 (N_7342,N_3797,N_5539);
or U7343 (N_7343,N_3895,N_4751);
nor U7344 (N_7344,N_4224,N_3739);
nand U7345 (N_7345,N_3718,N_5044);
xor U7346 (N_7346,N_3391,N_3823);
or U7347 (N_7347,N_4399,N_5340);
nand U7348 (N_7348,N_4059,N_3030);
nor U7349 (N_7349,N_4266,N_3019);
or U7350 (N_7350,N_5255,N_4401);
nand U7351 (N_7351,N_3462,N_4713);
and U7352 (N_7352,N_3485,N_4698);
and U7353 (N_7353,N_3494,N_3588);
nand U7354 (N_7354,N_5799,N_5243);
nor U7355 (N_7355,N_5465,N_3110);
nand U7356 (N_7356,N_5717,N_4933);
nand U7357 (N_7357,N_5842,N_3423);
nand U7358 (N_7358,N_3027,N_4117);
nand U7359 (N_7359,N_4199,N_3092);
nand U7360 (N_7360,N_5417,N_3411);
nand U7361 (N_7361,N_3066,N_3395);
xnor U7362 (N_7362,N_4406,N_5071);
and U7363 (N_7363,N_5580,N_5665);
or U7364 (N_7364,N_3700,N_4013);
nand U7365 (N_7365,N_5795,N_3513);
and U7366 (N_7366,N_3059,N_4111);
and U7367 (N_7367,N_3007,N_3338);
nand U7368 (N_7368,N_3165,N_3819);
and U7369 (N_7369,N_5908,N_3560);
and U7370 (N_7370,N_5073,N_5714);
or U7371 (N_7371,N_4110,N_3746);
nand U7372 (N_7372,N_5099,N_4096);
nand U7373 (N_7373,N_4112,N_4284);
nor U7374 (N_7374,N_4301,N_5179);
nand U7375 (N_7375,N_3587,N_5801);
nor U7376 (N_7376,N_5947,N_3146);
or U7377 (N_7377,N_4516,N_5637);
nand U7378 (N_7378,N_3720,N_4504);
nand U7379 (N_7379,N_4892,N_4089);
and U7380 (N_7380,N_4950,N_5246);
nor U7381 (N_7381,N_5096,N_3096);
nor U7382 (N_7382,N_5722,N_4917);
or U7383 (N_7383,N_4115,N_4856);
or U7384 (N_7384,N_5885,N_3289);
or U7385 (N_7385,N_4077,N_5130);
nor U7386 (N_7386,N_5237,N_4126);
nor U7387 (N_7387,N_3854,N_5691);
nand U7388 (N_7388,N_5599,N_3196);
nand U7389 (N_7389,N_4890,N_3612);
or U7390 (N_7390,N_3572,N_3370);
or U7391 (N_7391,N_5974,N_4348);
xnor U7392 (N_7392,N_5251,N_3336);
nand U7393 (N_7393,N_5253,N_5015);
and U7394 (N_7394,N_3291,N_3316);
or U7395 (N_7395,N_3904,N_4245);
nand U7396 (N_7396,N_5906,N_3573);
and U7397 (N_7397,N_3076,N_3668);
nand U7398 (N_7398,N_3266,N_5240);
nor U7399 (N_7399,N_3742,N_5365);
nand U7400 (N_7400,N_3525,N_4459);
or U7401 (N_7401,N_5018,N_5811);
nand U7402 (N_7402,N_3993,N_5281);
and U7403 (N_7403,N_4310,N_4575);
nand U7404 (N_7404,N_3726,N_3111);
nand U7405 (N_7405,N_4018,N_5514);
nand U7406 (N_7406,N_4557,N_4416);
nand U7407 (N_7407,N_5412,N_3491);
nor U7408 (N_7408,N_4275,N_4579);
or U7409 (N_7409,N_3828,N_3774);
nor U7410 (N_7410,N_4771,N_4246);
and U7411 (N_7411,N_4543,N_5005);
and U7412 (N_7412,N_5334,N_4678);
nand U7413 (N_7413,N_5287,N_4500);
nor U7414 (N_7414,N_3830,N_4478);
and U7415 (N_7415,N_4809,N_3670);
or U7416 (N_7416,N_3440,N_3189);
or U7417 (N_7417,N_4141,N_3524);
or U7418 (N_7418,N_4396,N_4193);
nor U7419 (N_7419,N_5278,N_4551);
or U7420 (N_7420,N_3859,N_3843);
or U7421 (N_7421,N_4213,N_3575);
nand U7422 (N_7422,N_3450,N_5077);
nand U7423 (N_7423,N_5087,N_4471);
or U7424 (N_7424,N_4586,N_3791);
xor U7425 (N_7425,N_3435,N_3399);
or U7426 (N_7426,N_5645,N_5214);
or U7427 (N_7427,N_5482,N_5076);
or U7428 (N_7428,N_4559,N_5352);
nand U7429 (N_7429,N_5311,N_3082);
nand U7430 (N_7430,N_5488,N_3698);
and U7431 (N_7431,N_4710,N_3400);
nand U7432 (N_7432,N_5663,N_3870);
nor U7433 (N_7433,N_5296,N_5895);
or U7434 (N_7434,N_4231,N_3927);
nand U7435 (N_7435,N_4610,N_4826);
or U7436 (N_7436,N_5878,N_4075);
or U7437 (N_7437,N_3982,N_5450);
or U7438 (N_7438,N_4048,N_3139);
or U7439 (N_7439,N_5940,N_4502);
nor U7440 (N_7440,N_4042,N_3891);
nor U7441 (N_7441,N_4997,N_3835);
or U7442 (N_7442,N_4796,N_4615);
xnor U7443 (N_7443,N_4131,N_3932);
nor U7444 (N_7444,N_3799,N_5150);
nor U7445 (N_7445,N_3486,N_4281);
and U7446 (N_7446,N_3793,N_3054);
nand U7447 (N_7447,N_3672,N_5268);
or U7448 (N_7448,N_4477,N_3384);
nor U7449 (N_7449,N_3340,N_5858);
nand U7450 (N_7450,N_4264,N_4499);
nor U7451 (N_7451,N_3887,N_5741);
and U7452 (N_7452,N_4379,N_4355);
and U7453 (N_7453,N_4962,N_4015);
or U7454 (N_7454,N_3427,N_5653);
or U7455 (N_7455,N_4501,N_3832);
nor U7456 (N_7456,N_5638,N_3813);
nor U7457 (N_7457,N_5486,N_5299);
nand U7458 (N_7458,N_4625,N_4481);
nand U7459 (N_7459,N_4718,N_5655);
or U7460 (N_7460,N_4635,N_5553);
nor U7461 (N_7461,N_3948,N_4243);
nand U7462 (N_7462,N_4681,N_5829);
or U7463 (N_7463,N_5584,N_4515);
or U7464 (N_7464,N_3766,N_3741);
nand U7465 (N_7465,N_3620,N_5241);
xor U7466 (N_7466,N_3817,N_3696);
nand U7467 (N_7467,N_5708,N_3725);
and U7468 (N_7468,N_5879,N_4137);
or U7469 (N_7469,N_3176,N_3892);
nand U7470 (N_7470,N_5232,N_5884);
nand U7471 (N_7471,N_4706,N_4510);
nor U7472 (N_7472,N_4216,N_3361);
and U7473 (N_7473,N_4685,N_4994);
xnor U7474 (N_7474,N_3262,N_5473);
nor U7475 (N_7475,N_5610,N_5806);
nand U7476 (N_7476,N_5565,N_4241);
and U7477 (N_7477,N_4726,N_3235);
and U7478 (N_7478,N_3767,N_4694);
and U7479 (N_7479,N_3656,N_3997);
or U7480 (N_7480,N_5033,N_5347);
nand U7481 (N_7481,N_5568,N_3592);
and U7482 (N_7482,N_4483,N_3593);
or U7483 (N_7483,N_4705,N_3822);
nor U7484 (N_7484,N_5724,N_3219);
nand U7485 (N_7485,N_4057,N_3737);
nor U7486 (N_7486,N_3995,N_5261);
nor U7487 (N_7487,N_3776,N_4358);
nand U7488 (N_7488,N_4540,N_4704);
nand U7489 (N_7489,N_3598,N_4739);
and U7490 (N_7490,N_5530,N_3992);
xor U7491 (N_7491,N_3298,N_5948);
or U7492 (N_7492,N_3708,N_4133);
nor U7493 (N_7493,N_4675,N_5006);
nand U7494 (N_7494,N_5113,N_3683);
nor U7495 (N_7495,N_3715,N_3642);
nand U7496 (N_7496,N_4674,N_5046);
or U7497 (N_7497,N_4524,N_4166);
xor U7498 (N_7498,N_4929,N_4341);
and U7499 (N_7499,N_3278,N_3712);
nand U7500 (N_7500,N_3554,N_3814);
or U7501 (N_7501,N_4764,N_5754);
nand U7502 (N_7502,N_5169,N_3177);
nor U7503 (N_7503,N_4834,N_4662);
and U7504 (N_7504,N_5183,N_4619);
or U7505 (N_7505,N_3660,N_5089);
nor U7506 (N_7506,N_4771,N_3537);
or U7507 (N_7507,N_4030,N_5244);
and U7508 (N_7508,N_3591,N_5681);
and U7509 (N_7509,N_3657,N_5687);
nand U7510 (N_7510,N_4200,N_3184);
or U7511 (N_7511,N_3258,N_3822);
nand U7512 (N_7512,N_5236,N_3319);
and U7513 (N_7513,N_3462,N_3162);
or U7514 (N_7514,N_5264,N_4956);
and U7515 (N_7515,N_4223,N_4016);
nand U7516 (N_7516,N_5556,N_4486);
or U7517 (N_7517,N_3878,N_5709);
nor U7518 (N_7518,N_4629,N_3819);
and U7519 (N_7519,N_4743,N_4237);
nand U7520 (N_7520,N_3442,N_3857);
xnor U7521 (N_7521,N_3496,N_4006);
or U7522 (N_7522,N_3091,N_4469);
and U7523 (N_7523,N_5655,N_3161);
and U7524 (N_7524,N_5650,N_4505);
or U7525 (N_7525,N_3728,N_3138);
nor U7526 (N_7526,N_4398,N_4617);
nand U7527 (N_7527,N_3970,N_3584);
or U7528 (N_7528,N_4667,N_5573);
or U7529 (N_7529,N_4860,N_3255);
nand U7530 (N_7530,N_4697,N_5410);
or U7531 (N_7531,N_4512,N_5468);
nor U7532 (N_7532,N_3908,N_4612);
nand U7533 (N_7533,N_3376,N_5594);
nor U7534 (N_7534,N_5420,N_4495);
or U7535 (N_7535,N_4854,N_5119);
or U7536 (N_7536,N_5434,N_3947);
or U7537 (N_7537,N_4402,N_3252);
nor U7538 (N_7538,N_4128,N_5324);
and U7539 (N_7539,N_3672,N_5440);
nor U7540 (N_7540,N_3397,N_5846);
nor U7541 (N_7541,N_4361,N_3044);
and U7542 (N_7542,N_3908,N_4161);
or U7543 (N_7543,N_4224,N_3360);
nor U7544 (N_7544,N_5496,N_5893);
and U7545 (N_7545,N_4110,N_3554);
nand U7546 (N_7546,N_3675,N_3552);
and U7547 (N_7547,N_5894,N_3278);
nor U7548 (N_7548,N_3844,N_3420);
and U7549 (N_7549,N_3967,N_4985);
or U7550 (N_7550,N_4653,N_3561);
or U7551 (N_7551,N_4065,N_3345);
nand U7552 (N_7552,N_5603,N_5557);
nor U7553 (N_7553,N_3605,N_4018);
and U7554 (N_7554,N_3025,N_4347);
or U7555 (N_7555,N_4470,N_3616);
or U7556 (N_7556,N_5162,N_5550);
and U7557 (N_7557,N_4318,N_5208);
nand U7558 (N_7558,N_3061,N_4263);
and U7559 (N_7559,N_5945,N_4911);
nand U7560 (N_7560,N_5581,N_3429);
nor U7561 (N_7561,N_5556,N_5642);
or U7562 (N_7562,N_4520,N_3292);
nand U7563 (N_7563,N_3603,N_4039);
nand U7564 (N_7564,N_3148,N_4301);
and U7565 (N_7565,N_3274,N_3207);
nor U7566 (N_7566,N_5208,N_3137);
nand U7567 (N_7567,N_4964,N_4199);
and U7568 (N_7568,N_3943,N_5605);
nand U7569 (N_7569,N_5507,N_3876);
or U7570 (N_7570,N_5400,N_3876);
xor U7571 (N_7571,N_3908,N_5889);
or U7572 (N_7572,N_4527,N_5301);
nor U7573 (N_7573,N_3371,N_5677);
nor U7574 (N_7574,N_3430,N_5943);
nand U7575 (N_7575,N_5397,N_4385);
or U7576 (N_7576,N_4279,N_4280);
nor U7577 (N_7577,N_3801,N_5337);
nand U7578 (N_7578,N_4839,N_4158);
or U7579 (N_7579,N_4546,N_4485);
nor U7580 (N_7580,N_4313,N_4725);
or U7581 (N_7581,N_3615,N_5946);
nand U7582 (N_7582,N_3011,N_3501);
nand U7583 (N_7583,N_4097,N_5278);
nand U7584 (N_7584,N_4988,N_3975);
or U7585 (N_7585,N_5492,N_5197);
nand U7586 (N_7586,N_5936,N_5634);
or U7587 (N_7587,N_3474,N_4828);
or U7588 (N_7588,N_3852,N_3252);
or U7589 (N_7589,N_3055,N_5063);
nor U7590 (N_7590,N_3468,N_5745);
nor U7591 (N_7591,N_5436,N_3173);
or U7592 (N_7592,N_5000,N_3207);
nand U7593 (N_7593,N_5247,N_4696);
and U7594 (N_7594,N_4162,N_4364);
nor U7595 (N_7595,N_5345,N_4451);
or U7596 (N_7596,N_4416,N_3612);
nor U7597 (N_7597,N_5186,N_4194);
and U7598 (N_7598,N_3930,N_4067);
and U7599 (N_7599,N_5639,N_4198);
and U7600 (N_7600,N_4995,N_3006);
nor U7601 (N_7601,N_5498,N_4253);
nand U7602 (N_7602,N_4932,N_4446);
nor U7603 (N_7603,N_5528,N_5076);
or U7604 (N_7604,N_4810,N_4427);
nand U7605 (N_7605,N_4836,N_4594);
or U7606 (N_7606,N_5397,N_4998);
or U7607 (N_7607,N_4030,N_5020);
and U7608 (N_7608,N_4499,N_4319);
nor U7609 (N_7609,N_5678,N_3010);
nor U7610 (N_7610,N_4345,N_4950);
nor U7611 (N_7611,N_4069,N_4419);
and U7612 (N_7612,N_4719,N_4040);
nand U7613 (N_7613,N_5885,N_4001);
and U7614 (N_7614,N_4614,N_5295);
or U7615 (N_7615,N_4899,N_3856);
nand U7616 (N_7616,N_4675,N_5552);
nor U7617 (N_7617,N_5997,N_3454);
or U7618 (N_7618,N_4960,N_4213);
nand U7619 (N_7619,N_4733,N_3686);
or U7620 (N_7620,N_3063,N_3388);
nand U7621 (N_7621,N_3653,N_5061);
and U7622 (N_7622,N_5433,N_3335);
nor U7623 (N_7623,N_4188,N_3615);
and U7624 (N_7624,N_5399,N_4753);
nor U7625 (N_7625,N_5712,N_4165);
xor U7626 (N_7626,N_3629,N_5823);
and U7627 (N_7627,N_5076,N_5721);
nand U7628 (N_7628,N_5783,N_4031);
nor U7629 (N_7629,N_3589,N_3808);
xor U7630 (N_7630,N_5930,N_5030);
or U7631 (N_7631,N_4472,N_3819);
or U7632 (N_7632,N_5595,N_4864);
nand U7633 (N_7633,N_4579,N_5244);
and U7634 (N_7634,N_5012,N_3956);
nor U7635 (N_7635,N_5098,N_5226);
or U7636 (N_7636,N_3219,N_4887);
nand U7637 (N_7637,N_3174,N_3711);
or U7638 (N_7638,N_4334,N_5705);
and U7639 (N_7639,N_5335,N_5212);
or U7640 (N_7640,N_5796,N_5068);
or U7641 (N_7641,N_5275,N_4123);
nor U7642 (N_7642,N_3904,N_5522);
nand U7643 (N_7643,N_4934,N_4492);
or U7644 (N_7644,N_5495,N_4796);
and U7645 (N_7645,N_5798,N_5068);
nor U7646 (N_7646,N_4068,N_4676);
nor U7647 (N_7647,N_3169,N_4120);
or U7648 (N_7648,N_4187,N_3913);
nand U7649 (N_7649,N_5682,N_5813);
nand U7650 (N_7650,N_3478,N_3714);
or U7651 (N_7651,N_3336,N_5978);
nand U7652 (N_7652,N_5047,N_3268);
or U7653 (N_7653,N_3300,N_3618);
and U7654 (N_7654,N_4939,N_3222);
nand U7655 (N_7655,N_4875,N_4148);
or U7656 (N_7656,N_3998,N_3588);
nor U7657 (N_7657,N_5431,N_4287);
or U7658 (N_7658,N_3370,N_3471);
nand U7659 (N_7659,N_5173,N_5232);
nor U7660 (N_7660,N_5028,N_4288);
nor U7661 (N_7661,N_5253,N_4574);
xnor U7662 (N_7662,N_5846,N_4752);
and U7663 (N_7663,N_5798,N_4987);
or U7664 (N_7664,N_4765,N_5542);
or U7665 (N_7665,N_3537,N_3769);
nor U7666 (N_7666,N_3204,N_5007);
nand U7667 (N_7667,N_4496,N_5456);
or U7668 (N_7668,N_4604,N_4442);
and U7669 (N_7669,N_4796,N_3519);
and U7670 (N_7670,N_4396,N_5667);
xnor U7671 (N_7671,N_5942,N_3763);
or U7672 (N_7672,N_5318,N_4835);
and U7673 (N_7673,N_3290,N_3378);
or U7674 (N_7674,N_5431,N_5708);
nand U7675 (N_7675,N_3197,N_4350);
and U7676 (N_7676,N_4752,N_3691);
or U7677 (N_7677,N_4337,N_3019);
nor U7678 (N_7678,N_4190,N_4435);
nor U7679 (N_7679,N_5319,N_4808);
nand U7680 (N_7680,N_3452,N_4369);
or U7681 (N_7681,N_4402,N_4793);
and U7682 (N_7682,N_5918,N_4273);
nor U7683 (N_7683,N_5742,N_5954);
or U7684 (N_7684,N_3744,N_5762);
or U7685 (N_7685,N_3089,N_4807);
xor U7686 (N_7686,N_4520,N_5092);
nand U7687 (N_7687,N_5011,N_4313);
nor U7688 (N_7688,N_4042,N_3499);
or U7689 (N_7689,N_4478,N_3566);
xnor U7690 (N_7690,N_4365,N_4815);
or U7691 (N_7691,N_5065,N_3881);
nand U7692 (N_7692,N_5793,N_3868);
and U7693 (N_7693,N_4028,N_5633);
and U7694 (N_7694,N_4482,N_5157);
and U7695 (N_7695,N_4624,N_5919);
nand U7696 (N_7696,N_5128,N_5556);
and U7697 (N_7697,N_5333,N_4680);
and U7698 (N_7698,N_5096,N_5904);
and U7699 (N_7699,N_3332,N_5257);
xor U7700 (N_7700,N_5881,N_3021);
or U7701 (N_7701,N_5837,N_5891);
nor U7702 (N_7702,N_4688,N_5531);
nor U7703 (N_7703,N_3675,N_4356);
xor U7704 (N_7704,N_5092,N_5131);
xor U7705 (N_7705,N_4752,N_3612);
nand U7706 (N_7706,N_5276,N_4874);
and U7707 (N_7707,N_5547,N_4932);
nor U7708 (N_7708,N_3323,N_5964);
nor U7709 (N_7709,N_4235,N_5818);
and U7710 (N_7710,N_5221,N_5826);
and U7711 (N_7711,N_5806,N_3571);
nand U7712 (N_7712,N_4212,N_3664);
nand U7713 (N_7713,N_3330,N_4497);
nor U7714 (N_7714,N_3214,N_3350);
nor U7715 (N_7715,N_3221,N_3040);
and U7716 (N_7716,N_4191,N_5286);
or U7717 (N_7717,N_5354,N_3922);
and U7718 (N_7718,N_4909,N_4440);
nand U7719 (N_7719,N_5722,N_5291);
and U7720 (N_7720,N_4711,N_4352);
nand U7721 (N_7721,N_3830,N_5811);
nand U7722 (N_7722,N_3809,N_4456);
nand U7723 (N_7723,N_3837,N_3074);
and U7724 (N_7724,N_4057,N_4480);
nand U7725 (N_7725,N_3453,N_3469);
and U7726 (N_7726,N_3085,N_4927);
nand U7727 (N_7727,N_3056,N_4537);
and U7728 (N_7728,N_4607,N_5590);
and U7729 (N_7729,N_5116,N_4668);
nor U7730 (N_7730,N_5365,N_4630);
nand U7731 (N_7731,N_3966,N_5745);
and U7732 (N_7732,N_4513,N_5392);
nor U7733 (N_7733,N_4490,N_4358);
nor U7734 (N_7734,N_3898,N_5563);
nand U7735 (N_7735,N_5440,N_5201);
nor U7736 (N_7736,N_4371,N_4657);
and U7737 (N_7737,N_3166,N_4137);
and U7738 (N_7738,N_5828,N_5338);
nand U7739 (N_7739,N_4198,N_5289);
and U7740 (N_7740,N_4454,N_5628);
xor U7741 (N_7741,N_3958,N_3095);
nor U7742 (N_7742,N_5641,N_5291);
or U7743 (N_7743,N_5340,N_5133);
nand U7744 (N_7744,N_4410,N_4203);
and U7745 (N_7745,N_5579,N_4108);
nand U7746 (N_7746,N_3803,N_4314);
nor U7747 (N_7747,N_5501,N_5517);
nand U7748 (N_7748,N_3259,N_4854);
and U7749 (N_7749,N_3429,N_3053);
nor U7750 (N_7750,N_5959,N_3556);
nand U7751 (N_7751,N_4374,N_4349);
nand U7752 (N_7752,N_3920,N_3610);
or U7753 (N_7753,N_3877,N_4574);
and U7754 (N_7754,N_3090,N_4494);
or U7755 (N_7755,N_5814,N_5377);
nor U7756 (N_7756,N_4524,N_5093);
nand U7757 (N_7757,N_4373,N_5608);
nor U7758 (N_7758,N_3401,N_5927);
nor U7759 (N_7759,N_5077,N_3759);
nor U7760 (N_7760,N_5780,N_3566);
nor U7761 (N_7761,N_4294,N_4499);
or U7762 (N_7762,N_5404,N_3282);
and U7763 (N_7763,N_5480,N_3690);
xnor U7764 (N_7764,N_5004,N_5311);
nand U7765 (N_7765,N_4088,N_4042);
nand U7766 (N_7766,N_3792,N_5400);
or U7767 (N_7767,N_5400,N_3715);
and U7768 (N_7768,N_4742,N_3344);
or U7769 (N_7769,N_4348,N_4347);
nor U7770 (N_7770,N_3303,N_5068);
and U7771 (N_7771,N_3781,N_5125);
or U7772 (N_7772,N_3557,N_3194);
xnor U7773 (N_7773,N_4188,N_3460);
nor U7774 (N_7774,N_3286,N_3815);
and U7775 (N_7775,N_3014,N_3280);
nor U7776 (N_7776,N_5841,N_5894);
nor U7777 (N_7777,N_4655,N_3479);
and U7778 (N_7778,N_5846,N_3886);
and U7779 (N_7779,N_5809,N_3425);
nand U7780 (N_7780,N_5356,N_4822);
and U7781 (N_7781,N_5712,N_4606);
nor U7782 (N_7782,N_3017,N_5652);
and U7783 (N_7783,N_4910,N_4198);
nor U7784 (N_7784,N_5939,N_4999);
and U7785 (N_7785,N_3827,N_4798);
nor U7786 (N_7786,N_5660,N_3868);
nor U7787 (N_7787,N_5295,N_4542);
nor U7788 (N_7788,N_5460,N_3630);
nand U7789 (N_7789,N_5035,N_3552);
and U7790 (N_7790,N_5873,N_5033);
nor U7791 (N_7791,N_3161,N_3724);
nor U7792 (N_7792,N_3025,N_5129);
nand U7793 (N_7793,N_4683,N_4440);
nor U7794 (N_7794,N_4724,N_5247);
or U7795 (N_7795,N_4849,N_3492);
nand U7796 (N_7796,N_3625,N_5324);
and U7797 (N_7797,N_5690,N_4212);
and U7798 (N_7798,N_5388,N_5992);
or U7799 (N_7799,N_4691,N_4798);
nor U7800 (N_7800,N_5241,N_3310);
and U7801 (N_7801,N_3321,N_4385);
and U7802 (N_7802,N_4286,N_5719);
or U7803 (N_7803,N_3559,N_3014);
or U7804 (N_7804,N_4727,N_5078);
nor U7805 (N_7805,N_3222,N_5926);
nor U7806 (N_7806,N_3678,N_4397);
nor U7807 (N_7807,N_4890,N_5162);
nor U7808 (N_7808,N_4534,N_4569);
nor U7809 (N_7809,N_4801,N_5095);
and U7810 (N_7810,N_5527,N_3834);
and U7811 (N_7811,N_5593,N_4457);
nor U7812 (N_7812,N_5301,N_4772);
and U7813 (N_7813,N_3206,N_5256);
and U7814 (N_7814,N_5662,N_4085);
and U7815 (N_7815,N_5749,N_4920);
nand U7816 (N_7816,N_3714,N_3695);
nor U7817 (N_7817,N_3767,N_3572);
and U7818 (N_7818,N_4775,N_4125);
and U7819 (N_7819,N_5247,N_3663);
nand U7820 (N_7820,N_3723,N_3318);
nor U7821 (N_7821,N_4354,N_3696);
nand U7822 (N_7822,N_4312,N_3699);
nand U7823 (N_7823,N_3651,N_4481);
nor U7824 (N_7824,N_3588,N_5827);
nand U7825 (N_7825,N_3757,N_5100);
nor U7826 (N_7826,N_4472,N_4516);
nor U7827 (N_7827,N_3121,N_4678);
nand U7828 (N_7828,N_4660,N_5041);
nand U7829 (N_7829,N_5815,N_5504);
nand U7830 (N_7830,N_3444,N_5862);
nand U7831 (N_7831,N_5134,N_4082);
nand U7832 (N_7832,N_5124,N_3841);
and U7833 (N_7833,N_3229,N_3111);
xnor U7834 (N_7834,N_3844,N_4620);
or U7835 (N_7835,N_5035,N_3079);
and U7836 (N_7836,N_3514,N_4758);
nand U7837 (N_7837,N_3124,N_3426);
and U7838 (N_7838,N_5579,N_4615);
and U7839 (N_7839,N_5419,N_5391);
nand U7840 (N_7840,N_3056,N_3717);
and U7841 (N_7841,N_3326,N_5481);
nor U7842 (N_7842,N_5668,N_3286);
and U7843 (N_7843,N_5407,N_4456);
nand U7844 (N_7844,N_3584,N_3654);
nand U7845 (N_7845,N_4349,N_5874);
and U7846 (N_7846,N_3919,N_4503);
and U7847 (N_7847,N_5028,N_3094);
or U7848 (N_7848,N_5338,N_4990);
nor U7849 (N_7849,N_5094,N_3057);
nand U7850 (N_7850,N_5508,N_5310);
nand U7851 (N_7851,N_3846,N_3812);
nor U7852 (N_7852,N_3972,N_3985);
and U7853 (N_7853,N_5998,N_4779);
and U7854 (N_7854,N_5324,N_5308);
and U7855 (N_7855,N_5404,N_5047);
nand U7856 (N_7856,N_3083,N_4530);
and U7857 (N_7857,N_3269,N_4258);
nand U7858 (N_7858,N_4912,N_3600);
and U7859 (N_7859,N_5673,N_3694);
nor U7860 (N_7860,N_3218,N_5463);
nand U7861 (N_7861,N_5467,N_5968);
and U7862 (N_7862,N_4326,N_4307);
nor U7863 (N_7863,N_5100,N_5270);
nor U7864 (N_7864,N_3302,N_3609);
or U7865 (N_7865,N_4771,N_3055);
or U7866 (N_7866,N_4612,N_5554);
or U7867 (N_7867,N_4409,N_5144);
and U7868 (N_7868,N_4909,N_4450);
or U7869 (N_7869,N_5490,N_5947);
or U7870 (N_7870,N_3493,N_4196);
nand U7871 (N_7871,N_3257,N_4766);
and U7872 (N_7872,N_3545,N_5836);
or U7873 (N_7873,N_3138,N_3812);
nand U7874 (N_7874,N_5842,N_4571);
or U7875 (N_7875,N_5732,N_4121);
or U7876 (N_7876,N_5536,N_3856);
and U7877 (N_7877,N_5845,N_5403);
and U7878 (N_7878,N_5328,N_4554);
xor U7879 (N_7879,N_5974,N_3468);
nor U7880 (N_7880,N_5698,N_4498);
and U7881 (N_7881,N_5481,N_4391);
nand U7882 (N_7882,N_5033,N_5917);
and U7883 (N_7883,N_4661,N_3943);
or U7884 (N_7884,N_4044,N_3698);
or U7885 (N_7885,N_3371,N_4239);
nand U7886 (N_7886,N_4166,N_3424);
nor U7887 (N_7887,N_5675,N_3807);
or U7888 (N_7888,N_4117,N_5539);
nor U7889 (N_7889,N_4162,N_3062);
or U7890 (N_7890,N_5144,N_3082);
and U7891 (N_7891,N_5596,N_4906);
nor U7892 (N_7892,N_4044,N_3013);
nor U7893 (N_7893,N_3629,N_4012);
or U7894 (N_7894,N_5587,N_4117);
nor U7895 (N_7895,N_4234,N_3677);
nor U7896 (N_7896,N_4926,N_3838);
or U7897 (N_7897,N_3400,N_5103);
nand U7898 (N_7898,N_4116,N_5397);
or U7899 (N_7899,N_5069,N_5632);
or U7900 (N_7900,N_4954,N_3637);
nor U7901 (N_7901,N_5316,N_5043);
or U7902 (N_7902,N_5369,N_3644);
nand U7903 (N_7903,N_5126,N_4218);
nand U7904 (N_7904,N_4197,N_3865);
nor U7905 (N_7905,N_3446,N_4930);
nand U7906 (N_7906,N_3366,N_4738);
nand U7907 (N_7907,N_4103,N_5739);
and U7908 (N_7908,N_5543,N_5802);
or U7909 (N_7909,N_5914,N_3238);
nand U7910 (N_7910,N_4285,N_5428);
or U7911 (N_7911,N_3821,N_4416);
and U7912 (N_7912,N_3484,N_4156);
or U7913 (N_7913,N_3083,N_4219);
or U7914 (N_7914,N_5894,N_5995);
nand U7915 (N_7915,N_5541,N_3589);
nor U7916 (N_7916,N_5464,N_3372);
nand U7917 (N_7917,N_5319,N_3448);
nor U7918 (N_7918,N_4076,N_3708);
and U7919 (N_7919,N_4469,N_5346);
or U7920 (N_7920,N_3603,N_5581);
nand U7921 (N_7921,N_3293,N_3094);
nor U7922 (N_7922,N_3810,N_5221);
nand U7923 (N_7923,N_3763,N_3429);
nand U7924 (N_7924,N_3843,N_3839);
or U7925 (N_7925,N_3487,N_3872);
nand U7926 (N_7926,N_4519,N_5140);
or U7927 (N_7927,N_4011,N_4192);
and U7928 (N_7928,N_3458,N_4279);
nor U7929 (N_7929,N_4973,N_4317);
and U7930 (N_7930,N_5870,N_3815);
or U7931 (N_7931,N_5293,N_3900);
or U7932 (N_7932,N_3308,N_4615);
nor U7933 (N_7933,N_5319,N_5662);
nor U7934 (N_7934,N_5685,N_4287);
and U7935 (N_7935,N_3689,N_3299);
and U7936 (N_7936,N_5438,N_4566);
and U7937 (N_7937,N_5567,N_3048);
nand U7938 (N_7938,N_5538,N_4015);
and U7939 (N_7939,N_3077,N_5390);
nor U7940 (N_7940,N_4602,N_3617);
and U7941 (N_7941,N_4629,N_5228);
or U7942 (N_7942,N_5112,N_3475);
nand U7943 (N_7943,N_5442,N_3022);
and U7944 (N_7944,N_4315,N_4932);
nand U7945 (N_7945,N_5268,N_3061);
nor U7946 (N_7946,N_5530,N_4146);
nand U7947 (N_7947,N_4435,N_3634);
and U7948 (N_7948,N_5446,N_4951);
or U7949 (N_7949,N_4933,N_3800);
or U7950 (N_7950,N_3658,N_3773);
nor U7951 (N_7951,N_5290,N_4651);
nand U7952 (N_7952,N_4187,N_4847);
and U7953 (N_7953,N_5309,N_4378);
nor U7954 (N_7954,N_5634,N_3931);
and U7955 (N_7955,N_3808,N_5035);
nand U7956 (N_7956,N_3110,N_4258);
and U7957 (N_7957,N_5733,N_4297);
or U7958 (N_7958,N_3132,N_5759);
nor U7959 (N_7959,N_5138,N_3317);
or U7960 (N_7960,N_4824,N_5978);
nor U7961 (N_7961,N_4234,N_5291);
or U7962 (N_7962,N_4391,N_5508);
or U7963 (N_7963,N_3410,N_4573);
or U7964 (N_7964,N_5721,N_4220);
or U7965 (N_7965,N_4794,N_5976);
or U7966 (N_7966,N_5285,N_5606);
and U7967 (N_7967,N_4487,N_3474);
nor U7968 (N_7968,N_3481,N_4030);
or U7969 (N_7969,N_4934,N_3776);
nor U7970 (N_7970,N_4540,N_5056);
or U7971 (N_7971,N_4398,N_3972);
and U7972 (N_7972,N_5706,N_4472);
nand U7973 (N_7973,N_3509,N_3865);
nor U7974 (N_7974,N_3681,N_3784);
nor U7975 (N_7975,N_4649,N_5300);
or U7976 (N_7976,N_4621,N_3528);
nor U7977 (N_7977,N_3047,N_4524);
and U7978 (N_7978,N_3860,N_5521);
xor U7979 (N_7979,N_5396,N_5961);
nor U7980 (N_7980,N_4579,N_4466);
nand U7981 (N_7981,N_5473,N_4709);
nor U7982 (N_7982,N_5904,N_3191);
or U7983 (N_7983,N_3037,N_4962);
nand U7984 (N_7984,N_4480,N_5627);
nand U7985 (N_7985,N_3601,N_3662);
nor U7986 (N_7986,N_5232,N_3385);
or U7987 (N_7987,N_3551,N_4131);
and U7988 (N_7988,N_5631,N_4275);
and U7989 (N_7989,N_5262,N_5645);
nand U7990 (N_7990,N_4317,N_3315);
xnor U7991 (N_7991,N_4743,N_3970);
xor U7992 (N_7992,N_4342,N_4664);
nor U7993 (N_7993,N_5466,N_5675);
or U7994 (N_7994,N_3042,N_4677);
nand U7995 (N_7995,N_5243,N_3368);
or U7996 (N_7996,N_4192,N_5215);
nor U7997 (N_7997,N_5255,N_5832);
or U7998 (N_7998,N_5028,N_4860);
and U7999 (N_7999,N_3441,N_4994);
and U8000 (N_8000,N_5893,N_4248);
nand U8001 (N_8001,N_3299,N_3874);
or U8002 (N_8002,N_4574,N_5917);
and U8003 (N_8003,N_4538,N_3647);
or U8004 (N_8004,N_4055,N_5658);
or U8005 (N_8005,N_3632,N_5151);
nand U8006 (N_8006,N_5150,N_3923);
and U8007 (N_8007,N_3372,N_5134);
nand U8008 (N_8008,N_3124,N_5720);
or U8009 (N_8009,N_3236,N_4035);
nand U8010 (N_8010,N_4891,N_4139);
nor U8011 (N_8011,N_3056,N_4254);
and U8012 (N_8012,N_4364,N_4777);
nor U8013 (N_8013,N_4360,N_5730);
or U8014 (N_8014,N_5698,N_4376);
nor U8015 (N_8015,N_3884,N_3633);
or U8016 (N_8016,N_4279,N_4305);
nor U8017 (N_8017,N_4123,N_4153);
xnor U8018 (N_8018,N_5509,N_5979);
nand U8019 (N_8019,N_5981,N_5688);
nand U8020 (N_8020,N_3732,N_5258);
and U8021 (N_8021,N_3103,N_3395);
nand U8022 (N_8022,N_4836,N_5718);
or U8023 (N_8023,N_5845,N_5211);
nand U8024 (N_8024,N_4701,N_3162);
and U8025 (N_8025,N_5399,N_3875);
or U8026 (N_8026,N_5111,N_4630);
nor U8027 (N_8027,N_4723,N_4748);
nand U8028 (N_8028,N_4751,N_4926);
or U8029 (N_8029,N_4375,N_4423);
or U8030 (N_8030,N_3561,N_5955);
and U8031 (N_8031,N_5459,N_3910);
nand U8032 (N_8032,N_4401,N_3380);
nand U8033 (N_8033,N_3622,N_3921);
nor U8034 (N_8034,N_3438,N_5423);
nor U8035 (N_8035,N_4946,N_5931);
or U8036 (N_8036,N_5679,N_4259);
nor U8037 (N_8037,N_4336,N_5809);
or U8038 (N_8038,N_4411,N_5753);
or U8039 (N_8039,N_4142,N_5814);
or U8040 (N_8040,N_4480,N_3466);
nor U8041 (N_8041,N_5856,N_5972);
nor U8042 (N_8042,N_3606,N_3386);
xnor U8043 (N_8043,N_4983,N_3199);
nand U8044 (N_8044,N_4806,N_3457);
nor U8045 (N_8045,N_4270,N_4474);
or U8046 (N_8046,N_3126,N_4674);
nor U8047 (N_8047,N_5952,N_4535);
nand U8048 (N_8048,N_3336,N_4957);
and U8049 (N_8049,N_4643,N_5336);
or U8050 (N_8050,N_5043,N_5239);
or U8051 (N_8051,N_4204,N_3532);
or U8052 (N_8052,N_3031,N_5093);
or U8053 (N_8053,N_4615,N_5457);
or U8054 (N_8054,N_3016,N_4751);
nor U8055 (N_8055,N_3458,N_3138);
nor U8056 (N_8056,N_4422,N_5902);
nand U8057 (N_8057,N_3346,N_3088);
nor U8058 (N_8058,N_5821,N_4027);
and U8059 (N_8059,N_5905,N_3360);
or U8060 (N_8060,N_3085,N_5654);
nor U8061 (N_8061,N_4003,N_5712);
nor U8062 (N_8062,N_4161,N_3901);
nand U8063 (N_8063,N_3319,N_5918);
nand U8064 (N_8064,N_5573,N_3065);
and U8065 (N_8065,N_5765,N_3008);
or U8066 (N_8066,N_3798,N_4923);
and U8067 (N_8067,N_4730,N_3697);
nor U8068 (N_8068,N_4885,N_5951);
nor U8069 (N_8069,N_3922,N_4074);
nor U8070 (N_8070,N_5334,N_3066);
and U8071 (N_8071,N_4415,N_4854);
or U8072 (N_8072,N_5721,N_3823);
or U8073 (N_8073,N_5873,N_5418);
nor U8074 (N_8074,N_3086,N_4206);
nand U8075 (N_8075,N_3195,N_5222);
and U8076 (N_8076,N_4993,N_3856);
nor U8077 (N_8077,N_5620,N_3011);
or U8078 (N_8078,N_4645,N_3344);
or U8079 (N_8079,N_4375,N_3692);
nand U8080 (N_8080,N_3647,N_4197);
nor U8081 (N_8081,N_3356,N_4044);
nand U8082 (N_8082,N_3707,N_5858);
and U8083 (N_8083,N_5369,N_5267);
or U8084 (N_8084,N_5341,N_4224);
or U8085 (N_8085,N_5453,N_3536);
or U8086 (N_8086,N_5358,N_4138);
nor U8087 (N_8087,N_3440,N_3457);
nor U8088 (N_8088,N_5524,N_5265);
nor U8089 (N_8089,N_4088,N_3544);
and U8090 (N_8090,N_4884,N_3186);
nand U8091 (N_8091,N_3658,N_5385);
or U8092 (N_8092,N_5967,N_3210);
or U8093 (N_8093,N_3322,N_3096);
nand U8094 (N_8094,N_3273,N_4575);
nor U8095 (N_8095,N_3201,N_5716);
and U8096 (N_8096,N_4798,N_3292);
and U8097 (N_8097,N_4699,N_5362);
nor U8098 (N_8098,N_4543,N_5638);
or U8099 (N_8099,N_5615,N_4603);
or U8100 (N_8100,N_4261,N_4571);
nor U8101 (N_8101,N_4529,N_3336);
nor U8102 (N_8102,N_5113,N_3444);
or U8103 (N_8103,N_4872,N_5353);
and U8104 (N_8104,N_5385,N_5024);
or U8105 (N_8105,N_5757,N_3634);
or U8106 (N_8106,N_4814,N_4673);
nor U8107 (N_8107,N_3964,N_4049);
and U8108 (N_8108,N_3452,N_3782);
nand U8109 (N_8109,N_3669,N_5854);
nor U8110 (N_8110,N_5268,N_4514);
or U8111 (N_8111,N_5405,N_3124);
xor U8112 (N_8112,N_3645,N_4969);
nor U8113 (N_8113,N_5433,N_5187);
and U8114 (N_8114,N_5895,N_5547);
nor U8115 (N_8115,N_4193,N_3702);
or U8116 (N_8116,N_4883,N_4149);
and U8117 (N_8117,N_3713,N_3063);
and U8118 (N_8118,N_3360,N_3321);
nand U8119 (N_8119,N_3964,N_4118);
nand U8120 (N_8120,N_3073,N_4504);
and U8121 (N_8121,N_5154,N_3922);
and U8122 (N_8122,N_5582,N_5074);
and U8123 (N_8123,N_4512,N_3622);
nor U8124 (N_8124,N_4149,N_4605);
nor U8125 (N_8125,N_4972,N_4199);
nand U8126 (N_8126,N_5955,N_3494);
nand U8127 (N_8127,N_5575,N_5092);
nand U8128 (N_8128,N_4673,N_3222);
and U8129 (N_8129,N_4812,N_3555);
nand U8130 (N_8130,N_4721,N_3334);
or U8131 (N_8131,N_3499,N_3476);
or U8132 (N_8132,N_4575,N_3102);
and U8133 (N_8133,N_5481,N_3640);
or U8134 (N_8134,N_5573,N_3824);
nor U8135 (N_8135,N_3058,N_5584);
or U8136 (N_8136,N_4024,N_4259);
or U8137 (N_8137,N_3162,N_4923);
nand U8138 (N_8138,N_5316,N_4554);
nor U8139 (N_8139,N_5387,N_5645);
xor U8140 (N_8140,N_3285,N_4009);
or U8141 (N_8141,N_3656,N_5682);
nand U8142 (N_8142,N_3448,N_4347);
and U8143 (N_8143,N_4927,N_5712);
nand U8144 (N_8144,N_5026,N_3506);
and U8145 (N_8145,N_3935,N_5156);
nor U8146 (N_8146,N_5340,N_5195);
xor U8147 (N_8147,N_4008,N_5235);
and U8148 (N_8148,N_4386,N_3033);
or U8149 (N_8149,N_3739,N_4072);
or U8150 (N_8150,N_5750,N_5998);
nand U8151 (N_8151,N_4970,N_3037);
nor U8152 (N_8152,N_5071,N_4126);
nor U8153 (N_8153,N_3484,N_3754);
nor U8154 (N_8154,N_3178,N_5306);
and U8155 (N_8155,N_5265,N_4748);
or U8156 (N_8156,N_3178,N_3574);
or U8157 (N_8157,N_5576,N_3245);
nor U8158 (N_8158,N_3653,N_5753);
nor U8159 (N_8159,N_3899,N_5389);
or U8160 (N_8160,N_4609,N_5555);
or U8161 (N_8161,N_3842,N_3884);
nand U8162 (N_8162,N_3893,N_5869);
nor U8163 (N_8163,N_5926,N_5340);
and U8164 (N_8164,N_3058,N_4511);
or U8165 (N_8165,N_4404,N_3078);
nor U8166 (N_8166,N_5458,N_5711);
or U8167 (N_8167,N_4581,N_4685);
or U8168 (N_8168,N_5686,N_3335);
or U8169 (N_8169,N_4049,N_3785);
or U8170 (N_8170,N_3086,N_4293);
or U8171 (N_8171,N_5980,N_5530);
nand U8172 (N_8172,N_3076,N_4792);
or U8173 (N_8173,N_3410,N_5910);
nor U8174 (N_8174,N_5496,N_5200);
or U8175 (N_8175,N_4086,N_4043);
xnor U8176 (N_8176,N_5340,N_5387);
nor U8177 (N_8177,N_5928,N_5250);
or U8178 (N_8178,N_3239,N_4442);
nor U8179 (N_8179,N_4621,N_4701);
nor U8180 (N_8180,N_5893,N_3077);
nor U8181 (N_8181,N_4278,N_4732);
nand U8182 (N_8182,N_4781,N_3853);
nand U8183 (N_8183,N_5631,N_3697);
and U8184 (N_8184,N_3536,N_4229);
nand U8185 (N_8185,N_5213,N_5418);
and U8186 (N_8186,N_3635,N_5491);
or U8187 (N_8187,N_3641,N_5546);
and U8188 (N_8188,N_4843,N_3666);
or U8189 (N_8189,N_5760,N_5769);
nor U8190 (N_8190,N_4155,N_4216);
nor U8191 (N_8191,N_5368,N_5132);
nand U8192 (N_8192,N_4498,N_4809);
nor U8193 (N_8193,N_3684,N_4519);
or U8194 (N_8194,N_3589,N_4343);
nor U8195 (N_8195,N_3864,N_5291);
xor U8196 (N_8196,N_5433,N_3372);
nand U8197 (N_8197,N_3597,N_5171);
or U8198 (N_8198,N_4955,N_3147);
or U8199 (N_8199,N_5778,N_4469);
nand U8200 (N_8200,N_5117,N_4180);
nor U8201 (N_8201,N_4473,N_4251);
nor U8202 (N_8202,N_5007,N_3338);
nand U8203 (N_8203,N_5171,N_3937);
and U8204 (N_8204,N_4679,N_4776);
nand U8205 (N_8205,N_4401,N_4641);
or U8206 (N_8206,N_4481,N_4759);
and U8207 (N_8207,N_5037,N_4985);
nand U8208 (N_8208,N_3200,N_4671);
nand U8209 (N_8209,N_3610,N_5909);
nand U8210 (N_8210,N_3263,N_4849);
or U8211 (N_8211,N_5489,N_4201);
and U8212 (N_8212,N_4612,N_3807);
nand U8213 (N_8213,N_5320,N_3391);
or U8214 (N_8214,N_5980,N_4899);
and U8215 (N_8215,N_4154,N_3086);
and U8216 (N_8216,N_4072,N_4631);
and U8217 (N_8217,N_5901,N_4498);
and U8218 (N_8218,N_3208,N_3730);
nand U8219 (N_8219,N_3272,N_4417);
and U8220 (N_8220,N_4673,N_5371);
nand U8221 (N_8221,N_3382,N_3590);
or U8222 (N_8222,N_3368,N_4296);
and U8223 (N_8223,N_4932,N_5820);
or U8224 (N_8224,N_3240,N_4154);
nor U8225 (N_8225,N_4632,N_3401);
and U8226 (N_8226,N_4746,N_3639);
nor U8227 (N_8227,N_3776,N_3011);
and U8228 (N_8228,N_3906,N_3659);
nand U8229 (N_8229,N_3266,N_4933);
xnor U8230 (N_8230,N_4730,N_4315);
and U8231 (N_8231,N_5531,N_3328);
and U8232 (N_8232,N_5570,N_3428);
nor U8233 (N_8233,N_4166,N_4710);
nor U8234 (N_8234,N_4436,N_4189);
nand U8235 (N_8235,N_4866,N_3135);
nand U8236 (N_8236,N_5907,N_5260);
and U8237 (N_8237,N_5459,N_3298);
and U8238 (N_8238,N_5323,N_3096);
nand U8239 (N_8239,N_5636,N_3446);
or U8240 (N_8240,N_5553,N_3027);
or U8241 (N_8241,N_5152,N_3200);
nand U8242 (N_8242,N_3513,N_5266);
nor U8243 (N_8243,N_3825,N_5396);
nand U8244 (N_8244,N_5765,N_3386);
and U8245 (N_8245,N_3860,N_4969);
nor U8246 (N_8246,N_4763,N_4631);
and U8247 (N_8247,N_5379,N_5345);
nand U8248 (N_8248,N_4587,N_5587);
or U8249 (N_8249,N_4379,N_5508);
or U8250 (N_8250,N_3259,N_3192);
nor U8251 (N_8251,N_5658,N_3064);
or U8252 (N_8252,N_4599,N_5396);
or U8253 (N_8253,N_3480,N_5582);
nand U8254 (N_8254,N_3632,N_3328);
nor U8255 (N_8255,N_4544,N_4511);
or U8256 (N_8256,N_3509,N_3868);
or U8257 (N_8257,N_3968,N_4768);
nor U8258 (N_8258,N_4565,N_4753);
nor U8259 (N_8259,N_5945,N_4287);
nand U8260 (N_8260,N_3871,N_3505);
and U8261 (N_8261,N_3231,N_3976);
and U8262 (N_8262,N_5687,N_5432);
nand U8263 (N_8263,N_3131,N_4021);
or U8264 (N_8264,N_4074,N_5278);
nand U8265 (N_8265,N_3286,N_3634);
nand U8266 (N_8266,N_3361,N_3724);
or U8267 (N_8267,N_4775,N_4874);
or U8268 (N_8268,N_5258,N_4582);
nor U8269 (N_8269,N_5455,N_5056);
nor U8270 (N_8270,N_5786,N_5591);
or U8271 (N_8271,N_4111,N_4537);
nor U8272 (N_8272,N_5081,N_3876);
and U8273 (N_8273,N_3355,N_5939);
nand U8274 (N_8274,N_4622,N_3364);
and U8275 (N_8275,N_4482,N_4411);
nor U8276 (N_8276,N_3722,N_3335);
nor U8277 (N_8277,N_3538,N_5352);
and U8278 (N_8278,N_3935,N_5676);
nand U8279 (N_8279,N_3527,N_5723);
nor U8280 (N_8280,N_3641,N_4658);
nor U8281 (N_8281,N_4860,N_5544);
nor U8282 (N_8282,N_4140,N_3323);
and U8283 (N_8283,N_3599,N_3544);
nor U8284 (N_8284,N_4677,N_4993);
nand U8285 (N_8285,N_5352,N_5777);
nor U8286 (N_8286,N_5760,N_5309);
and U8287 (N_8287,N_4851,N_5270);
and U8288 (N_8288,N_5439,N_5345);
and U8289 (N_8289,N_4054,N_3887);
nor U8290 (N_8290,N_3056,N_3011);
or U8291 (N_8291,N_3713,N_5802);
or U8292 (N_8292,N_3335,N_5572);
nand U8293 (N_8293,N_4546,N_3223);
and U8294 (N_8294,N_5059,N_4935);
and U8295 (N_8295,N_3148,N_5746);
nand U8296 (N_8296,N_4215,N_4598);
and U8297 (N_8297,N_4444,N_3263);
and U8298 (N_8298,N_5657,N_5323);
nor U8299 (N_8299,N_5779,N_4258);
or U8300 (N_8300,N_4111,N_3641);
and U8301 (N_8301,N_4865,N_5728);
or U8302 (N_8302,N_5903,N_3143);
nand U8303 (N_8303,N_4332,N_4954);
nor U8304 (N_8304,N_5204,N_4873);
or U8305 (N_8305,N_4692,N_5886);
nand U8306 (N_8306,N_3960,N_4776);
nor U8307 (N_8307,N_3213,N_5547);
nor U8308 (N_8308,N_5225,N_4682);
nand U8309 (N_8309,N_4717,N_3118);
nor U8310 (N_8310,N_5336,N_5861);
or U8311 (N_8311,N_3212,N_3289);
nand U8312 (N_8312,N_4205,N_4732);
and U8313 (N_8313,N_3614,N_4626);
nand U8314 (N_8314,N_3448,N_4297);
or U8315 (N_8315,N_4400,N_4274);
or U8316 (N_8316,N_4913,N_4410);
nor U8317 (N_8317,N_5799,N_4969);
nor U8318 (N_8318,N_3588,N_3332);
or U8319 (N_8319,N_3939,N_3911);
and U8320 (N_8320,N_5917,N_4749);
nor U8321 (N_8321,N_3229,N_5786);
nand U8322 (N_8322,N_3872,N_4218);
nor U8323 (N_8323,N_4999,N_4652);
nand U8324 (N_8324,N_3582,N_5859);
nor U8325 (N_8325,N_4769,N_4072);
nor U8326 (N_8326,N_5162,N_3962);
or U8327 (N_8327,N_4936,N_5520);
or U8328 (N_8328,N_4755,N_5148);
and U8329 (N_8329,N_3111,N_5752);
or U8330 (N_8330,N_4611,N_5365);
nand U8331 (N_8331,N_4227,N_5627);
nor U8332 (N_8332,N_3034,N_3952);
and U8333 (N_8333,N_4366,N_4305);
and U8334 (N_8334,N_4259,N_4146);
or U8335 (N_8335,N_3244,N_3015);
nand U8336 (N_8336,N_5632,N_3652);
and U8337 (N_8337,N_5142,N_3524);
and U8338 (N_8338,N_5752,N_5542);
xor U8339 (N_8339,N_5378,N_4382);
nor U8340 (N_8340,N_3045,N_5839);
nor U8341 (N_8341,N_4032,N_5962);
and U8342 (N_8342,N_3957,N_5460);
and U8343 (N_8343,N_4313,N_4194);
nand U8344 (N_8344,N_4020,N_4665);
nor U8345 (N_8345,N_5428,N_3090);
or U8346 (N_8346,N_4742,N_5973);
or U8347 (N_8347,N_3284,N_4556);
and U8348 (N_8348,N_4022,N_4654);
and U8349 (N_8349,N_3595,N_4974);
and U8350 (N_8350,N_5665,N_4658);
and U8351 (N_8351,N_4430,N_5595);
and U8352 (N_8352,N_3529,N_5961);
nand U8353 (N_8353,N_4112,N_5628);
nand U8354 (N_8354,N_5039,N_3997);
and U8355 (N_8355,N_5994,N_5275);
nor U8356 (N_8356,N_3778,N_5866);
or U8357 (N_8357,N_4895,N_3976);
nand U8358 (N_8358,N_4373,N_5433);
or U8359 (N_8359,N_5068,N_3954);
nand U8360 (N_8360,N_3430,N_5019);
nand U8361 (N_8361,N_5286,N_3345);
nand U8362 (N_8362,N_3423,N_3153);
and U8363 (N_8363,N_5078,N_3599);
nor U8364 (N_8364,N_4812,N_5273);
or U8365 (N_8365,N_5417,N_5741);
nor U8366 (N_8366,N_3673,N_5741);
nand U8367 (N_8367,N_3905,N_4032);
nand U8368 (N_8368,N_4780,N_3317);
nand U8369 (N_8369,N_3700,N_4850);
and U8370 (N_8370,N_5209,N_4688);
nand U8371 (N_8371,N_5372,N_3145);
or U8372 (N_8372,N_5205,N_3105);
nor U8373 (N_8373,N_5865,N_5449);
or U8374 (N_8374,N_4567,N_4514);
xnor U8375 (N_8375,N_5218,N_5723);
nand U8376 (N_8376,N_3863,N_3948);
nand U8377 (N_8377,N_5775,N_5734);
and U8378 (N_8378,N_5962,N_3671);
or U8379 (N_8379,N_5551,N_4743);
or U8380 (N_8380,N_3648,N_4098);
nand U8381 (N_8381,N_5608,N_5265);
and U8382 (N_8382,N_5413,N_3979);
or U8383 (N_8383,N_4906,N_5218);
nor U8384 (N_8384,N_4156,N_3561);
and U8385 (N_8385,N_3305,N_5684);
and U8386 (N_8386,N_5112,N_5595);
nor U8387 (N_8387,N_5951,N_3766);
or U8388 (N_8388,N_5286,N_3254);
and U8389 (N_8389,N_3885,N_5632);
and U8390 (N_8390,N_5670,N_4578);
or U8391 (N_8391,N_4240,N_3808);
and U8392 (N_8392,N_4974,N_3305);
nor U8393 (N_8393,N_5196,N_4378);
and U8394 (N_8394,N_3906,N_3745);
or U8395 (N_8395,N_4387,N_5493);
nor U8396 (N_8396,N_5540,N_5101);
nor U8397 (N_8397,N_5034,N_4413);
or U8398 (N_8398,N_4405,N_4974);
nand U8399 (N_8399,N_3777,N_5585);
or U8400 (N_8400,N_3266,N_4907);
nand U8401 (N_8401,N_4226,N_5106);
nor U8402 (N_8402,N_5677,N_5815);
nand U8403 (N_8403,N_3768,N_3260);
nand U8404 (N_8404,N_3312,N_3180);
nor U8405 (N_8405,N_5339,N_4415);
nor U8406 (N_8406,N_5996,N_4084);
or U8407 (N_8407,N_3082,N_3345);
or U8408 (N_8408,N_4681,N_5306);
or U8409 (N_8409,N_4024,N_5816);
or U8410 (N_8410,N_5174,N_5409);
and U8411 (N_8411,N_3092,N_4585);
or U8412 (N_8412,N_5720,N_5555);
or U8413 (N_8413,N_3006,N_4362);
nand U8414 (N_8414,N_3608,N_3569);
or U8415 (N_8415,N_5972,N_5931);
nand U8416 (N_8416,N_5531,N_5214);
nand U8417 (N_8417,N_4201,N_4389);
and U8418 (N_8418,N_3681,N_3755);
nor U8419 (N_8419,N_3296,N_3280);
or U8420 (N_8420,N_4481,N_5271);
or U8421 (N_8421,N_5884,N_5058);
and U8422 (N_8422,N_5618,N_5510);
nand U8423 (N_8423,N_5977,N_4289);
nand U8424 (N_8424,N_3002,N_4786);
or U8425 (N_8425,N_5849,N_4876);
nand U8426 (N_8426,N_4349,N_5402);
or U8427 (N_8427,N_4741,N_5294);
and U8428 (N_8428,N_5133,N_3920);
nand U8429 (N_8429,N_4113,N_4255);
nor U8430 (N_8430,N_3567,N_5615);
and U8431 (N_8431,N_5474,N_4110);
and U8432 (N_8432,N_4447,N_4073);
nand U8433 (N_8433,N_3774,N_5992);
nand U8434 (N_8434,N_5121,N_4514);
nor U8435 (N_8435,N_4710,N_3351);
and U8436 (N_8436,N_5174,N_4156);
nand U8437 (N_8437,N_4935,N_4227);
xor U8438 (N_8438,N_4409,N_3943);
and U8439 (N_8439,N_4082,N_3526);
or U8440 (N_8440,N_3977,N_5387);
or U8441 (N_8441,N_4548,N_5071);
nand U8442 (N_8442,N_5660,N_3005);
and U8443 (N_8443,N_3295,N_3818);
nand U8444 (N_8444,N_4778,N_4888);
or U8445 (N_8445,N_5366,N_4476);
xor U8446 (N_8446,N_4004,N_4228);
nor U8447 (N_8447,N_3844,N_5391);
nand U8448 (N_8448,N_5606,N_4225);
nand U8449 (N_8449,N_4123,N_5405);
nand U8450 (N_8450,N_3684,N_3619);
or U8451 (N_8451,N_4112,N_4708);
and U8452 (N_8452,N_3793,N_3154);
and U8453 (N_8453,N_3426,N_4054);
and U8454 (N_8454,N_3494,N_5108);
or U8455 (N_8455,N_3293,N_4328);
nand U8456 (N_8456,N_5967,N_5801);
nor U8457 (N_8457,N_3251,N_4951);
and U8458 (N_8458,N_4764,N_3324);
nand U8459 (N_8459,N_4849,N_5179);
and U8460 (N_8460,N_3212,N_5430);
nand U8461 (N_8461,N_4985,N_4434);
and U8462 (N_8462,N_3059,N_3845);
xor U8463 (N_8463,N_3677,N_5075);
xor U8464 (N_8464,N_5037,N_3193);
nor U8465 (N_8465,N_4726,N_3690);
and U8466 (N_8466,N_4706,N_4426);
nand U8467 (N_8467,N_3127,N_5547);
and U8468 (N_8468,N_5976,N_4106);
nor U8469 (N_8469,N_5077,N_5337);
xor U8470 (N_8470,N_4070,N_5818);
or U8471 (N_8471,N_5811,N_3202);
and U8472 (N_8472,N_5786,N_4830);
and U8473 (N_8473,N_5956,N_5550);
and U8474 (N_8474,N_5482,N_3929);
nor U8475 (N_8475,N_3802,N_4936);
nand U8476 (N_8476,N_4678,N_5362);
or U8477 (N_8477,N_3550,N_4810);
nand U8478 (N_8478,N_3280,N_5633);
nand U8479 (N_8479,N_4236,N_3690);
nor U8480 (N_8480,N_3503,N_3914);
nand U8481 (N_8481,N_3361,N_4631);
or U8482 (N_8482,N_3140,N_3253);
xor U8483 (N_8483,N_5187,N_3611);
or U8484 (N_8484,N_3826,N_5277);
and U8485 (N_8485,N_5804,N_5155);
or U8486 (N_8486,N_5920,N_5293);
and U8487 (N_8487,N_4608,N_5075);
or U8488 (N_8488,N_4126,N_3771);
and U8489 (N_8489,N_4667,N_5692);
and U8490 (N_8490,N_4850,N_3154);
nand U8491 (N_8491,N_3951,N_4645);
nand U8492 (N_8492,N_4113,N_4121);
and U8493 (N_8493,N_3934,N_5135);
nor U8494 (N_8494,N_3422,N_3923);
or U8495 (N_8495,N_4152,N_3873);
or U8496 (N_8496,N_3262,N_3900);
and U8497 (N_8497,N_3153,N_5024);
and U8498 (N_8498,N_4259,N_5786);
nand U8499 (N_8499,N_4508,N_3214);
nand U8500 (N_8500,N_3088,N_5871);
nand U8501 (N_8501,N_3975,N_5615);
and U8502 (N_8502,N_4319,N_4214);
and U8503 (N_8503,N_4894,N_3616);
and U8504 (N_8504,N_3002,N_3614);
or U8505 (N_8505,N_3611,N_3005);
nor U8506 (N_8506,N_5257,N_5576);
or U8507 (N_8507,N_5312,N_5686);
or U8508 (N_8508,N_3581,N_3955);
and U8509 (N_8509,N_4993,N_4157);
nand U8510 (N_8510,N_3068,N_3705);
and U8511 (N_8511,N_3132,N_4886);
nor U8512 (N_8512,N_5301,N_5827);
or U8513 (N_8513,N_5803,N_4756);
and U8514 (N_8514,N_3000,N_5831);
or U8515 (N_8515,N_5045,N_5642);
and U8516 (N_8516,N_3676,N_4977);
or U8517 (N_8517,N_4634,N_4892);
and U8518 (N_8518,N_3702,N_3752);
or U8519 (N_8519,N_5276,N_5961);
or U8520 (N_8520,N_4299,N_5303);
nor U8521 (N_8521,N_3042,N_5535);
or U8522 (N_8522,N_3320,N_3060);
nand U8523 (N_8523,N_3077,N_5285);
and U8524 (N_8524,N_3368,N_3935);
and U8525 (N_8525,N_3434,N_3208);
nand U8526 (N_8526,N_4787,N_4611);
and U8527 (N_8527,N_4106,N_3693);
nor U8528 (N_8528,N_5586,N_5277);
and U8529 (N_8529,N_4269,N_5577);
and U8530 (N_8530,N_4963,N_4511);
nand U8531 (N_8531,N_3261,N_5789);
nand U8532 (N_8532,N_3554,N_5965);
or U8533 (N_8533,N_4681,N_4456);
nand U8534 (N_8534,N_4309,N_5057);
nor U8535 (N_8535,N_5515,N_5276);
and U8536 (N_8536,N_5234,N_3625);
nand U8537 (N_8537,N_5841,N_3995);
and U8538 (N_8538,N_5626,N_5868);
nand U8539 (N_8539,N_5834,N_5664);
or U8540 (N_8540,N_3338,N_4184);
xnor U8541 (N_8541,N_4108,N_4891);
nand U8542 (N_8542,N_5980,N_3449);
and U8543 (N_8543,N_5269,N_3692);
nand U8544 (N_8544,N_3536,N_3854);
or U8545 (N_8545,N_4906,N_3082);
nor U8546 (N_8546,N_3427,N_4666);
or U8547 (N_8547,N_5907,N_3210);
or U8548 (N_8548,N_4178,N_3826);
or U8549 (N_8549,N_4655,N_3378);
xnor U8550 (N_8550,N_5074,N_5626);
xor U8551 (N_8551,N_3615,N_5088);
and U8552 (N_8552,N_3914,N_3957);
xor U8553 (N_8553,N_3090,N_5850);
nand U8554 (N_8554,N_4073,N_3410);
and U8555 (N_8555,N_4772,N_3127);
and U8556 (N_8556,N_3820,N_5105);
nor U8557 (N_8557,N_5039,N_3452);
and U8558 (N_8558,N_4378,N_4434);
and U8559 (N_8559,N_4283,N_3473);
and U8560 (N_8560,N_5920,N_4608);
nor U8561 (N_8561,N_3382,N_5657);
nor U8562 (N_8562,N_5281,N_3388);
nand U8563 (N_8563,N_5000,N_5967);
and U8564 (N_8564,N_5083,N_4581);
xor U8565 (N_8565,N_4291,N_4342);
nor U8566 (N_8566,N_3001,N_3106);
nand U8567 (N_8567,N_3177,N_5329);
nor U8568 (N_8568,N_5348,N_5409);
nand U8569 (N_8569,N_3209,N_4484);
nand U8570 (N_8570,N_5966,N_3078);
and U8571 (N_8571,N_5758,N_3452);
or U8572 (N_8572,N_5831,N_5147);
nor U8573 (N_8573,N_3985,N_3447);
nand U8574 (N_8574,N_4206,N_5491);
nand U8575 (N_8575,N_3150,N_5269);
or U8576 (N_8576,N_3925,N_5302);
nor U8577 (N_8577,N_3724,N_4587);
nor U8578 (N_8578,N_4810,N_3963);
and U8579 (N_8579,N_3350,N_4078);
or U8580 (N_8580,N_3797,N_4121);
and U8581 (N_8581,N_5420,N_3068);
or U8582 (N_8582,N_4136,N_4548);
nand U8583 (N_8583,N_3820,N_5674);
or U8584 (N_8584,N_4917,N_4456);
nor U8585 (N_8585,N_4217,N_5081);
or U8586 (N_8586,N_3410,N_3700);
or U8587 (N_8587,N_3773,N_5532);
or U8588 (N_8588,N_3655,N_5975);
nor U8589 (N_8589,N_5600,N_4077);
and U8590 (N_8590,N_3403,N_4789);
nand U8591 (N_8591,N_3849,N_4993);
nor U8592 (N_8592,N_5675,N_4362);
nand U8593 (N_8593,N_4650,N_5546);
nor U8594 (N_8594,N_4511,N_3168);
nand U8595 (N_8595,N_5024,N_5148);
nor U8596 (N_8596,N_4664,N_4804);
nor U8597 (N_8597,N_5813,N_4696);
xor U8598 (N_8598,N_3645,N_4887);
nand U8599 (N_8599,N_5746,N_5133);
nor U8600 (N_8600,N_3853,N_5629);
and U8601 (N_8601,N_4656,N_5965);
nor U8602 (N_8602,N_5039,N_5478);
and U8603 (N_8603,N_3284,N_5059);
and U8604 (N_8604,N_3821,N_4283);
and U8605 (N_8605,N_4783,N_3611);
nand U8606 (N_8606,N_4862,N_5733);
and U8607 (N_8607,N_4483,N_3272);
nor U8608 (N_8608,N_5008,N_3569);
nand U8609 (N_8609,N_4931,N_5283);
nand U8610 (N_8610,N_5239,N_4099);
nor U8611 (N_8611,N_4027,N_3959);
and U8612 (N_8612,N_5411,N_3065);
or U8613 (N_8613,N_4962,N_3602);
or U8614 (N_8614,N_4160,N_3773);
or U8615 (N_8615,N_4572,N_3848);
or U8616 (N_8616,N_4306,N_4641);
and U8617 (N_8617,N_4643,N_3211);
nand U8618 (N_8618,N_3780,N_3537);
nand U8619 (N_8619,N_3465,N_4136);
and U8620 (N_8620,N_5393,N_5408);
or U8621 (N_8621,N_5428,N_3086);
nand U8622 (N_8622,N_5165,N_5230);
xor U8623 (N_8623,N_3428,N_3162);
nand U8624 (N_8624,N_4914,N_4631);
xor U8625 (N_8625,N_3343,N_5732);
nand U8626 (N_8626,N_5388,N_4588);
or U8627 (N_8627,N_3781,N_3911);
nor U8628 (N_8628,N_4793,N_5432);
nor U8629 (N_8629,N_5284,N_5329);
nor U8630 (N_8630,N_3135,N_3092);
nand U8631 (N_8631,N_5778,N_3713);
nor U8632 (N_8632,N_4230,N_3353);
or U8633 (N_8633,N_3745,N_4002);
and U8634 (N_8634,N_4371,N_4530);
or U8635 (N_8635,N_3289,N_5276);
or U8636 (N_8636,N_5395,N_5107);
and U8637 (N_8637,N_5548,N_3983);
and U8638 (N_8638,N_4518,N_3390);
nor U8639 (N_8639,N_3276,N_3824);
or U8640 (N_8640,N_3439,N_5846);
nor U8641 (N_8641,N_4509,N_4208);
nor U8642 (N_8642,N_5979,N_4635);
or U8643 (N_8643,N_4971,N_4289);
and U8644 (N_8644,N_5896,N_5161);
nand U8645 (N_8645,N_5295,N_5786);
nand U8646 (N_8646,N_5841,N_5709);
or U8647 (N_8647,N_5126,N_5435);
nor U8648 (N_8648,N_3172,N_5287);
and U8649 (N_8649,N_5885,N_3014);
nor U8650 (N_8650,N_4315,N_5911);
or U8651 (N_8651,N_3313,N_5666);
and U8652 (N_8652,N_3026,N_5331);
nand U8653 (N_8653,N_3295,N_5870);
nand U8654 (N_8654,N_3624,N_5505);
nand U8655 (N_8655,N_5927,N_4141);
or U8656 (N_8656,N_5965,N_3163);
and U8657 (N_8657,N_5249,N_4607);
and U8658 (N_8658,N_3450,N_5314);
xnor U8659 (N_8659,N_4774,N_3181);
nand U8660 (N_8660,N_3456,N_5240);
and U8661 (N_8661,N_3994,N_5933);
or U8662 (N_8662,N_5337,N_5080);
nor U8663 (N_8663,N_5179,N_5092);
nand U8664 (N_8664,N_4838,N_4126);
nor U8665 (N_8665,N_4876,N_5970);
and U8666 (N_8666,N_4287,N_3428);
nor U8667 (N_8667,N_5433,N_5536);
or U8668 (N_8668,N_3093,N_4171);
nand U8669 (N_8669,N_4852,N_3670);
nand U8670 (N_8670,N_5088,N_4518);
nand U8671 (N_8671,N_5624,N_4836);
or U8672 (N_8672,N_4882,N_3393);
or U8673 (N_8673,N_5148,N_4565);
xnor U8674 (N_8674,N_4316,N_3933);
nand U8675 (N_8675,N_3103,N_5542);
or U8676 (N_8676,N_5211,N_3065);
and U8677 (N_8677,N_3439,N_3910);
nand U8678 (N_8678,N_5727,N_5761);
nor U8679 (N_8679,N_3474,N_4823);
nor U8680 (N_8680,N_3260,N_5911);
nand U8681 (N_8681,N_3482,N_5846);
or U8682 (N_8682,N_4044,N_3001);
nor U8683 (N_8683,N_3810,N_4455);
or U8684 (N_8684,N_5908,N_4943);
and U8685 (N_8685,N_4031,N_4922);
and U8686 (N_8686,N_4811,N_3066);
nor U8687 (N_8687,N_3282,N_4481);
nand U8688 (N_8688,N_4165,N_4559);
nand U8689 (N_8689,N_3649,N_3293);
nand U8690 (N_8690,N_3121,N_4977);
nor U8691 (N_8691,N_4609,N_3900);
nor U8692 (N_8692,N_4953,N_5065);
or U8693 (N_8693,N_5220,N_3668);
nand U8694 (N_8694,N_5834,N_3877);
or U8695 (N_8695,N_5051,N_3148);
nor U8696 (N_8696,N_3236,N_5950);
nand U8697 (N_8697,N_5255,N_3723);
or U8698 (N_8698,N_4681,N_5726);
and U8699 (N_8699,N_4810,N_3974);
and U8700 (N_8700,N_4599,N_5965);
nor U8701 (N_8701,N_4162,N_4409);
nand U8702 (N_8702,N_3914,N_3892);
nand U8703 (N_8703,N_5525,N_5948);
nor U8704 (N_8704,N_4035,N_4976);
xnor U8705 (N_8705,N_4116,N_3620);
nand U8706 (N_8706,N_5589,N_3981);
nor U8707 (N_8707,N_4756,N_3635);
nand U8708 (N_8708,N_3631,N_4055);
and U8709 (N_8709,N_4874,N_5710);
and U8710 (N_8710,N_3460,N_5983);
and U8711 (N_8711,N_5006,N_3801);
or U8712 (N_8712,N_4996,N_3748);
nor U8713 (N_8713,N_5635,N_3552);
or U8714 (N_8714,N_5694,N_5461);
nor U8715 (N_8715,N_3214,N_3993);
nor U8716 (N_8716,N_5532,N_4764);
or U8717 (N_8717,N_4002,N_3422);
xor U8718 (N_8718,N_4851,N_4448);
nand U8719 (N_8719,N_3508,N_4556);
nor U8720 (N_8720,N_3810,N_5675);
nand U8721 (N_8721,N_3560,N_4109);
nor U8722 (N_8722,N_3777,N_5526);
or U8723 (N_8723,N_3511,N_3388);
or U8724 (N_8724,N_3741,N_3411);
and U8725 (N_8725,N_4022,N_4031);
nand U8726 (N_8726,N_4644,N_3524);
or U8727 (N_8727,N_3233,N_4214);
nand U8728 (N_8728,N_5380,N_3981);
and U8729 (N_8729,N_5144,N_3948);
nand U8730 (N_8730,N_4830,N_4833);
and U8731 (N_8731,N_3535,N_5046);
and U8732 (N_8732,N_4796,N_4938);
and U8733 (N_8733,N_3451,N_3386);
or U8734 (N_8734,N_5374,N_4815);
or U8735 (N_8735,N_4442,N_4174);
or U8736 (N_8736,N_5311,N_4147);
nor U8737 (N_8737,N_5395,N_3564);
or U8738 (N_8738,N_3436,N_4977);
nor U8739 (N_8739,N_4257,N_5630);
nand U8740 (N_8740,N_5577,N_3375);
nor U8741 (N_8741,N_3005,N_5048);
and U8742 (N_8742,N_4128,N_5065);
nand U8743 (N_8743,N_4569,N_5039);
and U8744 (N_8744,N_3623,N_3042);
and U8745 (N_8745,N_4646,N_4655);
and U8746 (N_8746,N_3012,N_3582);
nor U8747 (N_8747,N_5845,N_5296);
xnor U8748 (N_8748,N_5577,N_5251);
nor U8749 (N_8749,N_3132,N_4884);
or U8750 (N_8750,N_3302,N_5629);
or U8751 (N_8751,N_5653,N_5955);
or U8752 (N_8752,N_4103,N_3313);
nand U8753 (N_8753,N_5006,N_4679);
or U8754 (N_8754,N_5033,N_3654);
and U8755 (N_8755,N_5339,N_4030);
nand U8756 (N_8756,N_4867,N_3801);
and U8757 (N_8757,N_4664,N_5147);
and U8758 (N_8758,N_4907,N_4539);
nor U8759 (N_8759,N_5078,N_5569);
and U8760 (N_8760,N_5947,N_5557);
or U8761 (N_8761,N_5831,N_4904);
nor U8762 (N_8762,N_3750,N_4224);
nand U8763 (N_8763,N_3786,N_3478);
or U8764 (N_8764,N_4589,N_4944);
nor U8765 (N_8765,N_3213,N_4508);
nor U8766 (N_8766,N_4367,N_5146);
and U8767 (N_8767,N_3715,N_3714);
and U8768 (N_8768,N_4147,N_4796);
nor U8769 (N_8769,N_5368,N_4850);
and U8770 (N_8770,N_3583,N_3993);
xnor U8771 (N_8771,N_4234,N_5840);
or U8772 (N_8772,N_5838,N_3648);
and U8773 (N_8773,N_5436,N_3541);
or U8774 (N_8774,N_4867,N_5474);
or U8775 (N_8775,N_4921,N_3308);
or U8776 (N_8776,N_3316,N_5254);
or U8777 (N_8777,N_3775,N_3293);
nor U8778 (N_8778,N_5526,N_4882);
nand U8779 (N_8779,N_3906,N_5631);
nor U8780 (N_8780,N_5391,N_5817);
nand U8781 (N_8781,N_3886,N_4072);
nor U8782 (N_8782,N_3145,N_5535);
nor U8783 (N_8783,N_5964,N_4495);
nand U8784 (N_8784,N_3824,N_5125);
or U8785 (N_8785,N_3003,N_5504);
and U8786 (N_8786,N_5402,N_5415);
and U8787 (N_8787,N_3093,N_5767);
nor U8788 (N_8788,N_3675,N_4693);
and U8789 (N_8789,N_3621,N_5904);
nand U8790 (N_8790,N_5790,N_3080);
or U8791 (N_8791,N_3981,N_4626);
nor U8792 (N_8792,N_4136,N_3538);
nand U8793 (N_8793,N_4303,N_3388);
nand U8794 (N_8794,N_3798,N_4380);
nand U8795 (N_8795,N_5941,N_3857);
or U8796 (N_8796,N_3882,N_5305);
nand U8797 (N_8797,N_3803,N_4665);
nor U8798 (N_8798,N_4101,N_4023);
or U8799 (N_8799,N_3148,N_3966);
or U8800 (N_8800,N_4375,N_3658);
nor U8801 (N_8801,N_5666,N_3883);
nor U8802 (N_8802,N_4399,N_5483);
or U8803 (N_8803,N_4168,N_4377);
nor U8804 (N_8804,N_3683,N_5876);
xnor U8805 (N_8805,N_4200,N_4030);
and U8806 (N_8806,N_4170,N_5068);
or U8807 (N_8807,N_3896,N_3246);
xnor U8808 (N_8808,N_4137,N_4902);
nor U8809 (N_8809,N_3035,N_4244);
nor U8810 (N_8810,N_3617,N_5612);
nor U8811 (N_8811,N_3447,N_3791);
and U8812 (N_8812,N_3034,N_5508);
nor U8813 (N_8813,N_3289,N_3395);
or U8814 (N_8814,N_3463,N_4405);
nand U8815 (N_8815,N_4902,N_4282);
nor U8816 (N_8816,N_3457,N_3666);
nand U8817 (N_8817,N_3983,N_3648);
and U8818 (N_8818,N_3745,N_5380);
nand U8819 (N_8819,N_3819,N_5438);
and U8820 (N_8820,N_5600,N_5884);
nor U8821 (N_8821,N_3361,N_4160);
nor U8822 (N_8822,N_3197,N_3131);
and U8823 (N_8823,N_4354,N_3387);
or U8824 (N_8824,N_4335,N_4988);
nand U8825 (N_8825,N_5216,N_5024);
or U8826 (N_8826,N_3618,N_4846);
xor U8827 (N_8827,N_4108,N_5472);
nand U8828 (N_8828,N_4171,N_3526);
or U8829 (N_8829,N_3001,N_5091);
or U8830 (N_8830,N_4766,N_4078);
nand U8831 (N_8831,N_4070,N_3770);
nor U8832 (N_8832,N_5152,N_4643);
nor U8833 (N_8833,N_5540,N_4910);
nor U8834 (N_8834,N_5294,N_5809);
nand U8835 (N_8835,N_3902,N_5633);
or U8836 (N_8836,N_5553,N_5673);
nand U8837 (N_8837,N_5498,N_5527);
or U8838 (N_8838,N_3351,N_5432);
and U8839 (N_8839,N_4484,N_5663);
nand U8840 (N_8840,N_3470,N_5969);
or U8841 (N_8841,N_4858,N_4879);
and U8842 (N_8842,N_5184,N_5272);
or U8843 (N_8843,N_4966,N_3685);
or U8844 (N_8844,N_3718,N_3840);
and U8845 (N_8845,N_3657,N_4096);
and U8846 (N_8846,N_3454,N_4268);
or U8847 (N_8847,N_3441,N_4298);
or U8848 (N_8848,N_5207,N_5863);
or U8849 (N_8849,N_3138,N_5893);
or U8850 (N_8850,N_3145,N_3273);
nor U8851 (N_8851,N_4581,N_3384);
or U8852 (N_8852,N_4054,N_4394);
nor U8853 (N_8853,N_3569,N_3325);
xnor U8854 (N_8854,N_5426,N_4175);
and U8855 (N_8855,N_4804,N_5092);
and U8856 (N_8856,N_5990,N_4959);
and U8857 (N_8857,N_4444,N_5475);
and U8858 (N_8858,N_4801,N_5854);
and U8859 (N_8859,N_3399,N_5586);
nor U8860 (N_8860,N_4118,N_4855);
or U8861 (N_8861,N_3259,N_4058);
nand U8862 (N_8862,N_4416,N_3865);
and U8863 (N_8863,N_5624,N_3121);
and U8864 (N_8864,N_5525,N_4608);
and U8865 (N_8865,N_4072,N_5780);
nor U8866 (N_8866,N_4997,N_5808);
nor U8867 (N_8867,N_3382,N_5214);
or U8868 (N_8868,N_4475,N_5001);
and U8869 (N_8869,N_4203,N_3760);
or U8870 (N_8870,N_5431,N_4460);
nor U8871 (N_8871,N_3415,N_3962);
xor U8872 (N_8872,N_4665,N_5707);
nor U8873 (N_8873,N_5075,N_4459);
and U8874 (N_8874,N_4422,N_4139);
and U8875 (N_8875,N_3370,N_5464);
xor U8876 (N_8876,N_5339,N_4587);
or U8877 (N_8877,N_3740,N_3789);
nand U8878 (N_8878,N_4490,N_3291);
and U8879 (N_8879,N_3847,N_4842);
nor U8880 (N_8880,N_4650,N_4711);
nor U8881 (N_8881,N_5777,N_4538);
or U8882 (N_8882,N_4367,N_5559);
or U8883 (N_8883,N_3400,N_4970);
and U8884 (N_8884,N_5947,N_4634);
xnor U8885 (N_8885,N_3109,N_5348);
and U8886 (N_8886,N_3104,N_4707);
and U8887 (N_8887,N_3254,N_3228);
or U8888 (N_8888,N_3792,N_5105);
or U8889 (N_8889,N_4183,N_3684);
and U8890 (N_8890,N_4110,N_5033);
or U8891 (N_8891,N_4752,N_3221);
or U8892 (N_8892,N_5419,N_4390);
and U8893 (N_8893,N_4877,N_3766);
and U8894 (N_8894,N_4913,N_4886);
and U8895 (N_8895,N_5400,N_5997);
or U8896 (N_8896,N_5989,N_5256);
nor U8897 (N_8897,N_5954,N_4263);
nor U8898 (N_8898,N_3268,N_3032);
xor U8899 (N_8899,N_4230,N_5521);
nand U8900 (N_8900,N_5831,N_5452);
nand U8901 (N_8901,N_4416,N_5592);
and U8902 (N_8902,N_3947,N_5860);
or U8903 (N_8903,N_3796,N_3080);
or U8904 (N_8904,N_4741,N_5268);
and U8905 (N_8905,N_5607,N_5316);
nand U8906 (N_8906,N_5058,N_5123);
nor U8907 (N_8907,N_3237,N_4836);
and U8908 (N_8908,N_5240,N_3689);
nand U8909 (N_8909,N_5227,N_3297);
nand U8910 (N_8910,N_5554,N_4136);
nand U8911 (N_8911,N_5423,N_4095);
or U8912 (N_8912,N_4662,N_5360);
nand U8913 (N_8913,N_5327,N_5142);
nor U8914 (N_8914,N_3577,N_4007);
nor U8915 (N_8915,N_3216,N_5513);
or U8916 (N_8916,N_4832,N_4830);
nand U8917 (N_8917,N_3031,N_3572);
or U8918 (N_8918,N_3581,N_3240);
or U8919 (N_8919,N_4745,N_5612);
and U8920 (N_8920,N_4954,N_5569);
nor U8921 (N_8921,N_4061,N_4763);
nand U8922 (N_8922,N_4060,N_5596);
nand U8923 (N_8923,N_3178,N_3025);
nor U8924 (N_8924,N_5212,N_3782);
or U8925 (N_8925,N_3644,N_4650);
nor U8926 (N_8926,N_5946,N_5973);
nor U8927 (N_8927,N_3345,N_4396);
or U8928 (N_8928,N_4060,N_5347);
or U8929 (N_8929,N_5229,N_5679);
or U8930 (N_8930,N_5522,N_5743);
nor U8931 (N_8931,N_3252,N_5594);
and U8932 (N_8932,N_3504,N_3927);
or U8933 (N_8933,N_5441,N_3242);
and U8934 (N_8934,N_5683,N_3301);
or U8935 (N_8935,N_4553,N_3917);
and U8936 (N_8936,N_4418,N_3715);
and U8937 (N_8937,N_4534,N_3623);
nand U8938 (N_8938,N_4725,N_3580);
and U8939 (N_8939,N_5446,N_4381);
and U8940 (N_8940,N_5979,N_5355);
nand U8941 (N_8941,N_4099,N_5660);
or U8942 (N_8942,N_5557,N_4906);
nor U8943 (N_8943,N_4243,N_4046);
or U8944 (N_8944,N_3904,N_5933);
and U8945 (N_8945,N_4468,N_3929);
xor U8946 (N_8946,N_5396,N_5244);
or U8947 (N_8947,N_4429,N_4106);
nor U8948 (N_8948,N_5479,N_4406);
nor U8949 (N_8949,N_5526,N_5908);
xor U8950 (N_8950,N_5978,N_4217);
nor U8951 (N_8951,N_4632,N_5086);
or U8952 (N_8952,N_4561,N_4325);
or U8953 (N_8953,N_5512,N_4383);
nor U8954 (N_8954,N_3884,N_4602);
and U8955 (N_8955,N_5354,N_3080);
or U8956 (N_8956,N_4016,N_4375);
nor U8957 (N_8957,N_3670,N_3411);
and U8958 (N_8958,N_4838,N_4478);
and U8959 (N_8959,N_4117,N_5313);
and U8960 (N_8960,N_3575,N_5708);
nor U8961 (N_8961,N_3644,N_5102);
nor U8962 (N_8962,N_4722,N_4996);
nor U8963 (N_8963,N_3064,N_3309);
or U8964 (N_8964,N_4577,N_5178);
xnor U8965 (N_8965,N_5649,N_3380);
nor U8966 (N_8966,N_5651,N_4944);
and U8967 (N_8967,N_3499,N_4207);
or U8968 (N_8968,N_3983,N_5404);
nand U8969 (N_8969,N_5945,N_3231);
nor U8970 (N_8970,N_3433,N_5141);
and U8971 (N_8971,N_4718,N_3771);
nor U8972 (N_8972,N_3089,N_5709);
or U8973 (N_8973,N_3614,N_4378);
nand U8974 (N_8974,N_3018,N_5551);
and U8975 (N_8975,N_5491,N_5304);
and U8976 (N_8976,N_4098,N_5846);
nor U8977 (N_8977,N_5259,N_3948);
nand U8978 (N_8978,N_4881,N_3169);
nand U8979 (N_8979,N_5090,N_3624);
or U8980 (N_8980,N_5419,N_3329);
and U8981 (N_8981,N_5748,N_4589);
and U8982 (N_8982,N_5623,N_3205);
or U8983 (N_8983,N_3062,N_4861);
and U8984 (N_8984,N_4446,N_3962);
nand U8985 (N_8985,N_5825,N_3872);
nand U8986 (N_8986,N_4237,N_3711);
nor U8987 (N_8987,N_4640,N_5381);
or U8988 (N_8988,N_5761,N_3423);
nor U8989 (N_8989,N_4378,N_5525);
or U8990 (N_8990,N_4980,N_3641);
or U8991 (N_8991,N_5199,N_4320);
and U8992 (N_8992,N_3868,N_3863);
nand U8993 (N_8993,N_4076,N_5966);
nand U8994 (N_8994,N_4207,N_3726);
or U8995 (N_8995,N_4594,N_5355);
nor U8996 (N_8996,N_3336,N_4537);
and U8997 (N_8997,N_4772,N_5630);
nor U8998 (N_8998,N_3499,N_5309);
or U8999 (N_8999,N_3949,N_4005);
and U9000 (N_9000,N_6224,N_6960);
and U9001 (N_9001,N_6728,N_8163);
nand U9002 (N_9002,N_7082,N_7371);
nand U9003 (N_9003,N_6695,N_8662);
nor U9004 (N_9004,N_6019,N_8739);
or U9005 (N_9005,N_8114,N_7592);
nor U9006 (N_9006,N_6394,N_8789);
or U9007 (N_9007,N_8217,N_6788);
and U9008 (N_9008,N_6818,N_7954);
nor U9009 (N_9009,N_6704,N_8246);
or U9010 (N_9010,N_6584,N_8266);
nor U9011 (N_9011,N_8263,N_6845);
nor U9012 (N_9012,N_8132,N_7616);
and U9013 (N_9013,N_6971,N_6794);
nor U9014 (N_9014,N_8883,N_6106);
or U9015 (N_9015,N_8095,N_6445);
or U9016 (N_9016,N_8866,N_7841);
and U9017 (N_9017,N_7631,N_7176);
nand U9018 (N_9018,N_8593,N_8735);
and U9019 (N_9019,N_7614,N_7063);
nand U9020 (N_9020,N_6828,N_8084);
or U9021 (N_9021,N_6824,N_6681);
and U9022 (N_9022,N_6316,N_6650);
and U9023 (N_9023,N_7333,N_6384);
nor U9024 (N_9024,N_7708,N_8365);
or U9025 (N_9025,N_7785,N_8340);
nor U9026 (N_9026,N_7925,N_6878);
or U9027 (N_9027,N_6022,N_7855);
nor U9028 (N_9028,N_6723,N_8526);
and U9029 (N_9029,N_8296,N_8403);
or U9030 (N_9030,N_8947,N_8093);
or U9031 (N_9031,N_8216,N_6899);
nor U9032 (N_9032,N_8142,N_8563);
or U9033 (N_9033,N_7237,N_8642);
nand U9034 (N_9034,N_7951,N_8130);
or U9035 (N_9035,N_6231,N_6443);
nand U9036 (N_9036,N_8439,N_8624);
nor U9037 (N_9037,N_6915,N_6377);
nand U9038 (N_9038,N_7780,N_8301);
or U9039 (N_9039,N_8727,N_6420);
nand U9040 (N_9040,N_6107,N_7573);
nor U9041 (N_9041,N_8887,N_8334);
nor U9042 (N_9042,N_7526,N_8074);
or U9043 (N_9043,N_6171,N_8945);
and U9044 (N_9044,N_6663,N_6177);
or U9045 (N_9045,N_6802,N_7190);
nor U9046 (N_9046,N_8949,N_8755);
nor U9047 (N_9047,N_8523,N_7759);
nor U9048 (N_9048,N_7239,N_7590);
nor U9049 (N_9049,N_6335,N_6843);
or U9050 (N_9050,N_8311,N_7873);
or U9051 (N_9051,N_7390,N_6626);
or U9052 (N_9052,N_6196,N_6905);
or U9053 (N_9053,N_8401,N_6199);
nor U9054 (N_9054,N_8864,N_7400);
xnor U9055 (N_9055,N_7787,N_7555);
nor U9056 (N_9056,N_6880,N_6313);
and U9057 (N_9057,N_6251,N_6396);
nor U9058 (N_9058,N_6853,N_7439);
and U9059 (N_9059,N_8753,N_7516);
nor U9060 (N_9060,N_8503,N_7952);
and U9061 (N_9061,N_7075,N_7721);
or U9062 (N_9062,N_7914,N_7202);
and U9063 (N_9063,N_6083,N_8494);
nand U9064 (N_9064,N_6285,N_7179);
and U9065 (N_9065,N_8536,N_6060);
or U9066 (N_9066,N_7680,N_7323);
nor U9067 (N_9067,N_7344,N_7603);
and U9068 (N_9068,N_7709,N_6413);
nor U9069 (N_9069,N_8912,N_6437);
nand U9070 (N_9070,N_8584,N_7950);
nor U9071 (N_9071,N_7277,N_7711);
or U9072 (N_9072,N_6137,N_6526);
or U9073 (N_9073,N_6797,N_7919);
or U9074 (N_9074,N_6261,N_8324);
or U9075 (N_9075,N_7114,N_7164);
and U9076 (N_9076,N_6616,N_8914);
nand U9077 (N_9077,N_8859,N_6169);
nand U9078 (N_9078,N_6987,N_7593);
nand U9079 (N_9079,N_6266,N_6719);
and U9080 (N_9080,N_6163,N_7405);
nand U9081 (N_9081,N_7985,N_7066);
nor U9082 (N_9082,N_7957,N_6622);
nor U9083 (N_9083,N_7550,N_6154);
nand U9084 (N_9084,N_8653,N_8366);
nand U9085 (N_9085,N_8221,N_7705);
or U9086 (N_9086,N_8414,N_7669);
or U9087 (N_9087,N_7067,N_7662);
or U9088 (N_9088,N_8353,N_7818);
nor U9089 (N_9089,N_7409,N_6844);
nand U9090 (N_9090,N_7672,N_8133);
or U9091 (N_9091,N_8853,N_6480);
nand U9092 (N_9092,N_7111,N_8666);
nand U9093 (N_9093,N_6867,N_7180);
or U9094 (N_9094,N_7304,N_6564);
and U9095 (N_9095,N_7949,N_6332);
or U9096 (N_9096,N_6061,N_6014);
nand U9097 (N_9097,N_8119,N_8239);
nand U9098 (N_9098,N_6576,N_6215);
and U9099 (N_9099,N_7487,N_8533);
and U9100 (N_9100,N_8919,N_8260);
nand U9101 (N_9101,N_8996,N_8169);
nand U9102 (N_9102,N_7702,N_8736);
xnor U9103 (N_9103,N_6525,N_6054);
nor U9104 (N_9104,N_8601,N_7094);
and U9105 (N_9105,N_8551,N_8514);
nor U9106 (N_9106,N_8223,N_7447);
nand U9107 (N_9107,N_7585,N_6995);
or U9108 (N_9108,N_7558,N_8137);
nand U9109 (N_9109,N_8147,N_8718);
xnor U9110 (N_9110,N_6263,N_7161);
or U9111 (N_9111,N_8261,N_6005);
or U9112 (N_9112,N_7532,N_7448);
and U9113 (N_9113,N_6479,N_7838);
nand U9114 (N_9114,N_7184,N_6382);
nand U9115 (N_9115,N_6557,N_6084);
or U9116 (N_9116,N_7658,N_6258);
nor U9117 (N_9117,N_6833,N_6721);
nand U9118 (N_9118,N_7046,N_6448);
nor U9119 (N_9119,N_7499,N_7695);
or U9120 (N_9120,N_6068,N_7188);
nand U9121 (N_9121,N_7820,N_8562);
and U9122 (N_9122,N_8175,N_6112);
or U9123 (N_9123,N_6315,N_7617);
or U9124 (N_9124,N_7621,N_6239);
or U9125 (N_9125,N_7494,N_7921);
nor U9126 (N_9126,N_6996,N_7481);
or U9127 (N_9127,N_7979,N_7297);
nand U9128 (N_9128,N_6892,N_8259);
nor U9129 (N_9129,N_7647,N_7264);
nor U9130 (N_9130,N_7927,N_8795);
nand U9131 (N_9131,N_6194,N_7163);
nor U9132 (N_9132,N_8884,N_6827);
nor U9133 (N_9133,N_8612,N_8599);
nand U9134 (N_9134,N_8959,N_8253);
nand U9135 (N_9135,N_6410,N_6111);
nand U9136 (N_9136,N_6545,N_6896);
nor U9137 (N_9137,N_8297,N_6297);
nand U9138 (N_9138,N_7977,N_7551);
and U9139 (N_9139,N_8452,N_7227);
nor U9140 (N_9140,N_8846,N_8487);
nor U9141 (N_9141,N_7899,N_8897);
nor U9142 (N_9142,N_8083,N_6729);
and U9143 (N_9143,N_8966,N_7769);
or U9144 (N_9144,N_7366,N_6730);
or U9145 (N_9145,N_8882,N_6539);
or U9146 (N_9146,N_6366,N_6898);
or U9147 (N_9147,N_7750,N_7113);
and U9148 (N_9148,N_7529,N_8788);
or U9149 (N_9149,N_7057,N_6524);
nor U9150 (N_9150,N_7348,N_8112);
or U9151 (N_9151,N_8549,N_6734);
or U9152 (N_9152,N_7345,N_8158);
or U9153 (N_9153,N_6162,N_8557);
xnor U9154 (N_9154,N_7588,N_8328);
nor U9155 (N_9155,N_7497,N_7714);
nand U9156 (N_9156,N_7607,N_8717);
nor U9157 (N_9157,N_8387,N_6758);
nand U9158 (N_9158,N_6087,N_6010);
nor U9159 (N_9159,N_7303,N_8850);
and U9160 (N_9160,N_8474,N_6974);
nand U9161 (N_9161,N_6837,N_7086);
or U9162 (N_9162,N_8757,N_8467);
and U9163 (N_9163,N_7410,N_7650);
nand U9164 (N_9164,N_8973,N_8363);
nand U9165 (N_9165,N_7801,N_8235);
nand U9166 (N_9166,N_6592,N_7065);
or U9167 (N_9167,N_6433,N_6213);
nor U9168 (N_9168,N_7562,N_8942);
nor U9169 (N_9169,N_8819,N_8111);
nor U9170 (N_9170,N_8288,N_8045);
and U9171 (N_9171,N_8576,N_8320);
nand U9172 (N_9172,N_7779,N_8185);
nand U9173 (N_9173,N_8779,N_7471);
or U9174 (N_9174,N_8139,N_6685);
nor U9175 (N_9175,N_6930,N_6478);
and U9176 (N_9176,N_7236,N_7147);
nor U9177 (N_9177,N_8929,N_8486);
nor U9178 (N_9178,N_7579,N_6630);
nand U9179 (N_9179,N_8034,N_6036);
or U9180 (N_9180,N_6246,N_7133);
nand U9181 (N_9181,N_6295,N_6588);
and U9182 (N_9182,N_6511,N_6652);
or U9183 (N_9183,N_6429,N_7538);
and U9184 (N_9184,N_8390,N_7268);
nor U9185 (N_9185,N_7634,N_7467);
nand U9186 (N_9186,N_6482,N_6464);
nand U9187 (N_9187,N_7933,N_6383);
or U9188 (N_9188,N_6737,N_7309);
or U9189 (N_9189,N_6970,N_8831);
nor U9190 (N_9190,N_7301,N_6795);
or U9191 (N_9191,N_6606,N_7070);
and U9192 (N_9192,N_6773,N_8454);
xnor U9193 (N_9193,N_6900,N_8247);
nor U9194 (N_9194,N_8315,N_8548);
nor U9195 (N_9195,N_8575,N_8763);
and U9196 (N_9196,N_6381,N_7477);
nand U9197 (N_9197,N_7924,N_6161);
nor U9198 (N_9198,N_8141,N_8432);
nor U9199 (N_9199,N_6854,N_7139);
nor U9200 (N_9200,N_6406,N_8103);
or U9201 (N_9201,N_8917,N_8607);
and U9202 (N_9202,N_8955,N_6253);
and U9203 (N_9203,N_8994,N_6062);
nor U9204 (N_9204,N_8314,N_6514);
and U9205 (N_9205,N_7817,N_6236);
and U9206 (N_9206,N_6641,N_7545);
and U9207 (N_9207,N_8344,N_6747);
and U9208 (N_9208,N_8146,N_8109);
and U9209 (N_9209,N_8043,N_8295);
xnor U9210 (N_9210,N_7974,N_8032);
or U9211 (N_9211,N_7503,N_6736);
or U9212 (N_9212,N_6400,N_8637);
nor U9213 (N_9213,N_6189,N_7570);
and U9214 (N_9214,N_8096,N_7712);
and U9215 (N_9215,N_7845,N_8944);
and U9216 (N_9216,N_6097,N_6959);
nor U9217 (N_9217,N_7868,N_8989);
nor U9218 (N_9218,N_6264,N_8086);
or U9219 (N_9219,N_8342,N_6373);
nor U9220 (N_9220,N_7866,N_7491);
or U9221 (N_9221,N_6484,N_7247);
or U9222 (N_9222,N_7825,N_7044);
and U9223 (N_9223,N_7001,N_8823);
or U9224 (N_9224,N_8206,N_7681);
and U9225 (N_9225,N_8335,N_6726);
nand U9226 (N_9226,N_6847,N_6368);
nor U9227 (N_9227,N_7772,N_7493);
nor U9228 (N_9228,N_6697,N_6459);
and U9229 (N_9229,N_7521,N_6079);
nand U9230 (N_9230,N_8911,N_7857);
and U9231 (N_9231,N_8535,N_6549);
and U9232 (N_9232,N_6160,N_7058);
nand U9233 (N_9233,N_8750,N_7666);
or U9234 (N_9234,N_7024,N_8257);
or U9235 (N_9235,N_8286,N_7288);
nand U9236 (N_9236,N_6846,N_7609);
and U9237 (N_9237,N_6598,N_6956);
nor U9238 (N_9238,N_7246,N_6658);
nor U9239 (N_9239,N_6753,N_7232);
or U9240 (N_9240,N_6746,N_6341);
nand U9241 (N_9241,N_6931,N_7639);
nand U9242 (N_9242,N_6318,N_6080);
nor U9243 (N_9243,N_7451,N_6447);
nand U9244 (N_9244,N_7733,N_6894);
nor U9245 (N_9245,N_6862,N_6345);
or U9246 (N_9246,N_8628,N_8180);
and U9247 (N_9247,N_8918,N_8079);
and U9248 (N_9248,N_6180,N_8786);
or U9249 (N_9249,N_7945,N_6041);
or U9250 (N_9250,N_7210,N_8571);
and U9251 (N_9251,N_8588,N_6259);
or U9252 (N_9252,N_8946,N_8409);
nor U9253 (N_9253,N_7206,N_7367);
or U9254 (N_9254,N_8159,N_8578);
nor U9255 (N_9255,N_7427,N_6967);
or U9256 (N_9256,N_7031,N_7221);
or U9257 (N_9257,N_8378,N_7556);
nand U9258 (N_9258,N_8639,N_7363);
and U9259 (N_9259,N_6324,N_6975);
nand U9260 (N_9260,N_6248,N_7698);
nand U9261 (N_9261,N_6372,N_7402);
and U9262 (N_9262,N_8025,N_6586);
nand U9263 (N_9263,N_8962,N_7765);
or U9264 (N_9264,N_8027,N_7986);
or U9265 (N_9265,N_7145,N_7880);
nand U9266 (N_9266,N_8954,N_6489);
nor U9267 (N_9267,N_7696,N_8981);
nor U9268 (N_9268,N_7960,N_7310);
nand U9269 (N_9269,N_7370,N_7198);
and U9270 (N_9270,N_7858,N_8650);
nand U9271 (N_9271,N_7178,N_8631);
and U9272 (N_9272,N_7170,N_6538);
nor U9273 (N_9273,N_6195,N_6810);
or U9274 (N_9274,N_6601,N_6895);
nand U9275 (N_9275,N_8670,N_7575);
nor U9276 (N_9276,N_6294,N_6317);
or U9277 (N_9277,N_7385,N_7963);
and U9278 (N_9278,N_8985,N_8657);
nand U9279 (N_9279,N_8177,N_8117);
nor U9280 (N_9280,N_7265,N_6289);
and U9281 (N_9281,N_7411,N_8292);
and U9282 (N_9282,N_8800,N_6943);
nor U9283 (N_9283,N_8188,N_8207);
and U9284 (N_9284,N_7229,N_8550);
nand U9285 (N_9285,N_7416,N_6809);
and U9286 (N_9286,N_7886,N_7527);
and U9287 (N_9287,N_7745,N_8015);
or U9288 (N_9288,N_8497,N_7946);
and U9289 (N_9289,N_6278,N_7701);
and U9290 (N_9290,N_6541,N_6490);
nand U9291 (N_9291,N_7119,N_8215);
or U9292 (N_9292,N_8513,N_6211);
and U9293 (N_9293,N_8965,N_6002);
or U9294 (N_9294,N_6638,N_6371);
and U9295 (N_9295,N_8026,N_7814);
nand U9296 (N_9296,N_7052,N_6945);
and U9297 (N_9297,N_7054,N_7916);
nor U9298 (N_9298,N_7665,N_6806);
nor U9299 (N_9299,N_8473,N_6679);
or U9300 (N_9300,N_8270,N_6268);
and U9301 (N_9301,N_8374,N_6825);
and U9302 (N_9302,N_6692,N_7177);
nand U9303 (N_9303,N_6811,N_8341);
nor U9304 (N_9304,N_6424,N_7428);
xnor U9305 (N_9305,N_8357,N_7536);
or U9306 (N_9306,N_7727,N_8860);
or U9307 (N_9307,N_8614,N_6861);
nor U9308 (N_9308,N_7498,N_8977);
and U9309 (N_9309,N_7822,N_8429);
xor U9310 (N_9310,N_7824,N_6548);
nand U9311 (N_9311,N_6343,N_8995);
and U9312 (N_9312,N_7235,N_6113);
nor U9313 (N_9313,N_6555,N_8056);
nand U9314 (N_9314,N_6863,N_6997);
and U9315 (N_9315,N_8245,N_7261);
nand U9316 (N_9316,N_7267,N_6375);
or U9317 (N_9317,N_7900,N_8988);
nor U9318 (N_9318,N_8048,N_8097);
nand U9319 (N_9319,N_7329,N_6059);
nor U9320 (N_9320,N_8833,N_7468);
and U9321 (N_9321,N_7327,N_8160);
nand U9322 (N_9322,N_7738,N_8230);
and U9323 (N_9323,N_6741,N_7112);
and U9324 (N_9324,N_6094,N_8101);
or U9325 (N_9325,N_6156,N_7852);
nor U9326 (N_9326,N_7150,N_6599);
and U9327 (N_9327,N_7968,N_6166);
nand U9328 (N_9328,N_6076,N_6286);
or U9329 (N_9329,N_7160,N_7656);
nand U9330 (N_9330,N_8665,N_8476);
nand U9331 (N_9331,N_8053,N_6201);
nand U9332 (N_9332,N_8457,N_8505);
nand U9333 (N_9333,N_8827,N_8771);
nand U9334 (N_9334,N_7175,N_6583);
or U9335 (N_9335,N_8219,N_6503);
and U9336 (N_9336,N_8225,N_7138);
and U9337 (N_9337,N_8004,N_8123);
xnor U9338 (N_9338,N_8325,N_6690);
or U9339 (N_9339,N_7223,N_6873);
and U9340 (N_9340,N_7988,N_7689);
nand U9341 (N_9341,N_6153,N_6104);
or U9342 (N_9342,N_8317,N_6150);
or U9343 (N_9343,N_6762,N_7287);
nand U9344 (N_9344,N_7445,N_6941);
nor U9345 (N_9345,N_7687,N_6405);
nand U9346 (N_9346,N_6040,N_6509);
or U9347 (N_9347,N_7074,N_8552);
or U9348 (N_9348,N_8029,N_6354);
nor U9349 (N_9349,N_8104,N_6561);
xnor U9350 (N_9350,N_8150,N_8449);
nor U9351 (N_9351,N_7426,N_8323);
nand U9352 (N_9352,N_8222,N_7980);
nand U9353 (N_9353,N_8404,N_6563);
nand U9354 (N_9354,N_7599,N_7399);
or U9355 (N_9355,N_6227,N_8463);
and U9356 (N_9356,N_8902,N_8051);
and U9357 (N_9357,N_6738,N_7002);
nor U9358 (N_9358,N_7196,N_8300);
nand U9359 (N_9359,N_6954,N_8226);
nor U9360 (N_9360,N_6742,N_8131);
nand U9361 (N_9361,N_8560,N_6401);
and U9362 (N_9362,N_6200,N_6502);
nor U9363 (N_9363,N_7099,N_8716);
and U9364 (N_9364,N_7574,N_7781);
nand U9365 (N_9365,N_8767,N_8544);
or U9366 (N_9366,N_7864,N_8368);
or U9367 (N_9367,N_7620,N_7887);
nand U9368 (N_9368,N_6929,N_6703);
or U9369 (N_9369,N_7697,N_7011);
and U9370 (N_9370,N_8021,N_6757);
and U9371 (N_9371,N_8237,N_7104);
nor U9372 (N_9372,N_8836,N_8367);
nor U9373 (N_9373,N_6216,N_6387);
nor U9374 (N_9374,N_6000,N_6591);
nand U9375 (N_9375,N_6691,N_7397);
or U9376 (N_9376,N_7973,N_8168);
nand U9377 (N_9377,N_8684,N_8790);
nor U9378 (N_9378,N_8446,N_6290);
nor U9379 (N_9379,N_7537,N_7379);
nor U9380 (N_9380,N_8932,N_7630);
or U9381 (N_9381,N_8754,N_8814);
and U9382 (N_9382,N_7463,N_8172);
and U9383 (N_9383,N_8891,N_7542);
nand U9384 (N_9384,N_7566,N_6888);
or U9385 (N_9385,N_6675,N_7600);
and U9386 (N_9386,N_6309,N_6336);
and U9387 (N_9387,N_7207,N_6562);
nand U9388 (N_9388,N_7719,N_6992);
nand U9389 (N_9389,N_6501,N_8766);
and U9390 (N_9390,N_6352,N_6980);
nand U9391 (N_9391,N_6467,N_6735);
nand U9392 (N_9392,N_8338,N_7107);
or U9393 (N_9393,N_6958,N_8153);
or U9394 (N_9394,N_6799,N_7464);
nand U9395 (N_9395,N_8213,N_7441);
nand U9396 (N_9396,N_7580,N_8254);
or U9397 (N_9397,N_7668,N_7736);
or U9398 (N_9398,N_8375,N_8746);
nand U9399 (N_9399,N_6395,N_7152);
nor U9400 (N_9400,N_7275,N_8858);
and U9401 (N_9401,N_6225,N_7671);
nor U9402 (N_9402,N_7096,N_7116);
nor U9403 (N_9403,N_8835,N_8256);
nor U9404 (N_9404,N_7211,N_7897);
or U9405 (N_9405,N_6287,N_7314);
nor U9406 (N_9406,N_6311,N_8499);
or U9407 (N_9407,N_7203,N_6350);
nor U9408 (N_9408,N_7611,N_7645);
and U9409 (N_9409,N_6934,N_7141);
nor U9410 (N_9410,N_8577,N_7742);
and U9411 (N_9411,N_6632,N_8354);
or U9412 (N_9412,N_8129,N_8033);
nor U9413 (N_9413,N_7557,N_8435);
and U9414 (N_9414,N_6303,N_8890);
nor U9415 (N_9415,N_7773,N_8616);
nor U9416 (N_9416,N_8915,N_8922);
or U9417 (N_9417,N_8234,N_6771);
and U9418 (N_9418,N_8258,N_7437);
nor U9419 (N_9419,N_8622,N_8098);
or U9420 (N_9420,N_6914,N_7515);
and U9421 (N_9421,N_8303,N_6506);
or U9422 (N_9422,N_7561,N_7601);
or U9423 (N_9423,N_6582,N_8149);
nor U9424 (N_9424,N_6038,N_8347);
nor U9425 (N_9425,N_7789,N_7757);
or U9426 (N_9426,N_8379,N_7081);
nand U9427 (N_9427,N_6370,N_8661);
and U9428 (N_9428,N_8880,N_8519);
or U9429 (N_9429,N_8595,N_8924);
and U9430 (N_9430,N_7512,N_8971);
nor U9431 (N_9431,N_7392,N_6450);
nand U9432 (N_9432,N_6380,N_7089);
and U9433 (N_9433,N_8696,N_8688);
or U9434 (N_9434,N_8695,N_8730);
nand U9435 (N_9435,N_6705,N_7528);
nor U9436 (N_9436,N_6714,N_6711);
or U9437 (N_9437,N_7241,N_8035);
nor U9438 (N_9438,N_8957,N_7364);
and U9439 (N_9439,N_7318,N_6026);
and U9440 (N_9440,N_7792,N_8385);
nor U9441 (N_9441,N_7505,N_6209);
nor U9442 (N_9442,N_6190,N_6042);
or U9443 (N_9443,N_8774,N_6296);
and U9444 (N_9444,N_8876,N_8849);
nand U9445 (N_9445,N_8009,N_7384);
nand U9446 (N_9446,N_7490,N_6300);
and U9447 (N_9447,N_6020,N_7679);
nor U9448 (N_9448,N_6487,N_6351);
and U9449 (N_9449,N_8841,N_7568);
nand U9450 (N_9450,N_6222,N_7930);
nand U9451 (N_9451,N_6206,N_7474);
or U9452 (N_9452,N_7425,N_7090);
or U9453 (N_9453,N_6120,N_7540);
nor U9454 (N_9454,N_6881,N_6666);
or U9455 (N_9455,N_7903,N_7577);
nand U9456 (N_9456,N_8472,N_6385);
nand U9457 (N_9457,N_8113,N_8214);
nor U9458 (N_9458,N_8444,N_8412);
nand U9459 (N_9459,N_7098,N_7084);
and U9460 (N_9460,N_8527,N_6938);
nor U9461 (N_9461,N_8842,N_7791);
and U9462 (N_9462,N_6440,N_8815);
nand U9463 (N_9463,N_8667,N_7943);
nand U9464 (N_9464,N_8050,N_6340);
nand U9465 (N_9465,N_7151,N_7643);
nand U9466 (N_9466,N_8834,N_6707);
nor U9467 (N_9467,N_8413,N_6173);
or U9468 (N_9468,N_7683,N_8676);
or U9469 (N_9469,N_7890,N_8282);
or U9470 (N_9470,N_8244,N_6720);
nor U9471 (N_9471,N_6271,N_6640);
and U9472 (N_9472,N_6800,N_7989);
or U9473 (N_9473,N_7118,N_8272);
or U9474 (N_9474,N_8729,N_8677);
nor U9475 (N_9475,N_7723,N_8006);
and U9476 (N_9476,N_8556,N_6320);
xor U9477 (N_9477,N_7522,N_7894);
nor U9478 (N_9478,N_7189,N_6789);
and U9479 (N_9479,N_8298,N_8904);
and U9480 (N_9480,N_7806,N_7608);
nor U9481 (N_9481,N_8496,N_8408);
and U9482 (N_9482,N_7173,N_8152);
nor U9483 (N_9483,N_6530,N_8352);
or U9484 (N_9484,N_7438,N_7535);
or U9485 (N_9485,N_6404,N_8801);
xnor U9486 (N_9486,N_6550,N_7828);
and U9487 (N_9487,N_7317,N_7214);
and U9488 (N_9488,N_6515,N_6617);
or U9489 (N_9489,N_8309,N_6593);
and U9490 (N_9490,N_6057,N_6744);
nand U9491 (N_9491,N_7569,N_6536);
xor U9492 (N_9492,N_6330,N_8743);
nand U9493 (N_9493,N_7225,N_8656);
or U9494 (N_9494,N_6835,N_6198);
nor U9495 (N_9495,N_8627,N_6454);
and U9496 (N_9496,N_6883,N_8632);
or U9497 (N_9497,N_6091,N_8406);
nor U9498 (N_9498,N_8640,N_7155);
nand U9499 (N_9499,N_7910,N_8212);
nor U9500 (N_9500,N_7250,N_8469);
or U9501 (N_9501,N_7774,N_8276);
or U9502 (N_9502,N_6684,N_6152);
nor U9503 (N_9503,N_7393,N_8313);
nor U9504 (N_9504,N_7230,N_7606);
nand U9505 (N_9505,N_6291,N_6043);
or U9506 (N_9506,N_6944,N_7166);
nand U9507 (N_9507,N_8384,N_6571);
or U9508 (N_9508,N_8377,N_7935);
nor U9509 (N_9509,N_6241,N_6155);
xnor U9510 (N_9510,N_7020,N_8392);
or U9511 (N_9511,N_6446,N_8895);
and U9512 (N_9512,N_7144,N_6612);
or U9513 (N_9513,N_8605,N_7129);
nand U9514 (N_9514,N_6783,N_6942);
or U9515 (N_9515,N_8787,N_7101);
nor U9516 (N_9516,N_8304,N_7183);
nor U9517 (N_9517,N_6618,N_6791);
and U9518 (N_9518,N_6966,N_6939);
nor U9519 (N_9519,N_6635,N_6803);
nand U9520 (N_9520,N_8450,N_6782);
or U9521 (N_9521,N_7953,N_7355);
nand U9522 (N_9522,N_7245,N_6553);
nand U9523 (N_9523,N_7055,N_6693);
or U9524 (N_9524,N_7661,N_6304);
or U9525 (N_9525,N_6532,N_7293);
or U9526 (N_9526,N_8005,N_6463);
or U9527 (N_9527,N_7934,N_8638);
or U9528 (N_9528,N_6269,N_6814);
nor U9529 (N_9529,N_7469,N_6776);
nor U9530 (N_9530,N_8003,N_8738);
nor U9531 (N_9531,N_8862,N_6767);
or U9532 (N_9532,N_6924,N_7324);
and U9533 (N_9533,N_8658,N_6860);
and U9534 (N_9534,N_8426,N_6476);
nor U9535 (N_9535,N_6416,N_7888);
and U9536 (N_9536,N_7716,N_6141);
and U9537 (N_9537,N_7395,N_6441);
nand U9538 (N_9538,N_6497,N_8979);
xnor U9539 (N_9539,N_6007,N_7169);
nor U9540 (N_9540,N_8067,N_6994);
nand U9541 (N_9541,N_7710,N_8916);
nor U9542 (N_9542,N_7386,N_8249);
nor U9543 (N_9543,N_6469,N_7812);
nor U9544 (N_9544,N_8105,N_8306);
or U9545 (N_9545,N_7137,N_7430);
and U9546 (N_9546,N_7215,N_6713);
and U9547 (N_9547,N_6848,N_6217);
or U9548 (N_9548,N_6534,N_6378);
or U9549 (N_9549,N_6918,N_7322);
nor U9550 (N_9550,N_7415,N_8453);
and U9551 (N_9551,N_8542,N_6969);
or U9552 (N_9552,N_8232,N_6024);
or U9553 (N_9553,N_8565,N_7388);
and U9554 (N_9554,N_6281,N_7642);
or U9555 (N_9555,N_8329,N_8719);
nor U9556 (N_9556,N_6388,N_7492);
nor U9557 (N_9557,N_6911,N_8706);
or U9558 (N_9558,N_8993,N_6893);
nor U9559 (N_9559,N_7008,N_8809);
or U9560 (N_9560,N_6698,N_6781);
nor U9561 (N_9561,N_6367,N_6573);
nand U9562 (N_9562,N_6552,N_8570);
or U9563 (N_9563,N_6168,N_8748);
nor U9564 (N_9564,N_7457,N_6882);
nor U9565 (N_9565,N_8307,N_8761);
and U9566 (N_9566,N_7511,N_6500);
or U9567 (N_9567,N_8115,N_6653);
nand U9568 (N_9568,N_6518,N_6499);
nor U9569 (N_9569,N_8961,N_8393);
nand U9570 (N_9570,N_6537,N_7793);
nor U9571 (N_9571,N_6355,N_7305);
or U9572 (N_9572,N_6566,N_6119);
or U9573 (N_9573,N_8346,N_7117);
or U9574 (N_9574,N_7290,N_7559);
nand U9575 (N_9575,N_6103,N_7100);
nand U9576 (N_9576,N_8875,N_7359);
xor U9577 (N_9577,N_7092,N_8553);
or U9578 (N_9578,N_6829,N_6282);
or U9579 (N_9579,N_6973,N_7983);
or U9580 (N_9580,N_8660,N_6871);
and U9581 (N_9581,N_8173,N_8921);
or U9582 (N_9582,N_6667,N_6035);
nand U9583 (N_9583,N_6504,N_6749);
nor U9584 (N_9584,N_6780,N_6718);
and U9585 (N_9585,N_7961,N_8590);
xor U9586 (N_9586,N_6648,N_6957);
or U9587 (N_9587,N_6556,N_6984);
nand U9588 (N_9588,N_8187,N_6838);
or U9589 (N_9589,N_7640,N_8524);
nor U9590 (N_9590,N_7744,N_6976);
nor U9591 (N_9591,N_6594,N_6977);
or U9592 (N_9592,N_7984,N_6046);
or U9593 (N_9593,N_7032,N_7051);
nor U9594 (N_9594,N_7720,N_7670);
or U9595 (N_9595,N_8863,N_8410);
nand U9596 (N_9596,N_6369,N_7784);
and U9597 (N_9597,N_7495,N_6347);
nor U9598 (N_9598,N_6620,N_8305);
and U9599 (N_9599,N_7717,N_7105);
and U9600 (N_9600,N_6540,N_6739);
nand U9601 (N_9601,N_8279,N_8539);
or U9602 (N_9602,N_7678,N_7216);
nand U9603 (N_9603,N_8913,N_8343);
nand U9604 (N_9604,N_7636,N_7990);
nor U9605 (N_9605,N_7586,N_6856);
nor U9606 (N_9606,N_8830,N_7480);
nand U9607 (N_9607,N_8415,N_8471);
nand U9608 (N_9608,N_7097,N_6875);
and U9609 (N_9609,N_7076,N_6218);
nand U9610 (N_9610,N_6004,N_8196);
nor U9611 (N_9611,N_6136,N_7053);
nor U9612 (N_9612,N_6823,N_7015);
nand U9613 (N_9613,N_7830,N_7767);
xor U9614 (N_9614,N_7021,N_7786);
or U9615 (N_9615,N_6634,N_7892);
nor U9616 (N_9616,N_6172,N_6132);
nand U9617 (N_9617,N_7604,N_8278);
nand U9618 (N_9618,N_6696,N_7654);
nand U9619 (N_9619,N_6358,N_8762);
or U9620 (N_9620,N_7509,N_6242);
and U9621 (N_9621,N_8070,N_6292);
nand U9622 (N_9622,N_8580,N_7417);
nor U9623 (N_9623,N_8844,N_6078);
nand U9624 (N_9624,N_7143,N_8047);
nor U9625 (N_9625,N_6146,N_6508);
nand U9626 (N_9626,N_8908,N_7724);
nor U9627 (N_9627,N_8990,N_7340);
or U9628 (N_9628,N_8610,N_7404);
nand U9629 (N_9629,N_8419,N_6466);
or U9630 (N_9630,N_6874,N_6774);
nand U9631 (N_9631,N_7077,N_6595);
nand U9632 (N_9632,N_6962,N_6683);
or U9633 (N_9633,N_6435,N_7186);
and U9634 (N_9634,N_8978,N_8772);
nor U9635 (N_9635,N_7228,N_8655);
or U9636 (N_9636,N_8975,N_8816);
nand U9637 (N_9637,N_6901,N_6661);
and U9638 (N_9638,N_6334,N_7270);
nand U9639 (N_9639,N_7664,N_8448);
nor U9640 (N_9640,N_7123,N_8933);
nand U9641 (N_9641,N_6775,N_7289);
or U9642 (N_9642,N_8195,N_7591);
nor U9643 (N_9643,N_7486,N_6625);
or U9644 (N_9644,N_6245,N_6948);
nand U9645 (N_9645,N_7976,N_6143);
nor U9646 (N_9646,N_7826,N_7244);
nand U9647 (N_9647,N_7504,N_6968);
or U9648 (N_9648,N_7014,N_8495);
and U9649 (N_9649,N_8792,N_6338);
and U9650 (N_9650,N_7254,N_7741);
or U9651 (N_9651,N_8956,N_8479);
and U9652 (N_9652,N_7859,N_6008);
or U9653 (N_9653,N_7939,N_6805);
nor U9654 (N_9654,N_8512,N_6165);
and U9655 (N_9655,N_7284,N_7506);
nand U9656 (N_9656,N_7917,N_7135);
nand U9657 (N_9657,N_8361,N_6305);
or U9658 (N_9658,N_8941,N_7839);
or U9659 (N_9659,N_7648,N_8869);
nand U9660 (N_9660,N_7338,N_8681);
nand U9661 (N_9661,N_8316,N_8905);
nor U9662 (N_9662,N_7583,N_8066);
nor U9663 (N_9663,N_6830,N_7737);
nor U9664 (N_9664,N_7320,N_6486);
or U9665 (N_9665,N_6275,N_7258);
or U9666 (N_9666,N_6072,N_7902);
or U9667 (N_9667,N_7154,N_7998);
nand U9668 (N_9668,N_8583,N_6682);
nor U9669 (N_9669,N_8573,N_8332);
and U9670 (N_9670,N_7534,N_8075);
and U9671 (N_9671,N_6769,N_8804);
or U9672 (N_9672,N_8466,N_7209);
nand U9673 (N_9673,N_8720,N_6284);
and U9674 (N_9674,N_7629,N_7004);
and U9675 (N_9675,N_6151,N_8651);
nand U9676 (N_9676,N_8355,N_7992);
nand U9677 (N_9677,N_8714,N_6578);
and U9678 (N_9678,N_7704,N_7408);
or U9679 (N_9679,N_7731,N_8724);
or U9680 (N_9680,N_7009,N_6523);
nand U9681 (N_9681,N_6114,N_7638);
and U9682 (N_9682,N_7282,N_7374);
and U9683 (N_9683,N_7013,N_8373);
nand U9684 (N_9684,N_7248,N_7418);
and U9685 (N_9685,N_8420,N_8485);
and U9686 (N_9686,N_8868,N_6786);
nor U9687 (N_9687,N_8893,N_6614);
nand U9688 (N_9688,N_6471,N_8889);
or U9689 (N_9689,N_7587,N_6922);
nand U9690 (N_9690,N_6346,N_6058);
and U9691 (N_9691,N_6483,N_7810);
nor U9692 (N_9692,N_6765,N_6928);
or U9693 (N_9693,N_6505,N_8591);
or U9694 (N_9694,N_6770,N_6865);
nand U9695 (N_9695,N_7676,N_8024);
and U9696 (N_9696,N_7429,N_7913);
and U9697 (N_9697,N_7667,N_7473);
and U9698 (N_9698,N_7078,N_8702);
nor U9699 (N_9699,N_7802,N_7308);
or U9700 (N_9700,N_8421,N_6003);
or U9701 (N_9701,N_7722,N_6221);
and U9702 (N_9702,N_7804,N_6917);
nand U9703 (N_9703,N_7928,N_6025);
or U9704 (N_9704,N_7931,N_8872);
and U9705 (N_9705,N_7028,N_7901);
and U9706 (N_9706,N_6023,N_7612);
xor U9707 (N_9707,N_7131,N_7860);
and U9708 (N_9708,N_8001,N_6621);
xnor U9709 (N_9709,N_7103,N_8707);
nor U9710 (N_9710,N_7728,N_8663);
or U9711 (N_9711,N_6034,N_7233);
and U9712 (N_9712,N_6686,N_8443);
nand U9713 (N_9713,N_8794,N_7337);
or U9714 (N_9714,N_8822,N_6531);
nand U9715 (N_9715,N_8156,N_8768);
and U9716 (N_9716,N_7549,N_6325);
xnor U9717 (N_9717,N_8821,N_7517);
nor U9718 (N_9718,N_6891,N_6302);
or U9719 (N_9719,N_7546,N_6270);
and U9720 (N_9720,N_7867,N_7905);
and U9721 (N_9721,N_8268,N_8972);
or U9722 (N_9722,N_8077,N_8685);
nor U9723 (N_9723,N_8515,N_7747);
or U9724 (N_9724,N_8782,N_8725);
nor U9725 (N_9725,N_8014,N_6529);
or U9726 (N_9726,N_6455,N_6589);
or U9727 (N_9727,N_7342,N_6585);
nor U9728 (N_9728,N_6575,N_8134);
nor U9729 (N_9729,N_8783,N_6596);
and U9730 (N_9730,N_6779,N_8319);
nand U9731 (N_9731,N_8991,N_8934);
or U9732 (N_9732,N_8732,N_7523);
or U9733 (N_9733,N_7302,N_6752);
nor U9734 (N_9734,N_8100,N_6086);
nand U9735 (N_9735,N_7414,N_7041);
and U9736 (N_9736,N_6065,N_7413);
and U9737 (N_9737,N_7891,N_8274);
and U9738 (N_9738,N_7513,N_6554);
nor U9739 (N_9739,N_7729,N_7657);
or U9740 (N_9740,N_6237,N_6460);
nand U9741 (N_9741,N_8262,N_8178);
and U9742 (N_9742,N_8857,N_6755);
nor U9743 (N_9743,N_6207,N_8348);
or U9744 (N_9744,N_8721,N_7039);
or U9745 (N_9745,N_8491,N_6133);
and U9746 (N_9746,N_6559,N_6050);
and U9747 (N_9747,N_6725,N_8776);
and U9748 (N_9748,N_8273,N_6045);
nor U9749 (N_9749,N_8484,N_6337);
nor U9750 (N_9750,N_8418,N_8252);
nand U9751 (N_9751,N_6826,N_7751);
nand U9752 (N_9752,N_7663,N_6952);
or U9753 (N_9753,N_8509,N_8224);
nor U9754 (N_9754,N_8986,N_6602);
nand U9755 (N_9755,N_8135,N_8892);
or U9756 (N_9756,N_8856,N_6047);
nor U9757 (N_9757,N_8510,N_6993);
or U9758 (N_9758,N_6465,N_6067);
nor U9759 (N_9759,N_8770,N_7313);
or U9760 (N_9760,N_6633,N_7191);
nor U9761 (N_9761,N_7850,N_6946);
nor U9762 (N_9762,N_8289,N_8094);
or U9763 (N_9763,N_8851,N_8861);
nor U9764 (N_9764,N_6990,N_8438);
nor U9765 (N_9765,N_6056,N_8391);
and U9766 (N_9766,N_8394,N_7208);
and U9767 (N_9767,N_8741,N_7800);
nand U9768 (N_9768,N_7699,N_6636);
and U9769 (N_9769,N_6363,N_7377);
and U9770 (N_9770,N_7042,N_8791);
nor U9771 (N_9771,N_6716,N_7768);
and U9772 (N_9772,N_6238,N_8626);
nor U9773 (N_9773,N_8960,N_6887);
or U9774 (N_9774,N_6669,N_8052);
and U9775 (N_9775,N_6105,N_8538);
or U9776 (N_9776,N_7613,N_8854);
or U9777 (N_9777,N_8669,N_8106);
nor U9778 (N_9778,N_6179,N_7813);
nor U9779 (N_9779,N_6603,N_8518);
nor U9780 (N_9780,N_8974,N_6414);
or U9781 (N_9781,N_8589,N_7655);
or U9782 (N_9782,N_8507,N_6963);
or U9783 (N_9783,N_6365,N_6127);
and U9784 (N_9784,N_6819,N_6676);
nor U9785 (N_9785,N_7893,N_6071);
nand U9786 (N_9786,N_6665,N_8061);
nand U9787 (N_9787,N_8810,N_7760);
and U9788 (N_9788,N_8264,N_7807);
nor U9789 (N_9789,N_8749,N_6581);
or U9790 (N_9790,N_8907,N_7281);
xnor U9791 (N_9791,N_8742,N_6998);
nand U9792 (N_9792,N_7996,N_8758);
nor U9793 (N_9793,N_8647,N_8759);
or U9794 (N_9794,N_8543,N_8407);
and U9795 (N_9795,N_8424,N_7286);
and U9796 (N_9796,N_7027,N_7446);
and U9797 (N_9797,N_7889,N_6089);
nand U9798 (N_9798,N_7115,N_8646);
or U9799 (N_9799,N_6671,N_6712);
nor U9800 (N_9800,N_7346,N_7273);
or U9801 (N_9801,N_8579,N_8508);
and U9802 (N_9802,N_6936,N_6768);
and U9803 (N_9803,N_6787,N_8308);
and U9804 (N_9804,N_7142,N_8958);
nand U9805 (N_9805,N_8874,N_8511);
nand U9806 (N_9806,N_8574,N_6680);
and U9807 (N_9807,N_7541,N_7253);
nor U9808 (N_9808,N_7162,N_6148);
or U9809 (N_9809,N_6462,N_7788);
or U9810 (N_9810,N_8364,N_7339);
nand U9811 (N_9811,N_6849,N_7251);
nand U9812 (N_9812,N_7279,N_8197);
nand U9813 (N_9813,N_6028,N_8039);
and U9814 (N_9814,N_7762,N_6474);
and U9815 (N_9815,N_8229,N_8405);
and U9816 (N_9816,N_6688,N_7632);
nor U9817 (N_9817,N_8397,N_6101);
and U9818 (N_9818,N_7605,N_6129);
or U9819 (N_9819,N_6909,N_8170);
or U9820 (N_9820,N_6280,N_7365);
and U9821 (N_9821,N_8561,N_8629);
and U9822 (N_9822,N_7688,N_6256);
nand U9823 (N_9823,N_6411,N_7923);
nor U9824 (N_9824,N_8906,N_8703);
and U9825 (N_9825,N_6999,N_7565);
or U9826 (N_9826,N_7874,N_6299);
and U9827 (N_9827,N_6235,N_8871);
or U9828 (N_9828,N_7444,N_8824);
nand U9829 (N_9829,N_6374,N_8431);
nand U9830 (N_9830,N_7256,N_7361);
and U9831 (N_9831,N_7006,N_8087);
or U9832 (N_9832,N_6247,N_6864);
and U9833 (N_9833,N_7962,N_6886);
xnor U9834 (N_9834,N_6274,N_6859);
nor U9835 (N_9835,N_8350,N_6750);
and U9836 (N_9836,N_8928,N_8200);
nor U9837 (N_9837,N_8619,N_8480);
nand U9838 (N_9838,N_6670,N_6955);
and U9839 (N_9839,N_7257,N_7476);
or U9840 (N_9840,N_7554,N_8498);
nor U9841 (N_9841,N_8275,N_8502);
xor U9842 (N_9842,N_8525,N_8672);
or U9843 (N_9843,N_8581,N_7982);
and U9844 (N_9844,N_8031,N_7120);
nand U9845 (N_9845,N_8602,N_7136);
and U9846 (N_9846,N_7501,N_8398);
or U9847 (N_9847,N_8243,N_6507);
nand U9848 (N_9848,N_6308,N_6597);
nand U9849 (N_9849,N_8948,N_7406);
or U9850 (N_9850,N_6813,N_6031);
or U9851 (N_9851,N_7706,N_7036);
nand U9852 (N_9852,N_8799,N_6815);
or U9853 (N_9853,N_7130,N_8812);
nand U9854 (N_9854,N_7823,N_7478);
or U9855 (N_9855,N_7334,N_6102);
or U9856 (N_9856,N_7997,N_7816);
nand U9857 (N_9857,N_8586,N_8594);
nand U9858 (N_9858,N_7651,N_8923);
nor U9859 (N_9859,N_8174,N_8829);
and U9860 (N_9860,N_6425,N_8002);
nand U9861 (N_9861,N_8012,N_7018);
and U9862 (N_9862,N_6044,N_7610);
or U9863 (N_9863,N_8192,N_7224);
and U9864 (N_9864,N_7912,N_8900);
or U9865 (N_9865,N_8694,N_8171);
nor U9866 (N_9866,N_8371,N_8028);
nor U9867 (N_9867,N_8982,N_6885);
nand U9868 (N_9868,N_7803,N_8643);
nand U9869 (N_9869,N_8673,N_8380);
nor U9870 (N_9870,N_7035,N_6778);
nand U9871 (N_9871,N_7624,N_8807);
or U9872 (N_9872,N_6699,N_7530);
or U9873 (N_9873,N_8395,N_7692);
nor U9874 (N_9874,N_7790,N_8964);
or U9875 (N_9875,N_7547,N_6098);
nand U9876 (N_9876,N_6988,N_7971);
nand U9877 (N_9877,N_7926,N_8675);
or U9878 (N_9878,N_8635,N_8072);
and U9879 (N_9879,N_8899,N_7396);
and U9880 (N_9880,N_7602,N_6700);
nand U9881 (N_9881,N_6100,N_8019);
and U9882 (N_9882,N_6131,N_8963);
or U9883 (N_9883,N_8726,N_8231);
nand U9884 (N_9884,N_7783,N_6426);
nand U9885 (N_9885,N_7622,N_8186);
and U9886 (N_9886,N_7856,N_7234);
nor U9887 (N_9887,N_7553,N_7970);
nand U9888 (N_9888,N_8678,N_6611);
or U9889 (N_9889,N_8569,N_6403);
xor U9890 (N_9890,N_7948,N_8011);
and U9891 (N_9891,N_6919,N_8765);
or U9892 (N_9892,N_8936,N_8447);
nor U9893 (N_9893,N_7691,N_6301);
nand U9894 (N_9894,N_8483,N_7403);
xor U9895 (N_9895,N_8558,N_7578);
and U9896 (N_9896,N_7332,N_7306);
nor U9897 (N_9897,N_7453,N_7192);
nand U9898 (N_9898,N_8680,N_8692);
or U9899 (N_9899,N_8587,N_7029);
nand U9900 (N_9900,N_7748,N_8878);
nor U9901 (N_9901,N_7898,N_8062);
nor U9902 (N_9902,N_6619,N_7037);
and U9903 (N_9903,N_8203,N_7165);
nand U9904 (N_9904,N_8671,N_7633);
nand U9905 (N_9905,N_7325,N_6985);
and U9906 (N_9906,N_8057,N_6764);
or U9907 (N_9907,N_8715,N_8522);
nand U9908 (N_9908,N_8068,N_7660);
nand U9909 (N_9909,N_7819,N_7628);
nand U9910 (N_9910,N_7007,N_7674);
and U9911 (N_9911,N_7644,N_6834);
nor U9912 (N_9912,N_6139,N_6283);
or U9913 (N_9913,N_8572,N_6857);
nor U9914 (N_9914,N_7091,N_6434);
nand U9915 (N_9915,N_7376,N_6668);
and U9916 (N_9916,N_6322,N_8608);
and U9917 (N_9917,N_8060,N_6812);
or U9918 (N_9918,N_6276,N_6254);
nor U9919 (N_9919,N_6850,N_8925);
nor U9920 (N_9920,N_6654,N_6841);
nor U9921 (N_9921,N_6432,N_8327);
nor U9922 (N_9922,N_6745,N_6851);
and U9923 (N_9923,N_6766,N_6333);
and U9924 (N_9924,N_7746,N_6037);
and U9925 (N_9925,N_8184,N_7576);
and U9926 (N_9926,N_8441,N_7981);
or U9927 (N_9927,N_7003,N_8036);
and U9928 (N_9928,N_6672,N_8952);
nor U9929 (N_9929,N_7594,N_7219);
nor U9930 (N_9930,N_8537,N_7703);
and U9931 (N_9931,N_6910,N_7878);
or U9932 (N_9932,N_6016,N_6751);
and U9933 (N_9933,N_8069,N_7947);
or U9934 (N_9934,N_8065,N_6232);
nand U9935 (N_9935,N_8910,N_7462);
nor U9936 (N_9936,N_8870,N_7753);
and U9937 (N_9937,N_6252,N_8205);
nor U9938 (N_9938,N_7739,N_8820);
nand U9939 (N_9939,N_7627,N_7127);
nand U9940 (N_9940,N_8909,N_6513);
or U9941 (N_9941,N_7083,N_7766);
and U9942 (N_9942,N_8896,N_7262);
or U9943 (N_9943,N_7936,N_8000);
and U9944 (N_9944,N_8930,N_7121);
nor U9945 (N_9945,N_6808,N_6923);
and U9946 (N_9946,N_6870,N_8118);
nor U9947 (N_9947,N_8847,N_7087);
nand U9948 (N_9948,N_8805,N_6831);
or U9949 (N_9949,N_8636,N_8227);
and U9950 (N_9950,N_7045,N_7016);
nor U9951 (N_9951,N_8073,N_6587);
or U9952 (N_9952,N_8359,N_8901);
nor U9953 (N_9953,N_8351,N_8712);
or U9954 (N_9954,N_7749,N_7357);
or U9955 (N_9955,N_8478,N_6470);
or U9956 (N_9956,N_8597,N_7756);
nor U9957 (N_9957,N_7686,N_8625);
nand U9958 (N_9958,N_7815,N_6468);
nor U9959 (N_9959,N_7375,N_8088);
xor U9960 (N_9960,N_6655,N_7799);
nor U9961 (N_9961,N_7204,N_7539);
or U9962 (N_9962,N_7932,N_8345);
and U9963 (N_9963,N_7863,N_7431);
or U9964 (N_9964,N_8310,N_8318);
nand U9965 (N_9965,N_6070,N_6109);
and U9966 (N_9966,N_7369,N_8269);
and U9967 (N_9967,N_6983,N_7102);
nand U9968 (N_9968,N_6339,N_8839);
and U9969 (N_9969,N_6021,N_6122);
or U9970 (N_9970,N_8778,N_6402);
and U9971 (N_9971,N_7966,N_7212);
nor U9972 (N_9972,N_7544,N_6701);
nor U9973 (N_9973,N_7877,N_8369);
or U9974 (N_9974,N_8654,N_7005);
nor U9975 (N_9975,N_8458,N_7071);
nor U9976 (N_9976,N_7626,N_6637);
or U9977 (N_9977,N_8120,N_7646);
and U9978 (N_9978,N_8641,N_6609);
and U9979 (N_9979,N_7489,N_8940);
or U9980 (N_9980,N_8837,N_7870);
nand U9981 (N_9981,N_6439,N_8144);
and U9982 (N_9982,N_6159,N_8490);
nor U9983 (N_9983,N_8293,N_6879);
and U9984 (N_9984,N_8183,N_6673);
or U9985 (N_9985,N_8999,N_7776);
nor U9986 (N_9986,N_8705,N_8585);
or U9987 (N_9987,N_8980,N_6642);
and U9988 (N_9988,N_7615,N_8634);
or U9989 (N_9989,N_7412,N_8201);
and U9990 (N_9990,N_7048,N_8248);
xnor U9991 (N_9991,N_6362,N_6937);
nor U9992 (N_9992,N_8204,N_6457);
and U9993 (N_9993,N_7775,N_7122);
and U9994 (N_9994,N_8110,N_8546);
nor U9995 (N_9995,N_8690,N_6255);
and U9996 (N_9996,N_6689,N_6391);
nand U9997 (N_9997,N_6306,N_8951);
or U9998 (N_9998,N_7435,N_8076);
nor U9999 (N_9999,N_7167,N_6674);
nand U10000 (N_10000,N_6422,N_8287);
or U10001 (N_10001,N_7572,N_7831);
xor U10002 (N_10002,N_6951,N_6314);
and U10003 (N_10003,N_7140,N_8145);
and U10004 (N_10004,N_7454,N_8664);
xnor U10005 (N_10005,N_6085,N_8194);
nand U10006 (N_10006,N_7064,N_7581);
and U10007 (N_10007,N_6134,N_7918);
nor U10008 (N_10008,N_8568,N_8058);
nand U10009 (N_10009,N_8531,N_7294);
and U10010 (N_10010,N_6989,N_6030);
nor U10011 (N_10011,N_6110,N_7059);
nand U10012 (N_10012,N_7743,N_7533);
and U10013 (N_10013,N_7335,N_7085);
or U10014 (N_10014,N_7146,N_7197);
or U10015 (N_10015,N_8683,N_7937);
or U10016 (N_10016,N_6197,N_7598);
or U10017 (N_10017,N_8049,N_7842);
nor U10018 (N_10018,N_8349,N_8336);
nor U10019 (N_10019,N_6590,N_6407);
or U10020 (N_10020,N_7422,N_6116);
nand U10021 (N_10021,N_6452,N_8283);
or U10022 (N_10022,N_6158,N_6574);
or U10023 (N_10023,N_7360,N_6412);
xnor U10024 (N_10024,N_8747,N_7571);
or U10025 (N_10025,N_8943,N_6978);
and U10026 (N_10026,N_6950,N_8843);
and U10027 (N_10027,N_8618,N_8157);
nand U10028 (N_10028,N_6228,N_8285);
nor U10029 (N_10029,N_7777,N_8456);
and U10030 (N_10030,N_6644,N_6226);
xor U10031 (N_10031,N_6233,N_6840);
nor U10032 (N_10032,N_7846,N_8042);
and U10033 (N_10033,N_6855,N_8617);
or U10034 (N_10034,N_7354,N_6516);
nor U10035 (N_10035,N_8442,N_8022);
nor U10036 (N_10036,N_7331,N_8976);
nor U10037 (N_10037,N_6890,N_6801);
and U10038 (N_10038,N_8488,N_7401);
or U10039 (N_10039,N_7482,N_7641);
nand U10040 (N_10040,N_8294,N_6210);
nor U10041 (N_10041,N_6063,N_8250);
or U10042 (N_10042,N_6702,N_7778);
and U10043 (N_10043,N_8793,N_8399);
and U10044 (N_10044,N_8489,N_8775);
xor U10045 (N_10045,N_6935,N_8040);
or U10046 (N_10046,N_8709,N_6419);
or U10047 (N_10047,N_7038,N_8504);
or U10048 (N_10048,N_6205,N_8529);
nor U10049 (N_10049,N_7735,N_8277);
nor U10050 (N_10050,N_6733,N_8455);
nor U10051 (N_10051,N_7682,N_6607);
nand U10052 (N_10052,N_8894,N_6551);
and U10053 (N_10053,N_7353,N_6722);
and U10054 (N_10054,N_6715,N_7222);
nor U10055 (N_10055,N_6149,N_7280);
and U10056 (N_10056,N_6535,N_6214);
or U10057 (N_10057,N_7524,N_7072);
nor U10058 (N_10058,N_8411,N_6009);
and U10059 (N_10059,N_7484,N_8240);
nor U10060 (N_10060,N_7069,N_8427);
xnor U10061 (N_10061,N_8189,N_6628);
nor U10062 (N_10062,N_6732,N_8818);
xor U10063 (N_10063,N_8796,N_8609);
nand U10064 (N_10064,N_8151,N_8462);
or U10065 (N_10065,N_8337,N_6662);
or U10066 (N_10066,N_8832,N_7840);
nand U10067 (N_10067,N_7126,N_7380);
nor U10068 (N_10068,N_8855,N_7421);
and U10069 (N_10069,N_7734,N_8482);
nand U10070 (N_10070,N_8434,N_7455);
xnor U10071 (N_10071,N_7752,N_7531);
and U10072 (N_10072,N_7715,N_6249);
or U10073 (N_10073,N_6986,N_6821);
nor U10074 (N_10074,N_8953,N_8803);
and U10075 (N_10075,N_6053,N_7758);
or U10076 (N_10076,N_7266,N_7879);
and U10077 (N_10077,N_7959,N_6376);
xnor U10078 (N_10078,N_8280,N_8785);
and U10079 (N_10079,N_6897,N_8698);
nor U10080 (N_10080,N_8825,N_8644);
or U10081 (N_10081,N_8090,N_7510);
nor U10082 (N_10082,N_8740,N_7195);
or U10083 (N_10083,N_7876,N_8037);
nand U10084 (N_10084,N_8127,N_6804);
nand U10085 (N_10085,N_6627,N_6512);
or U10086 (N_10086,N_6323,N_7836);
nand U10087 (N_10087,N_8210,N_6357);
and U10088 (N_10088,N_8689,N_7625);
and U10089 (N_10089,N_8506,N_8806);
or U10090 (N_10090,N_8648,N_7978);
nand U10091 (N_10091,N_6353,N_6615);
and U10092 (N_10092,N_8008,N_8358);
nand U10093 (N_10093,N_7149,N_8879);
nand U10094 (N_10094,N_7829,N_6493);
and U10095 (N_10095,N_8255,N_7040);
and U10096 (N_10096,N_7956,N_6092);
nand U10097 (N_10097,N_6390,N_8445);
and U10098 (N_10098,N_6144,N_6884);
or U10099 (N_10099,N_6444,N_6186);
and U10100 (N_10100,N_6074,N_6759);
or U10101 (N_10101,N_6442,N_6604);
or U10102 (N_10102,N_8089,N_7994);
nand U10103 (N_10103,N_6093,N_6051);
or U10104 (N_10104,N_8422,N_7259);
nand U10105 (N_10105,N_6415,N_8540);
nor U10106 (N_10106,N_6212,N_6082);
or U10107 (N_10107,N_7185,N_8400);
nor U10108 (N_10108,N_7049,N_7019);
or U10109 (N_10109,N_7659,N_7341);
and U10110 (N_10110,N_6889,N_8865);
nor U10111 (N_10111,N_8645,N_7809);
nand U10112 (N_10112,N_8430,N_6694);
or U10113 (N_10113,N_6664,N_7938);
nand U10114 (N_10114,N_8211,N_6138);
and U10115 (N_10115,N_7260,N_7881);
nand U10116 (N_10116,N_6754,N_6279);
or U10117 (N_10117,N_7922,N_6631);
and U10118 (N_10118,N_6312,N_8567);
or U10119 (N_10119,N_6418,N_6488);
or U10120 (N_10120,N_6932,N_8228);
or U10121 (N_10121,N_8532,N_6192);
nand U10122 (N_10122,N_8372,N_6451);
or U10123 (N_10123,N_7181,N_7187);
xor U10124 (N_10124,N_6836,N_8674);
or U10125 (N_10125,N_7470,N_6327);
nor U10126 (N_10126,N_8389,N_7022);
xor U10127 (N_10127,N_8382,N_6740);
nor U10128 (N_10128,N_7272,N_6784);
nor U10129 (N_10129,N_8284,N_6409);
nand U10130 (N_10130,N_8528,N_8970);
nand U10131 (N_10131,N_7479,N_7182);
nand U10132 (N_10132,N_7851,N_8756);
nor U10133 (N_10133,N_7466,N_7519);
nor U10134 (N_10134,N_6521,N_6906);
and U10135 (N_10135,N_6510,N_6203);
and U10136 (N_10136,N_6049,N_8290);
nor U10137 (N_10137,N_7732,N_7883);
nor U10138 (N_10138,N_8984,N_6230);
nor U10139 (N_10139,N_6128,N_8517);
or U10140 (N_10140,N_7394,N_6777);
nor U10141 (N_10141,N_6342,N_6743);
nor U10142 (N_10142,N_8138,N_6643);
or U10143 (N_10143,N_8402,N_6181);
or U10144 (N_10144,N_7316,N_6090);
and U10145 (N_10145,N_8808,N_8920);
nand U10146 (N_10146,N_7907,N_7862);
and U10147 (N_10147,N_7200,N_6145);
nor U10148 (N_10148,N_8198,N_8620);
nand U10149 (N_10149,N_6785,N_6257);
or U10150 (N_10150,N_8356,N_8939);
xor U10151 (N_10151,N_7226,N_6243);
or U10152 (N_10152,N_7964,N_6717);
nand U10153 (N_10153,N_6925,N_6048);
nor U10154 (N_10154,N_7958,N_8867);
nor U10155 (N_10155,N_7991,N_8708);
and U10156 (N_10156,N_8534,N_6250);
nand U10157 (N_10157,N_7043,N_7296);
or U10158 (N_10158,N_8555,N_8541);
and U10159 (N_10159,N_8623,N_8425);
nand U10160 (N_10160,N_7797,N_7068);
and U10161 (N_10161,N_7944,N_8633);
or U10162 (N_10162,N_8233,N_7158);
nor U10163 (N_10163,N_6579,N_6477);
and U10164 (N_10164,N_8668,N_7424);
or U10165 (N_10165,N_8148,N_7485);
nand U10166 (N_10166,N_8128,N_6117);
and U10167 (N_10167,N_6496,N_8046);
nor U10168 (N_10168,N_8802,N_7726);
nor U10169 (N_10169,N_6646,N_8191);
or U10170 (N_10170,N_8251,N_6329);
nor U10171 (N_10171,N_7995,N_7407);
nand U10172 (N_10172,N_8752,N_8099);
xor U10173 (N_10173,N_7419,N_7514);
nor U10174 (N_10174,N_6979,N_6678);
or U10175 (N_10175,N_8711,N_6560);
or U10176 (N_10176,N_7295,N_7502);
or U10177 (N_10177,N_8687,N_7373);
or U10178 (N_10178,N_7730,N_8700);
and U10179 (N_10179,N_7619,N_6124);
and U10180 (N_10180,N_8828,N_7560);
nand U10181 (N_10181,N_6868,N_7764);
and U10182 (N_10182,N_8362,N_6869);
or U10183 (N_10183,N_7194,N_7243);
nand U10184 (N_10184,N_7653,N_8998);
nand U10185 (N_10185,N_7056,N_6761);
and U10186 (N_10186,N_6972,N_8728);
and U10187 (N_10187,N_8360,N_6298);
and U10188 (N_10188,N_7132,N_7073);
or U10189 (N_10189,N_6519,N_6219);
or U10190 (N_10190,N_8501,N_7582);
and U10191 (N_10191,N_6167,N_6600);
or U10192 (N_10192,N_8764,N_8460);
nand U10193 (N_10193,N_8241,N_8416);
and U10194 (N_10194,N_6647,N_7263);
nor U10195 (N_10195,N_7201,N_6947);
and U10196 (N_10196,N_8388,N_7300);
or U10197 (N_10197,N_6796,N_7109);
or U10198 (N_10198,N_7915,N_6130);
nor U10199 (N_10199,N_6272,N_8167);
nand U10200 (N_10200,N_8521,N_6142);
nand U10201 (N_10201,N_8193,N_6544);
or U10202 (N_10202,N_6839,N_7010);
nand U10203 (N_10203,N_7034,N_6115);
and U10204 (N_10204,N_7171,N_6386);
and U10205 (N_10205,N_7134,N_7458);
nand U10206 (N_10206,N_6542,N_8547);
nor U10207 (N_10207,N_6533,N_7205);
or U10208 (N_10208,N_7854,N_6481);
and U10209 (N_10209,N_8630,N_6081);
or U10210 (N_10210,N_6260,N_7827);
nor U10211 (N_10211,N_6408,N_7770);
and U10212 (N_10212,N_7771,N_7378);
and U10213 (N_10213,N_8722,N_8697);
nand U10214 (N_10214,N_6639,N_8299);
or U10215 (N_10215,N_6399,N_6006);
and U10216 (N_10216,N_6820,N_8116);
nand U10217 (N_10217,N_7596,N_6326);
and U10218 (N_10218,N_6543,N_6027);
nor U10219 (N_10219,N_6965,N_7677);
or U10220 (N_10220,N_6727,N_7618);
or U10221 (N_10221,N_7326,N_7026);
nor U10222 (N_10222,N_7882,N_6423);
or U10223 (N_10223,N_7507,N_8383);
and U10224 (N_10224,N_6495,N_6017);
or U10225 (N_10225,N_8967,N_7442);
xor U10226 (N_10226,N_6822,N_7383);
nand U10227 (N_10227,N_8992,N_8852);
or U10228 (N_10228,N_7061,N_6629);
nand U10229 (N_10229,N_7319,N_8744);
and U10230 (N_10230,N_6349,N_7347);
nand U10231 (N_10231,N_7969,N_7832);
nor U10232 (N_10232,N_7623,N_6876);
nor U10233 (N_10233,N_8968,N_6018);
nor U10234 (N_10234,N_7153,N_6790);
and U10235 (N_10235,N_8236,N_8091);
and U10236 (N_10236,N_6677,N_7199);
or U10237 (N_10237,N_7285,N_7796);
nor U10238 (N_10238,N_6066,N_7871);
nor U10239 (N_10239,N_8603,N_6055);
nand U10240 (N_10240,N_8330,N_8107);
or U10241 (N_10241,N_7321,N_8840);
and U10242 (N_10242,N_7693,N_8092);
nand U10243 (N_10243,N_8433,N_6438);
and U10244 (N_10244,N_7909,N_8020);
nor U10245 (N_10245,N_8686,N_7238);
or U10246 (N_10246,N_7798,N_7754);
nand U10247 (N_10247,N_8493,N_8606);
nand U10248 (N_10248,N_6356,N_8898);
nand U10249 (N_10249,N_6760,N_6013);
nor U10250 (N_10250,N_6427,N_6069);
or U10251 (N_10251,N_7255,N_6546);
nand U10252 (N_10252,N_7050,N_8545);
or U10253 (N_10253,N_6547,N_8848);
or U10254 (N_10254,N_6073,N_7242);
nor U10255 (N_10255,N_7382,N_7564);
nand U10256 (N_10256,N_8126,N_6147);
nand U10257 (N_10257,N_7987,N_6182);
or U10258 (N_10258,N_7675,N_6075);
nor U10259 (N_10259,N_7835,N_8826);
or U10260 (N_10260,N_6184,N_8078);
and U10261 (N_10261,N_6907,N_6033);
and U10262 (N_10262,N_7389,N_8613);
or U10263 (N_10263,N_7387,N_6570);
and U10264 (N_10264,N_7794,N_8464);
nor U10265 (N_10265,N_7358,N_7352);
and U10266 (N_10266,N_7488,N_8023);
or U10267 (N_10267,N_6565,N_6393);
and U10268 (N_10268,N_8886,N_6389);
nand U10269 (N_10269,N_6307,N_7443);
nand U10270 (N_10270,N_6953,N_7496);
nor U10271 (N_10271,N_7292,N_6926);
nand U10272 (N_10272,N_8691,N_7108);
and U10273 (N_10273,N_6234,N_8220);
and U10274 (N_10274,N_7330,N_6392);
nor U10275 (N_10275,N_7595,N_7685);
nand U10276 (N_10276,N_8877,N_7834);
or U10277 (N_10277,N_6265,N_7000);
nor U10278 (N_10278,N_8481,N_7861);
nor U10279 (N_10279,N_7391,N_7763);
or U10280 (N_10280,N_8108,N_6916);
or U10281 (N_10281,N_7080,N_6262);
and U10282 (N_10282,N_6417,N_7213);
and U10283 (N_10283,N_7884,N_7351);
nor U10284 (N_10284,N_7483,N_7343);
nor U10285 (N_10285,N_6902,N_6458);
and U10286 (N_10286,N_8733,N_8208);
nand U10287 (N_10287,N_7159,N_8935);
and U10288 (N_10288,N_6852,N_6453);
and U10289 (N_10289,N_8082,N_6656);
or U10290 (N_10290,N_7423,N_7518);
nand U10291 (N_10291,N_8038,N_7725);
nor U10292 (N_10292,N_8370,N_6064);
nand U10293 (N_10293,N_8176,N_8181);
and U10294 (N_10294,N_6359,N_7252);
nand U10295 (N_10295,N_8165,N_8649);
nand U10296 (N_10296,N_7128,N_6187);
and U10297 (N_10297,N_6608,N_6651);
or U10298 (N_10298,N_7030,N_8161);
xor U10299 (N_10299,N_6927,N_6361);
or U10300 (N_10300,N_8339,N_6772);
nand U10301 (N_10301,N_7434,N_6572);
or U10302 (N_10302,N_7079,N_8085);
or U10303 (N_10303,N_6108,N_7869);
and U10304 (N_10304,N_6872,N_7124);
nand U10305 (N_10305,N_6473,N_7420);
nand U10306 (N_10306,N_7461,N_7906);
and U10307 (N_10307,N_8938,N_6981);
nor U10308 (N_10308,N_6421,N_6240);
nor U10309 (N_10309,N_8312,N_8166);
nand U10310 (N_10310,N_6001,N_7967);
or U10311 (N_10311,N_8751,N_7942);
or U10312 (N_10312,N_8154,N_8615);
nand U10313 (N_10313,N_8322,N_8773);
nor U10314 (N_10314,N_7563,N_6567);
nor U10315 (N_10315,N_7017,N_8016);
nand U10316 (N_10316,N_8013,N_8018);
nand U10317 (N_10317,N_6817,N_6475);
nand U10318 (N_10318,N_7755,N_6430);
and U10319 (N_10319,N_8559,N_6223);
nor U10320 (N_10320,N_8983,N_8218);
and U10321 (N_10321,N_6398,N_7999);
or U10322 (N_10322,N_7193,N_7298);
and U10323 (N_10323,N_6267,N_8199);
nand U10324 (N_10324,N_6052,N_8987);
nand U10325 (N_10325,N_8950,N_6118);
or U10326 (N_10326,N_7911,N_7436);
nor U10327 (N_10327,N_7362,N_7088);
or U10328 (N_10328,N_7449,N_6183);
or U10329 (N_10329,N_7452,N_7635);
and U10330 (N_10330,N_7972,N_8030);
nand U10331 (N_10331,N_6580,N_7895);
or U10332 (N_10332,N_6558,N_7356);
or U10333 (N_10333,N_6520,N_7398);
nor U10334 (N_10334,N_7472,N_7311);
nor U10335 (N_10335,N_8059,N_8931);
or U10336 (N_10336,N_8164,N_6792);
nor U10337 (N_10337,N_7168,N_8679);
or U10338 (N_10338,N_8659,N_6175);
and U10339 (N_10339,N_8423,N_7520);
and U10340 (N_10340,N_6908,N_8693);
or U10341 (N_10341,N_6095,N_8530);
nand U10342 (N_10342,N_8797,N_8604);
or U10343 (N_10343,N_6991,N_8784);
or U10344 (N_10344,N_7673,N_7567);
or U10345 (N_10345,N_6277,N_8155);
and U10346 (N_10346,N_6125,N_6178);
nand U10347 (N_10347,N_8926,N_6321);
nor U10348 (N_10348,N_7368,N_8461);
nor U10349 (N_10349,N_7217,N_8190);
nor U10350 (N_10350,N_7276,N_7350);
nand U10351 (N_10351,N_6472,N_8331);
nor U10352 (N_10352,N_8242,N_6135);
or U10353 (N_10353,N_8737,N_6461);
nand U10354 (N_10354,N_7157,N_6185);
or U10355 (N_10355,N_8817,N_6904);
nand U10356 (N_10356,N_7349,N_6710);
nor U10357 (N_10357,N_7649,N_7093);
or U10358 (N_10358,N_7174,N_6012);
xnor U10359 (N_10359,N_7110,N_8600);
nand U10360 (N_10360,N_7941,N_6706);
or U10361 (N_10361,N_7156,N_8888);
or U10362 (N_10362,N_8451,N_6517);
and U10363 (N_10363,N_8734,N_7062);
nor U10364 (N_10364,N_6348,N_6123);
nand U10365 (N_10365,N_8845,N_8798);
or U10366 (N_10366,N_7993,N_6649);
and U10367 (N_10367,N_7106,N_6659);
and U10368 (N_10368,N_7707,N_8179);
and U10369 (N_10369,N_7012,N_8271);
nand U10370 (N_10370,N_7885,N_6624);
nor U10371 (N_10371,N_7218,N_7459);
or U10372 (N_10372,N_8699,N_6793);
and U10373 (N_10373,N_6807,N_8281);
nor U10374 (N_10374,N_8682,N_6310);
and U10375 (N_10375,N_6498,N_7047);
or U10376 (N_10376,N_8723,N_8291);
nor U10377 (N_10377,N_8710,N_8396);
nor U10378 (N_10378,N_8302,N_8477);
xnor U10379 (N_10379,N_6176,N_8937);
nand U10380 (N_10380,N_8122,N_7312);
nor U10381 (N_10381,N_6748,N_6096);
nor U10382 (N_10382,N_7278,N_6933);
nand U10383 (N_10383,N_8500,N_7808);
or U10384 (N_10384,N_8386,N_8713);
or U10385 (N_10385,N_8745,N_7844);
nor U10386 (N_10386,N_8054,N_6088);
and U10387 (N_10387,N_6032,N_7908);
nor U10388 (N_10388,N_7543,N_6193);
nor U10389 (N_10389,N_8428,N_7456);
nand U10390 (N_10390,N_6982,N_6208);
xor U10391 (N_10391,N_8969,N_8475);
and U10392 (N_10392,N_7381,N_6328);
and U10393 (N_10393,N_7465,N_6645);
or U10394 (N_10394,N_6494,N_8598);
nor U10395 (N_10395,N_7548,N_6903);
nor U10396 (N_10396,N_7875,N_7291);
nor U10397 (N_10397,N_7718,N_7440);
nor U10398 (N_10398,N_6491,N_7848);
xor U10399 (N_10399,N_8564,N_7965);
and U10400 (N_10400,N_6029,N_6431);
and U10401 (N_10401,N_6436,N_8136);
or U10402 (N_10402,N_6816,N_8007);
nand U10403 (N_10403,N_8566,N_8516);
nand U10404 (N_10404,N_6961,N_6921);
and U10405 (N_10405,N_7837,N_7500);
nand U10406 (N_10406,N_7271,N_7372);
nand U10407 (N_10407,N_6157,N_7508);
nor U10408 (N_10408,N_6568,N_6724);
nor U10409 (N_10409,N_6528,N_7637);
nand U10410 (N_10410,N_7955,N_7849);
and U10411 (N_10411,N_6610,N_6687);
nand U10412 (N_10412,N_6121,N_8143);
nor U10413 (N_10413,N_8813,N_6039);
or U10414 (N_10414,N_8436,N_7821);
and U10415 (N_10415,N_6360,N_6449);
nor U10416 (N_10416,N_7694,N_8063);
or U10417 (N_10417,N_7172,N_8017);
and U10418 (N_10418,N_8041,N_7148);
and U10419 (N_10419,N_7525,N_7782);
nor U10420 (N_10420,N_6077,N_8182);
and U10421 (N_10421,N_7847,N_8592);
nor U10422 (N_10422,N_7552,N_8470);
or U10423 (N_10423,N_6011,N_7315);
or U10424 (N_10424,N_6293,N_7283);
or U10425 (N_10425,N_7975,N_8811);
nor U10426 (N_10426,N_7896,N_8124);
nor U10427 (N_10427,N_8492,N_6709);
nor U10428 (N_10428,N_7805,N_7940);
nor U10429 (N_10429,N_6613,N_6174);
nand U10430 (N_10430,N_6331,N_6866);
nor U10431 (N_10431,N_8652,N_7432);
or U10432 (N_10432,N_6456,N_8238);
nand U10433 (N_10433,N_6527,N_7811);
or U10434 (N_10434,N_7460,N_7249);
nor U10435 (N_10435,N_6344,N_6428);
or U10436 (N_10436,N_8381,N_7433);
nor U10437 (N_10437,N_6188,N_6842);
nor U10438 (N_10438,N_8326,N_7328);
or U10439 (N_10439,N_7450,N_8465);
nand U10440 (N_10440,N_8731,N_7843);
or U10441 (N_10441,N_6492,N_7095);
or U10442 (N_10442,N_6964,N_7700);
and U10443 (N_10443,N_8055,N_6220);
or U10444 (N_10444,N_6397,N_6569);
and U10445 (N_10445,N_6140,N_6204);
nor U10446 (N_10446,N_7795,N_6485);
nand U10447 (N_10447,N_6940,N_8596);
or U10448 (N_10448,N_8704,N_6657);
nand U10449 (N_10449,N_7125,N_7865);
nor U10450 (N_10450,N_8701,N_7690);
nor U10451 (N_10451,N_6605,N_7872);
and U10452 (N_10452,N_7060,N_8997);
and U10453 (N_10453,N_6877,N_8121);
nor U10454 (N_10454,N_8417,N_6912);
nor U10455 (N_10455,N_6913,N_7033);
nor U10456 (N_10456,N_8321,N_6126);
nand U10457 (N_10457,N_6731,N_6288);
nand U10458 (N_10458,N_7853,N_8780);
and U10459 (N_10459,N_6522,N_7274);
nor U10460 (N_10460,N_8081,N_8468);
and U10461 (N_10461,N_7220,N_6832);
or U10462 (N_10462,N_8162,N_8102);
nor U10463 (N_10463,N_8838,N_8554);
or U10464 (N_10464,N_8777,N_6191);
nor U10465 (N_10465,N_6623,N_7307);
or U10466 (N_10466,N_7920,N_8125);
nor U10467 (N_10467,N_8080,N_6229);
xnor U10468 (N_10468,N_8621,N_6379);
xnor U10469 (N_10469,N_7299,N_8885);
nor U10470 (N_10470,N_8927,N_6660);
nand U10471 (N_10471,N_6708,N_8209);
and U10472 (N_10472,N_8881,N_8520);
nor U10473 (N_10473,N_8781,N_7929);
and U10474 (N_10474,N_7833,N_8459);
or U10475 (N_10475,N_7684,N_8760);
nand U10476 (N_10476,N_8437,N_7740);
nand U10477 (N_10477,N_6920,N_6949);
nand U10478 (N_10478,N_8267,N_8769);
xnor U10479 (N_10479,N_6798,N_6364);
nor U10480 (N_10480,N_8064,N_6099);
nand U10481 (N_10481,N_6858,N_7652);
nand U10482 (N_10482,N_8265,N_7761);
nand U10483 (N_10483,N_6273,N_7240);
xor U10484 (N_10484,N_8873,N_8140);
nand U10485 (N_10485,N_6577,N_7475);
xnor U10486 (N_10486,N_7336,N_8582);
or U10487 (N_10487,N_6319,N_8044);
nand U10488 (N_10488,N_6756,N_6763);
and U10489 (N_10489,N_6202,N_6170);
or U10490 (N_10490,N_6164,N_8611);
nor U10491 (N_10491,N_7589,N_7597);
or U10492 (N_10492,N_6015,N_7713);
or U10493 (N_10493,N_8333,N_7231);
and U10494 (N_10494,N_7023,N_7269);
nand U10495 (N_10495,N_7904,N_7584);
nand U10496 (N_10496,N_8071,N_8903);
or U10497 (N_10497,N_8440,N_7025);
and U10498 (N_10498,N_8376,N_6244);
or U10499 (N_10499,N_8010,N_8202);
nand U10500 (N_10500,N_8357,N_6268);
nor U10501 (N_10501,N_8736,N_6093);
and U10502 (N_10502,N_6832,N_8651);
and U10503 (N_10503,N_6344,N_8022);
and U10504 (N_10504,N_6731,N_6341);
nor U10505 (N_10505,N_6777,N_6879);
nand U10506 (N_10506,N_6772,N_8833);
nand U10507 (N_10507,N_7075,N_7639);
xor U10508 (N_10508,N_6380,N_6291);
nor U10509 (N_10509,N_6638,N_8550);
nand U10510 (N_10510,N_8618,N_6186);
nand U10511 (N_10511,N_7429,N_8956);
nand U10512 (N_10512,N_6199,N_7339);
or U10513 (N_10513,N_7918,N_7400);
nand U10514 (N_10514,N_6810,N_7159);
nor U10515 (N_10515,N_7896,N_7969);
nand U10516 (N_10516,N_7863,N_7666);
nor U10517 (N_10517,N_6133,N_6348);
xor U10518 (N_10518,N_8183,N_8587);
nand U10519 (N_10519,N_7602,N_7888);
nand U10520 (N_10520,N_6308,N_6276);
nor U10521 (N_10521,N_6962,N_8283);
or U10522 (N_10522,N_6894,N_8973);
and U10523 (N_10523,N_8283,N_6541);
and U10524 (N_10524,N_8332,N_6705);
nand U10525 (N_10525,N_6755,N_6850);
xnor U10526 (N_10526,N_7992,N_6413);
nor U10527 (N_10527,N_8676,N_8506);
and U10528 (N_10528,N_8957,N_8148);
nor U10529 (N_10529,N_6659,N_7304);
nor U10530 (N_10530,N_8555,N_8651);
or U10531 (N_10531,N_7402,N_8061);
nand U10532 (N_10532,N_7136,N_6438);
and U10533 (N_10533,N_6524,N_6778);
xnor U10534 (N_10534,N_6423,N_6345);
nand U10535 (N_10535,N_6159,N_6330);
or U10536 (N_10536,N_8977,N_8399);
xnor U10537 (N_10537,N_7642,N_7623);
xor U10538 (N_10538,N_8020,N_8739);
or U10539 (N_10539,N_7102,N_8314);
nor U10540 (N_10540,N_7976,N_7250);
or U10541 (N_10541,N_8584,N_7577);
or U10542 (N_10542,N_6052,N_8738);
and U10543 (N_10543,N_7910,N_6998);
nand U10544 (N_10544,N_6286,N_7833);
and U10545 (N_10545,N_6219,N_8263);
nand U10546 (N_10546,N_6266,N_7104);
nor U10547 (N_10547,N_8472,N_8376);
and U10548 (N_10548,N_6275,N_6923);
nor U10549 (N_10549,N_8600,N_6491);
or U10550 (N_10550,N_6697,N_8592);
nor U10551 (N_10551,N_8709,N_7549);
nand U10552 (N_10552,N_6481,N_6618);
nor U10553 (N_10553,N_6961,N_6158);
nor U10554 (N_10554,N_6806,N_7158);
nand U10555 (N_10555,N_7206,N_7050);
nor U10556 (N_10556,N_6822,N_8863);
and U10557 (N_10557,N_6965,N_8558);
nand U10558 (N_10558,N_7003,N_8324);
and U10559 (N_10559,N_7733,N_8868);
and U10560 (N_10560,N_8900,N_7384);
nor U10561 (N_10561,N_8357,N_6158);
nand U10562 (N_10562,N_8153,N_8665);
nor U10563 (N_10563,N_6004,N_6374);
nor U10564 (N_10564,N_8132,N_6939);
and U10565 (N_10565,N_6413,N_7270);
nor U10566 (N_10566,N_6657,N_8011);
nor U10567 (N_10567,N_7201,N_7466);
or U10568 (N_10568,N_6886,N_7154);
nand U10569 (N_10569,N_8188,N_7311);
nor U10570 (N_10570,N_6747,N_8710);
nand U10571 (N_10571,N_6916,N_7617);
or U10572 (N_10572,N_6516,N_8076);
and U10573 (N_10573,N_6195,N_8098);
or U10574 (N_10574,N_8426,N_6259);
nand U10575 (N_10575,N_7577,N_8398);
or U10576 (N_10576,N_8504,N_6021);
or U10577 (N_10577,N_6120,N_6203);
and U10578 (N_10578,N_8412,N_7671);
nor U10579 (N_10579,N_8404,N_8748);
nand U10580 (N_10580,N_6521,N_7374);
xnor U10581 (N_10581,N_7590,N_6629);
nor U10582 (N_10582,N_8956,N_6803);
nand U10583 (N_10583,N_8734,N_8107);
xor U10584 (N_10584,N_8584,N_7716);
nand U10585 (N_10585,N_6993,N_8340);
or U10586 (N_10586,N_8593,N_7566);
nand U10587 (N_10587,N_7025,N_8439);
and U10588 (N_10588,N_7296,N_6168);
nor U10589 (N_10589,N_8499,N_8638);
nor U10590 (N_10590,N_7543,N_8933);
and U10591 (N_10591,N_8742,N_8289);
nor U10592 (N_10592,N_7190,N_6090);
or U10593 (N_10593,N_8175,N_8273);
nand U10594 (N_10594,N_6047,N_7719);
or U10595 (N_10595,N_8468,N_6459);
and U10596 (N_10596,N_6293,N_7044);
or U10597 (N_10597,N_6048,N_8170);
and U10598 (N_10598,N_7852,N_7337);
nand U10599 (N_10599,N_8682,N_6788);
nor U10600 (N_10600,N_6945,N_7473);
nor U10601 (N_10601,N_8158,N_6159);
and U10602 (N_10602,N_8078,N_6861);
or U10603 (N_10603,N_8727,N_7070);
nand U10604 (N_10604,N_8099,N_6612);
or U10605 (N_10605,N_8266,N_8240);
nand U10606 (N_10606,N_7431,N_6908);
nand U10607 (N_10607,N_7417,N_8433);
or U10608 (N_10608,N_7684,N_6426);
and U10609 (N_10609,N_7295,N_7692);
or U10610 (N_10610,N_8192,N_7135);
or U10611 (N_10611,N_7859,N_7135);
nor U10612 (N_10612,N_7909,N_8069);
or U10613 (N_10613,N_8297,N_8164);
nand U10614 (N_10614,N_6258,N_8166);
xor U10615 (N_10615,N_7275,N_7334);
nor U10616 (N_10616,N_8620,N_8968);
or U10617 (N_10617,N_7255,N_6769);
and U10618 (N_10618,N_8849,N_7441);
nand U10619 (N_10619,N_8041,N_6453);
or U10620 (N_10620,N_8839,N_8141);
and U10621 (N_10621,N_8720,N_7496);
nand U10622 (N_10622,N_8912,N_6225);
and U10623 (N_10623,N_7112,N_7698);
and U10624 (N_10624,N_6815,N_6869);
and U10625 (N_10625,N_6510,N_7572);
nor U10626 (N_10626,N_8202,N_6015);
nand U10627 (N_10627,N_8405,N_8003);
or U10628 (N_10628,N_8163,N_8028);
and U10629 (N_10629,N_7016,N_7586);
or U10630 (N_10630,N_6649,N_7573);
nor U10631 (N_10631,N_7343,N_6722);
or U10632 (N_10632,N_7235,N_6180);
or U10633 (N_10633,N_7131,N_7092);
and U10634 (N_10634,N_7412,N_7487);
and U10635 (N_10635,N_7343,N_7312);
or U10636 (N_10636,N_7115,N_8157);
nand U10637 (N_10637,N_6670,N_8407);
nor U10638 (N_10638,N_6340,N_8851);
nor U10639 (N_10639,N_6359,N_7382);
and U10640 (N_10640,N_8739,N_7918);
and U10641 (N_10641,N_8376,N_8922);
or U10642 (N_10642,N_6197,N_8394);
or U10643 (N_10643,N_6304,N_7426);
nand U10644 (N_10644,N_6836,N_7402);
and U10645 (N_10645,N_8659,N_8583);
or U10646 (N_10646,N_6175,N_7734);
xor U10647 (N_10647,N_6026,N_8701);
nor U10648 (N_10648,N_8805,N_8544);
nor U10649 (N_10649,N_8403,N_7524);
and U10650 (N_10650,N_8080,N_7777);
and U10651 (N_10651,N_8680,N_6842);
nand U10652 (N_10652,N_6316,N_8036);
and U10653 (N_10653,N_7766,N_8902);
nor U10654 (N_10654,N_6929,N_7427);
xnor U10655 (N_10655,N_8519,N_8918);
or U10656 (N_10656,N_8757,N_6521);
or U10657 (N_10657,N_7509,N_6099);
and U10658 (N_10658,N_7832,N_6036);
nor U10659 (N_10659,N_8192,N_6206);
and U10660 (N_10660,N_8957,N_8782);
nand U10661 (N_10661,N_6018,N_6868);
or U10662 (N_10662,N_8852,N_7389);
nor U10663 (N_10663,N_8158,N_8074);
nor U10664 (N_10664,N_6810,N_7887);
and U10665 (N_10665,N_6497,N_8841);
nor U10666 (N_10666,N_6423,N_6230);
or U10667 (N_10667,N_6425,N_8577);
nand U10668 (N_10668,N_8944,N_6076);
nand U10669 (N_10669,N_8440,N_7238);
nand U10670 (N_10670,N_8569,N_8609);
nand U10671 (N_10671,N_8269,N_7239);
nor U10672 (N_10672,N_8820,N_6910);
nand U10673 (N_10673,N_8259,N_6963);
nor U10674 (N_10674,N_6002,N_7023);
nand U10675 (N_10675,N_6469,N_7702);
nand U10676 (N_10676,N_8319,N_7199);
and U10677 (N_10677,N_7569,N_6767);
or U10678 (N_10678,N_7124,N_6043);
nor U10679 (N_10679,N_7426,N_6564);
or U10680 (N_10680,N_8975,N_7579);
and U10681 (N_10681,N_6142,N_7590);
nor U10682 (N_10682,N_6079,N_7627);
and U10683 (N_10683,N_8090,N_7576);
and U10684 (N_10684,N_6405,N_6433);
or U10685 (N_10685,N_7666,N_6998);
xnor U10686 (N_10686,N_8430,N_6488);
or U10687 (N_10687,N_6676,N_7133);
nor U10688 (N_10688,N_6326,N_6824);
nor U10689 (N_10689,N_7603,N_7038);
nor U10690 (N_10690,N_7980,N_7868);
or U10691 (N_10691,N_6205,N_8539);
nand U10692 (N_10692,N_7242,N_8605);
nand U10693 (N_10693,N_6239,N_8430);
and U10694 (N_10694,N_6685,N_7339);
nand U10695 (N_10695,N_6902,N_7806);
and U10696 (N_10696,N_6244,N_6935);
nand U10697 (N_10697,N_8876,N_7669);
and U10698 (N_10698,N_6266,N_8910);
nand U10699 (N_10699,N_8210,N_7842);
or U10700 (N_10700,N_8072,N_8748);
xor U10701 (N_10701,N_8304,N_8165);
nor U10702 (N_10702,N_6489,N_8890);
xnor U10703 (N_10703,N_6977,N_6818);
and U10704 (N_10704,N_8039,N_7781);
and U10705 (N_10705,N_8903,N_6194);
and U10706 (N_10706,N_6584,N_8348);
and U10707 (N_10707,N_6539,N_6367);
or U10708 (N_10708,N_7734,N_6427);
nand U10709 (N_10709,N_7303,N_7888);
nand U10710 (N_10710,N_6351,N_8303);
or U10711 (N_10711,N_6976,N_6756);
nor U10712 (N_10712,N_6929,N_6919);
nand U10713 (N_10713,N_7774,N_8488);
and U10714 (N_10714,N_7784,N_7005);
nor U10715 (N_10715,N_8128,N_8647);
nand U10716 (N_10716,N_8809,N_6890);
nor U10717 (N_10717,N_8817,N_8487);
or U10718 (N_10718,N_6134,N_7055);
and U10719 (N_10719,N_8856,N_8143);
and U10720 (N_10720,N_6796,N_8910);
and U10721 (N_10721,N_7155,N_8181);
nand U10722 (N_10722,N_7194,N_6168);
or U10723 (N_10723,N_6997,N_6262);
and U10724 (N_10724,N_7669,N_8058);
nor U10725 (N_10725,N_8902,N_7880);
nand U10726 (N_10726,N_7467,N_7882);
or U10727 (N_10727,N_6783,N_7376);
and U10728 (N_10728,N_7858,N_7499);
nor U10729 (N_10729,N_7886,N_6767);
nand U10730 (N_10730,N_8342,N_6005);
nand U10731 (N_10731,N_7654,N_6615);
nor U10732 (N_10732,N_7940,N_6075);
nand U10733 (N_10733,N_6081,N_8580);
nand U10734 (N_10734,N_6209,N_7456);
nor U10735 (N_10735,N_7124,N_8047);
or U10736 (N_10736,N_7715,N_6139);
or U10737 (N_10737,N_7307,N_7430);
and U10738 (N_10738,N_6366,N_7398);
or U10739 (N_10739,N_6366,N_8029);
nor U10740 (N_10740,N_7251,N_7424);
and U10741 (N_10741,N_8727,N_8832);
or U10742 (N_10742,N_7661,N_7377);
or U10743 (N_10743,N_6743,N_7489);
and U10744 (N_10744,N_8004,N_8586);
nor U10745 (N_10745,N_8744,N_7840);
and U10746 (N_10746,N_6789,N_7119);
and U10747 (N_10747,N_7529,N_8724);
and U10748 (N_10748,N_6820,N_8214);
nor U10749 (N_10749,N_8577,N_6388);
nor U10750 (N_10750,N_8526,N_6744);
nand U10751 (N_10751,N_7092,N_6129);
nand U10752 (N_10752,N_6214,N_7368);
and U10753 (N_10753,N_7436,N_8910);
nand U10754 (N_10754,N_6372,N_7961);
nand U10755 (N_10755,N_8931,N_8783);
and U10756 (N_10756,N_7775,N_7027);
nand U10757 (N_10757,N_7497,N_8806);
nor U10758 (N_10758,N_7343,N_6375);
and U10759 (N_10759,N_7558,N_8025);
nor U10760 (N_10760,N_8062,N_7188);
and U10761 (N_10761,N_8770,N_7930);
nand U10762 (N_10762,N_6931,N_6707);
nand U10763 (N_10763,N_8617,N_7976);
and U10764 (N_10764,N_8443,N_6384);
or U10765 (N_10765,N_8300,N_7544);
nand U10766 (N_10766,N_6621,N_8885);
nand U10767 (N_10767,N_7472,N_6423);
and U10768 (N_10768,N_8747,N_6946);
or U10769 (N_10769,N_7715,N_7972);
nand U10770 (N_10770,N_7684,N_6526);
or U10771 (N_10771,N_8451,N_7069);
nand U10772 (N_10772,N_7461,N_6634);
or U10773 (N_10773,N_6620,N_6409);
nor U10774 (N_10774,N_8521,N_7307);
and U10775 (N_10775,N_7472,N_6618);
nand U10776 (N_10776,N_7177,N_7614);
nor U10777 (N_10777,N_8564,N_7336);
nor U10778 (N_10778,N_6321,N_7769);
and U10779 (N_10779,N_8171,N_6882);
xor U10780 (N_10780,N_6867,N_8657);
nand U10781 (N_10781,N_7582,N_7678);
and U10782 (N_10782,N_6390,N_6046);
or U10783 (N_10783,N_8194,N_8960);
and U10784 (N_10784,N_8988,N_8941);
or U10785 (N_10785,N_6391,N_7127);
and U10786 (N_10786,N_6661,N_7928);
xnor U10787 (N_10787,N_8442,N_8811);
nor U10788 (N_10788,N_7113,N_6366);
nor U10789 (N_10789,N_8380,N_8121);
nor U10790 (N_10790,N_7867,N_7662);
nor U10791 (N_10791,N_8258,N_8577);
or U10792 (N_10792,N_7680,N_8397);
and U10793 (N_10793,N_7305,N_8646);
nand U10794 (N_10794,N_6814,N_7643);
and U10795 (N_10795,N_6533,N_7977);
and U10796 (N_10796,N_6103,N_8067);
nor U10797 (N_10797,N_6561,N_6089);
nand U10798 (N_10798,N_8666,N_6144);
or U10799 (N_10799,N_7977,N_7289);
nand U10800 (N_10800,N_8300,N_7715);
nand U10801 (N_10801,N_8537,N_7624);
nand U10802 (N_10802,N_7424,N_6197);
nand U10803 (N_10803,N_7897,N_7027);
nor U10804 (N_10804,N_6077,N_6282);
nand U10805 (N_10805,N_7686,N_6620);
or U10806 (N_10806,N_8567,N_8783);
and U10807 (N_10807,N_8784,N_8773);
and U10808 (N_10808,N_6308,N_7223);
or U10809 (N_10809,N_7557,N_8005);
nor U10810 (N_10810,N_7963,N_7622);
nand U10811 (N_10811,N_6270,N_8040);
nand U10812 (N_10812,N_6949,N_6049);
or U10813 (N_10813,N_6776,N_8514);
and U10814 (N_10814,N_6637,N_7975);
nand U10815 (N_10815,N_6717,N_6454);
and U10816 (N_10816,N_6370,N_8028);
and U10817 (N_10817,N_6309,N_7608);
or U10818 (N_10818,N_8393,N_8669);
and U10819 (N_10819,N_6544,N_7953);
or U10820 (N_10820,N_8083,N_8210);
nand U10821 (N_10821,N_8849,N_8685);
nor U10822 (N_10822,N_6767,N_7412);
and U10823 (N_10823,N_7170,N_8185);
nor U10824 (N_10824,N_8730,N_8888);
nor U10825 (N_10825,N_7148,N_7679);
and U10826 (N_10826,N_7808,N_7991);
and U10827 (N_10827,N_7953,N_7659);
nor U10828 (N_10828,N_7581,N_8192);
or U10829 (N_10829,N_6848,N_8669);
nor U10830 (N_10830,N_6977,N_7352);
nor U10831 (N_10831,N_7039,N_6601);
nand U10832 (N_10832,N_6886,N_6160);
or U10833 (N_10833,N_8283,N_8294);
and U10834 (N_10834,N_8487,N_8171);
nor U10835 (N_10835,N_6574,N_8818);
nand U10836 (N_10836,N_7015,N_8988);
and U10837 (N_10837,N_7180,N_8719);
nand U10838 (N_10838,N_6195,N_6859);
nand U10839 (N_10839,N_8710,N_7525);
and U10840 (N_10840,N_8205,N_7303);
and U10841 (N_10841,N_6940,N_7115);
and U10842 (N_10842,N_8858,N_6136);
nor U10843 (N_10843,N_6568,N_8478);
nor U10844 (N_10844,N_6170,N_8656);
or U10845 (N_10845,N_6048,N_7948);
or U10846 (N_10846,N_6040,N_7670);
xor U10847 (N_10847,N_6303,N_6599);
or U10848 (N_10848,N_8953,N_7448);
and U10849 (N_10849,N_6915,N_8354);
or U10850 (N_10850,N_8626,N_7396);
or U10851 (N_10851,N_8464,N_8259);
and U10852 (N_10852,N_7608,N_7447);
or U10853 (N_10853,N_8064,N_6333);
and U10854 (N_10854,N_8003,N_8770);
nor U10855 (N_10855,N_7308,N_8107);
nand U10856 (N_10856,N_6064,N_7662);
or U10857 (N_10857,N_8534,N_7591);
or U10858 (N_10858,N_7429,N_6217);
and U10859 (N_10859,N_7723,N_8005);
xor U10860 (N_10860,N_6383,N_7463);
nor U10861 (N_10861,N_6665,N_8130);
nand U10862 (N_10862,N_8604,N_7236);
nor U10863 (N_10863,N_8429,N_8477);
xnor U10864 (N_10864,N_6833,N_7829);
or U10865 (N_10865,N_8254,N_6372);
and U10866 (N_10866,N_6363,N_6154);
nand U10867 (N_10867,N_6197,N_6663);
nor U10868 (N_10868,N_7943,N_7571);
nor U10869 (N_10869,N_8521,N_8146);
nor U10870 (N_10870,N_6470,N_8426);
nor U10871 (N_10871,N_8354,N_8912);
and U10872 (N_10872,N_8061,N_7934);
xor U10873 (N_10873,N_8007,N_8364);
nand U10874 (N_10874,N_6761,N_6216);
nand U10875 (N_10875,N_7358,N_8066);
nand U10876 (N_10876,N_8226,N_7423);
or U10877 (N_10877,N_8419,N_7730);
nor U10878 (N_10878,N_8248,N_6297);
nand U10879 (N_10879,N_6268,N_6047);
nand U10880 (N_10880,N_7655,N_7268);
and U10881 (N_10881,N_7716,N_8858);
nor U10882 (N_10882,N_6104,N_6997);
nand U10883 (N_10883,N_8157,N_7959);
nand U10884 (N_10884,N_8135,N_6323);
nand U10885 (N_10885,N_8801,N_6761);
and U10886 (N_10886,N_8749,N_6052);
nor U10887 (N_10887,N_7155,N_7599);
or U10888 (N_10888,N_6502,N_6834);
nand U10889 (N_10889,N_8580,N_6100);
and U10890 (N_10890,N_6001,N_7549);
and U10891 (N_10891,N_7567,N_8564);
or U10892 (N_10892,N_8682,N_7247);
and U10893 (N_10893,N_7573,N_6083);
and U10894 (N_10894,N_6909,N_7878);
nor U10895 (N_10895,N_8745,N_8349);
nand U10896 (N_10896,N_8379,N_6207);
nand U10897 (N_10897,N_7364,N_7450);
and U10898 (N_10898,N_6252,N_8592);
xnor U10899 (N_10899,N_7486,N_8147);
and U10900 (N_10900,N_7495,N_7711);
nor U10901 (N_10901,N_7490,N_8119);
nand U10902 (N_10902,N_8605,N_8662);
and U10903 (N_10903,N_7912,N_6449);
and U10904 (N_10904,N_6839,N_6404);
and U10905 (N_10905,N_6066,N_6423);
and U10906 (N_10906,N_7774,N_7709);
nand U10907 (N_10907,N_6181,N_7775);
or U10908 (N_10908,N_7427,N_8070);
or U10909 (N_10909,N_6092,N_8901);
nand U10910 (N_10910,N_6864,N_6756);
or U10911 (N_10911,N_7978,N_8430);
nand U10912 (N_10912,N_6622,N_8393);
nor U10913 (N_10913,N_7761,N_6201);
nor U10914 (N_10914,N_7592,N_6799);
nand U10915 (N_10915,N_7224,N_6298);
or U10916 (N_10916,N_8922,N_6918);
nand U10917 (N_10917,N_6043,N_6868);
nand U10918 (N_10918,N_7477,N_7377);
nand U10919 (N_10919,N_6450,N_6481);
nor U10920 (N_10920,N_8729,N_7539);
nor U10921 (N_10921,N_8750,N_8696);
and U10922 (N_10922,N_6308,N_6179);
or U10923 (N_10923,N_6109,N_8588);
nor U10924 (N_10924,N_6424,N_6640);
or U10925 (N_10925,N_6542,N_7025);
and U10926 (N_10926,N_8053,N_7200);
and U10927 (N_10927,N_8348,N_7523);
or U10928 (N_10928,N_8566,N_6392);
nand U10929 (N_10929,N_8545,N_8559);
nor U10930 (N_10930,N_8285,N_8103);
nor U10931 (N_10931,N_6908,N_8928);
and U10932 (N_10932,N_6685,N_8430);
or U10933 (N_10933,N_8765,N_6730);
nor U10934 (N_10934,N_6484,N_7683);
nand U10935 (N_10935,N_7524,N_6845);
and U10936 (N_10936,N_7920,N_8521);
and U10937 (N_10937,N_6690,N_8994);
or U10938 (N_10938,N_8975,N_7869);
and U10939 (N_10939,N_8985,N_7708);
nand U10940 (N_10940,N_7814,N_7218);
nand U10941 (N_10941,N_7578,N_6031);
or U10942 (N_10942,N_7516,N_8499);
or U10943 (N_10943,N_8867,N_8918);
nor U10944 (N_10944,N_6644,N_7696);
or U10945 (N_10945,N_8755,N_8511);
and U10946 (N_10946,N_7298,N_7522);
nand U10947 (N_10947,N_8717,N_6781);
and U10948 (N_10948,N_7738,N_8546);
nand U10949 (N_10949,N_7568,N_7125);
nor U10950 (N_10950,N_8524,N_6494);
nor U10951 (N_10951,N_8422,N_7111);
nor U10952 (N_10952,N_8549,N_7391);
or U10953 (N_10953,N_7903,N_7527);
or U10954 (N_10954,N_8912,N_6627);
or U10955 (N_10955,N_6973,N_6795);
nor U10956 (N_10956,N_6791,N_6526);
and U10957 (N_10957,N_6662,N_7596);
nor U10958 (N_10958,N_6864,N_7494);
and U10959 (N_10959,N_6868,N_8121);
xor U10960 (N_10960,N_6564,N_7937);
nor U10961 (N_10961,N_6771,N_7483);
nand U10962 (N_10962,N_8775,N_8681);
and U10963 (N_10963,N_7491,N_7688);
nand U10964 (N_10964,N_8183,N_6227);
and U10965 (N_10965,N_8706,N_6905);
and U10966 (N_10966,N_7331,N_8728);
and U10967 (N_10967,N_6763,N_8078);
or U10968 (N_10968,N_8758,N_7187);
nor U10969 (N_10969,N_8937,N_8275);
or U10970 (N_10970,N_7009,N_6963);
and U10971 (N_10971,N_6144,N_7373);
or U10972 (N_10972,N_7699,N_6677);
nand U10973 (N_10973,N_8286,N_7504);
xor U10974 (N_10974,N_6413,N_6748);
nor U10975 (N_10975,N_6258,N_7513);
or U10976 (N_10976,N_6291,N_7761);
and U10977 (N_10977,N_6200,N_7906);
and U10978 (N_10978,N_6929,N_6624);
nor U10979 (N_10979,N_6045,N_8040);
and U10980 (N_10980,N_6635,N_6096);
nor U10981 (N_10981,N_7577,N_8393);
nand U10982 (N_10982,N_6742,N_7203);
nand U10983 (N_10983,N_6476,N_7938);
nor U10984 (N_10984,N_8081,N_7889);
or U10985 (N_10985,N_7519,N_6595);
and U10986 (N_10986,N_7717,N_6687);
nor U10987 (N_10987,N_8154,N_6526);
or U10988 (N_10988,N_8951,N_8412);
or U10989 (N_10989,N_8550,N_8442);
or U10990 (N_10990,N_7849,N_6395);
xor U10991 (N_10991,N_8841,N_6029);
nor U10992 (N_10992,N_7093,N_8711);
nor U10993 (N_10993,N_8243,N_7981);
and U10994 (N_10994,N_7139,N_8598);
and U10995 (N_10995,N_7750,N_6518);
nand U10996 (N_10996,N_6953,N_7069);
nor U10997 (N_10997,N_6657,N_6128);
and U10998 (N_10998,N_6505,N_8810);
nor U10999 (N_10999,N_6949,N_6985);
or U11000 (N_11000,N_8175,N_7949);
nor U11001 (N_11001,N_7401,N_8613);
nor U11002 (N_11002,N_8353,N_6013);
or U11003 (N_11003,N_8610,N_8661);
nor U11004 (N_11004,N_8563,N_7154);
or U11005 (N_11005,N_6500,N_7198);
xor U11006 (N_11006,N_8563,N_6719);
and U11007 (N_11007,N_8992,N_8632);
xor U11008 (N_11008,N_8874,N_8810);
and U11009 (N_11009,N_8874,N_7819);
nand U11010 (N_11010,N_7120,N_7504);
nor U11011 (N_11011,N_6581,N_8822);
nand U11012 (N_11012,N_7568,N_7363);
nor U11013 (N_11013,N_8896,N_7305);
xnor U11014 (N_11014,N_6687,N_7799);
nor U11015 (N_11015,N_8085,N_6921);
nand U11016 (N_11016,N_7418,N_7142);
nand U11017 (N_11017,N_7036,N_7107);
nand U11018 (N_11018,N_6669,N_8355);
and U11019 (N_11019,N_7972,N_7753);
nor U11020 (N_11020,N_7205,N_8888);
nor U11021 (N_11021,N_8252,N_7170);
or U11022 (N_11022,N_6814,N_8809);
and U11023 (N_11023,N_8665,N_7297);
nor U11024 (N_11024,N_7533,N_6630);
or U11025 (N_11025,N_6562,N_7395);
and U11026 (N_11026,N_6936,N_8819);
and U11027 (N_11027,N_6682,N_6444);
or U11028 (N_11028,N_8604,N_7631);
nand U11029 (N_11029,N_7373,N_7819);
nor U11030 (N_11030,N_8008,N_7732);
or U11031 (N_11031,N_8580,N_7102);
and U11032 (N_11032,N_8309,N_8847);
nand U11033 (N_11033,N_8210,N_7982);
or U11034 (N_11034,N_8303,N_7644);
and U11035 (N_11035,N_6031,N_8361);
or U11036 (N_11036,N_7704,N_8813);
and U11037 (N_11037,N_7972,N_6995);
and U11038 (N_11038,N_8294,N_8977);
nor U11039 (N_11039,N_7820,N_8477);
nand U11040 (N_11040,N_6181,N_8635);
nor U11041 (N_11041,N_8050,N_7481);
and U11042 (N_11042,N_6055,N_6624);
or U11043 (N_11043,N_8753,N_6321);
or U11044 (N_11044,N_7477,N_6349);
and U11045 (N_11045,N_6002,N_8658);
nor U11046 (N_11046,N_6311,N_8064);
nand U11047 (N_11047,N_8867,N_7466);
and U11048 (N_11048,N_7773,N_6174);
nor U11049 (N_11049,N_8833,N_7258);
nand U11050 (N_11050,N_6429,N_6071);
nor U11051 (N_11051,N_8062,N_6894);
or U11052 (N_11052,N_8966,N_6196);
or U11053 (N_11053,N_8806,N_7920);
and U11054 (N_11054,N_7801,N_6246);
and U11055 (N_11055,N_7050,N_7785);
and U11056 (N_11056,N_7473,N_6612);
nor U11057 (N_11057,N_8649,N_8920);
or U11058 (N_11058,N_8919,N_6632);
nand U11059 (N_11059,N_7926,N_6358);
and U11060 (N_11060,N_8441,N_7860);
and U11061 (N_11061,N_6014,N_8144);
nand U11062 (N_11062,N_8913,N_8467);
or U11063 (N_11063,N_8893,N_7661);
nor U11064 (N_11064,N_6720,N_6808);
nor U11065 (N_11065,N_6775,N_7665);
and U11066 (N_11066,N_7626,N_7432);
nor U11067 (N_11067,N_6143,N_6255);
nor U11068 (N_11068,N_7910,N_6040);
and U11069 (N_11069,N_6409,N_7017);
nand U11070 (N_11070,N_7355,N_7013);
and U11071 (N_11071,N_7376,N_8711);
and U11072 (N_11072,N_8115,N_6243);
nor U11073 (N_11073,N_6592,N_8928);
and U11074 (N_11074,N_8617,N_6376);
nor U11075 (N_11075,N_7012,N_8935);
nor U11076 (N_11076,N_6433,N_8385);
and U11077 (N_11077,N_6594,N_8554);
and U11078 (N_11078,N_7066,N_7409);
and U11079 (N_11079,N_8743,N_7121);
xnor U11080 (N_11080,N_8435,N_8424);
and U11081 (N_11081,N_8351,N_8526);
and U11082 (N_11082,N_7547,N_6137);
and U11083 (N_11083,N_8291,N_6052);
xnor U11084 (N_11084,N_8970,N_7046);
and U11085 (N_11085,N_6273,N_7445);
nor U11086 (N_11086,N_7304,N_7980);
or U11087 (N_11087,N_8168,N_6514);
and U11088 (N_11088,N_7788,N_8595);
xnor U11089 (N_11089,N_8453,N_6613);
nor U11090 (N_11090,N_8747,N_8425);
nand U11091 (N_11091,N_7380,N_8512);
nand U11092 (N_11092,N_7587,N_7684);
and U11093 (N_11093,N_6015,N_8807);
nor U11094 (N_11094,N_6860,N_6644);
or U11095 (N_11095,N_8300,N_8473);
and U11096 (N_11096,N_8243,N_6167);
or U11097 (N_11097,N_8042,N_7334);
or U11098 (N_11098,N_6807,N_6594);
nor U11099 (N_11099,N_6422,N_6896);
or U11100 (N_11100,N_6377,N_8805);
or U11101 (N_11101,N_8278,N_6667);
nand U11102 (N_11102,N_7634,N_6340);
nor U11103 (N_11103,N_6276,N_8713);
or U11104 (N_11104,N_7157,N_8112);
nand U11105 (N_11105,N_8534,N_8051);
nand U11106 (N_11106,N_7715,N_8015);
nor U11107 (N_11107,N_8583,N_7830);
nand U11108 (N_11108,N_7584,N_7050);
nand U11109 (N_11109,N_8250,N_6130);
or U11110 (N_11110,N_8690,N_6981);
nor U11111 (N_11111,N_6512,N_7178);
nor U11112 (N_11112,N_8515,N_7162);
nand U11113 (N_11113,N_8228,N_8376);
nand U11114 (N_11114,N_7017,N_7137);
or U11115 (N_11115,N_8142,N_6872);
nor U11116 (N_11116,N_8542,N_7749);
and U11117 (N_11117,N_7752,N_8801);
nand U11118 (N_11118,N_6938,N_8630);
nand U11119 (N_11119,N_7786,N_6821);
nand U11120 (N_11120,N_6693,N_7409);
nand U11121 (N_11121,N_8876,N_7574);
and U11122 (N_11122,N_7061,N_8806);
and U11123 (N_11123,N_7763,N_8459);
nor U11124 (N_11124,N_8776,N_6139);
nor U11125 (N_11125,N_8273,N_7334);
and U11126 (N_11126,N_7957,N_7000);
nor U11127 (N_11127,N_7406,N_6279);
nor U11128 (N_11128,N_8178,N_7586);
nand U11129 (N_11129,N_6177,N_6936);
or U11130 (N_11130,N_8567,N_8753);
nand U11131 (N_11131,N_8934,N_7184);
or U11132 (N_11132,N_6988,N_7099);
nor U11133 (N_11133,N_6533,N_8652);
xnor U11134 (N_11134,N_8233,N_8196);
or U11135 (N_11135,N_7247,N_8558);
or U11136 (N_11136,N_8431,N_8757);
or U11137 (N_11137,N_7368,N_6342);
and U11138 (N_11138,N_8340,N_6285);
nor U11139 (N_11139,N_7820,N_6925);
nand U11140 (N_11140,N_7735,N_7278);
nand U11141 (N_11141,N_8525,N_6246);
and U11142 (N_11142,N_8359,N_8807);
or U11143 (N_11143,N_6407,N_6592);
or U11144 (N_11144,N_7638,N_8559);
or U11145 (N_11145,N_7689,N_8188);
and U11146 (N_11146,N_7126,N_6615);
nand U11147 (N_11147,N_7134,N_6491);
or U11148 (N_11148,N_6488,N_8260);
nor U11149 (N_11149,N_7967,N_6203);
and U11150 (N_11150,N_8322,N_6703);
and U11151 (N_11151,N_7275,N_7828);
or U11152 (N_11152,N_7874,N_7391);
and U11153 (N_11153,N_8338,N_7979);
nand U11154 (N_11154,N_7805,N_6397);
nand U11155 (N_11155,N_7048,N_8761);
or U11156 (N_11156,N_6586,N_7636);
and U11157 (N_11157,N_8984,N_7805);
or U11158 (N_11158,N_7875,N_7673);
and U11159 (N_11159,N_8771,N_6266);
nor U11160 (N_11160,N_7669,N_8864);
nand U11161 (N_11161,N_7563,N_8437);
nor U11162 (N_11162,N_6835,N_6526);
and U11163 (N_11163,N_8232,N_7346);
and U11164 (N_11164,N_6663,N_7398);
or U11165 (N_11165,N_6764,N_8115);
nand U11166 (N_11166,N_6070,N_6657);
and U11167 (N_11167,N_7440,N_7795);
nor U11168 (N_11168,N_7878,N_7188);
nand U11169 (N_11169,N_6830,N_6386);
and U11170 (N_11170,N_6733,N_8218);
nand U11171 (N_11171,N_7017,N_8755);
nand U11172 (N_11172,N_8325,N_8458);
nand U11173 (N_11173,N_7464,N_8261);
nand U11174 (N_11174,N_8853,N_6222);
nor U11175 (N_11175,N_6076,N_6112);
and U11176 (N_11176,N_7055,N_7489);
and U11177 (N_11177,N_7817,N_7811);
and U11178 (N_11178,N_6383,N_6913);
nor U11179 (N_11179,N_7158,N_6379);
nor U11180 (N_11180,N_6455,N_6565);
nor U11181 (N_11181,N_6638,N_6997);
nor U11182 (N_11182,N_7762,N_7658);
nor U11183 (N_11183,N_8346,N_7469);
and U11184 (N_11184,N_6775,N_8343);
nand U11185 (N_11185,N_8938,N_8259);
nand U11186 (N_11186,N_8182,N_7311);
and U11187 (N_11187,N_8217,N_7283);
nand U11188 (N_11188,N_7892,N_8797);
or U11189 (N_11189,N_6577,N_8488);
or U11190 (N_11190,N_7209,N_6514);
and U11191 (N_11191,N_6439,N_7979);
or U11192 (N_11192,N_6197,N_7200);
nand U11193 (N_11193,N_8870,N_8896);
nor U11194 (N_11194,N_7821,N_7366);
nor U11195 (N_11195,N_8615,N_8722);
and U11196 (N_11196,N_7100,N_7243);
and U11197 (N_11197,N_8083,N_7026);
nor U11198 (N_11198,N_7639,N_8261);
and U11199 (N_11199,N_6599,N_6267);
or U11200 (N_11200,N_6224,N_6741);
nor U11201 (N_11201,N_7405,N_7710);
nor U11202 (N_11202,N_8295,N_6725);
and U11203 (N_11203,N_6008,N_8638);
and U11204 (N_11204,N_6962,N_7773);
nand U11205 (N_11205,N_6015,N_6280);
nor U11206 (N_11206,N_6203,N_7193);
nand U11207 (N_11207,N_7263,N_7907);
nor U11208 (N_11208,N_8812,N_7428);
nand U11209 (N_11209,N_6282,N_6817);
nand U11210 (N_11210,N_8763,N_7984);
nand U11211 (N_11211,N_6809,N_6439);
and U11212 (N_11212,N_7876,N_8290);
or U11213 (N_11213,N_8947,N_6745);
nor U11214 (N_11214,N_8770,N_6300);
and U11215 (N_11215,N_8299,N_6754);
or U11216 (N_11216,N_6788,N_6256);
and U11217 (N_11217,N_8973,N_6378);
nand U11218 (N_11218,N_8784,N_7354);
and U11219 (N_11219,N_6862,N_8925);
nand U11220 (N_11220,N_8453,N_8685);
or U11221 (N_11221,N_8947,N_7890);
nor U11222 (N_11222,N_8648,N_6710);
or U11223 (N_11223,N_8837,N_7910);
nor U11224 (N_11224,N_7163,N_6542);
nor U11225 (N_11225,N_6084,N_8016);
or U11226 (N_11226,N_8986,N_6493);
nand U11227 (N_11227,N_6117,N_7200);
nor U11228 (N_11228,N_6632,N_8177);
nor U11229 (N_11229,N_8000,N_8336);
and U11230 (N_11230,N_8607,N_7685);
nand U11231 (N_11231,N_7572,N_8688);
and U11232 (N_11232,N_8354,N_8826);
or U11233 (N_11233,N_6124,N_8926);
xor U11234 (N_11234,N_7201,N_6831);
and U11235 (N_11235,N_6461,N_6552);
and U11236 (N_11236,N_6861,N_7485);
or U11237 (N_11237,N_7428,N_8702);
nor U11238 (N_11238,N_6861,N_6871);
and U11239 (N_11239,N_6469,N_8021);
and U11240 (N_11240,N_8347,N_7968);
and U11241 (N_11241,N_6573,N_6393);
or U11242 (N_11242,N_7537,N_8439);
and U11243 (N_11243,N_8814,N_6784);
and U11244 (N_11244,N_8204,N_7126);
nor U11245 (N_11245,N_7343,N_7372);
nand U11246 (N_11246,N_6574,N_8753);
nand U11247 (N_11247,N_6272,N_8492);
and U11248 (N_11248,N_6845,N_7041);
or U11249 (N_11249,N_8621,N_6136);
nor U11250 (N_11250,N_6006,N_7297);
nand U11251 (N_11251,N_8026,N_7921);
or U11252 (N_11252,N_8461,N_6331);
nor U11253 (N_11253,N_6007,N_8792);
nand U11254 (N_11254,N_6015,N_7741);
or U11255 (N_11255,N_8334,N_8433);
nand U11256 (N_11256,N_8786,N_7100);
or U11257 (N_11257,N_8276,N_7452);
and U11258 (N_11258,N_8841,N_8915);
nor U11259 (N_11259,N_7143,N_7057);
nor U11260 (N_11260,N_7684,N_7073);
or U11261 (N_11261,N_8349,N_8063);
nor U11262 (N_11262,N_6542,N_6825);
and U11263 (N_11263,N_6241,N_8971);
nand U11264 (N_11264,N_7021,N_8933);
or U11265 (N_11265,N_6924,N_6629);
nor U11266 (N_11266,N_6573,N_6947);
or U11267 (N_11267,N_7491,N_8073);
and U11268 (N_11268,N_7585,N_7770);
nand U11269 (N_11269,N_6434,N_7835);
and U11270 (N_11270,N_7497,N_8820);
nor U11271 (N_11271,N_6291,N_6825);
nand U11272 (N_11272,N_6663,N_8797);
or U11273 (N_11273,N_8539,N_8460);
nor U11274 (N_11274,N_7151,N_7243);
and U11275 (N_11275,N_7653,N_6600);
and U11276 (N_11276,N_7273,N_7232);
and U11277 (N_11277,N_8499,N_6162);
nor U11278 (N_11278,N_7327,N_7867);
nor U11279 (N_11279,N_6540,N_8902);
and U11280 (N_11280,N_8644,N_6556);
and U11281 (N_11281,N_6073,N_7286);
nand U11282 (N_11282,N_8715,N_8270);
and U11283 (N_11283,N_6169,N_8116);
nand U11284 (N_11284,N_6441,N_6474);
nand U11285 (N_11285,N_8109,N_7109);
nor U11286 (N_11286,N_7270,N_7781);
and U11287 (N_11287,N_7965,N_6459);
nand U11288 (N_11288,N_8078,N_6512);
nor U11289 (N_11289,N_8575,N_7168);
nor U11290 (N_11290,N_7633,N_8083);
nand U11291 (N_11291,N_8754,N_8323);
and U11292 (N_11292,N_6046,N_7797);
or U11293 (N_11293,N_8404,N_8620);
or U11294 (N_11294,N_8355,N_7579);
nand U11295 (N_11295,N_8593,N_7607);
nand U11296 (N_11296,N_8058,N_6103);
or U11297 (N_11297,N_6278,N_6759);
and U11298 (N_11298,N_8196,N_7893);
and U11299 (N_11299,N_6837,N_7328);
nor U11300 (N_11300,N_7989,N_6512);
nand U11301 (N_11301,N_7976,N_8221);
nand U11302 (N_11302,N_6239,N_6332);
or U11303 (N_11303,N_8144,N_6540);
or U11304 (N_11304,N_6070,N_6271);
nand U11305 (N_11305,N_8362,N_6009);
and U11306 (N_11306,N_6272,N_6929);
nor U11307 (N_11307,N_8609,N_6240);
nor U11308 (N_11308,N_8097,N_6628);
xor U11309 (N_11309,N_7655,N_8309);
or U11310 (N_11310,N_7171,N_6740);
nor U11311 (N_11311,N_7378,N_6943);
and U11312 (N_11312,N_8808,N_7233);
xor U11313 (N_11313,N_8895,N_7011);
nor U11314 (N_11314,N_8172,N_6380);
nand U11315 (N_11315,N_7346,N_6736);
nor U11316 (N_11316,N_8512,N_7128);
or U11317 (N_11317,N_8593,N_7034);
and U11318 (N_11318,N_7304,N_6260);
nand U11319 (N_11319,N_7143,N_7691);
nand U11320 (N_11320,N_8794,N_6025);
nor U11321 (N_11321,N_6361,N_7448);
nand U11322 (N_11322,N_6210,N_6446);
nand U11323 (N_11323,N_8576,N_6637);
nand U11324 (N_11324,N_6852,N_8516);
and U11325 (N_11325,N_7435,N_7522);
or U11326 (N_11326,N_8030,N_8897);
and U11327 (N_11327,N_8051,N_7209);
nand U11328 (N_11328,N_8652,N_8354);
nor U11329 (N_11329,N_8332,N_6041);
nor U11330 (N_11330,N_7410,N_7131);
or U11331 (N_11331,N_8998,N_7751);
or U11332 (N_11332,N_6683,N_8201);
or U11333 (N_11333,N_7092,N_8757);
nor U11334 (N_11334,N_7544,N_7944);
and U11335 (N_11335,N_6208,N_8201);
xnor U11336 (N_11336,N_7590,N_7364);
nor U11337 (N_11337,N_7411,N_8956);
nor U11338 (N_11338,N_8528,N_7266);
nand U11339 (N_11339,N_6074,N_6766);
nand U11340 (N_11340,N_6906,N_6834);
nor U11341 (N_11341,N_6579,N_8118);
and U11342 (N_11342,N_6316,N_6923);
nand U11343 (N_11343,N_7113,N_6406);
and U11344 (N_11344,N_6501,N_7489);
xnor U11345 (N_11345,N_7875,N_6905);
or U11346 (N_11346,N_6465,N_7076);
nor U11347 (N_11347,N_6240,N_6786);
and U11348 (N_11348,N_8639,N_6961);
and U11349 (N_11349,N_8705,N_6879);
or U11350 (N_11350,N_6038,N_8861);
xor U11351 (N_11351,N_7429,N_8724);
and U11352 (N_11352,N_7461,N_7728);
nand U11353 (N_11353,N_6645,N_8083);
and U11354 (N_11354,N_6653,N_8920);
or U11355 (N_11355,N_6087,N_8584);
nand U11356 (N_11356,N_7506,N_6909);
nand U11357 (N_11357,N_7460,N_6601);
and U11358 (N_11358,N_8468,N_6690);
and U11359 (N_11359,N_6682,N_6990);
and U11360 (N_11360,N_7608,N_7495);
nor U11361 (N_11361,N_6637,N_6828);
or U11362 (N_11362,N_8273,N_8335);
nand U11363 (N_11363,N_8604,N_6379);
nand U11364 (N_11364,N_6747,N_6054);
or U11365 (N_11365,N_6327,N_8812);
nor U11366 (N_11366,N_6893,N_7428);
and U11367 (N_11367,N_7968,N_8431);
nor U11368 (N_11368,N_7374,N_8823);
or U11369 (N_11369,N_6478,N_8763);
and U11370 (N_11370,N_6578,N_6370);
nor U11371 (N_11371,N_7901,N_8988);
nor U11372 (N_11372,N_8028,N_6720);
nor U11373 (N_11373,N_7569,N_7143);
nand U11374 (N_11374,N_6612,N_7670);
nand U11375 (N_11375,N_7603,N_7362);
nand U11376 (N_11376,N_6684,N_7608);
nand U11377 (N_11377,N_6354,N_7411);
nand U11378 (N_11378,N_6147,N_6329);
nor U11379 (N_11379,N_8830,N_7305);
nand U11380 (N_11380,N_6733,N_6583);
nand U11381 (N_11381,N_8149,N_8395);
or U11382 (N_11382,N_7907,N_8377);
nor U11383 (N_11383,N_8521,N_8490);
nor U11384 (N_11384,N_7500,N_8142);
nor U11385 (N_11385,N_7786,N_7918);
xor U11386 (N_11386,N_8495,N_8078);
and U11387 (N_11387,N_6206,N_7520);
and U11388 (N_11388,N_7921,N_7075);
or U11389 (N_11389,N_6152,N_6060);
and U11390 (N_11390,N_8679,N_6860);
or U11391 (N_11391,N_7193,N_6780);
nor U11392 (N_11392,N_6307,N_6972);
nor U11393 (N_11393,N_8446,N_7559);
nand U11394 (N_11394,N_8320,N_6304);
nand U11395 (N_11395,N_6265,N_8433);
or U11396 (N_11396,N_6081,N_8983);
nor U11397 (N_11397,N_8231,N_7522);
nor U11398 (N_11398,N_6601,N_8641);
and U11399 (N_11399,N_8369,N_7203);
or U11400 (N_11400,N_6543,N_7926);
nand U11401 (N_11401,N_7805,N_7088);
or U11402 (N_11402,N_7638,N_6876);
and U11403 (N_11403,N_6890,N_8500);
or U11404 (N_11404,N_8762,N_8430);
or U11405 (N_11405,N_7961,N_8697);
or U11406 (N_11406,N_7686,N_8164);
and U11407 (N_11407,N_7539,N_6926);
nand U11408 (N_11408,N_7179,N_8052);
and U11409 (N_11409,N_8771,N_7040);
and U11410 (N_11410,N_7099,N_7875);
xor U11411 (N_11411,N_6032,N_7689);
or U11412 (N_11412,N_6101,N_8992);
and U11413 (N_11413,N_6578,N_7088);
nand U11414 (N_11414,N_8538,N_7339);
or U11415 (N_11415,N_7113,N_6512);
nand U11416 (N_11416,N_8022,N_8311);
nor U11417 (N_11417,N_7756,N_6519);
and U11418 (N_11418,N_6662,N_8700);
and U11419 (N_11419,N_8920,N_7849);
and U11420 (N_11420,N_6575,N_7998);
and U11421 (N_11421,N_7039,N_8120);
nand U11422 (N_11422,N_6482,N_6562);
nand U11423 (N_11423,N_8390,N_7515);
and U11424 (N_11424,N_8583,N_6269);
or U11425 (N_11425,N_7125,N_7147);
and U11426 (N_11426,N_8429,N_6041);
nor U11427 (N_11427,N_7759,N_7172);
nand U11428 (N_11428,N_6302,N_7658);
nor U11429 (N_11429,N_7494,N_6900);
nor U11430 (N_11430,N_6688,N_6517);
or U11431 (N_11431,N_8953,N_8496);
nand U11432 (N_11432,N_8279,N_8191);
nor U11433 (N_11433,N_8782,N_7183);
nor U11434 (N_11434,N_6208,N_7452);
nand U11435 (N_11435,N_8307,N_6484);
nor U11436 (N_11436,N_7850,N_7196);
or U11437 (N_11437,N_6602,N_6071);
and U11438 (N_11438,N_8825,N_6204);
or U11439 (N_11439,N_6358,N_8707);
nor U11440 (N_11440,N_7750,N_6945);
or U11441 (N_11441,N_7497,N_6701);
xor U11442 (N_11442,N_6122,N_7328);
and U11443 (N_11443,N_6285,N_8190);
nand U11444 (N_11444,N_6922,N_6973);
and U11445 (N_11445,N_7592,N_8063);
xor U11446 (N_11446,N_8075,N_8481);
nor U11447 (N_11447,N_7241,N_6119);
and U11448 (N_11448,N_6236,N_6504);
nor U11449 (N_11449,N_8626,N_8989);
nand U11450 (N_11450,N_6411,N_8322);
nand U11451 (N_11451,N_7455,N_7539);
nor U11452 (N_11452,N_8193,N_8055);
nand U11453 (N_11453,N_7496,N_8934);
or U11454 (N_11454,N_6132,N_7205);
nand U11455 (N_11455,N_8297,N_6697);
nand U11456 (N_11456,N_6418,N_7212);
nor U11457 (N_11457,N_8700,N_6962);
and U11458 (N_11458,N_7004,N_6763);
or U11459 (N_11459,N_6804,N_7844);
or U11460 (N_11460,N_6288,N_8034);
xnor U11461 (N_11461,N_6507,N_6565);
nor U11462 (N_11462,N_7887,N_7451);
and U11463 (N_11463,N_7259,N_7578);
nand U11464 (N_11464,N_6507,N_7624);
nor U11465 (N_11465,N_6350,N_8311);
and U11466 (N_11466,N_7714,N_7218);
or U11467 (N_11467,N_8702,N_6473);
or U11468 (N_11468,N_7709,N_6100);
or U11469 (N_11469,N_8559,N_7186);
nor U11470 (N_11470,N_6240,N_7189);
nand U11471 (N_11471,N_6649,N_7730);
nor U11472 (N_11472,N_7492,N_6745);
nor U11473 (N_11473,N_8516,N_6477);
nand U11474 (N_11474,N_6616,N_6861);
nand U11475 (N_11475,N_6106,N_6603);
and U11476 (N_11476,N_6097,N_8854);
nand U11477 (N_11477,N_8472,N_7472);
nand U11478 (N_11478,N_8256,N_7219);
nand U11479 (N_11479,N_8227,N_7004);
nor U11480 (N_11480,N_8644,N_7731);
and U11481 (N_11481,N_7666,N_7404);
nor U11482 (N_11482,N_6069,N_7662);
and U11483 (N_11483,N_8865,N_7055);
and U11484 (N_11484,N_7255,N_8698);
nor U11485 (N_11485,N_7041,N_6848);
nand U11486 (N_11486,N_6078,N_7145);
or U11487 (N_11487,N_6668,N_7568);
and U11488 (N_11488,N_8023,N_6438);
and U11489 (N_11489,N_6822,N_8900);
and U11490 (N_11490,N_7096,N_6813);
and U11491 (N_11491,N_8162,N_7714);
nand U11492 (N_11492,N_6315,N_6331);
nor U11493 (N_11493,N_7526,N_8150);
nor U11494 (N_11494,N_8690,N_7875);
nand U11495 (N_11495,N_6575,N_7762);
xor U11496 (N_11496,N_7625,N_7653);
nand U11497 (N_11497,N_6474,N_8900);
nor U11498 (N_11498,N_7271,N_8060);
or U11499 (N_11499,N_6210,N_8291);
and U11500 (N_11500,N_8833,N_8630);
and U11501 (N_11501,N_8717,N_7149);
nor U11502 (N_11502,N_8866,N_6288);
nor U11503 (N_11503,N_8565,N_7590);
and U11504 (N_11504,N_8642,N_6035);
nand U11505 (N_11505,N_7621,N_6509);
nand U11506 (N_11506,N_7677,N_7533);
nor U11507 (N_11507,N_8786,N_7161);
or U11508 (N_11508,N_8594,N_8918);
nor U11509 (N_11509,N_8126,N_8353);
nor U11510 (N_11510,N_8381,N_8382);
nand U11511 (N_11511,N_8420,N_6044);
or U11512 (N_11512,N_6291,N_7029);
nand U11513 (N_11513,N_8469,N_7983);
nor U11514 (N_11514,N_8979,N_7420);
nand U11515 (N_11515,N_6216,N_7128);
or U11516 (N_11516,N_7255,N_6094);
or U11517 (N_11517,N_7941,N_6819);
or U11518 (N_11518,N_6064,N_6073);
and U11519 (N_11519,N_8751,N_8508);
nand U11520 (N_11520,N_7142,N_8903);
or U11521 (N_11521,N_7234,N_7062);
or U11522 (N_11522,N_7586,N_6795);
or U11523 (N_11523,N_6592,N_8930);
nor U11524 (N_11524,N_7436,N_7655);
nor U11525 (N_11525,N_7504,N_8163);
nand U11526 (N_11526,N_8149,N_8407);
and U11527 (N_11527,N_8480,N_8025);
nand U11528 (N_11528,N_6556,N_6137);
nor U11529 (N_11529,N_8527,N_7834);
and U11530 (N_11530,N_6126,N_7433);
and U11531 (N_11531,N_7810,N_7117);
nor U11532 (N_11532,N_6504,N_7999);
and U11533 (N_11533,N_6031,N_6242);
and U11534 (N_11534,N_6231,N_8678);
or U11535 (N_11535,N_8176,N_6100);
nand U11536 (N_11536,N_6115,N_8367);
or U11537 (N_11537,N_6081,N_6765);
nor U11538 (N_11538,N_6291,N_8115);
nand U11539 (N_11539,N_8030,N_8035);
nand U11540 (N_11540,N_8494,N_6071);
nand U11541 (N_11541,N_7524,N_8769);
and U11542 (N_11542,N_7521,N_8770);
and U11543 (N_11543,N_6316,N_7465);
nand U11544 (N_11544,N_7693,N_8642);
nor U11545 (N_11545,N_6882,N_8872);
nand U11546 (N_11546,N_8893,N_6873);
and U11547 (N_11547,N_7731,N_6758);
or U11548 (N_11548,N_8496,N_8712);
or U11549 (N_11549,N_7218,N_6411);
or U11550 (N_11550,N_7723,N_8633);
nor U11551 (N_11551,N_8460,N_7928);
or U11552 (N_11552,N_7507,N_8305);
nor U11553 (N_11553,N_7257,N_7709);
or U11554 (N_11554,N_7700,N_7506);
xnor U11555 (N_11555,N_8750,N_6436);
nand U11556 (N_11556,N_7275,N_6548);
nand U11557 (N_11557,N_7837,N_8054);
nor U11558 (N_11558,N_7191,N_8288);
nor U11559 (N_11559,N_6860,N_7010);
and U11560 (N_11560,N_6267,N_8201);
nor U11561 (N_11561,N_7271,N_6777);
nor U11562 (N_11562,N_8449,N_8311);
or U11563 (N_11563,N_7617,N_6524);
nand U11564 (N_11564,N_7620,N_8384);
and U11565 (N_11565,N_7007,N_6271);
nor U11566 (N_11566,N_8748,N_8249);
nand U11567 (N_11567,N_8585,N_7995);
or U11568 (N_11568,N_7957,N_6870);
nand U11569 (N_11569,N_6042,N_7756);
nor U11570 (N_11570,N_6324,N_6707);
or U11571 (N_11571,N_8756,N_7340);
nor U11572 (N_11572,N_7422,N_6304);
or U11573 (N_11573,N_6773,N_7454);
or U11574 (N_11574,N_6521,N_7690);
and U11575 (N_11575,N_7607,N_7966);
nor U11576 (N_11576,N_6168,N_8572);
nor U11577 (N_11577,N_7343,N_6529);
or U11578 (N_11578,N_7447,N_6309);
or U11579 (N_11579,N_8380,N_8060);
or U11580 (N_11580,N_8074,N_7185);
and U11581 (N_11581,N_6755,N_6202);
nor U11582 (N_11582,N_6851,N_7051);
nor U11583 (N_11583,N_7038,N_8891);
nor U11584 (N_11584,N_6701,N_7916);
or U11585 (N_11585,N_8148,N_8109);
and U11586 (N_11586,N_8475,N_7079);
and U11587 (N_11587,N_6912,N_6060);
nand U11588 (N_11588,N_7659,N_7028);
nor U11589 (N_11589,N_7341,N_8003);
nor U11590 (N_11590,N_7245,N_7350);
nor U11591 (N_11591,N_8424,N_7888);
nor U11592 (N_11592,N_7115,N_8262);
and U11593 (N_11593,N_6360,N_6832);
and U11594 (N_11594,N_7632,N_7542);
nand U11595 (N_11595,N_7791,N_7792);
nand U11596 (N_11596,N_6484,N_8076);
and U11597 (N_11597,N_8291,N_7688);
and U11598 (N_11598,N_7645,N_6228);
xnor U11599 (N_11599,N_7736,N_7382);
nor U11600 (N_11600,N_8755,N_7439);
nor U11601 (N_11601,N_7106,N_6490);
nor U11602 (N_11602,N_6089,N_6313);
and U11603 (N_11603,N_6073,N_6332);
nand U11604 (N_11604,N_8534,N_6884);
or U11605 (N_11605,N_7135,N_8790);
or U11606 (N_11606,N_7158,N_7526);
nand U11607 (N_11607,N_8248,N_6852);
nand U11608 (N_11608,N_7042,N_6489);
and U11609 (N_11609,N_7861,N_7716);
and U11610 (N_11610,N_7544,N_7835);
or U11611 (N_11611,N_8570,N_7032);
nand U11612 (N_11612,N_6541,N_8046);
and U11613 (N_11613,N_7180,N_8595);
nor U11614 (N_11614,N_6648,N_7237);
nor U11615 (N_11615,N_8163,N_6627);
or U11616 (N_11616,N_7457,N_7747);
nand U11617 (N_11617,N_7026,N_7736);
nor U11618 (N_11618,N_7300,N_8204);
or U11619 (N_11619,N_7484,N_7943);
nand U11620 (N_11620,N_6638,N_8887);
nor U11621 (N_11621,N_8270,N_8346);
nand U11622 (N_11622,N_7020,N_8602);
nand U11623 (N_11623,N_6405,N_8010);
or U11624 (N_11624,N_8221,N_6495);
or U11625 (N_11625,N_6075,N_6531);
nand U11626 (N_11626,N_8756,N_6613);
and U11627 (N_11627,N_7850,N_8121);
nand U11628 (N_11628,N_7152,N_6986);
nand U11629 (N_11629,N_8522,N_7574);
nand U11630 (N_11630,N_8606,N_7458);
nor U11631 (N_11631,N_7005,N_6105);
nor U11632 (N_11632,N_6506,N_6993);
and U11633 (N_11633,N_7091,N_7340);
or U11634 (N_11634,N_7865,N_6387);
nor U11635 (N_11635,N_6404,N_8554);
or U11636 (N_11636,N_7330,N_8443);
and U11637 (N_11637,N_7885,N_7032);
and U11638 (N_11638,N_8015,N_7081);
nand U11639 (N_11639,N_6304,N_6679);
and U11640 (N_11640,N_7147,N_7193);
nor U11641 (N_11641,N_8653,N_8008);
nor U11642 (N_11642,N_8292,N_6616);
nand U11643 (N_11643,N_7435,N_8895);
nand U11644 (N_11644,N_6267,N_6318);
nand U11645 (N_11645,N_7621,N_6137);
or U11646 (N_11646,N_8582,N_6880);
or U11647 (N_11647,N_7586,N_8951);
xnor U11648 (N_11648,N_6373,N_7416);
or U11649 (N_11649,N_7589,N_6700);
or U11650 (N_11650,N_7644,N_7255);
nor U11651 (N_11651,N_7682,N_6781);
and U11652 (N_11652,N_8942,N_6948);
nor U11653 (N_11653,N_8300,N_8440);
nand U11654 (N_11654,N_6330,N_6637);
and U11655 (N_11655,N_7025,N_7169);
nand U11656 (N_11656,N_6330,N_7213);
xor U11657 (N_11657,N_6440,N_7357);
nor U11658 (N_11658,N_6541,N_8834);
nand U11659 (N_11659,N_7629,N_7402);
or U11660 (N_11660,N_8601,N_6386);
or U11661 (N_11661,N_7915,N_7429);
or U11662 (N_11662,N_6051,N_6258);
or U11663 (N_11663,N_6624,N_7325);
and U11664 (N_11664,N_6946,N_6454);
nand U11665 (N_11665,N_6742,N_8472);
and U11666 (N_11666,N_7557,N_6263);
and U11667 (N_11667,N_6764,N_6840);
or U11668 (N_11668,N_7733,N_6883);
nand U11669 (N_11669,N_6499,N_8105);
nor U11670 (N_11670,N_7256,N_6563);
and U11671 (N_11671,N_8659,N_7991);
nor U11672 (N_11672,N_7807,N_6546);
nand U11673 (N_11673,N_6768,N_8824);
xor U11674 (N_11674,N_8732,N_7581);
or U11675 (N_11675,N_8365,N_8289);
nand U11676 (N_11676,N_8561,N_8594);
or U11677 (N_11677,N_7364,N_6520);
or U11678 (N_11678,N_8507,N_7247);
nor U11679 (N_11679,N_6002,N_8505);
nor U11680 (N_11680,N_6106,N_7828);
or U11681 (N_11681,N_7083,N_6498);
and U11682 (N_11682,N_7595,N_8225);
and U11683 (N_11683,N_6834,N_7052);
or U11684 (N_11684,N_8702,N_8669);
and U11685 (N_11685,N_8473,N_8732);
nor U11686 (N_11686,N_6258,N_7883);
and U11687 (N_11687,N_7182,N_8858);
nor U11688 (N_11688,N_6438,N_8327);
nand U11689 (N_11689,N_7140,N_6009);
and U11690 (N_11690,N_8566,N_6420);
and U11691 (N_11691,N_8944,N_7952);
nand U11692 (N_11692,N_7818,N_8647);
and U11693 (N_11693,N_7250,N_8779);
or U11694 (N_11694,N_8005,N_8446);
or U11695 (N_11695,N_8187,N_7280);
and U11696 (N_11696,N_7734,N_8204);
or U11697 (N_11697,N_6234,N_7400);
nor U11698 (N_11698,N_7931,N_6177);
and U11699 (N_11699,N_8383,N_7614);
or U11700 (N_11700,N_7829,N_7605);
nor U11701 (N_11701,N_6343,N_6295);
or U11702 (N_11702,N_6634,N_7052);
or U11703 (N_11703,N_7060,N_6906);
nand U11704 (N_11704,N_7369,N_7939);
nor U11705 (N_11705,N_8858,N_7297);
and U11706 (N_11706,N_8284,N_8854);
and U11707 (N_11707,N_7373,N_8783);
nor U11708 (N_11708,N_8689,N_7411);
and U11709 (N_11709,N_6006,N_6858);
and U11710 (N_11710,N_8705,N_7772);
or U11711 (N_11711,N_8844,N_6268);
or U11712 (N_11712,N_7385,N_6148);
or U11713 (N_11713,N_8079,N_7977);
nor U11714 (N_11714,N_8423,N_7830);
nor U11715 (N_11715,N_8208,N_6363);
nor U11716 (N_11716,N_8133,N_6454);
nand U11717 (N_11717,N_7782,N_6057);
nor U11718 (N_11718,N_8456,N_6354);
or U11719 (N_11719,N_7564,N_6912);
and U11720 (N_11720,N_8249,N_7333);
or U11721 (N_11721,N_6584,N_7903);
nor U11722 (N_11722,N_6210,N_7977);
nor U11723 (N_11723,N_6719,N_8236);
or U11724 (N_11724,N_7352,N_7556);
xnor U11725 (N_11725,N_8211,N_6759);
or U11726 (N_11726,N_8337,N_7450);
nor U11727 (N_11727,N_7330,N_6125);
and U11728 (N_11728,N_6375,N_8267);
and U11729 (N_11729,N_8364,N_7751);
nor U11730 (N_11730,N_6409,N_6416);
nand U11731 (N_11731,N_7965,N_8662);
and U11732 (N_11732,N_8159,N_8618);
nand U11733 (N_11733,N_8870,N_8407);
nand U11734 (N_11734,N_6225,N_8004);
and U11735 (N_11735,N_8073,N_8693);
nand U11736 (N_11736,N_6054,N_8108);
nor U11737 (N_11737,N_6890,N_8787);
nand U11738 (N_11738,N_6723,N_7287);
nor U11739 (N_11739,N_7353,N_8302);
nor U11740 (N_11740,N_6498,N_8889);
and U11741 (N_11741,N_7971,N_8522);
and U11742 (N_11742,N_7785,N_6918);
nand U11743 (N_11743,N_6164,N_6300);
nor U11744 (N_11744,N_8156,N_8004);
and U11745 (N_11745,N_6326,N_6920);
or U11746 (N_11746,N_6546,N_6784);
nor U11747 (N_11747,N_6456,N_6592);
nand U11748 (N_11748,N_6039,N_6337);
or U11749 (N_11749,N_6533,N_7757);
or U11750 (N_11750,N_8220,N_6726);
and U11751 (N_11751,N_8987,N_7793);
nor U11752 (N_11752,N_8537,N_6843);
nor U11753 (N_11753,N_7619,N_7865);
or U11754 (N_11754,N_7800,N_6774);
nor U11755 (N_11755,N_6811,N_6652);
xor U11756 (N_11756,N_6363,N_6694);
or U11757 (N_11757,N_8652,N_8457);
or U11758 (N_11758,N_6912,N_8255);
or U11759 (N_11759,N_8415,N_6379);
xnor U11760 (N_11760,N_6832,N_8988);
nor U11761 (N_11761,N_8473,N_6048);
or U11762 (N_11762,N_7019,N_6027);
nand U11763 (N_11763,N_7434,N_8709);
nand U11764 (N_11764,N_6130,N_8500);
or U11765 (N_11765,N_7513,N_6487);
nand U11766 (N_11766,N_6767,N_6073);
or U11767 (N_11767,N_8653,N_7055);
nand U11768 (N_11768,N_6835,N_6227);
or U11769 (N_11769,N_6026,N_7533);
or U11770 (N_11770,N_8179,N_8582);
or U11771 (N_11771,N_6662,N_8655);
and U11772 (N_11772,N_7866,N_8698);
and U11773 (N_11773,N_6915,N_6663);
nor U11774 (N_11774,N_6405,N_7780);
nand U11775 (N_11775,N_6044,N_8582);
and U11776 (N_11776,N_6873,N_6644);
and U11777 (N_11777,N_6764,N_7368);
nand U11778 (N_11778,N_7803,N_6278);
nor U11779 (N_11779,N_8173,N_8077);
nor U11780 (N_11780,N_7636,N_8200);
nor U11781 (N_11781,N_7914,N_7936);
nand U11782 (N_11782,N_7256,N_6735);
nor U11783 (N_11783,N_7351,N_7252);
or U11784 (N_11784,N_6409,N_8652);
or U11785 (N_11785,N_8905,N_7423);
or U11786 (N_11786,N_6482,N_6368);
nand U11787 (N_11787,N_8100,N_6871);
and U11788 (N_11788,N_6663,N_7231);
and U11789 (N_11789,N_8640,N_6425);
and U11790 (N_11790,N_6538,N_7262);
nand U11791 (N_11791,N_6008,N_7808);
nand U11792 (N_11792,N_7869,N_8225);
or U11793 (N_11793,N_6107,N_7141);
nand U11794 (N_11794,N_6980,N_7946);
nand U11795 (N_11795,N_8412,N_8935);
and U11796 (N_11796,N_6397,N_8767);
or U11797 (N_11797,N_7041,N_7236);
or U11798 (N_11798,N_6495,N_6485);
or U11799 (N_11799,N_6386,N_6790);
nand U11800 (N_11800,N_7053,N_8776);
nor U11801 (N_11801,N_7165,N_6699);
or U11802 (N_11802,N_8711,N_8478);
or U11803 (N_11803,N_7965,N_6416);
nor U11804 (N_11804,N_7224,N_7780);
and U11805 (N_11805,N_8227,N_7836);
and U11806 (N_11806,N_8678,N_7468);
and U11807 (N_11807,N_6041,N_6236);
xor U11808 (N_11808,N_8140,N_8259);
and U11809 (N_11809,N_8954,N_8414);
nor U11810 (N_11810,N_7944,N_8112);
nor U11811 (N_11811,N_6775,N_7198);
nor U11812 (N_11812,N_6027,N_6555);
and U11813 (N_11813,N_6424,N_8280);
or U11814 (N_11814,N_7912,N_6336);
and U11815 (N_11815,N_8859,N_6768);
nand U11816 (N_11816,N_7297,N_7831);
nand U11817 (N_11817,N_7588,N_7396);
nand U11818 (N_11818,N_6941,N_6294);
and U11819 (N_11819,N_6049,N_7761);
or U11820 (N_11820,N_6842,N_8776);
nor U11821 (N_11821,N_8093,N_8228);
and U11822 (N_11822,N_7441,N_8415);
or U11823 (N_11823,N_6590,N_6228);
or U11824 (N_11824,N_8398,N_8169);
nand U11825 (N_11825,N_8342,N_7287);
nand U11826 (N_11826,N_6381,N_8656);
nor U11827 (N_11827,N_6730,N_8784);
or U11828 (N_11828,N_7985,N_8177);
nor U11829 (N_11829,N_8513,N_6176);
or U11830 (N_11830,N_8843,N_7965);
xor U11831 (N_11831,N_6240,N_8228);
nor U11832 (N_11832,N_7435,N_8199);
nor U11833 (N_11833,N_7903,N_7859);
or U11834 (N_11834,N_8005,N_7934);
or U11835 (N_11835,N_6957,N_6379);
or U11836 (N_11836,N_8064,N_8841);
nand U11837 (N_11837,N_8831,N_8224);
nor U11838 (N_11838,N_8042,N_7929);
and U11839 (N_11839,N_8690,N_7205);
nor U11840 (N_11840,N_6744,N_6370);
or U11841 (N_11841,N_8734,N_7479);
or U11842 (N_11842,N_8193,N_7510);
or U11843 (N_11843,N_6899,N_6503);
and U11844 (N_11844,N_7378,N_6408);
nand U11845 (N_11845,N_6155,N_8999);
and U11846 (N_11846,N_8867,N_8258);
and U11847 (N_11847,N_6416,N_7184);
nand U11848 (N_11848,N_6350,N_8800);
nand U11849 (N_11849,N_7904,N_7295);
or U11850 (N_11850,N_7018,N_7419);
xnor U11851 (N_11851,N_7586,N_7353);
nand U11852 (N_11852,N_7170,N_7901);
and U11853 (N_11853,N_6914,N_6001);
nor U11854 (N_11854,N_8335,N_7698);
and U11855 (N_11855,N_8100,N_8044);
nand U11856 (N_11856,N_7830,N_6411);
nand U11857 (N_11857,N_6952,N_6102);
and U11858 (N_11858,N_6594,N_6906);
and U11859 (N_11859,N_8943,N_8086);
and U11860 (N_11860,N_6392,N_8562);
nand U11861 (N_11861,N_7476,N_7447);
nand U11862 (N_11862,N_7547,N_7624);
nand U11863 (N_11863,N_7993,N_8551);
nor U11864 (N_11864,N_7653,N_8517);
nand U11865 (N_11865,N_8418,N_8207);
and U11866 (N_11866,N_8145,N_6926);
or U11867 (N_11867,N_8573,N_6438);
nand U11868 (N_11868,N_8167,N_6784);
or U11869 (N_11869,N_7908,N_8131);
and U11870 (N_11870,N_7888,N_8901);
and U11871 (N_11871,N_6038,N_6977);
nor U11872 (N_11872,N_6323,N_8516);
nor U11873 (N_11873,N_8962,N_7913);
nand U11874 (N_11874,N_7983,N_6109);
nor U11875 (N_11875,N_7231,N_8866);
and U11876 (N_11876,N_6483,N_7447);
nand U11877 (N_11877,N_7220,N_7896);
nor U11878 (N_11878,N_6811,N_8335);
nand U11879 (N_11879,N_8402,N_8220);
nand U11880 (N_11880,N_6296,N_7821);
nand U11881 (N_11881,N_8629,N_8914);
xnor U11882 (N_11882,N_7493,N_8797);
or U11883 (N_11883,N_8550,N_7424);
nor U11884 (N_11884,N_7143,N_6278);
nand U11885 (N_11885,N_6141,N_7848);
nand U11886 (N_11886,N_6765,N_7471);
nor U11887 (N_11887,N_6367,N_7200);
xor U11888 (N_11888,N_7592,N_8976);
and U11889 (N_11889,N_6375,N_8989);
or U11890 (N_11890,N_7060,N_8378);
nand U11891 (N_11891,N_7768,N_8893);
and U11892 (N_11892,N_8508,N_7234);
or U11893 (N_11893,N_7984,N_7807);
and U11894 (N_11894,N_7635,N_7318);
xor U11895 (N_11895,N_7056,N_6519);
or U11896 (N_11896,N_8719,N_6918);
xor U11897 (N_11897,N_6581,N_7009);
and U11898 (N_11898,N_6421,N_8588);
nand U11899 (N_11899,N_8991,N_8842);
nor U11900 (N_11900,N_6753,N_6525);
nand U11901 (N_11901,N_6972,N_7691);
nor U11902 (N_11902,N_6250,N_6866);
and U11903 (N_11903,N_6047,N_6717);
nor U11904 (N_11904,N_6335,N_6620);
nor U11905 (N_11905,N_7378,N_7560);
and U11906 (N_11906,N_7285,N_6290);
nand U11907 (N_11907,N_7238,N_6615);
nand U11908 (N_11908,N_8611,N_7826);
or U11909 (N_11909,N_8199,N_8733);
nor U11910 (N_11910,N_7205,N_6331);
or U11911 (N_11911,N_7687,N_8520);
or U11912 (N_11912,N_6922,N_7565);
nor U11913 (N_11913,N_6247,N_8896);
and U11914 (N_11914,N_8198,N_6960);
nand U11915 (N_11915,N_8342,N_8776);
nor U11916 (N_11916,N_7053,N_6080);
nor U11917 (N_11917,N_7096,N_8446);
nand U11918 (N_11918,N_7171,N_7568);
and U11919 (N_11919,N_6835,N_8560);
or U11920 (N_11920,N_7736,N_6874);
nor U11921 (N_11921,N_7262,N_7264);
or U11922 (N_11922,N_6894,N_8976);
or U11923 (N_11923,N_8045,N_7070);
and U11924 (N_11924,N_8370,N_7068);
nor U11925 (N_11925,N_7685,N_6328);
and U11926 (N_11926,N_8672,N_8167);
nor U11927 (N_11927,N_6001,N_8832);
nand U11928 (N_11928,N_8182,N_7833);
and U11929 (N_11929,N_7003,N_7521);
and U11930 (N_11930,N_7877,N_7276);
xor U11931 (N_11931,N_6627,N_8164);
and U11932 (N_11932,N_8960,N_7488);
or U11933 (N_11933,N_7991,N_7008);
and U11934 (N_11934,N_8270,N_7256);
or U11935 (N_11935,N_7167,N_7451);
and U11936 (N_11936,N_7815,N_7188);
or U11937 (N_11937,N_6607,N_8459);
and U11938 (N_11938,N_6140,N_8697);
nand U11939 (N_11939,N_7046,N_8994);
nor U11940 (N_11940,N_7041,N_8628);
xor U11941 (N_11941,N_6330,N_7441);
nor U11942 (N_11942,N_6650,N_8998);
nand U11943 (N_11943,N_6133,N_7058);
or U11944 (N_11944,N_7206,N_7427);
nand U11945 (N_11945,N_8217,N_7453);
nand U11946 (N_11946,N_8831,N_6331);
nor U11947 (N_11947,N_6471,N_8710);
or U11948 (N_11948,N_6119,N_7002);
and U11949 (N_11949,N_8687,N_8187);
nand U11950 (N_11950,N_6100,N_6174);
nor U11951 (N_11951,N_8261,N_7659);
nand U11952 (N_11952,N_8364,N_7371);
nor U11953 (N_11953,N_7973,N_8649);
nand U11954 (N_11954,N_8640,N_7037);
nor U11955 (N_11955,N_8597,N_8332);
and U11956 (N_11956,N_8133,N_6960);
nor U11957 (N_11957,N_6229,N_8799);
or U11958 (N_11958,N_6261,N_6303);
nand U11959 (N_11959,N_7431,N_7630);
xor U11960 (N_11960,N_8686,N_7858);
and U11961 (N_11961,N_7812,N_7015);
or U11962 (N_11962,N_6497,N_8665);
or U11963 (N_11963,N_7107,N_8215);
and U11964 (N_11964,N_7601,N_8969);
nor U11965 (N_11965,N_8611,N_7628);
or U11966 (N_11966,N_8614,N_8671);
nor U11967 (N_11967,N_7425,N_8550);
or U11968 (N_11968,N_6909,N_6051);
and U11969 (N_11969,N_8154,N_6312);
and U11970 (N_11970,N_7690,N_8566);
and U11971 (N_11971,N_7914,N_6411);
xnor U11972 (N_11972,N_7001,N_6002);
and U11973 (N_11973,N_8124,N_6016);
nand U11974 (N_11974,N_8224,N_7863);
nand U11975 (N_11975,N_6042,N_8928);
and U11976 (N_11976,N_7336,N_6636);
or U11977 (N_11977,N_6512,N_6732);
or U11978 (N_11978,N_8127,N_8521);
nand U11979 (N_11979,N_8325,N_7059);
and U11980 (N_11980,N_8879,N_6400);
and U11981 (N_11981,N_6370,N_6262);
nor U11982 (N_11982,N_6931,N_8408);
or U11983 (N_11983,N_7301,N_8761);
nand U11984 (N_11984,N_8246,N_8100);
or U11985 (N_11985,N_7493,N_7581);
or U11986 (N_11986,N_6178,N_6342);
nor U11987 (N_11987,N_7762,N_8562);
and U11988 (N_11988,N_7069,N_8982);
xor U11989 (N_11989,N_6543,N_8516);
nand U11990 (N_11990,N_6313,N_6333);
nand U11991 (N_11991,N_6891,N_7046);
nor U11992 (N_11992,N_8467,N_7680);
nor U11993 (N_11993,N_8043,N_8423);
nor U11994 (N_11994,N_7406,N_7805);
nand U11995 (N_11995,N_6648,N_7856);
nor U11996 (N_11996,N_6664,N_8830);
nor U11997 (N_11997,N_6703,N_7101);
nand U11998 (N_11998,N_8480,N_7283);
nand U11999 (N_11999,N_7276,N_7419);
nor U12000 (N_12000,N_11982,N_10429);
nand U12001 (N_12001,N_10888,N_9566);
nand U12002 (N_12002,N_11954,N_11064);
or U12003 (N_12003,N_10372,N_11917);
nor U12004 (N_12004,N_9239,N_11183);
and U12005 (N_12005,N_9131,N_9297);
and U12006 (N_12006,N_11358,N_11531);
nand U12007 (N_12007,N_10725,N_9611);
or U12008 (N_12008,N_10179,N_10420);
xnor U12009 (N_12009,N_11411,N_11245);
and U12010 (N_12010,N_10640,N_11243);
and U12011 (N_12011,N_11153,N_9561);
nand U12012 (N_12012,N_9232,N_9456);
xnor U12013 (N_12013,N_9783,N_9903);
nor U12014 (N_12014,N_9393,N_11686);
nor U12015 (N_12015,N_11990,N_9021);
or U12016 (N_12016,N_9996,N_9159);
and U12017 (N_12017,N_11994,N_11258);
and U12018 (N_12018,N_11928,N_9374);
nand U12019 (N_12019,N_11360,N_9137);
or U12020 (N_12020,N_10434,N_10439);
or U12021 (N_12021,N_9043,N_10245);
or U12022 (N_12022,N_11938,N_11627);
or U12023 (N_12023,N_9258,N_11577);
nor U12024 (N_12024,N_10384,N_10298);
nand U12025 (N_12025,N_11366,N_11875);
nand U12026 (N_12026,N_9375,N_11911);
nor U12027 (N_12027,N_9099,N_11563);
and U12028 (N_12028,N_9146,N_10403);
nor U12029 (N_12029,N_11225,N_10806);
nor U12030 (N_12030,N_11675,N_11651);
and U12031 (N_12031,N_11777,N_9116);
or U12032 (N_12032,N_10023,N_11302);
and U12033 (N_12033,N_9005,N_9169);
or U12034 (N_12034,N_9778,N_9488);
nor U12035 (N_12035,N_10927,N_9390);
nand U12036 (N_12036,N_9040,N_10968);
or U12037 (N_12037,N_11019,N_11043);
nand U12038 (N_12038,N_10648,N_10087);
nand U12039 (N_12039,N_9529,N_11680);
nand U12040 (N_12040,N_11771,N_9802);
nand U12041 (N_12041,N_11658,N_9145);
nor U12042 (N_12042,N_11539,N_10558);
nor U12043 (N_12043,N_9072,N_11461);
xor U12044 (N_12044,N_9753,N_10543);
and U12045 (N_12045,N_9752,N_10870);
nand U12046 (N_12046,N_11889,N_11780);
or U12047 (N_12047,N_11620,N_9853);
or U12048 (N_12048,N_10821,N_11697);
and U12049 (N_12049,N_10180,N_11608);
nand U12050 (N_12050,N_9787,N_9246);
nand U12051 (N_12051,N_11858,N_10122);
nand U12052 (N_12052,N_9054,N_10794);
nor U12053 (N_12053,N_10526,N_9893);
nor U12054 (N_12054,N_11457,N_9167);
nand U12055 (N_12055,N_10534,N_11552);
nor U12056 (N_12056,N_11405,N_10528);
or U12057 (N_12057,N_11262,N_10343);
or U12058 (N_12058,N_11960,N_9846);
or U12059 (N_12059,N_9793,N_11385);
nor U12060 (N_12060,N_11321,N_11486);
and U12061 (N_12061,N_10547,N_10132);
nand U12062 (N_12062,N_10818,N_9245);
nor U12063 (N_12063,N_9217,N_11103);
nor U12064 (N_12064,N_9707,N_9823);
nor U12065 (N_12065,N_11499,N_11713);
and U12066 (N_12066,N_11930,N_11794);
nor U12067 (N_12067,N_10017,N_10746);
nand U12068 (N_12068,N_9838,N_11547);
or U12069 (N_12069,N_11899,N_9808);
or U12070 (N_12070,N_11284,N_10684);
or U12071 (N_12071,N_10586,N_9209);
nand U12072 (N_12072,N_9990,N_10082);
or U12073 (N_12073,N_10771,N_11348);
or U12074 (N_12074,N_9000,N_10931);
or U12075 (N_12075,N_9182,N_10598);
or U12076 (N_12076,N_9136,N_11801);
nor U12077 (N_12077,N_11334,N_10871);
nand U12078 (N_12078,N_9966,N_11255);
and U12079 (N_12079,N_11747,N_11033);
or U12080 (N_12080,N_11212,N_11710);
or U12081 (N_12081,N_11407,N_10109);
nor U12082 (N_12082,N_9337,N_11687);
nand U12083 (N_12083,N_10945,N_11134);
or U12084 (N_12084,N_11616,N_10016);
or U12085 (N_12085,N_11751,N_11571);
nand U12086 (N_12086,N_9888,N_11646);
nand U12087 (N_12087,N_10444,N_10233);
and U12088 (N_12088,N_10290,N_10212);
nand U12089 (N_12089,N_10568,N_9304);
nand U12090 (N_12090,N_9833,N_9979);
nand U12091 (N_12091,N_11736,N_10786);
nor U12092 (N_12092,N_9497,N_10501);
nor U12093 (N_12093,N_10302,N_11685);
xnor U12094 (N_12094,N_10916,N_9770);
nor U12095 (N_12095,N_11723,N_11410);
or U12096 (N_12096,N_11108,N_11843);
or U12097 (N_12097,N_9100,N_10485);
nand U12098 (N_12098,N_10912,N_10032);
or U12099 (N_12099,N_9719,N_9762);
or U12100 (N_12100,N_9689,N_9178);
nor U12101 (N_12101,N_9960,N_10317);
xor U12102 (N_12102,N_10440,N_11576);
nor U12103 (N_12103,N_11980,N_10637);
nand U12104 (N_12104,N_10563,N_9621);
nand U12105 (N_12105,N_9610,N_11691);
nor U12106 (N_12106,N_10597,N_10987);
and U12107 (N_12107,N_11196,N_11223);
and U12108 (N_12108,N_9803,N_9494);
nor U12109 (N_12109,N_9103,N_11417);
or U12110 (N_12110,N_9053,N_9475);
or U12111 (N_12111,N_10483,N_10405);
nand U12112 (N_12112,N_9837,N_9505);
or U12113 (N_12113,N_11080,N_11684);
and U12114 (N_12114,N_11682,N_9491);
and U12115 (N_12115,N_10837,N_9757);
nor U12116 (N_12116,N_11762,N_10276);
and U12117 (N_12117,N_11944,N_10866);
or U12118 (N_12118,N_10634,N_11275);
nor U12119 (N_12119,N_10116,N_9037);
and U12120 (N_12120,N_9588,N_10519);
nand U12121 (N_12121,N_10129,N_10283);
nand U12122 (N_12122,N_9578,N_9076);
and U12123 (N_12123,N_11190,N_9704);
nor U12124 (N_12124,N_9740,N_10869);
and U12125 (N_12125,N_9210,N_11048);
nand U12126 (N_12126,N_10636,N_10432);
nand U12127 (N_12127,N_9344,N_9300);
nor U12128 (N_12128,N_9222,N_9089);
or U12129 (N_12129,N_11449,N_10120);
nor U12130 (N_12130,N_11227,N_9556);
nor U12131 (N_12131,N_10450,N_10578);
nand U12132 (N_12132,N_9627,N_11157);
or U12133 (N_12133,N_9964,N_10537);
nand U12134 (N_12134,N_11289,N_9503);
nor U12135 (N_12135,N_9788,N_11343);
or U12136 (N_12136,N_10493,N_9568);
or U12137 (N_12137,N_10666,N_11003);
or U12138 (N_12138,N_11965,N_9854);
or U12139 (N_12139,N_11995,N_10781);
nand U12140 (N_12140,N_9359,N_11611);
or U12141 (N_12141,N_10565,N_11543);
or U12142 (N_12142,N_9316,N_10386);
xor U12143 (N_12143,N_10264,N_10961);
or U12144 (N_12144,N_10373,N_10995);
nand U12145 (N_12145,N_10095,N_10754);
or U12146 (N_12146,N_11739,N_11176);
nand U12147 (N_12147,N_10893,N_11708);
and U12148 (N_12148,N_10123,N_9800);
or U12149 (N_12149,N_10426,N_10993);
and U12150 (N_12150,N_11919,N_11890);
and U12151 (N_12151,N_10166,N_10335);
nand U12152 (N_12152,N_9512,N_10353);
xnor U12153 (N_12153,N_10988,N_9867);
or U12154 (N_12154,N_10554,N_9738);
or U12155 (N_12155,N_9332,N_10864);
nor U12156 (N_12156,N_9051,N_10235);
nor U12157 (N_12157,N_9306,N_9825);
nand U12158 (N_12158,N_10887,N_9420);
nor U12159 (N_12159,N_10607,N_11783);
or U12160 (N_12160,N_10813,N_11831);
xor U12161 (N_12161,N_9013,N_9114);
nor U12162 (N_12162,N_10058,N_11955);
and U12163 (N_12163,N_10532,N_9541);
or U12164 (N_12164,N_10329,N_11841);
nand U12165 (N_12165,N_10203,N_10530);
nand U12166 (N_12166,N_11718,N_11342);
nand U12167 (N_12167,N_11291,N_9220);
and U12168 (N_12168,N_11396,N_10743);
nor U12169 (N_12169,N_9642,N_11894);
or U12170 (N_12170,N_9913,N_11098);
and U12171 (N_12171,N_11162,N_9672);
or U12172 (N_12172,N_9955,N_9458);
or U12173 (N_12173,N_9731,N_11614);
nor U12174 (N_12174,N_11453,N_9322);
nand U12175 (N_12175,N_9083,N_11881);
or U12176 (N_12176,N_9760,N_10117);
or U12177 (N_12177,N_9668,N_9171);
or U12178 (N_12178,N_11170,N_11617);
and U12179 (N_12179,N_10655,N_9685);
or U12180 (N_12180,N_10936,N_11720);
and U12181 (N_12181,N_10823,N_10567);
or U12182 (N_12182,N_9267,N_11203);
or U12183 (N_12183,N_9292,N_10632);
nand U12184 (N_12184,N_10847,N_10728);
or U12185 (N_12185,N_9408,N_11250);
and U12186 (N_12186,N_10822,N_10247);
and U12187 (N_12187,N_9001,N_11025);
or U12188 (N_12188,N_10121,N_9038);
nand U12189 (N_12189,N_10748,N_10992);
or U12190 (N_12190,N_11529,N_11676);
nand U12191 (N_12191,N_10240,N_11032);
or U12192 (N_12192,N_10625,N_10659);
and U12193 (N_12193,N_10626,N_10839);
nand U12194 (N_12194,N_9667,N_11042);
or U12195 (N_12195,N_9724,N_9057);
or U12196 (N_12196,N_9933,N_10348);
or U12197 (N_12197,N_11905,N_9922);
nand U12198 (N_12198,N_10792,N_10587);
nand U12199 (N_12199,N_11422,N_9864);
nand U12200 (N_12200,N_9695,N_9443);
nand U12201 (N_12201,N_11288,N_9563);
nand U12202 (N_12202,N_11404,N_10480);
nand U12203 (N_12203,N_11705,N_11711);
or U12204 (N_12204,N_10722,N_9533);
nand U12205 (N_12205,N_10727,N_9781);
and U12206 (N_12206,N_9474,N_9774);
or U12207 (N_12207,N_11068,N_9839);
nand U12208 (N_12208,N_10478,N_11833);
nor U12209 (N_12209,N_10257,N_10422);
nor U12210 (N_12210,N_11013,N_9127);
or U12211 (N_12211,N_9354,N_11824);
nand U12212 (N_12212,N_11773,N_10458);
nor U12213 (N_12213,N_11607,N_10631);
nor U12214 (N_12214,N_10555,N_10072);
or U12215 (N_12215,N_9438,N_10843);
nand U12216 (N_12216,N_9799,N_10063);
or U12217 (N_12217,N_10454,N_9550);
nand U12218 (N_12218,N_11029,N_9705);
or U12219 (N_12219,N_11659,N_10374);
nand U12220 (N_12220,N_10521,N_11173);
and U12221 (N_12221,N_10595,N_10499);
nand U12222 (N_12222,N_9382,N_11765);
and U12223 (N_12223,N_9652,N_9489);
and U12224 (N_12224,N_11985,N_9660);
and U12225 (N_12225,N_10889,N_9834);
nand U12226 (N_12226,N_11340,N_11163);
nand U12227 (N_12227,N_11290,N_9993);
and U12228 (N_12228,N_10341,N_10160);
or U12229 (N_12229,N_10602,N_9502);
nand U12230 (N_12230,N_11946,N_9930);
nor U12231 (N_12231,N_11267,N_11998);
nor U12232 (N_12232,N_9792,N_10211);
or U12233 (N_12233,N_9714,N_9938);
nor U12234 (N_12234,N_9481,N_9397);
nor U12235 (N_12235,N_9727,N_10327);
or U12236 (N_12236,N_9863,N_9650);
nand U12237 (N_12237,N_11696,N_11601);
nor U12238 (N_12238,N_10672,N_9543);
or U12239 (N_12239,N_9994,N_10738);
nor U12240 (N_12240,N_10114,N_10919);
and U12241 (N_12241,N_11778,N_11933);
xor U12242 (N_12242,N_11512,N_9343);
xor U12243 (N_12243,N_9284,N_10219);
and U12244 (N_12244,N_11505,N_9177);
or U12245 (N_12245,N_9634,N_9873);
nand U12246 (N_12246,N_10879,N_11363);
xnor U12247 (N_12247,N_9790,N_11692);
or U12248 (N_12248,N_11187,N_9936);
and U12249 (N_12249,N_10783,N_11528);
or U12250 (N_12250,N_9969,N_10028);
and U12251 (N_12251,N_9765,N_10278);
nor U12252 (N_12252,N_9551,N_10724);
nor U12253 (N_12253,N_11690,N_9624);
and U12254 (N_12254,N_9287,N_9965);
or U12255 (N_12255,N_9951,N_10868);
nand U12256 (N_12256,N_10394,N_9391);
nor U12257 (N_12257,N_9142,N_9882);
or U12258 (N_12258,N_10577,N_11230);
or U12259 (N_12259,N_11594,N_10898);
nor U12260 (N_12260,N_10044,N_10065);
nand U12261 (N_12261,N_9646,N_9439);
nand U12262 (N_12262,N_11509,N_11458);
and U12263 (N_12263,N_10662,N_9315);
and U12264 (N_12264,N_9927,N_9449);
or U12265 (N_12265,N_10030,N_10717);
and U12266 (N_12266,N_9579,N_9835);
nor U12267 (N_12267,N_11981,N_9176);
nand U12268 (N_12268,N_11179,N_10610);
or U12269 (N_12269,N_10891,N_11737);
or U12270 (N_12270,N_9451,N_10934);
nor U12271 (N_12271,N_11660,N_10046);
nor U12272 (N_12272,N_11971,N_10024);
nand U12273 (N_12273,N_10875,N_11122);
and U12274 (N_12274,N_9797,N_9776);
nor U12275 (N_12275,N_10273,N_11090);
nand U12276 (N_12276,N_9892,N_11439);
nand U12277 (N_12277,N_10294,N_10066);
or U12278 (N_12278,N_9971,N_11605);
or U12279 (N_12279,N_10098,N_11525);
and U12280 (N_12280,N_10050,N_11425);
and U12281 (N_12281,N_11236,N_9656);
nand U12282 (N_12282,N_9891,N_9036);
nor U12283 (N_12283,N_9164,N_10291);
and U12284 (N_12284,N_11118,N_9047);
nor U12285 (N_12285,N_11319,N_9592);
or U12286 (N_12286,N_9278,N_11473);
or U12287 (N_12287,N_9694,N_10107);
or U12288 (N_12288,N_9952,N_9745);
and U12289 (N_12289,N_10943,N_9432);
and U12290 (N_12290,N_10108,N_9985);
and U12291 (N_12291,N_11888,N_11333);
and U12292 (N_12292,N_9218,N_9252);
nor U12293 (N_12293,N_11560,N_9128);
and U12294 (N_12294,N_11892,N_10979);
nand U12295 (N_12295,N_10363,N_10141);
and U12296 (N_12296,N_11202,N_11146);
and U12297 (N_12297,N_11572,N_10209);
or U12298 (N_12298,N_10337,N_9593);
or U12299 (N_12299,N_10126,N_10999);
nor U12300 (N_12300,N_11991,N_10653);
nor U12301 (N_12301,N_11872,N_9004);
nand U12302 (N_12302,N_10364,N_9415);
nor U12303 (N_12303,N_11311,N_10709);
nand U12304 (N_12304,N_11306,N_9862);
nor U12305 (N_12305,N_10917,N_11785);
nand U12306 (N_12306,N_10315,N_10125);
or U12307 (N_12307,N_10884,N_9605);
nor U12308 (N_12308,N_11372,N_9812);
nand U12309 (N_12309,N_10789,N_11533);
and U12310 (N_12310,N_11564,N_9842);
nor U12311 (N_12311,N_10639,N_11702);
nand U12312 (N_12312,N_11735,N_10407);
xnor U12313 (N_12313,N_9305,N_9470);
nand U12314 (N_12314,N_9747,N_10347);
or U12315 (N_12315,N_10608,N_11167);
and U12316 (N_12316,N_10649,N_11078);
nor U12317 (N_12317,N_10835,N_10881);
nand U12318 (N_12318,N_10520,N_11062);
and U12319 (N_12319,N_11506,N_9299);
and U12320 (N_12320,N_11770,N_11796);
and U12321 (N_12321,N_11234,N_10859);
nor U12322 (N_12322,N_10241,N_11352);
and U12323 (N_12323,N_11790,N_10045);
or U12324 (N_12324,N_11268,N_9381);
xor U12325 (N_12325,N_9373,N_11839);
and U12326 (N_12326,N_11624,N_10712);
and U12327 (N_12327,N_11272,N_10707);
nand U12328 (N_12328,N_11757,N_9016);
nor U12329 (N_12329,N_10105,N_9437);
nor U12330 (N_12330,N_11959,N_10047);
or U12331 (N_12331,N_9830,N_9338);
and U12332 (N_12332,N_9163,N_9919);
or U12333 (N_12333,N_10756,N_11475);
nand U12334 (N_12334,N_10720,N_9982);
and U12335 (N_12335,N_10198,N_9582);
nand U12336 (N_12336,N_11656,N_9251);
nand U12337 (N_12337,N_10067,N_9387);
xnor U12338 (N_12338,N_10338,N_9386);
nand U12339 (N_12339,N_10675,N_11084);
nand U12340 (N_12340,N_9763,N_10162);
nor U12341 (N_12341,N_9257,N_9378);
and U12342 (N_12342,N_9355,N_11591);
and U12343 (N_12343,N_9150,N_10421);
xnor U12344 (N_12344,N_9670,N_11004);
nor U12345 (N_12345,N_9786,N_10400);
nor U12346 (N_12346,N_11018,N_9976);
xor U12347 (N_12347,N_10767,N_11421);
and U12348 (N_12348,N_11077,N_9754);
or U12349 (N_12349,N_11148,N_9447);
nand U12350 (N_12350,N_11673,N_11805);
and U12351 (N_12351,N_10031,N_9268);
nand U12352 (N_12352,N_10591,N_9463);
nor U12353 (N_12353,N_10310,N_11063);
nand U12354 (N_12354,N_9585,N_11443);
or U12355 (N_12355,N_11244,N_9140);
or U12356 (N_12356,N_9755,N_11559);
nand U12357 (N_12357,N_10115,N_10185);
or U12358 (N_12358,N_9430,N_10011);
nor U12359 (N_12359,N_10583,N_11054);
or U12360 (N_12360,N_9603,N_11067);
or U12361 (N_12361,N_11393,N_10303);
nand U12362 (N_12362,N_10124,N_11432);
nor U12363 (N_12363,N_9874,N_11436);
or U12364 (N_12364,N_9682,N_10680);
nor U12365 (N_12365,N_11768,N_11040);
or U12366 (N_12366,N_9241,N_11482);
and U12367 (N_12367,N_9347,N_10503);
or U12368 (N_12368,N_11200,N_10167);
nor U12369 (N_12369,N_11679,N_9207);
and U12370 (N_12370,N_11265,N_11039);
nand U12371 (N_12371,N_10852,N_9195);
or U12372 (N_12372,N_9225,N_11451);
and U12373 (N_12373,N_10260,N_10950);
xor U12374 (N_12374,N_10330,N_9017);
nor U12375 (N_12375,N_11270,N_10603);
and U12376 (N_12376,N_9926,N_11117);
and U12377 (N_12377,N_11566,N_9581);
nand U12378 (N_12378,N_9523,N_10252);
or U12379 (N_12379,N_10571,N_9819);
or U12380 (N_12380,N_10614,N_9844);
or U12381 (N_12381,N_9698,N_10234);
or U12382 (N_12382,N_9120,N_10404);
or U12383 (N_12383,N_9484,N_9352);
nor U12384 (N_12384,N_10750,N_9622);
or U12385 (N_12385,N_10790,N_9206);
and U12386 (N_12386,N_10208,N_10361);
or U12387 (N_12387,N_10763,N_9690);
nand U12388 (N_12388,N_10923,N_11584);
or U12389 (N_12389,N_9925,N_9877);
nor U12390 (N_12390,N_11815,N_11469);
nor U12391 (N_12391,N_11222,N_9791);
and U12392 (N_12392,N_10542,N_10736);
and U12393 (N_12393,N_9730,N_10305);
and U12394 (N_12394,N_9321,N_11631);
nor U12395 (N_12395,N_9018,N_11415);
nor U12396 (N_12396,N_9875,N_9843);
or U12397 (N_12397,N_9370,N_11721);
or U12398 (N_12398,N_10101,N_9905);
or U12399 (N_12399,N_11857,N_11695);
and U12400 (N_12400,N_11851,N_10815);
or U12401 (N_12401,N_9483,N_9006);
nand U12402 (N_12402,N_11859,N_9441);
nand U12403 (N_12403,N_10076,N_10069);
xor U12404 (N_12404,N_10388,N_10183);
and U12405 (N_12405,N_10716,N_10894);
or U12406 (N_12406,N_10304,N_9202);
nor U12407 (N_12407,N_11688,N_10991);
or U12408 (N_12408,N_11021,N_11279);
and U12409 (N_12409,N_9594,N_10617);
or U12410 (N_12410,N_10104,N_9186);
and U12411 (N_12411,N_10863,N_10842);
nand U12412 (N_12412,N_10490,N_11915);
nand U12413 (N_12413,N_10702,N_10787);
or U12414 (N_12414,N_10187,N_9900);
and U12415 (N_12415,N_9193,N_10773);
and U12416 (N_12416,N_9166,N_10110);
nand U12417 (N_12417,N_9115,N_11388);
and U12418 (N_12418,N_11952,N_10477);
and U12419 (N_12419,N_10090,N_9860);
and U12420 (N_12420,N_10574,N_11072);
nand U12421 (N_12421,N_10119,N_11112);
nor U12422 (N_12422,N_10594,N_10535);
or U12423 (N_12423,N_10230,N_10883);
or U12424 (N_12424,N_9733,N_10522);
nor U12425 (N_12425,N_11782,N_11105);
or U12426 (N_12426,N_9263,N_11536);
or U12427 (N_12427,N_11438,N_11485);
or U12428 (N_12428,N_11286,N_11207);
nor U12429 (N_12429,N_10370,N_11650);
nor U12430 (N_12430,N_11570,N_9535);
nand U12431 (N_12431,N_11500,N_11440);
xor U12432 (N_12432,N_11958,N_10573);
and U12433 (N_12433,N_11487,N_9929);
nand U12434 (N_12434,N_9924,N_9644);
nor U12435 (N_12435,N_10819,N_11184);
nand U12436 (N_12436,N_9619,N_11725);
and U12437 (N_12437,N_9673,N_11802);
nand U12438 (N_12438,N_11391,N_11376);
nand U12439 (N_12439,N_10612,N_10003);
and U12440 (N_12440,N_11037,N_9199);
nand U12441 (N_12441,N_10613,N_10645);
nand U12442 (N_12442,N_11256,N_10137);
nand U12443 (N_12443,N_10825,N_9172);
nand U12444 (N_12444,N_11337,N_10469);
or U12445 (N_12445,N_11086,N_9360);
or U12446 (N_12446,N_10643,N_9857);
nor U12447 (N_12447,N_11674,N_11807);
nand U12448 (N_12448,N_9628,N_9106);
nand U12449 (N_12449,N_10502,N_9970);
nand U12450 (N_12450,N_9935,N_10377);
or U12451 (N_12451,N_10663,N_10733);
nand U12452 (N_12452,N_9967,N_11527);
or U12453 (N_12453,N_9383,N_9680);
nor U12454 (N_12454,N_11093,N_10557);
or U12455 (N_12455,N_11502,N_11942);
nand U12456 (N_12456,N_9009,N_10606);
nand U12457 (N_12457,N_9155,N_11830);
nor U12458 (N_12458,N_11215,N_9804);
nand U12459 (N_12459,N_10641,N_10669);
and U12460 (N_12460,N_9423,N_10500);
nor U12461 (N_12461,N_10697,N_10147);
nor U12462 (N_12462,N_11515,N_11192);
nor U12463 (N_12463,N_11643,N_9950);
nand U12464 (N_12464,N_9637,N_10286);
nand U12465 (N_12465,N_9462,N_11082);
nor U12466 (N_12466,N_11992,N_9912);
nor U12467 (N_12467,N_11657,N_10957);
and U12468 (N_12468,N_11392,N_9840);
nand U12469 (N_12469,N_9596,N_9324);
and U12470 (N_12470,N_9331,N_11495);
and U12471 (N_12471,N_10168,N_10100);
nand U12472 (N_12472,N_11494,N_9358);
and U12473 (N_12473,N_9460,N_9191);
and U12474 (N_12474,N_10638,N_10963);
and U12475 (N_12475,N_10599,N_10904);
nor U12476 (N_12476,N_11140,N_9767);
and U12477 (N_12477,N_10425,N_9020);
nand U12478 (N_12478,N_9384,N_9564);
nor U12479 (N_12479,N_11518,N_10517);
or U12480 (N_12480,N_10080,N_10473);
or U12481 (N_12481,N_11767,N_11452);
and U12482 (N_12482,N_11367,N_11371);
or U12483 (N_12483,N_9998,N_10250);
or U12484 (N_12484,N_11497,N_11836);
or U12485 (N_12485,N_9417,N_9785);
and U12486 (N_12486,N_11613,N_10505);
and U12487 (N_12487,N_9075,N_10552);
nor U12488 (N_12488,N_11544,N_10106);
or U12489 (N_12489,N_10002,N_10415);
nor U12490 (N_12490,N_10958,N_9519);
nand U12491 (N_12491,N_10062,N_9796);
and U12492 (N_12492,N_9144,N_9188);
or U12493 (N_12493,N_10512,N_11488);
nand U12494 (N_12494,N_9729,N_11984);
nor U12495 (N_12495,N_9546,N_10188);
or U12496 (N_12496,N_10464,N_9537);
or U12497 (N_12497,N_10296,N_10381);
and U12498 (N_12498,N_10651,N_11731);
and U12499 (N_12499,N_11310,N_10757);
nand U12500 (N_12500,N_10671,N_11678);
or U12501 (N_12501,N_10205,N_11556);
nor U12502 (N_12502,N_9118,N_11041);
or U12503 (N_12503,N_10022,N_11880);
nor U12504 (N_12504,N_11891,N_11640);
nor U12505 (N_12505,N_11354,N_11848);
nor U12506 (N_12506,N_9279,N_9577);
or U12507 (N_12507,N_9722,N_10686);
and U12508 (N_12508,N_11280,N_10548);
and U12509 (N_12509,N_11699,N_11939);
nor U12510 (N_12510,N_11182,N_11530);
nand U12511 (N_12511,N_9702,N_10545);
xnor U12512 (N_12512,N_11951,N_10202);
nor U12513 (N_12513,N_9055,N_11592);
nand U12514 (N_12514,N_9229,N_11877);
or U12515 (N_12515,N_9431,N_11430);
nor U12516 (N_12516,N_10433,N_10592);
nand U12517 (N_12517,N_11171,N_9542);
nand U12518 (N_12518,N_11408,N_9204);
nor U12519 (N_12519,N_10165,N_11997);
nand U12520 (N_12520,N_11524,N_9356);
nand U12521 (N_12521,N_9265,N_10383);
xor U12522 (N_12522,N_11621,N_10497);
and U12523 (N_12523,N_11743,N_11057);
and U12524 (N_12524,N_10518,N_11921);
or U12525 (N_12525,N_11373,N_11361);
or U12526 (N_12526,N_10744,N_11826);
nand U12527 (N_12527,N_11870,N_11323);
nand U12528 (N_12528,N_10081,N_9310);
and U12529 (N_12529,N_9986,N_9440);
xnor U12530 (N_12530,N_10035,N_11834);
nand U12531 (N_12531,N_9398,N_11844);
and U12532 (N_12532,N_10873,N_10449);
nor U12533 (N_12533,N_9631,N_10997);
nor U12534 (N_12534,N_9389,N_11719);
and U12535 (N_12535,N_9980,N_11876);
or U12536 (N_12536,N_9269,N_10368);
and U12537 (N_12537,N_10005,N_11867);
and U12538 (N_12538,N_10354,N_11299);
and U12539 (N_12539,N_11812,N_11233);
or U12540 (N_12540,N_9410,N_11305);
nor U12541 (N_12541,N_9732,N_10325);
and U12542 (N_12542,N_9699,N_9671);
nand U12543 (N_12543,N_11160,N_11823);
nand U12544 (N_12544,N_10804,N_11626);
and U12545 (N_12545,N_10134,N_11759);
nor U12546 (N_12546,N_9200,N_11186);
nand U12547 (N_12547,N_11353,N_9034);
and U12548 (N_12548,N_9330,N_10516);
or U12549 (N_12549,N_11419,N_11308);
and U12550 (N_12550,N_11869,N_9666);
nor U12551 (N_12551,N_10914,N_9810);
and U12552 (N_12552,N_9108,N_9189);
nor U12553 (N_12553,N_10805,N_9879);
or U12554 (N_12554,N_9769,N_11989);
and U12555 (N_12555,N_9649,N_9062);
nand U12556 (N_12556,N_9836,N_10776);
nor U12557 (N_12557,N_11000,N_9028);
and U12558 (N_12558,N_9651,N_10424);
and U12559 (N_12559,N_11508,N_11450);
nor U12560 (N_12560,N_9445,N_10828);
and U12561 (N_12561,N_10360,N_11047);
nor U12562 (N_12562,N_10091,N_9019);
and U12563 (N_12563,N_9538,N_10416);
xor U12564 (N_12564,N_11456,N_9107);
or U12565 (N_12565,N_9805,N_10689);
xnor U12566 (N_12566,N_9586,N_11498);
nor U12567 (N_12567,N_11689,N_10605);
nand U12568 (N_12568,N_10172,N_10920);
nand U12569 (N_12569,N_10986,N_9015);
nand U12570 (N_12570,N_9342,N_11465);
nand U12571 (N_12571,N_11197,N_10048);
or U12572 (N_12572,N_11724,N_11618);
and U12573 (N_12573,N_9414,N_10741);
nor U12574 (N_12574,N_9553,N_10054);
nor U12575 (N_12575,N_11517,N_9726);
and U12576 (N_12576,N_10840,N_10948);
nor U12577 (N_12577,N_9663,N_10349);
xnor U12578 (N_12578,N_9088,N_9850);
and U12579 (N_12579,N_9196,N_9064);
nor U12580 (N_12580,N_11198,N_11774);
nor U12581 (N_12581,N_11259,N_11503);
or U12582 (N_12582,N_11328,N_10816);
and U12583 (N_12583,N_11429,N_9334);
nand U12584 (N_12584,N_10718,N_11389);
nand U12585 (N_12585,N_10693,N_10486);
xor U12586 (N_12586,N_10149,N_11254);
or U12587 (N_12587,N_11322,N_11753);
or U12588 (N_12588,N_11546,N_10527);
and U12589 (N_12589,N_9855,N_9710);
nand U12590 (N_12590,N_9676,N_9490);
nand U12591 (N_12591,N_9655,N_10947);
or U12592 (N_12592,N_11740,N_11855);
or U12593 (N_12593,N_11251,N_9276);
or U12594 (N_12594,N_9831,N_10907);
and U12595 (N_12595,N_11164,N_9240);
or U12596 (N_12596,N_11789,N_11115);
and U12597 (N_12597,N_9248,N_11069);
and U12598 (N_12598,N_9498,N_10471);
and U12599 (N_12599,N_9285,N_11507);
or U12600 (N_12600,N_11304,N_11957);
and U12601 (N_12601,N_9401,N_10309);
and U12602 (N_12602,N_10414,N_9149);
or U12603 (N_12603,N_11116,N_11011);
or U12604 (N_12604,N_11007,N_9224);
nand U12605 (N_12605,N_10488,N_9711);
nand U12606 (N_12606,N_10779,N_10903);
nor U12607 (N_12607,N_9205,N_11175);
nor U12608 (N_12608,N_9625,N_10419);
nand U12609 (N_12609,N_10312,N_11448);
and U12610 (N_12610,N_9509,N_11159);
or U12611 (N_12611,N_10214,N_10004);
nand U12612 (N_12612,N_11941,N_9758);
and U12613 (N_12613,N_10282,N_11142);
or U12614 (N_12614,N_10299,N_9198);
xnor U12615 (N_12615,N_10367,N_9908);
nand U12616 (N_12616,N_9534,N_10758);
nor U12617 (N_12617,N_9528,N_10411);
nor U12618 (N_12618,N_11271,N_9943);
or U12619 (N_12619,N_10268,N_9328);
nand U12620 (N_12620,N_10026,N_9852);
or U12621 (N_12621,N_10146,N_9858);
nand U12622 (N_12622,N_9824,N_9049);
xor U12623 (N_12623,N_9527,N_11800);
or U12624 (N_12624,N_11028,N_9348);
or U12625 (N_12625,N_10267,N_9794);
or U12626 (N_12626,N_9633,N_9454);
nor U12627 (N_12627,N_11523,N_9084);
or U12628 (N_12628,N_10013,N_10646);
xnor U12629 (N_12629,N_11811,N_9288);
and U12630 (N_12630,N_9190,N_10319);
and U12631 (N_12631,N_9436,N_10284);
and U12632 (N_12632,N_9898,N_10199);
nand U12633 (N_12633,N_11455,N_10695);
nor U12634 (N_12634,N_9761,N_9866);
or U12635 (N_12635,N_11799,N_11378);
nor U12636 (N_12636,N_9237,N_11065);
nand U12637 (N_12637,N_11492,N_11386);
or U12638 (N_12638,N_9095,N_9455);
or U12639 (N_12639,N_11155,N_10142);
or U12640 (N_12640,N_9350,N_11125);
nand U12641 (N_12641,N_11850,N_9464);
and U12642 (N_12642,N_10445,N_11402);
nor U12643 (N_12643,N_9030,N_11803);
nand U12644 (N_12644,N_10706,N_9657);
and U12645 (N_12645,N_10911,N_11472);
and U12646 (N_12646,N_10487,N_11968);
nand U12647 (N_12647,N_10242,N_9896);
nor U12648 (N_12648,N_9870,N_10376);
and U12649 (N_12649,N_9147,N_9968);
nor U12650 (N_12650,N_9399,N_11882);
or U12651 (N_12651,N_11295,N_10551);
and U12652 (N_12652,N_11583,N_10937);
or U12653 (N_12653,N_10877,N_11630);
nor U12654 (N_12654,N_9789,N_11015);
and U12655 (N_12655,N_10222,N_9235);
nor U12656 (N_12656,N_9664,N_9482);
or U12657 (N_12657,N_10323,N_10569);
or U12658 (N_12658,N_10099,N_11347);
or U12659 (N_12659,N_11329,N_9442);
and U12660 (N_12660,N_9692,N_9405);
nor U12661 (N_12661,N_9063,N_11504);
or U12662 (N_12662,N_9567,N_10431);
or U12663 (N_12663,N_10393,N_10392);
nor U12664 (N_12664,N_10451,N_10495);
nand U12665 (N_12665,N_9275,N_9409);
and U12666 (N_12666,N_10784,N_10094);
and U12667 (N_12667,N_9845,N_10467);
and U12668 (N_12668,N_9478,N_10581);
and U12669 (N_12669,N_10719,N_10865);
nand U12670 (N_12670,N_10007,N_11586);
or U12671 (N_12671,N_11961,N_9944);
and U12672 (N_12672,N_11338,N_11587);
nor U12673 (N_12673,N_10135,N_10862);
nor U12674 (N_12674,N_10845,N_10075);
xor U12675 (N_12675,N_10674,N_10078);
nor U12676 (N_12676,N_10892,N_10229);
and U12677 (N_12677,N_10764,N_11351);
nand U12678 (N_12678,N_10882,N_11479);
and U12679 (N_12679,N_10714,N_9881);
or U12680 (N_12680,N_9094,N_9932);
or U12681 (N_12681,N_11217,N_9764);
or U12682 (N_12682,N_9571,N_10955);
nand U12683 (N_12683,N_9515,N_10308);
and U12684 (N_12684,N_9156,N_9890);
or U12685 (N_12685,N_11139,N_10153);
and U12686 (N_12686,N_11099,N_11061);
or U12687 (N_12687,N_11845,N_11964);
nand U12688 (N_12688,N_10766,N_11726);
and U12689 (N_12689,N_9325,N_10753);
and U12690 (N_12690,N_11936,N_9557);
nand U12691 (N_12691,N_11672,N_11248);
nand U12692 (N_12692,N_10807,N_10694);
nand U12693 (N_12693,N_11931,N_9572);
nand U12694 (N_12694,N_9376,N_9085);
nor U12695 (N_12695,N_11383,N_10140);
xor U12696 (N_12696,N_9914,N_9876);
or U12697 (N_12697,N_11706,N_9223);
or U12698 (N_12698,N_10658,N_10696);
nand U12699 (N_12699,N_11535,N_10523);
and U12700 (N_12700,N_10836,N_10878);
and U12701 (N_12701,N_10885,N_11748);
nand U12702 (N_12702,N_9638,N_9807);
and U12703 (N_12703,N_11477,N_11932);
and U12704 (N_12704,N_9700,N_9366);
and U12705 (N_12705,N_9766,N_9126);
and U12706 (N_12706,N_11355,N_9684);
or U12707 (N_12707,N_11849,N_10895);
nor U12708 (N_12708,N_11252,N_10726);
or U12709 (N_12709,N_11763,N_9152);
nor U12710 (N_12710,N_11606,N_11044);
and U12711 (N_12711,N_11318,N_10735);
nor U12712 (N_12712,N_11050,N_10676);
and U12713 (N_12713,N_9999,N_10390);
and U12714 (N_12714,N_9717,N_9995);
nand U12715 (N_12715,N_9192,N_10043);
or U12716 (N_12716,N_9165,N_9402);
and U12717 (N_12717,N_9939,N_10721);
and U12718 (N_12718,N_10611,N_10742);
or U12719 (N_12719,N_11575,N_11459);
and U12720 (N_12720,N_9427,N_11454);
or U12721 (N_12721,N_11493,N_11734);
nor U12722 (N_12722,N_9056,N_9514);
nand U12723 (N_12723,N_9031,N_9214);
and U12724 (N_12724,N_10089,N_9050);
and U12725 (N_12725,N_11463,N_11131);
nor U12726 (N_12726,N_10618,N_11677);
nor U12727 (N_12727,N_11609,N_9364);
nand U12728 (N_12728,N_10929,N_11829);
and U12729 (N_12729,N_9082,N_11387);
nor U12730 (N_12730,N_9079,N_11119);
and U12731 (N_12731,N_10018,N_11636);
nand U12732 (N_12732,N_9012,N_11798);
and U12733 (N_12733,N_10009,N_9477);
and U12734 (N_12734,N_11483,N_9466);
nand U12735 (N_12735,N_9307,N_11052);
and U12736 (N_12736,N_9749,N_9404);
and U12737 (N_12737,N_11827,N_9506);
nand U12738 (N_12738,N_9661,N_11754);
nor U12739 (N_12739,N_10566,N_11722);
nand U12740 (N_12740,N_10430,N_10679);
nor U12741 (N_12741,N_10759,N_9308);
nand U12742 (N_12742,N_10496,N_10791);
nand U12743 (N_12743,N_10899,N_10301);
nand U12744 (N_12744,N_11335,N_9916);
and U12745 (N_12745,N_9286,N_9097);
nand U12746 (N_12746,N_11365,N_9066);
or U12747 (N_12747,N_10668,N_9113);
and U12748 (N_12748,N_10041,N_10848);
or U12749 (N_12749,N_11910,N_9598);
nand U12750 (N_12750,N_11423,N_9314);
or U12751 (N_12751,N_11394,N_10243);
and U12752 (N_12752,N_9024,N_11792);
and U12753 (N_12753,N_10322,N_9910);
nand U12754 (N_12754,N_9161,N_9403);
nand U12755 (N_12755,N_9215,N_9868);
and U12756 (N_12756,N_10856,N_11610);
xor U12757 (N_12757,N_10596,N_9620);
nand U12758 (N_12758,N_9238,N_10036);
nand U12759 (N_12759,N_10051,N_11445);
nor U12760 (N_12760,N_9254,N_9138);
or U12761 (N_12761,N_11350,N_11934);
or U12762 (N_12762,N_10025,N_9829);
nor U12763 (N_12763,N_10984,N_10113);
nor U12764 (N_12764,N_9061,N_11426);
nand U12765 (N_12765,N_9872,N_11810);
and U12766 (N_12766,N_10514,N_9453);
nor U12767 (N_12767,N_9984,N_10174);
nand U12768 (N_12768,N_10782,N_9045);
and U12769 (N_12769,N_9608,N_10918);
nor U12770 (N_12770,N_11970,N_9904);
nand U12771 (N_12771,N_10533,N_9869);
nor U12772 (N_12772,N_11441,N_11639);
or U12773 (N_12773,N_11593,N_9226);
nand U12774 (N_12774,N_11242,N_11226);
or U12775 (N_12775,N_9434,N_11274);
nand U12776 (N_12776,N_11300,N_11433);
nor U12777 (N_12777,N_10306,N_11622);
and U12778 (N_12778,N_11149,N_11832);
or U12779 (N_12779,N_10930,N_11094);
and U12780 (N_12780,N_10000,N_11924);
xnor U12781 (N_12781,N_9230,N_10210);
nand U12782 (N_12782,N_9435,N_10985);
nand U12783 (N_12783,N_10867,N_10924);
or U12784 (N_12784,N_9849,N_11374);
nand U12785 (N_12785,N_11169,N_9947);
nor U12786 (N_12786,N_9591,N_10084);
nand U12787 (N_12787,N_9419,N_9816);
nor U12788 (N_12788,N_10086,N_9516);
nand U12789 (N_12789,N_10788,N_10982);
nor U12790 (N_12790,N_9496,N_10096);
nand U12791 (N_12791,N_11199,N_9975);
or U12792 (N_12792,N_9521,N_11144);
or U12793 (N_12793,N_11681,N_11549);
or U12794 (N_12794,N_9713,N_11861);
nor U12795 (N_12795,N_11126,N_9813);
nor U12796 (N_12796,N_10307,N_11447);
and U12797 (N_12797,N_10795,N_11413);
or U12798 (N_12798,N_9119,N_10144);
and U12799 (N_12799,N_10197,N_11956);
or U12800 (N_12800,N_10670,N_11014);
nor U12801 (N_12801,N_11795,N_9388);
nand U12802 (N_12802,N_10777,N_9162);
xor U12803 (N_12803,N_9558,N_9906);
and U12804 (N_12804,N_11793,N_9632);
and U12805 (N_12805,N_10316,N_9302);
nor U12806 (N_12806,N_9277,N_11652);
and U12807 (N_12807,N_10761,N_9185);
nor U12808 (N_12808,N_11293,N_9720);
or U12809 (N_12809,N_11886,N_11249);
nor U12810 (N_12810,N_9957,N_10810);
nand U12811 (N_12811,N_11406,N_10796);
or U12812 (N_12812,N_9654,N_11545);
nor U12813 (N_12813,N_11862,N_11693);
and U12814 (N_12814,N_10295,N_10256);
and U12815 (N_12815,N_10227,N_11903);
nor U12816 (N_12816,N_9327,N_9674);
and U12817 (N_12817,N_11835,N_10561);
nand U12818 (N_12818,N_9878,N_11058);
or U12819 (N_12819,N_10270,N_10579);
nand U12820 (N_12820,N_10262,N_10770);
and U12821 (N_12821,N_10366,N_10340);
nor U12822 (N_12822,N_11156,N_11653);
and U12823 (N_12823,N_10752,N_10708);
nand U12824 (N_12824,N_9884,N_10660);
nor U12825 (N_12825,N_9067,N_10279);
nand U12826 (N_12826,N_10681,N_10745);
or U12827 (N_12827,N_11764,N_9723);
and U12828 (N_12828,N_11009,N_11316);
and U12829 (N_12829,N_11522,N_9525);
xnor U12830 (N_12830,N_9228,N_10624);
or U12831 (N_12831,N_9725,N_11649);
nor U12832 (N_12832,N_11893,N_11555);
or U12833 (N_12833,N_11097,N_11579);
nand U12834 (N_12834,N_11853,N_9549);
nor U12835 (N_12835,N_10111,N_10311);
and U12836 (N_12836,N_11641,N_9678);
and U12837 (N_12837,N_10699,N_11978);
and U12838 (N_12838,N_9087,N_9261);
nor U12839 (N_12839,N_10616,N_10131);
and U12840 (N_12840,N_10192,N_11444);
nand U12841 (N_12841,N_9597,N_10077);
and U12842 (N_12842,N_10820,N_10409);
or U12843 (N_12843,N_9981,N_10944);
and U12844 (N_12844,N_9911,N_11664);
nor U12845 (N_12845,N_9552,N_11049);
or U12846 (N_12846,N_9974,N_11056);
or U12847 (N_12847,N_10691,N_10774);
nor U12848 (N_12848,N_9122,N_9479);
nand U12849 (N_12849,N_9715,N_10900);
nor U12850 (N_12850,N_10127,N_11788);
and U12851 (N_12851,N_9227,N_9212);
nand U12852 (N_12852,N_10940,N_11420);
nor U12853 (N_12853,N_11260,N_10959);
or U12854 (N_12854,N_10941,N_10378);
or U12855 (N_12855,N_10628,N_11277);
nand U12856 (N_12856,N_9187,N_10176);
and U12857 (N_12857,N_11776,N_9272);
xor U12858 (N_12858,N_11478,N_9121);
xnor U12859 (N_12859,N_9428,N_10402);
xor U12860 (N_12860,N_9111,N_11220);
nor U12861 (N_12861,N_10328,N_10217);
nor U12862 (N_12862,N_10970,N_11038);
or U12863 (N_12863,N_10336,N_9003);
xor U12864 (N_12864,N_9978,N_9335);
or U12865 (N_12865,N_10466,N_10186);
or U12866 (N_12866,N_9025,N_10513);
nor U12867 (N_12867,N_9313,N_10181);
nor U12868 (N_12868,N_10396,N_9452);
nor U12869 (N_12869,N_11842,N_11602);
nor U12870 (N_12870,N_11424,N_9626);
or U12871 (N_12871,N_10749,N_11362);
and U12872 (N_12872,N_11666,N_9706);
nand U12873 (N_12873,N_11231,N_11879);
or U12874 (N_12874,N_9117,N_11809);
nand U12875 (N_12875,N_9069,N_10644);
nand U12876 (N_12876,N_11562,N_11694);
nand U12877 (N_12877,N_10401,N_11416);
nor U12878 (N_12878,N_11818,N_10972);
nand U12879 (N_12879,N_9081,N_10287);
or U12880 (N_12880,N_11246,N_10705);
and U12881 (N_12881,N_10275,N_11481);
nor U12882 (N_12882,N_10128,N_9059);
or U12883 (N_12883,N_11923,N_9168);
nand U12884 (N_12884,N_10442,N_11020);
or U12885 (N_12885,N_9320,N_9317);
and U12886 (N_12886,N_10196,N_11177);
nor U12887 (N_12887,N_10980,N_11446);
nor U12888 (N_12888,N_11434,N_10410);
nor U12889 (N_12889,N_10798,N_11412);
or U12890 (N_12890,N_11296,N_11005);
and U12891 (N_12891,N_10826,N_11814);
nor U12892 (N_12892,N_10647,N_9485);
or U12893 (N_12893,N_10604,N_10161);
nand U12894 (N_12894,N_9539,N_9473);
and U12895 (N_12895,N_10318,N_10905);
and U12896 (N_12896,N_11661,N_10504);
nor U12897 (N_12897,N_10463,N_10849);
nor U12898 (N_12898,N_11669,N_11307);
nor U12899 (N_12899,N_10482,N_9262);
and U12900 (N_12900,N_11906,N_9822);
or U12901 (N_12901,N_9080,N_11568);
nor U12902 (N_12902,N_9861,N_11635);
nand U12903 (N_12903,N_11887,N_10371);
or U12904 (N_12904,N_11247,N_9413);
nand U12905 (N_12905,N_11026,N_9153);
or U12906 (N_12906,N_11476,N_9894);
nand U12907 (N_12907,N_10375,N_10288);
nor U12908 (N_12908,N_11654,N_11969);
and U12909 (N_12909,N_10880,N_9526);
nor U12910 (N_12910,N_10932,N_11902);
nand U12911 (N_12911,N_9777,N_11313);
nor U12912 (N_12912,N_11781,N_10896);
nor U12913 (N_12913,N_11914,N_10369);
nor U12914 (N_12914,N_11399,N_9283);
nand U12915 (N_12915,N_10178,N_11377);
and U12916 (N_12916,N_9221,N_9326);
nand U12917 (N_12917,N_11428,N_11519);
nand U12918 (N_12918,N_9469,N_11273);
nand U12919 (N_12919,N_11996,N_11466);
nor U12920 (N_12920,N_9920,N_9630);
nand U12921 (N_12921,N_9942,N_11238);
and U12922 (N_12922,N_11937,N_9883);
nor U12923 (N_12923,N_10436,N_10145);
and U12924 (N_12924,N_10218,N_9587);
nor U12925 (N_12925,N_11281,N_9989);
nor U12926 (N_12926,N_9959,N_10012);
nor U12927 (N_12927,N_10713,N_10964);
or U12928 (N_12928,N_10395,N_9180);
or U12929 (N_12929,N_11435,N_10739);
and U12930 (N_12930,N_9231,N_9683);
and U12931 (N_12931,N_9595,N_11821);
and U12932 (N_12932,N_9739,N_9022);
and U12933 (N_12933,N_10978,N_11541);
or U12934 (N_12934,N_11988,N_9008);
and U12935 (N_12935,N_10935,N_11534);
nor U12936 (N_12936,N_11569,N_9203);
nand U12937 (N_12937,N_11766,N_11211);
and U12938 (N_12938,N_11229,N_9480);
and U12939 (N_12939,N_9500,N_10755);
or U12940 (N_12940,N_9213,N_9851);
nor U12941 (N_12941,N_9341,N_10824);
nand U12942 (N_12942,N_10010,N_10232);
nor U12943 (N_12943,N_10507,N_9487);
nor U12944 (N_12944,N_9886,N_11398);
nor U12945 (N_12945,N_10762,N_11683);
nand U12946 (N_12946,N_9618,N_9677);
and U12947 (N_12947,N_10580,N_9923);
and U12948 (N_12948,N_10258,N_9102);
nand U12949 (N_12949,N_11106,N_9425);
or U12950 (N_12950,N_10812,N_11489);
nand U12951 (N_12951,N_11194,N_9179);
or U12952 (N_12952,N_9532,N_11644);
nand U12953 (N_12953,N_9697,N_9058);
and U12954 (N_12954,N_11102,N_9817);
nand U12955 (N_12955,N_10452,N_9918);
or U12956 (N_12956,N_11925,N_9183);
nand U12957 (N_12957,N_9728,N_9645);
and U12958 (N_12958,N_11110,N_11897);
and U12959 (N_12959,N_11979,N_11967);
or U12960 (N_12960,N_9345,N_10215);
nor U12961 (N_12961,N_9418,N_10479);
nor U12962 (N_12962,N_10817,N_10182);
nor U12963 (N_12963,N_10983,N_11375);
nor U12964 (N_12964,N_10772,N_11087);
nor U12965 (N_12965,N_10620,N_10476);
and U12966 (N_12966,N_9461,N_10623);
or U12967 (N_12967,N_10491,N_11918);
nand U12968 (N_12968,N_9820,N_11532);
or U12969 (N_12969,N_11161,N_10965);
or U12970 (N_12970,N_9495,N_11330);
nand U12971 (N_12971,N_11120,N_10814);
nor U12972 (N_12972,N_10539,N_11257);
xnor U12973 (N_12973,N_9421,N_10073);
and U12974 (N_12974,N_10802,N_9601);
or U12975 (N_12975,N_9686,N_11667);
or U12976 (N_12976,N_9784,N_11059);
or U12977 (N_12977,N_10266,N_9827);
nand U12978 (N_12978,N_11467,N_9065);
nor U12979 (N_12979,N_9014,N_10391);
nor U12980 (N_12980,N_10472,N_10831);
or U12981 (N_12981,N_10969,N_10803);
nand U12982 (N_12982,N_11993,N_9092);
and U12983 (N_12983,N_11213,N_10590);
nor U12984 (N_12984,N_9590,N_9243);
and U12985 (N_12985,N_10701,N_11885);
xnor U12986 (N_12986,N_11595,N_10910);
or U12987 (N_12987,N_11612,N_11581);
nand U12988 (N_12988,N_11317,N_10356);
nor U12989 (N_12989,N_10037,N_9899);
nor U12990 (N_12990,N_10342,N_9319);
or U12991 (N_12991,N_11219,N_10418);
nor U12992 (N_12992,N_10254,N_10536);
nor U12993 (N_12993,N_9041,N_9973);
or U12994 (N_12994,N_11741,N_10692);
nor U12995 (N_12995,N_11553,N_9318);
nand U12996 (N_12996,N_9296,N_10346);
or U12997 (N_12997,N_9741,N_11195);
and U12998 (N_12998,N_11847,N_10582);
nor U12999 (N_12999,N_9696,N_10915);
xnor U13000 (N_13000,N_11221,N_10710);
or U13001 (N_13001,N_11582,N_11130);
nor U13002 (N_13002,N_11027,N_10635);
xnor U13003 (N_13003,N_10630,N_10506);
and U13004 (N_13004,N_10191,N_10494);
nand U13005 (N_13005,N_10800,N_10633);
and U13006 (N_13006,N_11401,N_9639);
nand U13007 (N_13007,N_10621,N_10155);
or U13008 (N_13008,N_10339,N_10443);
and U13009 (N_13009,N_9901,N_11261);
or U13010 (N_13010,N_11285,N_11036);
xor U13011 (N_13011,N_10171,N_11819);
or U13012 (N_13012,N_11158,N_10775);
nand U13013 (N_13013,N_9157,N_9782);
nand U13014 (N_13014,N_9885,N_9963);
nand U13015 (N_13015,N_10261,N_10093);
nor U13016 (N_13016,N_9365,N_9493);
nor U13017 (N_13017,N_11390,N_11382);
or U13018 (N_13018,N_10345,N_9395);
nor U13019 (N_13019,N_11174,N_11501);
nand U13020 (N_13020,N_11101,N_10564);
or U13021 (N_13021,N_11943,N_11282);
nand U13022 (N_13022,N_10546,N_9609);
nor U13023 (N_13023,N_10236,N_10475);
or U13024 (N_13024,N_11700,N_11662);
and U13025 (N_13025,N_10874,N_10350);
and U13026 (N_13026,N_10698,N_9104);
or U13027 (N_13027,N_11703,N_9736);
and U13028 (N_13028,N_11729,N_10459);
nor U13029 (N_13029,N_9547,N_11707);
nand U13030 (N_13030,N_9492,N_10332);
and U13031 (N_13031,N_9613,N_11292);
nand U13032 (N_13032,N_9143,N_11239);
and U13033 (N_13033,N_11484,N_11597);
nand U13034 (N_13034,N_11071,N_11218);
nor U13035 (N_13035,N_11983,N_11898);
nor U13036 (N_13036,N_10677,N_11141);
and U13037 (N_13037,N_10562,N_9972);
nand U13038 (N_13038,N_11797,N_10006);
and U13039 (N_13039,N_10690,N_11369);
nor U13040 (N_13040,N_11873,N_9139);
nor U13041 (N_13041,N_10946,N_11580);
nand U13042 (N_13042,N_11017,N_11520);
or U13043 (N_13043,N_11840,N_11091);
nor U13044 (N_13044,N_10263,N_10531);
and U13045 (N_13045,N_11128,N_11418);
nor U13046 (N_13046,N_9636,N_11976);
and U13047 (N_13047,N_10423,N_11806);
or U13048 (N_13048,N_11346,N_9756);
nand U13049 (N_13049,N_11301,N_9992);
and U13050 (N_13050,N_9216,N_10949);
nor U13051 (N_13051,N_10994,N_11822);
or U13052 (N_13052,N_9259,N_10977);
and U13053 (N_13053,N_9653,N_10246);
nor U13054 (N_13054,N_11963,N_10385);
or U13055 (N_13055,N_10901,N_10223);
and U13056 (N_13056,N_11585,N_9540);
or U13057 (N_13057,N_10785,N_11066);
nor U13058 (N_13058,N_10938,N_9576);
and U13059 (N_13059,N_11866,N_10297);
or U13060 (N_13060,N_9599,N_11111);
nor U13061 (N_13061,N_11331,N_10971);
nor U13062 (N_13062,N_10962,N_11326);
xnor U13063 (N_13063,N_10292,N_10834);
or U13064 (N_13064,N_9801,N_9815);
and U13065 (N_13065,N_11540,N_10221);
nand U13066 (N_13066,N_10830,N_11309);
or U13067 (N_13067,N_10177,N_9775);
nor U13068 (N_13068,N_11266,N_9499);
or U13069 (N_13069,N_9333,N_11325);
nand U13070 (N_13070,N_11947,N_9472);
and U13071 (N_13071,N_11619,N_9281);
and U13072 (N_13072,N_9446,N_9060);
or U13073 (N_13073,N_10333,N_11085);
and U13074 (N_13074,N_10715,N_11002);
or U13075 (N_13075,N_10664,N_11276);
nand U13076 (N_13076,N_10428,N_10928);
nand U13077 (N_13077,N_9721,N_10151);
or U13078 (N_13078,N_11884,N_10461);
nand U13079 (N_13079,N_11332,N_9368);
nor U13080 (N_13080,N_10549,N_9510);
nand U13081 (N_13081,N_9174,N_9665);
nor U13082 (N_13082,N_9513,N_11868);
and U13083 (N_13083,N_10427,N_11414);
or U13084 (N_13084,N_10244,N_9011);
nor U13085 (N_13085,N_11095,N_10049);
nand U13086 (N_13086,N_10584,N_10886);
or U13087 (N_13087,N_10737,N_11395);
nand U13088 (N_13088,N_11647,N_11838);
nand U13089 (N_13089,N_9616,N_10352);
and U13090 (N_13090,N_10974,N_10358);
or U13091 (N_13091,N_9735,N_11750);
and U13092 (N_13092,N_9669,N_9607);
and U13093 (N_13093,N_10102,N_10996);
nand U13094 (N_13094,N_9931,N_10509);
nor U13095 (N_13095,N_10642,N_9135);
and U13096 (N_13096,N_9508,N_11973);
nand U13097 (N_13097,N_11828,N_10169);
or U13098 (N_13098,N_10960,N_11339);
nand U13099 (N_13099,N_10492,N_9052);
nand U13100 (N_13100,N_9407,N_10600);
and U13101 (N_13101,N_10966,N_11253);
or U13102 (N_13102,N_9841,N_9486);
or U13103 (N_13103,N_10470,N_9809);
nor U13104 (N_13104,N_11565,N_10231);
nand U13105 (N_13105,N_9309,N_11024);
and U13106 (N_13106,N_10059,N_11900);
nand U13107 (N_13107,N_11871,N_10300);
and U13108 (N_13108,N_10083,N_9954);
nor U13109 (N_13109,N_11860,N_10926);
or U13110 (N_13110,N_10158,N_10344);
and U13111 (N_13111,N_11949,N_9915);
xnor U13112 (N_13112,N_10194,N_11092);
nor U13113 (N_13113,N_9520,N_9909);
nor U13114 (N_13114,N_9048,N_11045);
nor U13115 (N_13115,N_11341,N_11548);
and U13116 (N_13116,N_9336,N_9429);
nand U13117 (N_13117,N_11188,N_11468);
nand U13118 (N_13118,N_10685,N_10976);
or U13119 (N_13119,N_10170,N_10841);
and U13120 (N_13120,N_9141,N_9007);
or U13121 (N_13121,N_10173,N_9569);
nor U13122 (N_13122,N_11055,N_9134);
and U13123 (N_13123,N_10855,N_9880);
or U13124 (N_13124,N_11837,N_10057);
nor U13125 (N_13125,N_11016,N_9468);
and U13126 (N_13126,N_11775,N_10237);
and U13127 (N_13127,N_10204,N_10097);
nor U13128 (N_13128,N_9411,N_9531);
and U13129 (N_13129,N_9125,N_9583);
or U13130 (N_13130,N_9255,N_11874);
nand U13131 (N_13131,N_9750,N_9379);
and U13132 (N_13132,N_11240,N_11856);
nand U13133 (N_13133,N_10846,N_11846);
or U13134 (N_13134,N_9253,N_11926);
or U13135 (N_13135,N_10020,N_10481);
nor U13136 (N_13136,N_10975,N_10998);
xnor U13137 (N_13137,N_11629,N_9614);
nand U13138 (N_13138,N_9112,N_11133);
nor U13139 (N_13139,N_11096,N_9961);
nor U13140 (N_13140,N_11235,N_11283);
and U13141 (N_13141,N_11804,N_9400);
nand U13142 (N_13142,N_11716,N_9606);
and U13143 (N_13143,N_11916,N_11312);
or U13144 (N_13144,N_11634,N_9175);
and U13145 (N_13145,N_11034,N_10760);
nand U13146 (N_13146,N_11588,N_9600);
xnor U13147 (N_13147,N_10362,N_9291);
nor U13148 (N_13148,N_10220,N_10437);
or U13149 (N_13149,N_9536,N_9105);
nand U13150 (N_13150,N_10939,N_11908);
or U13151 (N_13151,N_10967,N_9412);
and U13152 (N_13152,N_10667,N_10320);
or U13153 (N_13153,N_11491,N_11715);
nor U13154 (N_13154,N_10585,N_10541);
or U13155 (N_13155,N_9298,N_11403);
nor U13156 (N_13156,N_9748,N_10154);
or U13157 (N_13157,N_11554,N_10446);
or U13158 (N_13158,N_10524,N_11349);
nor U13159 (N_13159,N_10053,N_11264);
or U13160 (N_13160,N_9070,N_11904);
nor U13161 (N_13161,N_10038,N_9832);
nor U13162 (N_13162,N_9948,N_9987);
or U13163 (N_13163,N_9385,N_9703);
or U13164 (N_13164,N_9795,N_11100);
and U13165 (N_13165,N_9737,N_10164);
nand U13166 (N_13166,N_10008,N_9662);
nor U13167 (N_13167,N_11008,N_11076);
nand U13168 (N_13168,N_11237,N_10324);
nand U13169 (N_13169,N_11589,N_10441);
xnor U13170 (N_13170,N_9351,N_11574);
and U13171 (N_13171,N_11670,N_10732);
or U13172 (N_13172,N_9363,N_10768);
and U13173 (N_13173,N_9042,N_11883);
nor U13174 (N_13174,N_9071,N_9361);
nor U13175 (N_13175,N_9396,N_9476);
or U13176 (N_13176,N_9362,N_10277);
or U13177 (N_13177,N_10953,N_11538);
or U13178 (N_13178,N_9589,N_9573);
nor U13179 (N_13179,N_10765,N_11204);
nor U13180 (N_13180,N_9371,N_9623);
nor U13181 (N_13181,N_10453,N_11384);
or U13182 (N_13182,N_10797,N_11185);
xor U13183 (N_13183,N_9643,N_9814);
nor U13184 (N_13184,N_9629,N_9865);
and U13185 (N_13185,N_9035,N_9545);
and U13186 (N_13186,N_9687,N_10853);
or U13187 (N_13187,N_9716,N_9002);
nor U13188 (N_13188,N_9124,N_10313);
or U13189 (N_13189,N_9701,N_10661);
or U13190 (N_13190,N_10876,N_10071);
and U13191 (N_13191,N_10462,N_11755);
nor U13192 (N_13192,N_11269,N_11030);
or U13193 (N_13193,N_11945,N_9945);
and U13194 (N_13194,N_10902,N_9023);
nor U13195 (N_13195,N_11511,N_9236);
or U13196 (N_13196,N_10039,N_10515);
nor U13197 (N_13197,N_11698,N_9917);
nor U13198 (N_13198,N_11913,N_9856);
or U13199 (N_13199,N_9078,N_10159);
nor U13200 (N_13200,N_9339,N_9584);
nand U13201 (N_13201,N_9293,N_9201);
or U13202 (N_13202,N_9271,N_11922);
nor U13203 (N_13203,N_10239,N_10990);
or U13204 (N_13204,N_9270,N_9129);
nor U13205 (N_13205,N_11191,N_10351);
nor U13206 (N_13206,N_9098,N_9093);
and U13207 (N_13207,N_9219,N_10665);
nor U13208 (N_13208,N_10942,N_11053);
nand U13209 (N_13209,N_10854,N_11336);
nand U13210 (N_13210,N_9635,N_10615);
nor U13211 (N_13211,N_9602,N_9282);
or U13212 (N_13212,N_11490,N_10556);
nand U13213 (N_13213,N_11733,N_11940);
or U13214 (N_13214,N_9518,N_11999);
nand U13215 (N_13215,N_9648,N_11645);
nor U13216 (N_13216,N_10269,N_11550);
nand U13217 (N_13217,N_10455,N_10811);
and U13218 (N_13218,N_11180,N_9090);
nor U13219 (N_13219,N_11012,N_11948);
nand U13220 (N_13220,N_11600,N_10656);
or U13221 (N_13221,N_11745,N_10801);
or U13222 (N_13222,N_11127,N_9380);
nand U13223 (N_13223,N_9295,N_9559);
and U13224 (N_13224,N_10379,N_9151);
nand U13225 (N_13225,N_9962,N_10833);
nor U13226 (N_13226,N_11909,N_9329);
nand U13227 (N_13227,N_10224,N_9895);
nor U13228 (N_13228,N_11717,N_11166);
and U13229 (N_13229,N_10559,N_10055);
and U13230 (N_13230,N_9471,N_10112);
nand U13231 (N_13231,N_10019,N_10731);
nand U13232 (N_13232,N_9340,N_10255);
nor U13233 (N_13233,N_9290,N_9511);
nor U13234 (N_13234,N_10225,N_11738);
xor U13235 (N_13235,N_11145,N_9289);
or U13236 (N_13236,N_10359,N_11114);
nand U13237 (N_13237,N_11124,N_10678);
nor U13238 (N_13238,N_11514,N_11214);
or U13239 (N_13239,N_10629,N_10355);
and U13240 (N_13240,N_9467,N_11209);
or U13241 (N_13241,N_9132,N_11368);
nor U13242 (N_13242,N_11379,N_11712);
and U13243 (N_13243,N_9280,N_10150);
nand U13244 (N_13244,N_9154,N_10525);
or U13245 (N_13245,N_10827,N_11625);
nor U13246 (N_13246,N_9312,N_10184);
nor U13247 (N_13247,N_11912,N_9956);
or U13248 (N_13248,N_9148,N_11542);
nor U13249 (N_13249,N_9771,N_11232);
nor U13250 (N_13250,N_10118,N_10397);
nand U13251 (N_13251,N_10809,N_9826);
nor U13252 (N_13252,N_10474,N_11817);
nor U13253 (N_13253,N_9160,N_10570);
nor U13254 (N_13254,N_10711,N_11521);
nor U13255 (N_13255,N_10723,N_10175);
nand U13256 (N_13256,N_10465,N_10703);
and U13257 (N_13257,N_9369,N_11787);
nor U13258 (N_13258,N_10575,N_11864);
or U13259 (N_13259,N_11756,N_9433);
nor U13260 (N_13260,N_11278,N_10860);
or U13261 (N_13261,N_11427,N_11381);
or U13262 (N_13262,N_10601,N_9517);
nand U13263 (N_13263,N_9264,N_11287);
nor U13264 (N_13264,N_11590,N_10925);
nand U13265 (N_13265,N_11320,N_9273);
and U13266 (N_13266,N_9772,N_10157);
nand U13267 (N_13267,N_10627,N_11442);
nor U13268 (N_13268,N_10331,N_10654);
and U13269 (N_13269,N_11599,N_9907);
nand U13270 (N_13270,N_11663,N_9507);
or U13271 (N_13271,N_11357,N_9091);
xnor U13272 (N_13272,N_10956,N_11121);
xnor U13273 (N_13273,N_11972,N_10001);
and U13274 (N_13274,N_9247,N_10769);
nand U13275 (N_13275,N_10778,N_11137);
nand U13276 (N_13276,N_11022,N_10133);
or U13277 (N_13277,N_9086,N_9242);
or U13278 (N_13278,N_10700,N_10954);
and U13279 (N_13279,N_10560,N_11070);
nand U13280 (N_13280,N_9170,N_11437);
nor U13281 (N_13281,N_11727,N_9575);
nor U13282 (N_13282,N_9459,N_11154);
nor U13283 (N_13283,N_11551,N_9311);
or U13284 (N_13284,N_11604,N_10468);
and U13285 (N_13285,N_11324,N_11852);
and U13286 (N_13286,N_10435,N_10265);
nor U13287 (N_13287,N_10538,N_9934);
nand U13288 (N_13288,N_9392,N_10056);
and U13289 (N_13289,N_10190,N_11006);
nand U13290 (N_13290,N_10657,N_11303);
nor U13291 (N_13291,N_11558,N_10829);
or U13292 (N_13292,N_10228,N_10249);
nor U13293 (N_13293,N_10042,N_9773);
or U13294 (N_13294,N_10040,N_11907);
nor U13295 (N_13295,N_10314,N_10688);
nand U13296 (N_13296,N_11950,N_9555);
xnor U13297 (N_13297,N_11714,N_9416);
or U13298 (N_13298,N_11642,N_9301);
nor U13299 (N_13299,N_9033,N_10248);
nor U13300 (N_13300,N_10085,N_10593);
or U13301 (N_13301,N_10274,N_11107);
or U13302 (N_13302,N_10489,N_9953);
nor U13303 (N_13303,N_10070,N_11470);
nor U13304 (N_13304,N_11808,N_10740);
nor U13305 (N_13305,N_11138,N_10682);
and U13306 (N_13306,N_11147,N_9806);
nor U13307 (N_13307,N_9073,N_9928);
and U13308 (N_13308,N_9612,N_10851);
or U13309 (N_13309,N_11758,N_10973);
or U13310 (N_13310,N_9158,N_10730);
xnor U13311 (N_13311,N_11083,N_9615);
nor U13312 (N_13312,N_11193,N_11671);
nor U13313 (N_13313,N_11668,N_11854);
nand U13314 (N_13314,N_11074,N_10189);
nand U13315 (N_13315,N_9346,N_10382);
nor U13316 (N_13316,N_10079,N_10021);
or U13317 (N_13317,N_10857,N_11132);
or U13318 (N_13318,N_11129,N_11878);
and U13319 (N_13319,N_11813,N_10399);
or U13320 (N_13320,N_11263,N_11462);
and U13321 (N_13321,N_9422,N_9184);
nor U13322 (N_13322,N_9691,N_11327);
nor U13323 (N_13323,N_11863,N_10380);
nor U13324 (N_13324,N_10321,N_9504);
or U13325 (N_13325,N_11359,N_11730);
and U13326 (N_13326,N_11820,N_10897);
nor U13327 (N_13327,N_9530,N_11772);
nor U13328 (N_13328,N_11637,N_11966);
nand U13329 (N_13329,N_10139,N_9798);
nand U13330 (N_13330,N_10460,N_9641);
and U13331 (N_13331,N_10408,N_10872);
nor U13332 (N_13332,N_9889,N_9570);
and U13333 (N_13333,N_10389,N_9746);
and U13334 (N_13334,N_10457,N_10068);
and U13335 (N_13335,N_11977,N_10251);
or U13336 (N_13336,N_11962,N_10357);
nand U13337 (N_13337,N_9708,N_11927);
or U13338 (N_13338,N_9208,N_9997);
and U13339 (N_13339,N_10540,N_10015);
nor U13340 (N_13340,N_10406,N_11431);
or U13341 (N_13341,N_11865,N_10448);
xnor U13342 (N_13342,N_9372,N_9709);
or U13343 (N_13343,N_10906,N_10951);
xor U13344 (N_13344,N_11561,N_11113);
and U13345 (N_13345,N_11031,N_10061);
or U13346 (N_13346,N_11896,N_10989);
nor U13347 (N_13347,N_11573,N_9640);
nor U13348 (N_13348,N_11051,N_11749);
and U13349 (N_13349,N_9780,N_11471);
or U13350 (N_13350,N_11060,N_9249);
and U13351 (N_13351,N_9110,N_10908);
or U13352 (N_13352,N_11123,N_11496);
nor U13353 (N_13353,N_11935,N_11975);
nand U13354 (N_13354,N_11046,N_11152);
and U13355 (N_13355,N_9074,N_10687);
or U13356 (N_13356,N_10729,N_11023);
or U13357 (N_13357,N_10387,N_10734);
or U13358 (N_13358,N_11205,N_9133);
nor U13359 (N_13359,N_10484,N_11181);
and U13360 (N_13360,N_9941,N_11010);
and U13361 (N_13361,N_11345,N_11001);
nand U13362 (N_13362,N_9130,N_9759);
nor U13363 (N_13363,N_11079,N_11628);
nor U13364 (N_13364,N_10588,N_11895);
nand U13365 (N_13365,N_9424,N_10259);
nor U13366 (N_13366,N_9027,N_9444);
nor U13367 (N_13367,N_10027,N_11578);
nor U13368 (N_13368,N_9751,N_11073);
and U13369 (N_13369,N_9940,N_9406);
nand U13370 (N_13370,N_10201,N_9983);
nor U13371 (N_13371,N_11143,N_10544);
and U13372 (N_13372,N_11557,N_9294);
and U13373 (N_13373,N_11224,N_10014);
nor U13374 (N_13374,N_10130,N_10412);
and U13375 (N_13375,N_9991,N_9659);
and U13376 (N_13376,N_10033,N_9897);
nand U13377 (N_13377,N_11241,N_10365);
nand U13378 (N_13378,N_11742,N_10334);
xor U13379 (N_13379,N_9096,N_11825);
xnor U13380 (N_13380,N_9958,N_9921);
xnor U13381 (N_13381,N_11035,N_10293);
xnor U13382 (N_13382,N_11665,N_11464);
nand U13383 (N_13383,N_10751,N_10074);
nand U13384 (N_13384,N_10921,N_10511);
nand U13385 (N_13385,N_11208,N_9693);
or U13386 (N_13386,N_9077,N_10456);
or U13387 (N_13387,N_11732,N_9688);
and U13388 (N_13388,N_11297,N_11623);
nor U13389 (N_13389,N_11526,N_10417);
nand U13390 (N_13390,N_9811,N_11779);
or U13391 (N_13391,N_10780,N_9256);
xor U13392 (N_13392,N_9554,N_11344);
and U13393 (N_13393,N_11648,N_11075);
and U13394 (N_13394,N_9250,N_10034);
and U13395 (N_13395,N_10226,N_11974);
and U13396 (N_13396,N_9197,N_10832);
or U13397 (N_13397,N_9977,N_11603);
nor U13398 (N_13398,N_10398,N_10092);
or U13399 (N_13399,N_10704,N_11480);
and U13400 (N_13400,N_9173,N_10193);
and U13401 (N_13401,N_11920,N_11769);
nor U13402 (N_13402,N_9266,N_10850);
or U13403 (N_13403,N_9821,N_10281);
nand U13404 (N_13404,N_10858,N_10981);
or U13405 (N_13405,N_11088,N_11510);
nor U13406 (N_13406,N_10029,N_10673);
and U13407 (N_13407,N_10808,N_10064);
nand U13408 (N_13408,N_9029,N_11460);
nand U13409 (N_13409,N_10438,N_9548);
and U13410 (N_13410,N_10152,N_9871);
or U13411 (N_13411,N_9560,N_11210);
nand U13412 (N_13412,N_11615,N_9260);
or U13413 (N_13413,N_11704,N_9244);
nor U13414 (N_13414,N_9039,N_11987);
and U13415 (N_13415,N_10508,N_10838);
nand U13416 (N_13416,N_9887,N_10747);
nor U13417 (N_13417,N_10861,N_11986);
nor U13418 (N_13418,N_10622,N_11701);
nor U13419 (N_13419,N_9742,N_9679);
nand U13420 (N_13420,N_11516,N_10060);
nor U13421 (N_13421,N_10206,N_11633);
nand U13422 (N_13422,N_10576,N_9580);
or U13423 (N_13423,N_9026,N_10195);
nor U13424 (N_13424,N_10498,N_9522);
or U13425 (N_13425,N_11356,N_10650);
and U13426 (N_13426,N_9818,N_10909);
and U13427 (N_13427,N_11567,N_11598);
or U13428 (N_13428,N_9949,N_9046);
nand U13429 (N_13429,N_11632,N_11400);
nor U13430 (N_13430,N_10844,N_11761);
nand U13431 (N_13431,N_9744,N_11206);
nor U13432 (N_13432,N_9743,N_11165);
nor U13433 (N_13433,N_9658,N_11172);
xnor U13434 (N_13434,N_9604,N_10799);
and U13435 (N_13435,N_10272,N_9501);
or U13436 (N_13436,N_10553,N_10529);
and U13437 (N_13437,N_9946,N_11901);
or U13438 (N_13438,N_11135,N_11189);
nor U13439 (N_13439,N_9274,N_11089);
or U13440 (N_13440,N_10890,N_10285);
and U13441 (N_13441,N_11816,N_10156);
or U13442 (N_13442,N_9068,N_10148);
or U13443 (N_13443,N_11104,N_9712);
or U13444 (N_13444,N_11150,N_10052);
nand U13445 (N_13445,N_9828,N_9448);
or U13446 (N_13446,N_10103,N_11109);
and U13447 (N_13447,N_11409,N_9859);
and U13448 (N_13448,N_9647,N_10447);
nand U13449 (N_13449,N_10289,N_9617);
or U13450 (N_13450,N_10619,N_9109);
and U13451 (N_13451,N_9323,N_11784);
or U13452 (N_13452,N_9465,N_10238);
nor U13453 (N_13453,N_11314,N_11178);
and U13454 (N_13454,N_9426,N_10609);
nand U13455 (N_13455,N_11216,N_11081);
and U13456 (N_13456,N_9123,N_9988);
or U13457 (N_13457,N_9848,N_9181);
and U13458 (N_13458,N_9718,N_10413);
or U13459 (N_13459,N_11655,N_11228);
nor U13460 (N_13460,N_11168,N_9010);
nand U13461 (N_13461,N_9847,N_10683);
and U13462 (N_13462,N_9357,N_11744);
and U13463 (N_13463,N_10207,N_9574);
nand U13464 (N_13464,N_10216,N_9353);
and U13465 (N_13465,N_11786,N_11364);
and U13466 (N_13466,N_9562,N_9937);
nor U13467 (N_13467,N_9681,N_11537);
nor U13468 (N_13468,N_11298,N_9450);
xnor U13469 (N_13469,N_10088,N_10589);
nand U13470 (N_13470,N_11791,N_10213);
nand U13471 (N_13471,N_9234,N_9394);
nand U13472 (N_13472,N_9377,N_9734);
nand U13473 (N_13473,N_9303,N_10550);
nand U13474 (N_13474,N_10326,N_11929);
nor U13475 (N_13475,N_11397,N_9032);
nor U13476 (N_13476,N_11760,N_10143);
nor U13477 (N_13477,N_11596,N_11201);
and U13478 (N_13478,N_9233,N_11380);
and U13479 (N_13479,N_10913,N_11953);
and U13480 (N_13480,N_10200,N_11752);
nand U13481 (N_13481,N_11151,N_9565);
and U13482 (N_13482,N_9367,N_10253);
nor U13483 (N_13483,N_9902,N_9044);
or U13484 (N_13484,N_11474,N_10280);
and U13485 (N_13485,N_11294,N_10136);
nor U13486 (N_13486,N_9779,N_9544);
nand U13487 (N_13487,N_9194,N_10652);
nor U13488 (N_13488,N_9349,N_9675);
nand U13489 (N_13489,N_11709,N_10952);
or U13490 (N_13490,N_10572,N_10271);
or U13491 (N_13491,N_10163,N_9101);
or U13492 (N_13492,N_9211,N_9524);
nor U13493 (N_13493,N_11513,N_11136);
or U13494 (N_13494,N_10922,N_10510);
or U13495 (N_13495,N_11728,N_10793);
or U13496 (N_13496,N_11315,N_11638);
nand U13497 (N_13497,N_10933,N_9457);
nor U13498 (N_13498,N_11746,N_9768);
nand U13499 (N_13499,N_11370,N_10138);
nor U13500 (N_13500,N_11863,N_11806);
nor U13501 (N_13501,N_11439,N_10553);
and U13502 (N_13502,N_10339,N_9627);
nand U13503 (N_13503,N_10453,N_11242);
nand U13504 (N_13504,N_11099,N_9174);
nor U13505 (N_13505,N_11048,N_11043);
nor U13506 (N_13506,N_11471,N_11591);
nor U13507 (N_13507,N_10334,N_11517);
and U13508 (N_13508,N_11694,N_10958);
or U13509 (N_13509,N_10107,N_11011);
nor U13510 (N_13510,N_10453,N_9815);
nand U13511 (N_13511,N_9929,N_11238);
nand U13512 (N_13512,N_11994,N_10349);
or U13513 (N_13513,N_10867,N_9140);
nand U13514 (N_13514,N_9357,N_10363);
or U13515 (N_13515,N_10470,N_9481);
nand U13516 (N_13516,N_10062,N_10702);
or U13517 (N_13517,N_11155,N_9893);
nor U13518 (N_13518,N_10570,N_10150);
nor U13519 (N_13519,N_9486,N_9333);
nor U13520 (N_13520,N_11072,N_9243);
or U13521 (N_13521,N_9377,N_9342);
or U13522 (N_13522,N_10016,N_9791);
and U13523 (N_13523,N_11900,N_10889);
nor U13524 (N_13524,N_11306,N_11957);
nand U13525 (N_13525,N_9851,N_10829);
nor U13526 (N_13526,N_11318,N_10844);
or U13527 (N_13527,N_9966,N_11573);
nor U13528 (N_13528,N_11980,N_11389);
nor U13529 (N_13529,N_11469,N_11237);
and U13530 (N_13530,N_11349,N_11071);
nand U13531 (N_13531,N_10085,N_9944);
or U13532 (N_13532,N_10239,N_10102);
nand U13533 (N_13533,N_10578,N_10692);
and U13534 (N_13534,N_10128,N_9038);
or U13535 (N_13535,N_10673,N_9989);
and U13536 (N_13536,N_9217,N_10154);
and U13537 (N_13537,N_11266,N_10785);
and U13538 (N_13538,N_11108,N_9426);
nand U13539 (N_13539,N_9445,N_10832);
and U13540 (N_13540,N_11753,N_11228);
and U13541 (N_13541,N_9879,N_10970);
or U13542 (N_13542,N_11499,N_9163);
and U13543 (N_13543,N_11076,N_10114);
and U13544 (N_13544,N_10155,N_11514);
nand U13545 (N_13545,N_10008,N_11403);
and U13546 (N_13546,N_10778,N_10122);
nor U13547 (N_13547,N_9632,N_10528);
or U13548 (N_13548,N_10694,N_9517);
or U13549 (N_13549,N_10930,N_11765);
nor U13550 (N_13550,N_10877,N_9387);
nand U13551 (N_13551,N_10353,N_11382);
nand U13552 (N_13552,N_11210,N_10292);
nor U13553 (N_13553,N_11069,N_10236);
nor U13554 (N_13554,N_10420,N_9231);
nor U13555 (N_13555,N_10948,N_9247);
nor U13556 (N_13556,N_10272,N_10780);
nand U13557 (N_13557,N_11161,N_10581);
xnor U13558 (N_13558,N_11276,N_9373);
and U13559 (N_13559,N_10775,N_10643);
and U13560 (N_13560,N_10556,N_11103);
and U13561 (N_13561,N_10098,N_9017);
nor U13562 (N_13562,N_11028,N_9292);
and U13563 (N_13563,N_10117,N_11940);
or U13564 (N_13564,N_10875,N_11365);
nor U13565 (N_13565,N_9523,N_9291);
and U13566 (N_13566,N_11466,N_10836);
or U13567 (N_13567,N_9743,N_11597);
nand U13568 (N_13568,N_9646,N_11467);
and U13569 (N_13569,N_9665,N_9951);
nand U13570 (N_13570,N_11666,N_9901);
or U13571 (N_13571,N_9054,N_9515);
nand U13572 (N_13572,N_9390,N_9538);
nor U13573 (N_13573,N_9141,N_10897);
and U13574 (N_13574,N_9930,N_10799);
nor U13575 (N_13575,N_9967,N_9814);
or U13576 (N_13576,N_10959,N_10717);
and U13577 (N_13577,N_10240,N_10399);
nand U13578 (N_13578,N_11965,N_11309);
or U13579 (N_13579,N_10605,N_9361);
or U13580 (N_13580,N_9734,N_10688);
nand U13581 (N_13581,N_11188,N_9950);
nand U13582 (N_13582,N_10596,N_10886);
or U13583 (N_13583,N_10926,N_11076);
nor U13584 (N_13584,N_10561,N_11205);
nand U13585 (N_13585,N_11407,N_9133);
or U13586 (N_13586,N_10629,N_11621);
or U13587 (N_13587,N_9637,N_10942);
and U13588 (N_13588,N_11291,N_11453);
or U13589 (N_13589,N_10931,N_9099);
nor U13590 (N_13590,N_11539,N_10322);
and U13591 (N_13591,N_9684,N_9875);
nand U13592 (N_13592,N_10944,N_9911);
or U13593 (N_13593,N_10490,N_11589);
or U13594 (N_13594,N_9753,N_11114);
nand U13595 (N_13595,N_11240,N_10100);
nand U13596 (N_13596,N_11157,N_10443);
or U13597 (N_13597,N_10862,N_11835);
and U13598 (N_13598,N_10053,N_11845);
nand U13599 (N_13599,N_10237,N_11310);
nor U13600 (N_13600,N_9993,N_10665);
nand U13601 (N_13601,N_10503,N_10050);
and U13602 (N_13602,N_9097,N_11990);
nand U13603 (N_13603,N_9156,N_9558);
and U13604 (N_13604,N_9147,N_9579);
nand U13605 (N_13605,N_11189,N_11160);
nand U13606 (N_13606,N_11196,N_11321);
nand U13607 (N_13607,N_9008,N_11307);
or U13608 (N_13608,N_9988,N_11250);
nand U13609 (N_13609,N_9223,N_11669);
nand U13610 (N_13610,N_10038,N_11439);
and U13611 (N_13611,N_11876,N_11110);
or U13612 (N_13612,N_10144,N_10887);
or U13613 (N_13613,N_9625,N_11707);
nor U13614 (N_13614,N_10657,N_10689);
nand U13615 (N_13615,N_11963,N_10229);
or U13616 (N_13616,N_10208,N_11992);
or U13617 (N_13617,N_10550,N_9210);
nor U13618 (N_13618,N_11740,N_9891);
nor U13619 (N_13619,N_10901,N_9068);
nand U13620 (N_13620,N_10642,N_10968);
and U13621 (N_13621,N_9428,N_11240);
nor U13622 (N_13622,N_9264,N_9113);
nand U13623 (N_13623,N_11897,N_11082);
nor U13624 (N_13624,N_10428,N_11252);
or U13625 (N_13625,N_9479,N_9051);
xnor U13626 (N_13626,N_10107,N_11715);
and U13627 (N_13627,N_9410,N_10982);
and U13628 (N_13628,N_10356,N_11759);
and U13629 (N_13629,N_10979,N_10753);
or U13630 (N_13630,N_9986,N_9382);
or U13631 (N_13631,N_9231,N_9339);
and U13632 (N_13632,N_9167,N_11166);
nor U13633 (N_13633,N_11486,N_10339);
nand U13634 (N_13634,N_9168,N_10112);
and U13635 (N_13635,N_9124,N_9496);
and U13636 (N_13636,N_11450,N_11984);
nand U13637 (N_13637,N_9765,N_9266);
and U13638 (N_13638,N_9953,N_9807);
and U13639 (N_13639,N_11095,N_9405);
nor U13640 (N_13640,N_10059,N_11365);
and U13641 (N_13641,N_9282,N_10617);
nand U13642 (N_13642,N_10927,N_10891);
and U13643 (N_13643,N_10436,N_9201);
nor U13644 (N_13644,N_10977,N_11459);
or U13645 (N_13645,N_9208,N_9776);
and U13646 (N_13646,N_10134,N_11955);
nand U13647 (N_13647,N_11303,N_11849);
nand U13648 (N_13648,N_10916,N_9808);
or U13649 (N_13649,N_9836,N_10780);
and U13650 (N_13650,N_9474,N_11861);
and U13651 (N_13651,N_10719,N_9375);
or U13652 (N_13652,N_9590,N_10010);
nand U13653 (N_13653,N_11345,N_11838);
nand U13654 (N_13654,N_9391,N_9102);
nand U13655 (N_13655,N_11193,N_9405);
and U13656 (N_13656,N_11151,N_9507);
or U13657 (N_13657,N_9543,N_10634);
nand U13658 (N_13658,N_10527,N_11559);
and U13659 (N_13659,N_10379,N_9202);
nand U13660 (N_13660,N_11487,N_11489);
nand U13661 (N_13661,N_9540,N_9376);
nand U13662 (N_13662,N_9633,N_11832);
nor U13663 (N_13663,N_9774,N_9581);
nor U13664 (N_13664,N_10159,N_9969);
nor U13665 (N_13665,N_10869,N_9626);
and U13666 (N_13666,N_10396,N_9449);
nor U13667 (N_13667,N_10069,N_9650);
nor U13668 (N_13668,N_10131,N_10172);
nand U13669 (N_13669,N_10009,N_10086);
and U13670 (N_13670,N_11793,N_9010);
nor U13671 (N_13671,N_10868,N_11319);
and U13672 (N_13672,N_11805,N_9997);
or U13673 (N_13673,N_10217,N_11489);
nand U13674 (N_13674,N_10983,N_10824);
or U13675 (N_13675,N_10255,N_10121);
or U13676 (N_13676,N_10805,N_9723);
and U13677 (N_13677,N_10218,N_9193);
nor U13678 (N_13678,N_11765,N_11464);
nor U13679 (N_13679,N_11882,N_11749);
nand U13680 (N_13680,N_10582,N_11692);
or U13681 (N_13681,N_9493,N_11611);
or U13682 (N_13682,N_9498,N_11603);
nor U13683 (N_13683,N_11523,N_11298);
nor U13684 (N_13684,N_9160,N_9597);
and U13685 (N_13685,N_9047,N_9901);
or U13686 (N_13686,N_11210,N_11867);
or U13687 (N_13687,N_10473,N_11916);
and U13688 (N_13688,N_9875,N_10241);
nor U13689 (N_13689,N_10008,N_11560);
nand U13690 (N_13690,N_9593,N_10012);
nor U13691 (N_13691,N_9132,N_9080);
nor U13692 (N_13692,N_11323,N_10141);
or U13693 (N_13693,N_11381,N_11986);
nand U13694 (N_13694,N_9751,N_10222);
nand U13695 (N_13695,N_10237,N_9083);
and U13696 (N_13696,N_9464,N_11502);
or U13697 (N_13697,N_9856,N_10927);
or U13698 (N_13698,N_11719,N_11965);
and U13699 (N_13699,N_10515,N_10730);
and U13700 (N_13700,N_10939,N_10369);
or U13701 (N_13701,N_10806,N_11737);
nor U13702 (N_13702,N_9991,N_9161);
or U13703 (N_13703,N_11172,N_10555);
and U13704 (N_13704,N_11386,N_11176);
or U13705 (N_13705,N_9473,N_9510);
and U13706 (N_13706,N_10404,N_9319);
nand U13707 (N_13707,N_10567,N_9223);
nor U13708 (N_13708,N_11177,N_9074);
nand U13709 (N_13709,N_11800,N_11011);
and U13710 (N_13710,N_9201,N_11532);
and U13711 (N_13711,N_9135,N_10466);
or U13712 (N_13712,N_10338,N_10470);
or U13713 (N_13713,N_10159,N_11910);
or U13714 (N_13714,N_11891,N_9634);
nor U13715 (N_13715,N_10372,N_11191);
nand U13716 (N_13716,N_10567,N_11132);
or U13717 (N_13717,N_9905,N_11980);
nand U13718 (N_13718,N_9156,N_11685);
and U13719 (N_13719,N_10438,N_10676);
nor U13720 (N_13720,N_10410,N_9134);
nand U13721 (N_13721,N_10881,N_10334);
nand U13722 (N_13722,N_11296,N_11779);
and U13723 (N_13723,N_9467,N_9302);
and U13724 (N_13724,N_9586,N_9243);
nor U13725 (N_13725,N_11166,N_11056);
nor U13726 (N_13726,N_9712,N_9128);
or U13727 (N_13727,N_9016,N_9823);
and U13728 (N_13728,N_10440,N_11379);
and U13729 (N_13729,N_9260,N_11113);
or U13730 (N_13730,N_11171,N_11273);
nor U13731 (N_13731,N_11422,N_10440);
nand U13732 (N_13732,N_9071,N_9738);
nor U13733 (N_13733,N_11536,N_10804);
nand U13734 (N_13734,N_9265,N_9458);
or U13735 (N_13735,N_10937,N_9382);
nor U13736 (N_13736,N_11441,N_9022);
or U13737 (N_13737,N_11022,N_10512);
and U13738 (N_13738,N_9180,N_10902);
nand U13739 (N_13739,N_11660,N_11760);
nand U13740 (N_13740,N_10829,N_10932);
and U13741 (N_13741,N_11291,N_10683);
nor U13742 (N_13742,N_10554,N_9362);
and U13743 (N_13743,N_10554,N_10988);
or U13744 (N_13744,N_11411,N_9151);
and U13745 (N_13745,N_11938,N_10778);
nor U13746 (N_13746,N_9256,N_9872);
or U13747 (N_13747,N_11532,N_11317);
or U13748 (N_13748,N_10313,N_9380);
nor U13749 (N_13749,N_10920,N_10687);
and U13750 (N_13750,N_10513,N_10231);
nand U13751 (N_13751,N_11801,N_11785);
nand U13752 (N_13752,N_9693,N_9487);
and U13753 (N_13753,N_10641,N_9843);
nand U13754 (N_13754,N_11150,N_9409);
or U13755 (N_13755,N_10138,N_10028);
and U13756 (N_13756,N_11417,N_11017);
and U13757 (N_13757,N_11044,N_11911);
nor U13758 (N_13758,N_9082,N_9672);
nor U13759 (N_13759,N_10599,N_9038);
nand U13760 (N_13760,N_11861,N_9710);
nand U13761 (N_13761,N_9005,N_10214);
nand U13762 (N_13762,N_11093,N_11102);
and U13763 (N_13763,N_10447,N_11606);
nor U13764 (N_13764,N_10367,N_10336);
or U13765 (N_13765,N_11520,N_11172);
or U13766 (N_13766,N_10577,N_10168);
and U13767 (N_13767,N_10347,N_9258);
nor U13768 (N_13768,N_11111,N_11112);
nor U13769 (N_13769,N_11177,N_11120);
nor U13770 (N_13770,N_9488,N_10485);
and U13771 (N_13771,N_10863,N_10209);
nor U13772 (N_13772,N_11630,N_10026);
nand U13773 (N_13773,N_9171,N_10230);
nor U13774 (N_13774,N_10668,N_9151);
or U13775 (N_13775,N_9223,N_9441);
nand U13776 (N_13776,N_9386,N_10900);
or U13777 (N_13777,N_11968,N_11206);
or U13778 (N_13778,N_9797,N_9937);
xnor U13779 (N_13779,N_10477,N_10532);
and U13780 (N_13780,N_10695,N_9006);
nor U13781 (N_13781,N_10561,N_11257);
nand U13782 (N_13782,N_9771,N_11883);
nor U13783 (N_13783,N_10414,N_10469);
or U13784 (N_13784,N_9667,N_9813);
and U13785 (N_13785,N_11526,N_10188);
nand U13786 (N_13786,N_9680,N_11923);
and U13787 (N_13787,N_9433,N_9752);
nand U13788 (N_13788,N_11122,N_9000);
or U13789 (N_13789,N_11961,N_10587);
nand U13790 (N_13790,N_10239,N_10966);
and U13791 (N_13791,N_10375,N_11062);
nor U13792 (N_13792,N_9178,N_9646);
or U13793 (N_13793,N_11401,N_9710);
nand U13794 (N_13794,N_10248,N_10329);
nor U13795 (N_13795,N_11566,N_10227);
nand U13796 (N_13796,N_11115,N_11023);
nor U13797 (N_13797,N_9947,N_9653);
nand U13798 (N_13798,N_9204,N_11583);
or U13799 (N_13799,N_11782,N_11745);
nand U13800 (N_13800,N_9364,N_10647);
nor U13801 (N_13801,N_9964,N_10733);
xor U13802 (N_13802,N_11370,N_11793);
nor U13803 (N_13803,N_10254,N_9227);
or U13804 (N_13804,N_10580,N_11401);
and U13805 (N_13805,N_10444,N_11870);
nand U13806 (N_13806,N_10078,N_9133);
or U13807 (N_13807,N_9661,N_9005);
nor U13808 (N_13808,N_10299,N_9771);
and U13809 (N_13809,N_11465,N_11596);
or U13810 (N_13810,N_11337,N_11317);
or U13811 (N_13811,N_9838,N_9222);
nand U13812 (N_13812,N_11954,N_11509);
nand U13813 (N_13813,N_10401,N_9695);
nor U13814 (N_13814,N_11563,N_9397);
nand U13815 (N_13815,N_11582,N_11306);
nand U13816 (N_13816,N_9291,N_10284);
nor U13817 (N_13817,N_10711,N_9451);
nor U13818 (N_13818,N_10615,N_9135);
and U13819 (N_13819,N_9110,N_11033);
or U13820 (N_13820,N_11821,N_11093);
or U13821 (N_13821,N_11710,N_9494);
and U13822 (N_13822,N_10659,N_9317);
nor U13823 (N_13823,N_9222,N_11283);
nor U13824 (N_13824,N_9402,N_9814);
nand U13825 (N_13825,N_10435,N_10505);
nor U13826 (N_13826,N_10965,N_9963);
nand U13827 (N_13827,N_10281,N_11699);
nand U13828 (N_13828,N_9104,N_9515);
or U13829 (N_13829,N_9701,N_11401);
or U13830 (N_13830,N_9860,N_11564);
nand U13831 (N_13831,N_9748,N_11989);
and U13832 (N_13832,N_10157,N_10958);
nand U13833 (N_13833,N_11452,N_10351);
nor U13834 (N_13834,N_10656,N_9989);
nand U13835 (N_13835,N_11661,N_11779);
and U13836 (N_13836,N_9027,N_11115);
nand U13837 (N_13837,N_9514,N_10410);
or U13838 (N_13838,N_10756,N_10657);
nor U13839 (N_13839,N_9199,N_9520);
xnor U13840 (N_13840,N_11156,N_11157);
or U13841 (N_13841,N_10985,N_10957);
nor U13842 (N_13842,N_11012,N_11969);
nand U13843 (N_13843,N_11167,N_10045);
and U13844 (N_13844,N_10257,N_10523);
and U13845 (N_13845,N_10425,N_9235);
and U13846 (N_13846,N_11023,N_11357);
nor U13847 (N_13847,N_11129,N_10947);
nand U13848 (N_13848,N_11465,N_11356);
or U13849 (N_13849,N_10638,N_11595);
xnor U13850 (N_13850,N_9045,N_9716);
or U13851 (N_13851,N_10728,N_10998);
or U13852 (N_13852,N_10329,N_11461);
nand U13853 (N_13853,N_9246,N_11942);
nand U13854 (N_13854,N_9540,N_9793);
nor U13855 (N_13855,N_11657,N_9752);
or U13856 (N_13856,N_10379,N_9669);
and U13857 (N_13857,N_9144,N_10761);
and U13858 (N_13858,N_11644,N_10055);
nand U13859 (N_13859,N_11281,N_11980);
or U13860 (N_13860,N_9708,N_10866);
nor U13861 (N_13861,N_9234,N_9931);
or U13862 (N_13862,N_11279,N_9076);
or U13863 (N_13863,N_9178,N_10364);
nand U13864 (N_13864,N_11111,N_10786);
and U13865 (N_13865,N_10388,N_10870);
or U13866 (N_13866,N_10088,N_9568);
nor U13867 (N_13867,N_11941,N_11230);
and U13868 (N_13868,N_11617,N_9361);
nand U13869 (N_13869,N_10342,N_11866);
or U13870 (N_13870,N_10681,N_10649);
or U13871 (N_13871,N_11453,N_10148);
or U13872 (N_13872,N_10094,N_10497);
or U13873 (N_13873,N_11161,N_10045);
nand U13874 (N_13874,N_10326,N_10565);
nor U13875 (N_13875,N_10632,N_9754);
or U13876 (N_13876,N_10267,N_10071);
or U13877 (N_13877,N_11618,N_11901);
nor U13878 (N_13878,N_10998,N_11640);
nor U13879 (N_13879,N_9113,N_9230);
or U13880 (N_13880,N_9133,N_9287);
and U13881 (N_13881,N_9159,N_11923);
xor U13882 (N_13882,N_10161,N_11608);
nand U13883 (N_13883,N_11810,N_10294);
or U13884 (N_13884,N_10724,N_11449);
nand U13885 (N_13885,N_9084,N_11774);
and U13886 (N_13886,N_11880,N_10024);
xor U13887 (N_13887,N_9615,N_11666);
or U13888 (N_13888,N_10567,N_10029);
or U13889 (N_13889,N_9185,N_10248);
nand U13890 (N_13890,N_11018,N_10496);
and U13891 (N_13891,N_10686,N_11358);
nor U13892 (N_13892,N_11569,N_10979);
nor U13893 (N_13893,N_11077,N_10148);
nor U13894 (N_13894,N_10107,N_11741);
nand U13895 (N_13895,N_10703,N_10725);
or U13896 (N_13896,N_10897,N_9493);
nand U13897 (N_13897,N_9015,N_10888);
or U13898 (N_13898,N_11233,N_10507);
or U13899 (N_13899,N_10655,N_9404);
or U13900 (N_13900,N_10139,N_10874);
or U13901 (N_13901,N_9668,N_9660);
nor U13902 (N_13902,N_9195,N_9467);
nand U13903 (N_13903,N_10805,N_9100);
or U13904 (N_13904,N_9327,N_9391);
nand U13905 (N_13905,N_11469,N_11882);
or U13906 (N_13906,N_9163,N_10861);
or U13907 (N_13907,N_9160,N_11270);
nor U13908 (N_13908,N_10063,N_10879);
nor U13909 (N_13909,N_11254,N_9054);
or U13910 (N_13910,N_11519,N_10410);
xnor U13911 (N_13911,N_10838,N_11646);
or U13912 (N_13912,N_11517,N_9122);
or U13913 (N_13913,N_10842,N_11124);
and U13914 (N_13914,N_9567,N_11242);
and U13915 (N_13915,N_9158,N_10732);
nand U13916 (N_13916,N_10238,N_9999);
nand U13917 (N_13917,N_11135,N_10206);
or U13918 (N_13918,N_10402,N_9411);
and U13919 (N_13919,N_10606,N_9243);
and U13920 (N_13920,N_11649,N_10535);
nor U13921 (N_13921,N_9204,N_10084);
and U13922 (N_13922,N_10448,N_9307);
nor U13923 (N_13923,N_9462,N_10020);
and U13924 (N_13924,N_11848,N_9555);
and U13925 (N_13925,N_9246,N_11026);
nor U13926 (N_13926,N_10548,N_10481);
nand U13927 (N_13927,N_11935,N_11377);
and U13928 (N_13928,N_11464,N_11231);
nand U13929 (N_13929,N_11313,N_10033);
or U13930 (N_13930,N_10875,N_9725);
nand U13931 (N_13931,N_11378,N_10929);
or U13932 (N_13932,N_10730,N_9490);
or U13933 (N_13933,N_11033,N_9216);
nor U13934 (N_13934,N_10960,N_11525);
and U13935 (N_13935,N_10040,N_11793);
or U13936 (N_13936,N_9862,N_11160);
nor U13937 (N_13937,N_11493,N_10129);
or U13938 (N_13938,N_11351,N_10934);
nor U13939 (N_13939,N_11044,N_11861);
or U13940 (N_13940,N_10326,N_10803);
nor U13941 (N_13941,N_9953,N_11344);
nand U13942 (N_13942,N_11441,N_10303);
and U13943 (N_13943,N_9977,N_9085);
and U13944 (N_13944,N_11189,N_9901);
nand U13945 (N_13945,N_10525,N_11768);
nor U13946 (N_13946,N_9212,N_10276);
nand U13947 (N_13947,N_11391,N_9194);
and U13948 (N_13948,N_9911,N_9316);
or U13949 (N_13949,N_9004,N_10574);
nor U13950 (N_13950,N_10307,N_11923);
and U13951 (N_13951,N_9638,N_9817);
and U13952 (N_13952,N_11899,N_9272);
nor U13953 (N_13953,N_11121,N_9416);
or U13954 (N_13954,N_9790,N_11589);
nor U13955 (N_13955,N_10964,N_10536);
or U13956 (N_13956,N_10970,N_9507);
nor U13957 (N_13957,N_9096,N_10310);
nor U13958 (N_13958,N_9768,N_9177);
nor U13959 (N_13959,N_10165,N_11991);
and U13960 (N_13960,N_10616,N_11666);
nand U13961 (N_13961,N_10160,N_10218);
and U13962 (N_13962,N_10525,N_9310);
nand U13963 (N_13963,N_11418,N_11083);
or U13964 (N_13964,N_9634,N_9845);
nor U13965 (N_13965,N_9593,N_9520);
xor U13966 (N_13966,N_9017,N_9684);
or U13967 (N_13967,N_11882,N_9812);
nand U13968 (N_13968,N_11440,N_11941);
and U13969 (N_13969,N_10673,N_10040);
and U13970 (N_13970,N_10055,N_9330);
xor U13971 (N_13971,N_10209,N_11412);
xnor U13972 (N_13972,N_10072,N_10675);
or U13973 (N_13973,N_9398,N_10921);
and U13974 (N_13974,N_10099,N_10100);
nand U13975 (N_13975,N_11278,N_10211);
and U13976 (N_13976,N_11955,N_9329);
or U13977 (N_13977,N_9496,N_11632);
nand U13978 (N_13978,N_11045,N_10834);
or U13979 (N_13979,N_10100,N_11780);
xor U13980 (N_13980,N_9299,N_11315);
nand U13981 (N_13981,N_10766,N_9605);
nor U13982 (N_13982,N_9887,N_9042);
nand U13983 (N_13983,N_11618,N_11799);
nor U13984 (N_13984,N_9048,N_9797);
nand U13985 (N_13985,N_11791,N_9302);
nor U13986 (N_13986,N_9549,N_9315);
and U13987 (N_13987,N_10609,N_10287);
and U13988 (N_13988,N_11695,N_10737);
and U13989 (N_13989,N_9442,N_9918);
or U13990 (N_13990,N_11710,N_9175);
nand U13991 (N_13991,N_11383,N_9083);
and U13992 (N_13992,N_9345,N_11680);
nor U13993 (N_13993,N_10875,N_9767);
and U13994 (N_13994,N_10232,N_10115);
nand U13995 (N_13995,N_11272,N_11964);
or U13996 (N_13996,N_10020,N_11172);
or U13997 (N_13997,N_9316,N_11181);
nand U13998 (N_13998,N_11985,N_10774);
nand U13999 (N_13999,N_9927,N_11695);
and U14000 (N_14000,N_9609,N_9937);
nand U14001 (N_14001,N_11352,N_11518);
and U14002 (N_14002,N_11135,N_9156);
nor U14003 (N_14003,N_10561,N_9432);
and U14004 (N_14004,N_9563,N_10277);
nand U14005 (N_14005,N_10711,N_10405);
and U14006 (N_14006,N_10731,N_9417);
or U14007 (N_14007,N_11901,N_9570);
and U14008 (N_14008,N_10512,N_11499);
nor U14009 (N_14009,N_9088,N_10593);
or U14010 (N_14010,N_11844,N_10863);
or U14011 (N_14011,N_10836,N_10269);
and U14012 (N_14012,N_11932,N_9496);
and U14013 (N_14013,N_11898,N_10389);
and U14014 (N_14014,N_9107,N_10414);
and U14015 (N_14015,N_11324,N_9337);
or U14016 (N_14016,N_11901,N_9124);
nor U14017 (N_14017,N_10732,N_9575);
nand U14018 (N_14018,N_11859,N_9277);
nand U14019 (N_14019,N_9813,N_11603);
nand U14020 (N_14020,N_9893,N_10541);
nand U14021 (N_14021,N_10530,N_10648);
and U14022 (N_14022,N_10332,N_11412);
and U14023 (N_14023,N_10203,N_11470);
nand U14024 (N_14024,N_10679,N_9647);
or U14025 (N_14025,N_9896,N_10171);
and U14026 (N_14026,N_11071,N_9032);
and U14027 (N_14027,N_11742,N_10518);
or U14028 (N_14028,N_10291,N_9656);
nor U14029 (N_14029,N_10619,N_11430);
and U14030 (N_14030,N_10822,N_10976);
nor U14031 (N_14031,N_10860,N_9761);
nor U14032 (N_14032,N_9260,N_11158);
or U14033 (N_14033,N_11649,N_11308);
nor U14034 (N_14034,N_10093,N_11300);
and U14035 (N_14035,N_10736,N_10094);
nand U14036 (N_14036,N_10630,N_11315);
and U14037 (N_14037,N_10385,N_9330);
nor U14038 (N_14038,N_9498,N_10486);
and U14039 (N_14039,N_10254,N_10196);
and U14040 (N_14040,N_11571,N_11365);
nand U14041 (N_14041,N_10403,N_9552);
nand U14042 (N_14042,N_9520,N_11713);
and U14043 (N_14043,N_10269,N_9343);
or U14044 (N_14044,N_10315,N_9525);
nor U14045 (N_14045,N_9708,N_9974);
or U14046 (N_14046,N_10968,N_10013);
nor U14047 (N_14047,N_10544,N_9686);
nor U14048 (N_14048,N_11545,N_11869);
or U14049 (N_14049,N_11296,N_10082);
and U14050 (N_14050,N_9342,N_10922);
nand U14051 (N_14051,N_10201,N_11922);
and U14052 (N_14052,N_11705,N_11950);
nor U14053 (N_14053,N_9660,N_10766);
or U14054 (N_14054,N_11206,N_11290);
nand U14055 (N_14055,N_9799,N_9363);
and U14056 (N_14056,N_11681,N_10164);
xnor U14057 (N_14057,N_9471,N_10740);
nand U14058 (N_14058,N_11880,N_9999);
nand U14059 (N_14059,N_10063,N_11448);
nor U14060 (N_14060,N_10202,N_9232);
nand U14061 (N_14061,N_9504,N_11369);
nor U14062 (N_14062,N_10317,N_11511);
nor U14063 (N_14063,N_11312,N_9002);
nor U14064 (N_14064,N_9936,N_11866);
nand U14065 (N_14065,N_9096,N_11779);
and U14066 (N_14066,N_11075,N_11124);
nor U14067 (N_14067,N_10271,N_9363);
and U14068 (N_14068,N_10800,N_11027);
nor U14069 (N_14069,N_9486,N_11822);
or U14070 (N_14070,N_10208,N_9258);
and U14071 (N_14071,N_11841,N_9321);
and U14072 (N_14072,N_10464,N_9962);
or U14073 (N_14073,N_10472,N_10093);
or U14074 (N_14074,N_11768,N_9409);
or U14075 (N_14075,N_11854,N_10829);
nand U14076 (N_14076,N_11626,N_11955);
nor U14077 (N_14077,N_9920,N_10475);
nor U14078 (N_14078,N_11846,N_10633);
nor U14079 (N_14079,N_10726,N_9122);
nand U14080 (N_14080,N_11875,N_9446);
and U14081 (N_14081,N_9991,N_9181);
and U14082 (N_14082,N_10506,N_11597);
nand U14083 (N_14083,N_10487,N_9529);
nor U14084 (N_14084,N_11380,N_10622);
and U14085 (N_14085,N_10793,N_9443);
or U14086 (N_14086,N_11620,N_11667);
nand U14087 (N_14087,N_11454,N_11271);
and U14088 (N_14088,N_11078,N_9223);
xor U14089 (N_14089,N_10511,N_9214);
nand U14090 (N_14090,N_11033,N_9666);
or U14091 (N_14091,N_11778,N_9704);
and U14092 (N_14092,N_10780,N_11093);
and U14093 (N_14093,N_10637,N_11377);
nand U14094 (N_14094,N_10128,N_10177);
nor U14095 (N_14095,N_10406,N_9393);
or U14096 (N_14096,N_10443,N_11831);
and U14097 (N_14097,N_10076,N_9411);
nand U14098 (N_14098,N_10077,N_11857);
nor U14099 (N_14099,N_11293,N_10555);
or U14100 (N_14100,N_10876,N_11092);
and U14101 (N_14101,N_9720,N_11004);
nand U14102 (N_14102,N_9869,N_11471);
nand U14103 (N_14103,N_9452,N_10771);
nand U14104 (N_14104,N_11963,N_10388);
and U14105 (N_14105,N_11573,N_11835);
or U14106 (N_14106,N_9127,N_9370);
xor U14107 (N_14107,N_11091,N_11165);
xor U14108 (N_14108,N_10478,N_11767);
nor U14109 (N_14109,N_11371,N_9957);
nand U14110 (N_14110,N_11657,N_11155);
and U14111 (N_14111,N_11380,N_10936);
nand U14112 (N_14112,N_9763,N_9311);
nand U14113 (N_14113,N_10048,N_9067);
xnor U14114 (N_14114,N_10104,N_10336);
or U14115 (N_14115,N_9558,N_10258);
and U14116 (N_14116,N_9589,N_11575);
or U14117 (N_14117,N_10311,N_9062);
or U14118 (N_14118,N_9996,N_11067);
nand U14119 (N_14119,N_10682,N_9135);
nor U14120 (N_14120,N_10964,N_11204);
nand U14121 (N_14121,N_11377,N_10673);
and U14122 (N_14122,N_10470,N_11282);
and U14123 (N_14123,N_9400,N_9473);
and U14124 (N_14124,N_10726,N_9944);
and U14125 (N_14125,N_9962,N_10425);
nor U14126 (N_14126,N_11113,N_11036);
or U14127 (N_14127,N_11972,N_11206);
and U14128 (N_14128,N_11984,N_9580);
nand U14129 (N_14129,N_10858,N_9955);
and U14130 (N_14130,N_11739,N_10986);
nand U14131 (N_14131,N_9526,N_9113);
nand U14132 (N_14132,N_9277,N_9357);
or U14133 (N_14133,N_9559,N_10312);
or U14134 (N_14134,N_9133,N_10546);
nor U14135 (N_14135,N_9551,N_11460);
nor U14136 (N_14136,N_11003,N_9543);
and U14137 (N_14137,N_9999,N_9703);
nand U14138 (N_14138,N_11732,N_11691);
nand U14139 (N_14139,N_9878,N_10002);
or U14140 (N_14140,N_9807,N_11662);
nor U14141 (N_14141,N_10896,N_9517);
nor U14142 (N_14142,N_11609,N_11732);
or U14143 (N_14143,N_10378,N_9112);
or U14144 (N_14144,N_11683,N_10430);
or U14145 (N_14145,N_11423,N_9927);
and U14146 (N_14146,N_11319,N_9462);
nor U14147 (N_14147,N_9962,N_9570);
nand U14148 (N_14148,N_11260,N_11763);
nand U14149 (N_14149,N_9803,N_11199);
and U14150 (N_14150,N_10218,N_10038);
and U14151 (N_14151,N_11890,N_10175);
and U14152 (N_14152,N_10421,N_9357);
nand U14153 (N_14153,N_11458,N_11120);
nand U14154 (N_14154,N_10411,N_11011);
and U14155 (N_14155,N_11766,N_10805);
or U14156 (N_14156,N_10946,N_11496);
nor U14157 (N_14157,N_11198,N_9169);
or U14158 (N_14158,N_9634,N_9956);
xor U14159 (N_14159,N_10783,N_9471);
and U14160 (N_14160,N_9757,N_10358);
or U14161 (N_14161,N_10167,N_9870);
and U14162 (N_14162,N_9666,N_9195);
nor U14163 (N_14163,N_9278,N_9504);
or U14164 (N_14164,N_10557,N_11614);
and U14165 (N_14165,N_9450,N_11192);
nand U14166 (N_14166,N_10830,N_11436);
and U14167 (N_14167,N_11887,N_11795);
and U14168 (N_14168,N_10024,N_10739);
or U14169 (N_14169,N_11524,N_11066);
or U14170 (N_14170,N_11098,N_9132);
or U14171 (N_14171,N_9294,N_9396);
nand U14172 (N_14172,N_10846,N_11148);
nor U14173 (N_14173,N_10637,N_11027);
and U14174 (N_14174,N_9418,N_9452);
and U14175 (N_14175,N_11543,N_9521);
or U14176 (N_14176,N_10872,N_10626);
or U14177 (N_14177,N_11831,N_9970);
and U14178 (N_14178,N_11092,N_11659);
nor U14179 (N_14179,N_10615,N_11589);
and U14180 (N_14180,N_10672,N_9159);
and U14181 (N_14181,N_10684,N_11745);
or U14182 (N_14182,N_10062,N_11754);
nand U14183 (N_14183,N_10007,N_9568);
or U14184 (N_14184,N_11822,N_10859);
or U14185 (N_14185,N_10051,N_9005);
nand U14186 (N_14186,N_9306,N_10695);
or U14187 (N_14187,N_9113,N_9687);
or U14188 (N_14188,N_10816,N_10664);
nand U14189 (N_14189,N_10563,N_10609);
xnor U14190 (N_14190,N_9332,N_10902);
or U14191 (N_14191,N_10113,N_10175);
nor U14192 (N_14192,N_9186,N_9119);
and U14193 (N_14193,N_11928,N_9757);
nand U14194 (N_14194,N_11982,N_10912);
nor U14195 (N_14195,N_11657,N_10871);
nor U14196 (N_14196,N_11079,N_9472);
xnor U14197 (N_14197,N_10312,N_10558);
nor U14198 (N_14198,N_11952,N_9392);
and U14199 (N_14199,N_10795,N_9035);
or U14200 (N_14200,N_10492,N_9056);
and U14201 (N_14201,N_11248,N_9535);
and U14202 (N_14202,N_10680,N_9210);
nor U14203 (N_14203,N_10791,N_9061);
nand U14204 (N_14204,N_11866,N_11819);
nand U14205 (N_14205,N_10199,N_11192);
and U14206 (N_14206,N_9596,N_11259);
nand U14207 (N_14207,N_11543,N_9312);
or U14208 (N_14208,N_11254,N_10510);
nand U14209 (N_14209,N_10782,N_9971);
nor U14210 (N_14210,N_10643,N_10417);
and U14211 (N_14211,N_10865,N_11737);
nand U14212 (N_14212,N_9582,N_11071);
nand U14213 (N_14213,N_9298,N_10386);
nor U14214 (N_14214,N_9024,N_11508);
nor U14215 (N_14215,N_11732,N_11044);
and U14216 (N_14216,N_11353,N_11983);
or U14217 (N_14217,N_10323,N_9328);
nand U14218 (N_14218,N_9878,N_9216);
and U14219 (N_14219,N_9718,N_9303);
nand U14220 (N_14220,N_9555,N_11597);
or U14221 (N_14221,N_10859,N_9400);
nand U14222 (N_14222,N_9823,N_9554);
nand U14223 (N_14223,N_10053,N_9989);
nand U14224 (N_14224,N_9062,N_10090);
nor U14225 (N_14225,N_9816,N_9997);
nor U14226 (N_14226,N_11297,N_11853);
nor U14227 (N_14227,N_10304,N_11496);
nor U14228 (N_14228,N_11236,N_11398);
nor U14229 (N_14229,N_11490,N_10721);
and U14230 (N_14230,N_11664,N_10280);
or U14231 (N_14231,N_9284,N_9158);
nand U14232 (N_14232,N_9893,N_9172);
nor U14233 (N_14233,N_11369,N_10279);
and U14234 (N_14234,N_9979,N_9814);
nand U14235 (N_14235,N_9720,N_11221);
or U14236 (N_14236,N_9758,N_9620);
nor U14237 (N_14237,N_10228,N_11230);
nor U14238 (N_14238,N_11323,N_10661);
or U14239 (N_14239,N_10368,N_11391);
or U14240 (N_14240,N_9343,N_11622);
nand U14241 (N_14241,N_9570,N_9564);
nand U14242 (N_14242,N_9111,N_10318);
and U14243 (N_14243,N_10532,N_9167);
nand U14244 (N_14244,N_11929,N_9610);
or U14245 (N_14245,N_11941,N_11468);
or U14246 (N_14246,N_11565,N_10516);
or U14247 (N_14247,N_10683,N_9805);
nor U14248 (N_14248,N_11802,N_11996);
nor U14249 (N_14249,N_11006,N_10912);
nor U14250 (N_14250,N_11281,N_10198);
and U14251 (N_14251,N_10123,N_9761);
or U14252 (N_14252,N_11959,N_9456);
nand U14253 (N_14253,N_10601,N_9537);
nor U14254 (N_14254,N_10870,N_11858);
xnor U14255 (N_14255,N_10406,N_11136);
nand U14256 (N_14256,N_10111,N_9792);
and U14257 (N_14257,N_9115,N_10379);
nor U14258 (N_14258,N_10931,N_9374);
nor U14259 (N_14259,N_11328,N_10116);
nor U14260 (N_14260,N_9258,N_9118);
or U14261 (N_14261,N_9861,N_10824);
nand U14262 (N_14262,N_10332,N_9823);
and U14263 (N_14263,N_11286,N_11719);
and U14264 (N_14264,N_10147,N_11639);
nand U14265 (N_14265,N_11798,N_10738);
or U14266 (N_14266,N_11143,N_10258);
or U14267 (N_14267,N_9727,N_10932);
and U14268 (N_14268,N_11285,N_10137);
nand U14269 (N_14269,N_9056,N_11880);
nand U14270 (N_14270,N_11026,N_11588);
and U14271 (N_14271,N_10249,N_11775);
nand U14272 (N_14272,N_11529,N_10903);
nand U14273 (N_14273,N_9292,N_9672);
nor U14274 (N_14274,N_11262,N_11877);
nor U14275 (N_14275,N_11082,N_10217);
or U14276 (N_14276,N_11928,N_9683);
and U14277 (N_14277,N_9708,N_9764);
or U14278 (N_14278,N_10891,N_9303);
or U14279 (N_14279,N_11443,N_11041);
nand U14280 (N_14280,N_10162,N_11473);
and U14281 (N_14281,N_10712,N_11205);
nand U14282 (N_14282,N_9140,N_10833);
and U14283 (N_14283,N_9541,N_10714);
and U14284 (N_14284,N_10197,N_10651);
and U14285 (N_14285,N_11114,N_9671);
nand U14286 (N_14286,N_11064,N_11372);
nand U14287 (N_14287,N_10400,N_10192);
nand U14288 (N_14288,N_9679,N_11701);
and U14289 (N_14289,N_10306,N_9549);
xor U14290 (N_14290,N_11729,N_11372);
and U14291 (N_14291,N_9699,N_11790);
nor U14292 (N_14292,N_11114,N_10851);
and U14293 (N_14293,N_9069,N_10600);
nand U14294 (N_14294,N_10236,N_9290);
or U14295 (N_14295,N_11125,N_10156);
nand U14296 (N_14296,N_11013,N_10196);
and U14297 (N_14297,N_11012,N_11195);
and U14298 (N_14298,N_9374,N_11938);
nand U14299 (N_14299,N_9789,N_11124);
xor U14300 (N_14300,N_10268,N_10719);
or U14301 (N_14301,N_11696,N_9414);
nor U14302 (N_14302,N_10183,N_9651);
nor U14303 (N_14303,N_10224,N_10732);
nand U14304 (N_14304,N_9970,N_9617);
nand U14305 (N_14305,N_11075,N_11056);
or U14306 (N_14306,N_9315,N_10600);
or U14307 (N_14307,N_10586,N_9969);
and U14308 (N_14308,N_11628,N_11144);
nand U14309 (N_14309,N_11544,N_10739);
and U14310 (N_14310,N_11053,N_11993);
nor U14311 (N_14311,N_11125,N_9339);
and U14312 (N_14312,N_10556,N_10142);
nor U14313 (N_14313,N_11905,N_11716);
nor U14314 (N_14314,N_9422,N_9467);
nand U14315 (N_14315,N_9984,N_11971);
and U14316 (N_14316,N_11623,N_11617);
and U14317 (N_14317,N_11345,N_10483);
or U14318 (N_14318,N_10782,N_10785);
or U14319 (N_14319,N_11185,N_10968);
or U14320 (N_14320,N_11362,N_10098);
nor U14321 (N_14321,N_11177,N_9995);
nor U14322 (N_14322,N_10103,N_10055);
or U14323 (N_14323,N_11450,N_9006);
nand U14324 (N_14324,N_10202,N_10244);
nor U14325 (N_14325,N_9571,N_11125);
nor U14326 (N_14326,N_10927,N_11538);
nor U14327 (N_14327,N_9876,N_11135);
or U14328 (N_14328,N_11682,N_11856);
nor U14329 (N_14329,N_9262,N_9228);
or U14330 (N_14330,N_10997,N_10646);
nand U14331 (N_14331,N_11443,N_9025);
nor U14332 (N_14332,N_11478,N_9088);
and U14333 (N_14333,N_11347,N_9657);
nand U14334 (N_14334,N_10412,N_11121);
nor U14335 (N_14335,N_11013,N_11548);
nor U14336 (N_14336,N_11536,N_11841);
nand U14337 (N_14337,N_10857,N_11942);
nand U14338 (N_14338,N_11767,N_10870);
nor U14339 (N_14339,N_11058,N_10681);
nor U14340 (N_14340,N_11502,N_11538);
nand U14341 (N_14341,N_10970,N_11130);
nand U14342 (N_14342,N_11896,N_11062);
nand U14343 (N_14343,N_11007,N_10825);
or U14344 (N_14344,N_10105,N_11958);
nand U14345 (N_14345,N_10630,N_10598);
or U14346 (N_14346,N_11880,N_10773);
and U14347 (N_14347,N_9005,N_10703);
nand U14348 (N_14348,N_10720,N_10823);
or U14349 (N_14349,N_9821,N_9250);
nor U14350 (N_14350,N_10782,N_10477);
or U14351 (N_14351,N_11222,N_9643);
or U14352 (N_14352,N_10667,N_10414);
and U14353 (N_14353,N_9778,N_11152);
nor U14354 (N_14354,N_11028,N_10160);
nor U14355 (N_14355,N_9736,N_11788);
and U14356 (N_14356,N_9617,N_9678);
nand U14357 (N_14357,N_9714,N_9120);
nand U14358 (N_14358,N_11876,N_10209);
or U14359 (N_14359,N_9498,N_11727);
and U14360 (N_14360,N_9613,N_11859);
or U14361 (N_14361,N_9451,N_11916);
nand U14362 (N_14362,N_11713,N_9860);
nand U14363 (N_14363,N_11721,N_9785);
and U14364 (N_14364,N_9363,N_10913);
and U14365 (N_14365,N_10089,N_11150);
xor U14366 (N_14366,N_11600,N_11774);
or U14367 (N_14367,N_10176,N_10445);
or U14368 (N_14368,N_10360,N_9359);
or U14369 (N_14369,N_11425,N_11416);
nand U14370 (N_14370,N_9274,N_9889);
and U14371 (N_14371,N_10558,N_9090);
and U14372 (N_14372,N_11089,N_9676);
nand U14373 (N_14373,N_10435,N_9137);
nor U14374 (N_14374,N_9856,N_11247);
nor U14375 (N_14375,N_10316,N_11836);
nand U14376 (N_14376,N_11347,N_10480);
or U14377 (N_14377,N_9921,N_11731);
or U14378 (N_14378,N_10822,N_10236);
nand U14379 (N_14379,N_11529,N_10799);
nor U14380 (N_14380,N_9522,N_10280);
and U14381 (N_14381,N_10078,N_11946);
or U14382 (N_14382,N_10653,N_9247);
nor U14383 (N_14383,N_9688,N_9870);
nor U14384 (N_14384,N_9867,N_10926);
or U14385 (N_14385,N_9882,N_9579);
xnor U14386 (N_14386,N_10523,N_10181);
nand U14387 (N_14387,N_10996,N_11611);
or U14388 (N_14388,N_10705,N_9025);
nor U14389 (N_14389,N_9362,N_9404);
or U14390 (N_14390,N_10804,N_10537);
nor U14391 (N_14391,N_10431,N_11915);
nor U14392 (N_14392,N_10602,N_11117);
and U14393 (N_14393,N_10836,N_10869);
or U14394 (N_14394,N_9748,N_9787);
nor U14395 (N_14395,N_9158,N_10171);
nand U14396 (N_14396,N_11285,N_11024);
nand U14397 (N_14397,N_9201,N_9353);
and U14398 (N_14398,N_9174,N_11412);
nor U14399 (N_14399,N_9423,N_10139);
or U14400 (N_14400,N_9805,N_11375);
and U14401 (N_14401,N_11995,N_9532);
nor U14402 (N_14402,N_10543,N_10978);
and U14403 (N_14403,N_10251,N_10260);
nor U14404 (N_14404,N_9363,N_11719);
nor U14405 (N_14405,N_10634,N_9612);
nand U14406 (N_14406,N_9409,N_10860);
nor U14407 (N_14407,N_11627,N_11186);
or U14408 (N_14408,N_10162,N_9739);
or U14409 (N_14409,N_9522,N_10672);
nand U14410 (N_14410,N_9732,N_10477);
or U14411 (N_14411,N_10326,N_10254);
nand U14412 (N_14412,N_10469,N_11322);
or U14413 (N_14413,N_9991,N_9080);
and U14414 (N_14414,N_10387,N_10613);
nor U14415 (N_14415,N_11056,N_10693);
or U14416 (N_14416,N_9491,N_10821);
nor U14417 (N_14417,N_11238,N_9998);
and U14418 (N_14418,N_10903,N_10774);
nor U14419 (N_14419,N_11640,N_10911);
nor U14420 (N_14420,N_10733,N_9135);
and U14421 (N_14421,N_11081,N_11871);
or U14422 (N_14422,N_10572,N_11906);
nand U14423 (N_14423,N_10020,N_11728);
nand U14424 (N_14424,N_9021,N_9675);
nand U14425 (N_14425,N_9502,N_9904);
and U14426 (N_14426,N_10619,N_11622);
and U14427 (N_14427,N_11661,N_11969);
and U14428 (N_14428,N_9589,N_11553);
nand U14429 (N_14429,N_9207,N_10266);
or U14430 (N_14430,N_11358,N_9083);
nand U14431 (N_14431,N_11118,N_11058);
nor U14432 (N_14432,N_11617,N_10678);
or U14433 (N_14433,N_9411,N_10436);
nand U14434 (N_14434,N_10954,N_9982);
nor U14435 (N_14435,N_9763,N_11008);
nor U14436 (N_14436,N_9423,N_10712);
nand U14437 (N_14437,N_9145,N_9938);
and U14438 (N_14438,N_9115,N_11010);
and U14439 (N_14439,N_9914,N_11702);
or U14440 (N_14440,N_9052,N_10310);
or U14441 (N_14441,N_9552,N_11146);
and U14442 (N_14442,N_9165,N_9649);
nor U14443 (N_14443,N_9309,N_11967);
nand U14444 (N_14444,N_10030,N_11762);
and U14445 (N_14445,N_9290,N_11745);
nor U14446 (N_14446,N_9601,N_10052);
nor U14447 (N_14447,N_10310,N_9764);
nor U14448 (N_14448,N_10306,N_10618);
nand U14449 (N_14449,N_11267,N_10034);
nor U14450 (N_14450,N_10778,N_11280);
or U14451 (N_14451,N_10378,N_10737);
nand U14452 (N_14452,N_11458,N_9942);
nand U14453 (N_14453,N_10289,N_11452);
nor U14454 (N_14454,N_9650,N_11228);
or U14455 (N_14455,N_11908,N_11915);
nand U14456 (N_14456,N_11011,N_9469);
nand U14457 (N_14457,N_11848,N_10050);
or U14458 (N_14458,N_11924,N_10756);
or U14459 (N_14459,N_11488,N_10032);
or U14460 (N_14460,N_11921,N_11533);
nor U14461 (N_14461,N_9081,N_9782);
xor U14462 (N_14462,N_11716,N_11682);
nand U14463 (N_14463,N_11267,N_11259);
nand U14464 (N_14464,N_10829,N_9262);
and U14465 (N_14465,N_10130,N_9967);
nor U14466 (N_14466,N_10064,N_10153);
and U14467 (N_14467,N_9387,N_11101);
nand U14468 (N_14468,N_11727,N_11991);
nor U14469 (N_14469,N_9584,N_9069);
nor U14470 (N_14470,N_9118,N_11858);
and U14471 (N_14471,N_11459,N_10913);
and U14472 (N_14472,N_10931,N_9925);
nor U14473 (N_14473,N_9316,N_10108);
and U14474 (N_14474,N_9993,N_9233);
and U14475 (N_14475,N_9645,N_10177);
nor U14476 (N_14476,N_9172,N_10385);
nand U14477 (N_14477,N_11606,N_11324);
nand U14478 (N_14478,N_10937,N_9259);
and U14479 (N_14479,N_9368,N_10224);
nor U14480 (N_14480,N_9148,N_11208);
nor U14481 (N_14481,N_10029,N_9115);
or U14482 (N_14482,N_11109,N_9183);
nor U14483 (N_14483,N_10790,N_10434);
or U14484 (N_14484,N_10093,N_10124);
nor U14485 (N_14485,N_10236,N_10649);
nand U14486 (N_14486,N_10134,N_9877);
nor U14487 (N_14487,N_9058,N_9134);
and U14488 (N_14488,N_10540,N_9491);
or U14489 (N_14489,N_11387,N_11424);
and U14490 (N_14490,N_9700,N_9513);
nor U14491 (N_14491,N_9574,N_10536);
nor U14492 (N_14492,N_10104,N_9522);
nor U14493 (N_14493,N_11939,N_9051);
nor U14494 (N_14494,N_9273,N_10988);
nand U14495 (N_14495,N_11832,N_10472);
and U14496 (N_14496,N_11278,N_11019);
and U14497 (N_14497,N_11203,N_10555);
and U14498 (N_14498,N_11696,N_10445);
nor U14499 (N_14499,N_10960,N_11246);
and U14500 (N_14500,N_11165,N_11377);
nand U14501 (N_14501,N_11041,N_11994);
or U14502 (N_14502,N_11677,N_11609);
and U14503 (N_14503,N_10515,N_11370);
and U14504 (N_14504,N_11435,N_10953);
or U14505 (N_14505,N_9273,N_11351);
nand U14506 (N_14506,N_11761,N_9635);
nand U14507 (N_14507,N_10503,N_11724);
and U14508 (N_14508,N_9724,N_11905);
nand U14509 (N_14509,N_10165,N_11290);
nand U14510 (N_14510,N_10528,N_11064);
and U14511 (N_14511,N_10558,N_11458);
nor U14512 (N_14512,N_10749,N_9625);
nand U14513 (N_14513,N_10109,N_10350);
nand U14514 (N_14514,N_10762,N_11096);
or U14515 (N_14515,N_10235,N_11248);
nor U14516 (N_14516,N_9671,N_10405);
and U14517 (N_14517,N_9493,N_10011);
nor U14518 (N_14518,N_10227,N_10230);
nand U14519 (N_14519,N_10195,N_11822);
nand U14520 (N_14520,N_9221,N_9337);
and U14521 (N_14521,N_10548,N_9866);
and U14522 (N_14522,N_9433,N_11978);
or U14523 (N_14523,N_10389,N_11737);
or U14524 (N_14524,N_11124,N_11183);
nor U14525 (N_14525,N_9069,N_10386);
nand U14526 (N_14526,N_9965,N_9683);
or U14527 (N_14527,N_9634,N_9915);
or U14528 (N_14528,N_9758,N_11712);
nor U14529 (N_14529,N_10714,N_11563);
or U14530 (N_14530,N_9468,N_10164);
nor U14531 (N_14531,N_11304,N_9395);
and U14532 (N_14532,N_10747,N_10289);
nand U14533 (N_14533,N_9295,N_10430);
or U14534 (N_14534,N_10717,N_10827);
nand U14535 (N_14535,N_11197,N_11511);
nand U14536 (N_14536,N_10376,N_9985);
and U14537 (N_14537,N_10933,N_11122);
or U14538 (N_14538,N_9386,N_10821);
nand U14539 (N_14539,N_10668,N_11577);
nor U14540 (N_14540,N_9966,N_9266);
or U14541 (N_14541,N_10203,N_10401);
nor U14542 (N_14542,N_9534,N_10795);
and U14543 (N_14543,N_11574,N_9625);
and U14544 (N_14544,N_9352,N_9637);
nor U14545 (N_14545,N_9467,N_11121);
or U14546 (N_14546,N_10493,N_11570);
nor U14547 (N_14547,N_11899,N_11903);
and U14548 (N_14548,N_9051,N_9415);
xnor U14549 (N_14549,N_9222,N_9932);
or U14550 (N_14550,N_10018,N_11691);
xnor U14551 (N_14551,N_10483,N_11933);
nor U14552 (N_14552,N_11071,N_9241);
and U14553 (N_14553,N_9198,N_9300);
nand U14554 (N_14554,N_9040,N_11152);
nand U14555 (N_14555,N_10418,N_9168);
nand U14556 (N_14556,N_11660,N_11964);
or U14557 (N_14557,N_10818,N_11364);
nand U14558 (N_14558,N_9738,N_9029);
nand U14559 (N_14559,N_9044,N_11467);
and U14560 (N_14560,N_9194,N_10051);
nor U14561 (N_14561,N_10563,N_10392);
or U14562 (N_14562,N_10490,N_11652);
nor U14563 (N_14563,N_10706,N_9559);
nand U14564 (N_14564,N_11459,N_10496);
nand U14565 (N_14565,N_9198,N_10261);
and U14566 (N_14566,N_11798,N_10270);
nand U14567 (N_14567,N_10044,N_9356);
and U14568 (N_14568,N_11519,N_11009);
and U14569 (N_14569,N_9656,N_9620);
nor U14570 (N_14570,N_11962,N_9560);
and U14571 (N_14571,N_11695,N_9140);
nor U14572 (N_14572,N_9630,N_10796);
or U14573 (N_14573,N_11338,N_9943);
nor U14574 (N_14574,N_11963,N_9454);
and U14575 (N_14575,N_10910,N_10420);
and U14576 (N_14576,N_9326,N_11475);
and U14577 (N_14577,N_9267,N_10794);
or U14578 (N_14578,N_10633,N_9313);
nor U14579 (N_14579,N_10046,N_11520);
nand U14580 (N_14580,N_11976,N_10767);
nand U14581 (N_14581,N_10070,N_11594);
or U14582 (N_14582,N_10395,N_11906);
or U14583 (N_14583,N_11213,N_9301);
and U14584 (N_14584,N_11792,N_9689);
and U14585 (N_14585,N_10568,N_11340);
or U14586 (N_14586,N_10127,N_9782);
nor U14587 (N_14587,N_10283,N_9529);
and U14588 (N_14588,N_9658,N_9376);
nand U14589 (N_14589,N_11666,N_9046);
nor U14590 (N_14590,N_9434,N_10784);
nand U14591 (N_14591,N_10465,N_10510);
and U14592 (N_14592,N_9880,N_9025);
xnor U14593 (N_14593,N_9471,N_11297);
or U14594 (N_14594,N_9250,N_10856);
nand U14595 (N_14595,N_10948,N_10490);
nand U14596 (N_14596,N_9754,N_10196);
nor U14597 (N_14597,N_10634,N_11518);
nand U14598 (N_14598,N_9742,N_10834);
nor U14599 (N_14599,N_9788,N_10535);
nor U14600 (N_14600,N_9986,N_9000);
or U14601 (N_14601,N_11896,N_9852);
or U14602 (N_14602,N_9109,N_10350);
and U14603 (N_14603,N_11637,N_11248);
or U14604 (N_14604,N_9588,N_10746);
and U14605 (N_14605,N_11469,N_11100);
and U14606 (N_14606,N_11819,N_9877);
or U14607 (N_14607,N_9973,N_9961);
and U14608 (N_14608,N_11170,N_9152);
and U14609 (N_14609,N_11793,N_11849);
and U14610 (N_14610,N_11338,N_11708);
nor U14611 (N_14611,N_9220,N_10406);
nor U14612 (N_14612,N_9742,N_11257);
nand U14613 (N_14613,N_11766,N_11971);
nor U14614 (N_14614,N_10304,N_10660);
and U14615 (N_14615,N_9820,N_9429);
and U14616 (N_14616,N_9245,N_11929);
and U14617 (N_14617,N_10889,N_11175);
or U14618 (N_14618,N_11088,N_9411);
or U14619 (N_14619,N_10204,N_9250);
nor U14620 (N_14620,N_10356,N_9627);
nor U14621 (N_14621,N_11452,N_11822);
nand U14622 (N_14622,N_10854,N_10005);
and U14623 (N_14623,N_10088,N_10117);
or U14624 (N_14624,N_9142,N_10581);
nor U14625 (N_14625,N_10494,N_9992);
and U14626 (N_14626,N_10166,N_9759);
and U14627 (N_14627,N_10027,N_10486);
or U14628 (N_14628,N_10630,N_11397);
or U14629 (N_14629,N_9361,N_10270);
nor U14630 (N_14630,N_10263,N_9773);
nor U14631 (N_14631,N_10827,N_9504);
or U14632 (N_14632,N_11557,N_10197);
nor U14633 (N_14633,N_10520,N_10914);
and U14634 (N_14634,N_9133,N_11270);
or U14635 (N_14635,N_11538,N_9187);
or U14636 (N_14636,N_9390,N_11845);
and U14637 (N_14637,N_10596,N_10111);
and U14638 (N_14638,N_10715,N_9519);
nor U14639 (N_14639,N_10272,N_11803);
nor U14640 (N_14640,N_11074,N_10547);
nand U14641 (N_14641,N_9991,N_10195);
or U14642 (N_14642,N_10772,N_9808);
nor U14643 (N_14643,N_10458,N_9044);
nand U14644 (N_14644,N_10142,N_9512);
and U14645 (N_14645,N_9045,N_10908);
nor U14646 (N_14646,N_11936,N_10058);
or U14647 (N_14647,N_9368,N_11292);
and U14648 (N_14648,N_11597,N_9639);
and U14649 (N_14649,N_11769,N_11371);
and U14650 (N_14650,N_9689,N_9976);
nand U14651 (N_14651,N_11184,N_10725);
and U14652 (N_14652,N_10743,N_10706);
and U14653 (N_14653,N_9130,N_11028);
nor U14654 (N_14654,N_10046,N_9414);
nor U14655 (N_14655,N_11058,N_11626);
or U14656 (N_14656,N_9370,N_9252);
nand U14657 (N_14657,N_9275,N_10147);
or U14658 (N_14658,N_11127,N_11939);
nand U14659 (N_14659,N_9299,N_11671);
nor U14660 (N_14660,N_10324,N_11790);
or U14661 (N_14661,N_9042,N_10643);
xnor U14662 (N_14662,N_9720,N_9659);
nand U14663 (N_14663,N_10957,N_10340);
and U14664 (N_14664,N_10415,N_11318);
and U14665 (N_14665,N_11031,N_9504);
nor U14666 (N_14666,N_9010,N_9857);
or U14667 (N_14667,N_11663,N_10023);
nand U14668 (N_14668,N_10116,N_11831);
nand U14669 (N_14669,N_11933,N_10450);
nor U14670 (N_14670,N_11074,N_9114);
xnor U14671 (N_14671,N_10716,N_10254);
or U14672 (N_14672,N_9045,N_10792);
or U14673 (N_14673,N_10404,N_11682);
or U14674 (N_14674,N_11972,N_9583);
nor U14675 (N_14675,N_10629,N_10922);
or U14676 (N_14676,N_10839,N_9606);
nor U14677 (N_14677,N_10905,N_10472);
nand U14678 (N_14678,N_9825,N_10228);
or U14679 (N_14679,N_11479,N_9308);
nor U14680 (N_14680,N_9155,N_11279);
nor U14681 (N_14681,N_9428,N_11451);
and U14682 (N_14682,N_9464,N_10027);
and U14683 (N_14683,N_10509,N_10501);
xnor U14684 (N_14684,N_9380,N_10751);
or U14685 (N_14685,N_10976,N_10560);
nor U14686 (N_14686,N_9919,N_9567);
nand U14687 (N_14687,N_11841,N_11522);
nor U14688 (N_14688,N_11439,N_9665);
or U14689 (N_14689,N_9794,N_10412);
or U14690 (N_14690,N_10459,N_9630);
nor U14691 (N_14691,N_9228,N_11722);
nand U14692 (N_14692,N_9884,N_9883);
and U14693 (N_14693,N_10671,N_9267);
and U14694 (N_14694,N_9637,N_11898);
and U14695 (N_14695,N_10618,N_9182);
or U14696 (N_14696,N_11458,N_9459);
nor U14697 (N_14697,N_9757,N_11724);
nand U14698 (N_14698,N_10836,N_9214);
or U14699 (N_14699,N_9817,N_9443);
nand U14700 (N_14700,N_10593,N_9896);
nor U14701 (N_14701,N_10836,N_9698);
or U14702 (N_14702,N_9760,N_10241);
or U14703 (N_14703,N_11226,N_9702);
or U14704 (N_14704,N_11424,N_11601);
or U14705 (N_14705,N_10825,N_11552);
nand U14706 (N_14706,N_10966,N_11080);
xor U14707 (N_14707,N_9369,N_11597);
nand U14708 (N_14708,N_11915,N_9541);
or U14709 (N_14709,N_11230,N_10194);
or U14710 (N_14710,N_10705,N_11410);
nor U14711 (N_14711,N_10638,N_11577);
nand U14712 (N_14712,N_9405,N_10516);
and U14713 (N_14713,N_11191,N_9469);
and U14714 (N_14714,N_9102,N_10943);
and U14715 (N_14715,N_11718,N_9272);
or U14716 (N_14716,N_9397,N_11130);
or U14717 (N_14717,N_10135,N_10992);
nand U14718 (N_14718,N_10439,N_9858);
nand U14719 (N_14719,N_11893,N_10669);
nand U14720 (N_14720,N_10376,N_9836);
and U14721 (N_14721,N_10714,N_9004);
and U14722 (N_14722,N_10231,N_10290);
or U14723 (N_14723,N_11972,N_9150);
nand U14724 (N_14724,N_11396,N_11381);
or U14725 (N_14725,N_9987,N_11888);
nand U14726 (N_14726,N_9491,N_10681);
or U14727 (N_14727,N_11964,N_10612);
and U14728 (N_14728,N_10990,N_10923);
nor U14729 (N_14729,N_9469,N_11951);
nor U14730 (N_14730,N_9483,N_11732);
nor U14731 (N_14731,N_11162,N_10237);
and U14732 (N_14732,N_10458,N_9038);
or U14733 (N_14733,N_10069,N_9757);
nor U14734 (N_14734,N_10291,N_9583);
xnor U14735 (N_14735,N_9831,N_9016);
or U14736 (N_14736,N_9137,N_9838);
and U14737 (N_14737,N_9769,N_10150);
nand U14738 (N_14738,N_11310,N_11052);
and U14739 (N_14739,N_9822,N_10716);
nand U14740 (N_14740,N_9039,N_10068);
nor U14741 (N_14741,N_11517,N_10080);
and U14742 (N_14742,N_10418,N_11514);
nor U14743 (N_14743,N_9843,N_9666);
and U14744 (N_14744,N_10116,N_10686);
or U14745 (N_14745,N_9901,N_9555);
or U14746 (N_14746,N_11000,N_11474);
and U14747 (N_14747,N_10059,N_9173);
and U14748 (N_14748,N_11928,N_10846);
or U14749 (N_14749,N_9468,N_9112);
and U14750 (N_14750,N_10353,N_9224);
nor U14751 (N_14751,N_10109,N_9263);
nand U14752 (N_14752,N_10285,N_9555);
or U14753 (N_14753,N_11441,N_11609);
nand U14754 (N_14754,N_11974,N_10691);
nor U14755 (N_14755,N_11401,N_10699);
nor U14756 (N_14756,N_9107,N_11492);
nor U14757 (N_14757,N_10352,N_11302);
and U14758 (N_14758,N_10344,N_11878);
and U14759 (N_14759,N_9450,N_11461);
or U14760 (N_14760,N_10221,N_10974);
nor U14761 (N_14761,N_10233,N_9056);
nor U14762 (N_14762,N_9895,N_10214);
nand U14763 (N_14763,N_9321,N_9578);
nor U14764 (N_14764,N_9495,N_11328);
and U14765 (N_14765,N_11762,N_9550);
nand U14766 (N_14766,N_9303,N_9206);
nand U14767 (N_14767,N_10262,N_11826);
nor U14768 (N_14768,N_9545,N_11694);
nor U14769 (N_14769,N_9349,N_10945);
nand U14770 (N_14770,N_11032,N_9945);
and U14771 (N_14771,N_9743,N_10247);
nor U14772 (N_14772,N_10473,N_10185);
nor U14773 (N_14773,N_9096,N_9363);
nor U14774 (N_14774,N_9234,N_10282);
or U14775 (N_14775,N_10591,N_10974);
and U14776 (N_14776,N_9293,N_9085);
nand U14777 (N_14777,N_11403,N_9773);
and U14778 (N_14778,N_11263,N_11609);
xor U14779 (N_14779,N_11956,N_9890);
and U14780 (N_14780,N_9798,N_9319);
and U14781 (N_14781,N_9107,N_10476);
and U14782 (N_14782,N_9363,N_10395);
and U14783 (N_14783,N_11662,N_10932);
and U14784 (N_14784,N_9834,N_9957);
and U14785 (N_14785,N_10138,N_9068);
nand U14786 (N_14786,N_10645,N_11479);
and U14787 (N_14787,N_11703,N_10762);
nor U14788 (N_14788,N_11348,N_11141);
nand U14789 (N_14789,N_10928,N_11870);
and U14790 (N_14790,N_10381,N_9622);
nand U14791 (N_14791,N_9966,N_9519);
nor U14792 (N_14792,N_11541,N_10991);
or U14793 (N_14793,N_10427,N_10654);
nand U14794 (N_14794,N_11787,N_11035);
nor U14795 (N_14795,N_10845,N_10105);
and U14796 (N_14796,N_9354,N_10205);
nor U14797 (N_14797,N_9052,N_11886);
nand U14798 (N_14798,N_10052,N_9977);
nand U14799 (N_14799,N_11319,N_10804);
and U14800 (N_14800,N_11877,N_9932);
nor U14801 (N_14801,N_10535,N_10345);
nand U14802 (N_14802,N_11959,N_11235);
and U14803 (N_14803,N_11243,N_9516);
nor U14804 (N_14804,N_9795,N_9686);
or U14805 (N_14805,N_10464,N_11474);
or U14806 (N_14806,N_9946,N_9310);
nor U14807 (N_14807,N_11646,N_11261);
nor U14808 (N_14808,N_11825,N_10216);
nand U14809 (N_14809,N_9844,N_11488);
nor U14810 (N_14810,N_10276,N_11868);
and U14811 (N_14811,N_11148,N_10902);
nor U14812 (N_14812,N_9818,N_10819);
or U14813 (N_14813,N_10440,N_11998);
nand U14814 (N_14814,N_9542,N_10703);
nand U14815 (N_14815,N_9790,N_9547);
xor U14816 (N_14816,N_9707,N_11502);
nor U14817 (N_14817,N_10983,N_9988);
nand U14818 (N_14818,N_11123,N_9487);
and U14819 (N_14819,N_11590,N_10352);
and U14820 (N_14820,N_11953,N_10837);
or U14821 (N_14821,N_9020,N_9365);
nand U14822 (N_14822,N_9896,N_10392);
xnor U14823 (N_14823,N_11981,N_10737);
nor U14824 (N_14824,N_9689,N_9673);
and U14825 (N_14825,N_9231,N_9662);
nand U14826 (N_14826,N_10885,N_10427);
nand U14827 (N_14827,N_11095,N_11151);
or U14828 (N_14828,N_11180,N_9475);
or U14829 (N_14829,N_10196,N_9300);
or U14830 (N_14830,N_11313,N_9166);
nand U14831 (N_14831,N_9524,N_10464);
nand U14832 (N_14832,N_11179,N_11158);
nor U14833 (N_14833,N_9194,N_11620);
nor U14834 (N_14834,N_10300,N_9877);
nor U14835 (N_14835,N_11769,N_11017);
xor U14836 (N_14836,N_9838,N_9141);
or U14837 (N_14837,N_10167,N_9231);
or U14838 (N_14838,N_10890,N_10697);
nor U14839 (N_14839,N_11049,N_10077);
or U14840 (N_14840,N_11274,N_9316);
or U14841 (N_14841,N_11611,N_11357);
nor U14842 (N_14842,N_11886,N_9835);
or U14843 (N_14843,N_10155,N_10800);
and U14844 (N_14844,N_10952,N_10848);
and U14845 (N_14845,N_9714,N_11657);
or U14846 (N_14846,N_11031,N_9178);
nor U14847 (N_14847,N_11626,N_10783);
or U14848 (N_14848,N_11089,N_9698);
nor U14849 (N_14849,N_9842,N_9453);
nand U14850 (N_14850,N_11584,N_11394);
nand U14851 (N_14851,N_11512,N_11411);
or U14852 (N_14852,N_9925,N_10661);
or U14853 (N_14853,N_11073,N_11932);
nand U14854 (N_14854,N_11804,N_11383);
nor U14855 (N_14855,N_10555,N_10801);
nor U14856 (N_14856,N_10887,N_9629);
nand U14857 (N_14857,N_11597,N_11820);
or U14858 (N_14858,N_11035,N_9599);
or U14859 (N_14859,N_11230,N_9959);
or U14860 (N_14860,N_10279,N_10885);
or U14861 (N_14861,N_11396,N_9438);
and U14862 (N_14862,N_9498,N_11747);
and U14863 (N_14863,N_11559,N_10066);
and U14864 (N_14864,N_10117,N_11240);
and U14865 (N_14865,N_9962,N_10804);
and U14866 (N_14866,N_9836,N_10987);
or U14867 (N_14867,N_10113,N_9585);
or U14868 (N_14868,N_9438,N_9366);
and U14869 (N_14869,N_10756,N_11632);
nor U14870 (N_14870,N_9486,N_9699);
and U14871 (N_14871,N_10291,N_10448);
and U14872 (N_14872,N_11896,N_10011);
nand U14873 (N_14873,N_11190,N_10090);
and U14874 (N_14874,N_9545,N_9136);
nor U14875 (N_14875,N_10663,N_11453);
nand U14876 (N_14876,N_11046,N_9933);
and U14877 (N_14877,N_10951,N_10841);
nand U14878 (N_14878,N_11445,N_9018);
and U14879 (N_14879,N_10464,N_10834);
and U14880 (N_14880,N_11881,N_11707);
and U14881 (N_14881,N_11004,N_9428);
and U14882 (N_14882,N_9220,N_9114);
nor U14883 (N_14883,N_10137,N_11074);
or U14884 (N_14884,N_11152,N_9221);
and U14885 (N_14885,N_11390,N_10564);
nand U14886 (N_14886,N_11732,N_10679);
nor U14887 (N_14887,N_11453,N_9552);
or U14888 (N_14888,N_10993,N_9022);
and U14889 (N_14889,N_11020,N_11753);
and U14890 (N_14890,N_9360,N_11724);
and U14891 (N_14891,N_10393,N_9393);
or U14892 (N_14892,N_11141,N_10788);
nor U14893 (N_14893,N_11119,N_10339);
or U14894 (N_14894,N_9828,N_10061);
nor U14895 (N_14895,N_11253,N_10720);
and U14896 (N_14896,N_9029,N_11761);
nand U14897 (N_14897,N_10156,N_10019);
nand U14898 (N_14898,N_10890,N_9772);
and U14899 (N_14899,N_10777,N_11028);
or U14900 (N_14900,N_11021,N_11936);
and U14901 (N_14901,N_10575,N_9347);
or U14902 (N_14902,N_10668,N_10572);
nand U14903 (N_14903,N_11347,N_11384);
and U14904 (N_14904,N_10392,N_10018);
nand U14905 (N_14905,N_10535,N_11750);
nand U14906 (N_14906,N_11422,N_10775);
nand U14907 (N_14907,N_9897,N_9274);
nand U14908 (N_14908,N_10545,N_10712);
or U14909 (N_14909,N_10224,N_10357);
nand U14910 (N_14910,N_10708,N_10113);
xnor U14911 (N_14911,N_9848,N_11747);
and U14912 (N_14912,N_9645,N_11619);
nor U14913 (N_14913,N_9701,N_11083);
nor U14914 (N_14914,N_11002,N_10344);
and U14915 (N_14915,N_11268,N_10613);
and U14916 (N_14916,N_11272,N_9202);
or U14917 (N_14917,N_10140,N_9539);
and U14918 (N_14918,N_11194,N_11656);
nor U14919 (N_14919,N_10180,N_11867);
nor U14920 (N_14920,N_10098,N_10615);
and U14921 (N_14921,N_11178,N_9824);
and U14922 (N_14922,N_9962,N_10279);
or U14923 (N_14923,N_9467,N_9855);
nor U14924 (N_14924,N_9280,N_9863);
or U14925 (N_14925,N_10291,N_10798);
and U14926 (N_14926,N_10613,N_11139);
nor U14927 (N_14927,N_10093,N_10134);
nand U14928 (N_14928,N_10360,N_11747);
and U14929 (N_14929,N_9674,N_11976);
or U14930 (N_14930,N_10768,N_10397);
nor U14931 (N_14931,N_11178,N_10987);
nand U14932 (N_14932,N_10004,N_11224);
and U14933 (N_14933,N_10855,N_9384);
or U14934 (N_14934,N_10915,N_11592);
nor U14935 (N_14935,N_9774,N_10126);
nand U14936 (N_14936,N_9893,N_11448);
xor U14937 (N_14937,N_9289,N_9302);
and U14938 (N_14938,N_10272,N_9079);
nor U14939 (N_14939,N_11897,N_9731);
or U14940 (N_14940,N_11403,N_9203);
and U14941 (N_14941,N_11251,N_9703);
nand U14942 (N_14942,N_10612,N_11623);
and U14943 (N_14943,N_10108,N_11822);
nand U14944 (N_14944,N_11155,N_9657);
nand U14945 (N_14945,N_10050,N_11241);
or U14946 (N_14946,N_11863,N_11652);
and U14947 (N_14947,N_10441,N_10580);
or U14948 (N_14948,N_11701,N_9589);
nand U14949 (N_14949,N_11145,N_11150);
nand U14950 (N_14950,N_9199,N_11849);
nand U14951 (N_14951,N_9996,N_11294);
nand U14952 (N_14952,N_10835,N_10180);
nor U14953 (N_14953,N_9353,N_9338);
nor U14954 (N_14954,N_9884,N_10222);
and U14955 (N_14955,N_11241,N_9183);
or U14956 (N_14956,N_9935,N_11701);
nor U14957 (N_14957,N_11911,N_11685);
and U14958 (N_14958,N_10462,N_9029);
and U14959 (N_14959,N_10109,N_9187);
nor U14960 (N_14960,N_9809,N_11414);
nor U14961 (N_14961,N_11069,N_11905);
or U14962 (N_14962,N_10006,N_11780);
and U14963 (N_14963,N_10361,N_11308);
nand U14964 (N_14964,N_9294,N_10536);
nand U14965 (N_14965,N_9048,N_11025);
nand U14966 (N_14966,N_11718,N_9131);
nand U14967 (N_14967,N_11350,N_10299);
and U14968 (N_14968,N_11630,N_10470);
or U14969 (N_14969,N_11141,N_10422);
nor U14970 (N_14970,N_11036,N_9169);
and U14971 (N_14971,N_11994,N_11453);
nand U14972 (N_14972,N_11948,N_11204);
nand U14973 (N_14973,N_11614,N_10198);
and U14974 (N_14974,N_11620,N_10185);
or U14975 (N_14975,N_11289,N_10834);
nand U14976 (N_14976,N_9467,N_11746);
nor U14977 (N_14977,N_9250,N_10178);
nor U14978 (N_14978,N_10184,N_11976);
nand U14979 (N_14979,N_11853,N_9134);
or U14980 (N_14980,N_10476,N_9539);
nand U14981 (N_14981,N_9340,N_9742);
nor U14982 (N_14982,N_11494,N_10587);
nor U14983 (N_14983,N_11972,N_11797);
and U14984 (N_14984,N_11412,N_10307);
or U14985 (N_14985,N_10492,N_11458);
or U14986 (N_14986,N_9135,N_11253);
or U14987 (N_14987,N_9193,N_11543);
xor U14988 (N_14988,N_10695,N_9021);
or U14989 (N_14989,N_11657,N_9230);
nor U14990 (N_14990,N_11498,N_11796);
or U14991 (N_14991,N_10974,N_10716);
nor U14992 (N_14992,N_11297,N_9036);
and U14993 (N_14993,N_10585,N_10267);
nand U14994 (N_14994,N_9165,N_10909);
and U14995 (N_14995,N_11352,N_11836);
and U14996 (N_14996,N_10277,N_11249);
and U14997 (N_14997,N_10449,N_10773);
nor U14998 (N_14998,N_9648,N_10145);
and U14999 (N_14999,N_9974,N_11287);
nor UO_0 (O_0,N_14658,N_14755);
nand UO_1 (O_1,N_12445,N_14621);
nor UO_2 (O_2,N_14500,N_12175);
or UO_3 (O_3,N_14217,N_14937);
nor UO_4 (O_4,N_14593,N_14764);
nor UO_5 (O_5,N_12106,N_14030);
nand UO_6 (O_6,N_12991,N_13277);
nor UO_7 (O_7,N_14638,N_13384);
and UO_8 (O_8,N_14125,N_14919);
xnor UO_9 (O_9,N_12505,N_14670);
and UO_10 (O_10,N_12479,N_14724);
nand UO_11 (O_11,N_14324,N_12005);
or UO_12 (O_12,N_12184,N_13713);
nand UO_13 (O_13,N_13619,N_14843);
xor UO_14 (O_14,N_13921,N_12302);
or UO_15 (O_15,N_14995,N_14808);
or UO_16 (O_16,N_13784,N_14429);
or UO_17 (O_17,N_14941,N_14795);
nor UO_18 (O_18,N_12921,N_14944);
or UO_19 (O_19,N_12665,N_14985);
nand UO_20 (O_20,N_14409,N_12997);
nand UO_21 (O_21,N_13284,N_14283);
or UO_22 (O_22,N_13190,N_14394);
nand UO_23 (O_23,N_13483,N_12103);
and UO_24 (O_24,N_12200,N_13388);
xnor UO_25 (O_25,N_14158,N_14149);
or UO_26 (O_26,N_12903,N_13746);
nor UO_27 (O_27,N_13426,N_12180);
or UO_28 (O_28,N_14488,N_13392);
and UO_29 (O_29,N_14981,N_14450);
nand UO_30 (O_30,N_13677,N_12700);
or UO_31 (O_31,N_12518,N_14544);
or UO_32 (O_32,N_12246,N_13592);
nand UO_33 (O_33,N_12710,N_13067);
nand UO_34 (O_34,N_14424,N_12026);
nor UO_35 (O_35,N_13706,N_12699);
nor UO_36 (O_36,N_13791,N_12872);
or UO_37 (O_37,N_12559,N_12449);
nand UO_38 (O_38,N_12863,N_12399);
or UO_39 (O_39,N_13969,N_13587);
nor UO_40 (O_40,N_12645,N_14165);
nor UO_41 (O_41,N_12545,N_12962);
or UO_42 (O_42,N_13006,N_13894);
xnor UO_43 (O_43,N_12671,N_12318);
and UO_44 (O_44,N_14470,N_12050);
xor UO_45 (O_45,N_12355,N_14066);
nor UO_46 (O_46,N_13280,N_14820);
and UO_47 (O_47,N_14940,N_14655);
or UO_48 (O_48,N_14922,N_13108);
nor UO_49 (O_49,N_14004,N_12868);
or UO_50 (O_50,N_14784,N_12380);
and UO_51 (O_51,N_14061,N_13538);
or UO_52 (O_52,N_14825,N_13232);
or UO_53 (O_53,N_14587,N_12929);
nand UO_54 (O_54,N_14953,N_14802);
xnor UO_55 (O_55,N_12810,N_14617);
or UO_56 (O_56,N_13263,N_13795);
nand UO_57 (O_57,N_12766,N_12476);
or UO_58 (O_58,N_13368,N_14659);
and UO_59 (O_59,N_12874,N_12031);
or UO_60 (O_60,N_14269,N_13663);
xnor UO_61 (O_61,N_13912,N_13193);
and UO_62 (O_62,N_12970,N_13009);
or UO_63 (O_63,N_14657,N_14276);
xor UO_64 (O_64,N_13617,N_14636);
nand UO_65 (O_65,N_12781,N_14917);
or UO_66 (O_66,N_12188,N_12178);
nor UO_67 (O_67,N_13700,N_12080);
and UO_68 (O_68,N_12247,N_14601);
and UO_69 (O_69,N_14069,N_12713);
and UO_70 (O_70,N_13983,N_13524);
nand UO_71 (O_71,N_12167,N_13900);
nor UO_72 (O_72,N_14093,N_12931);
nand UO_73 (O_73,N_13680,N_12585);
and UO_74 (O_74,N_13201,N_13371);
nand UO_75 (O_75,N_13712,N_12564);
nand UO_76 (O_76,N_13597,N_14739);
or UO_77 (O_77,N_12692,N_12331);
and UO_78 (O_78,N_13025,N_13080);
or UO_79 (O_79,N_14199,N_13157);
or UO_80 (O_80,N_12177,N_14564);
nor UO_81 (O_81,N_14455,N_13393);
nor UO_82 (O_82,N_12697,N_13906);
nand UO_83 (O_83,N_13824,N_13938);
nor UO_84 (O_84,N_12631,N_12539);
nor UO_85 (O_85,N_14014,N_12373);
and UO_86 (O_86,N_14759,N_13576);
nand UO_87 (O_87,N_13817,N_13955);
or UO_88 (O_88,N_13116,N_14619);
or UO_89 (O_89,N_14926,N_14547);
and UO_90 (O_90,N_14725,N_14958);
nor UO_91 (O_91,N_13716,N_12638);
nor UO_92 (O_92,N_13069,N_14967);
and UO_93 (O_93,N_12329,N_13585);
nor UO_94 (O_94,N_14748,N_12403);
and UO_95 (O_95,N_13419,N_14119);
nor UO_96 (O_96,N_14310,N_14452);
or UO_97 (O_97,N_13366,N_13763);
nand UO_98 (O_98,N_12846,N_14572);
nand UO_99 (O_99,N_14960,N_14205);
and UO_100 (O_100,N_14107,N_13998);
nor UO_101 (O_101,N_12947,N_12450);
or UO_102 (O_102,N_14718,N_13101);
nor UO_103 (O_103,N_14542,N_13302);
nand UO_104 (O_104,N_14242,N_12214);
or UO_105 (O_105,N_12864,N_14989);
nor UO_106 (O_106,N_12704,N_12624);
and UO_107 (O_107,N_13059,N_14528);
and UO_108 (O_108,N_14527,N_13612);
and UO_109 (O_109,N_14524,N_12590);
nand UO_110 (O_110,N_14975,N_12012);
and UO_111 (O_111,N_13406,N_12208);
and UO_112 (O_112,N_12532,N_14910);
nand UO_113 (O_113,N_14584,N_12800);
nand UO_114 (O_114,N_12058,N_13249);
nor UO_115 (O_115,N_14523,N_13654);
xor UO_116 (O_116,N_12357,N_12547);
nor UO_117 (O_117,N_14647,N_13153);
or UO_118 (O_118,N_14315,N_12609);
nand UO_119 (O_119,N_12428,N_14151);
nor UO_120 (O_120,N_13110,N_12375);
or UO_121 (O_121,N_12642,N_13724);
or UO_122 (O_122,N_14024,N_12739);
and UO_123 (O_123,N_12988,N_13409);
and UO_124 (O_124,N_14566,N_14537);
and UO_125 (O_125,N_13527,N_12897);
nand UO_126 (O_126,N_12360,N_12848);
and UO_127 (O_127,N_13287,N_13556);
and UO_128 (O_128,N_12575,N_14189);
or UO_129 (O_129,N_13016,N_12880);
nor UO_130 (O_130,N_13273,N_13567);
nor UO_131 (O_131,N_14682,N_14195);
nor UO_132 (O_132,N_13013,N_13057);
and UO_133 (O_133,N_14899,N_14738);
or UO_134 (O_134,N_13467,N_14824);
nor UO_135 (O_135,N_12010,N_12675);
nand UO_136 (O_136,N_13689,N_14309);
nor UO_137 (O_137,N_14322,N_12322);
and UO_138 (O_138,N_13181,N_13865);
and UO_139 (O_139,N_14717,N_13781);
nand UO_140 (O_140,N_14698,N_12119);
nand UO_141 (O_141,N_12827,N_12224);
nor UO_142 (O_142,N_14260,N_13365);
or UO_143 (O_143,N_14270,N_13687);
nand UO_144 (O_144,N_12153,N_14951);
or UO_145 (O_145,N_12840,N_14391);
nor UO_146 (O_146,N_14762,N_12557);
nand UO_147 (O_147,N_14290,N_12716);
and UO_148 (O_148,N_12714,N_13884);
nor UO_149 (O_149,N_13186,N_12459);
or UO_150 (O_150,N_14306,N_13997);
nand UO_151 (O_151,N_12035,N_12682);
nand UO_152 (O_152,N_14763,N_12552);
nand UO_153 (O_153,N_14463,N_13091);
and UO_154 (O_154,N_14422,N_13143);
or UO_155 (O_155,N_12796,N_13604);
nor UO_156 (O_156,N_14461,N_13326);
nor UO_157 (O_157,N_12218,N_12454);
or UO_158 (O_158,N_14861,N_12820);
nor UO_159 (O_159,N_13550,N_12952);
nor UO_160 (O_160,N_12297,N_12905);
or UO_161 (O_161,N_14479,N_14635);
nor UO_162 (O_162,N_14325,N_12724);
or UO_163 (O_163,N_13657,N_13098);
nor UO_164 (O_164,N_14374,N_12548);
nand UO_165 (O_165,N_13065,N_14673);
or UO_166 (O_166,N_13564,N_12812);
nor UO_167 (O_167,N_14174,N_12460);
xnor UO_168 (O_168,N_14384,N_12654);
nand UO_169 (O_169,N_14320,N_14774);
or UO_170 (O_170,N_13047,N_12625);
nand UO_171 (O_171,N_13103,N_13942);
xor UO_172 (O_172,N_14513,N_12251);
and UO_173 (O_173,N_14331,N_13507);
or UO_174 (O_174,N_12081,N_13805);
or UO_175 (O_175,N_12274,N_13624);
or UO_176 (O_176,N_14776,N_13199);
nand UO_177 (O_177,N_14538,N_12029);
and UO_178 (O_178,N_13140,N_12299);
and UO_179 (O_179,N_12345,N_13215);
nand UO_180 (O_180,N_14058,N_13329);
or UO_181 (O_181,N_13749,N_13463);
nor UO_182 (O_182,N_12105,N_13794);
nor UO_183 (O_183,N_14109,N_13470);
or UO_184 (O_184,N_12752,N_12022);
or UO_185 (O_185,N_12678,N_12294);
nor UO_186 (O_186,N_13875,N_13328);
or UO_187 (O_187,N_12183,N_12668);
and UO_188 (O_188,N_12364,N_12596);
and UO_189 (O_189,N_14811,N_13142);
or UO_190 (O_190,N_12254,N_13734);
or UO_191 (O_191,N_12530,N_14906);
and UO_192 (O_192,N_12501,N_13165);
nor UO_193 (O_193,N_14730,N_14801);
nand UO_194 (O_194,N_14462,N_12225);
nand UO_195 (O_195,N_12475,N_12870);
nand UO_196 (O_196,N_14531,N_13346);
nor UO_197 (O_197,N_12976,N_14023);
nor UO_198 (O_198,N_13899,N_12579);
or UO_199 (O_199,N_12451,N_12803);
and UO_200 (O_200,N_14842,N_13078);
and UO_201 (O_201,N_13084,N_12664);
nor UO_202 (O_202,N_14339,N_13980);
and UO_203 (O_203,N_13603,N_13373);
nor UO_204 (O_204,N_12157,N_14075);
xor UO_205 (O_205,N_14247,N_14857);
nand UO_206 (O_206,N_12582,N_14907);
or UO_207 (O_207,N_12356,N_14240);
nand UO_208 (O_208,N_12835,N_14336);
xor UO_209 (O_209,N_12444,N_13885);
nand UO_210 (O_210,N_12107,N_14577);
and UO_211 (O_211,N_14961,N_14299);
xnor UO_212 (O_212,N_13648,N_13396);
and UO_213 (O_213,N_14929,N_13382);
nand UO_214 (O_214,N_13656,N_12317);
nor UO_215 (O_215,N_12577,N_13231);
nand UO_216 (O_216,N_12676,N_13639);
or UO_217 (O_217,N_12956,N_13503);
or UO_218 (O_218,N_12269,N_14752);
or UO_219 (O_219,N_13695,N_12199);
nand UO_220 (O_220,N_13905,N_14472);
nand UO_221 (O_221,N_12712,N_12937);
xor UO_222 (O_222,N_14445,N_14925);
or UO_223 (O_223,N_13693,N_14948);
or UO_224 (O_224,N_12448,N_12101);
nor UO_225 (O_225,N_14859,N_14273);
or UO_226 (O_226,N_12967,N_12759);
nand UO_227 (O_227,N_14311,N_12938);
nand UO_228 (O_228,N_12071,N_12566);
nor UO_229 (O_229,N_12737,N_13423);
or UO_230 (O_230,N_14565,N_12011);
or UO_231 (O_231,N_13094,N_12984);
nand UO_232 (O_232,N_13130,N_14142);
and UO_233 (O_233,N_12788,N_12162);
nand UO_234 (O_234,N_14794,N_13523);
nand UO_235 (O_235,N_12535,N_14560);
and UO_236 (O_236,N_12075,N_12472);
or UO_237 (O_237,N_14683,N_13278);
xor UO_238 (O_238,N_12248,N_13721);
and UO_239 (O_239,N_14049,N_12122);
or UO_240 (O_240,N_13407,N_13888);
and UO_241 (O_241,N_14459,N_13886);
or UO_242 (O_242,N_14353,N_12068);
nand UO_243 (O_243,N_12016,N_13126);
or UO_244 (O_244,N_14979,N_13953);
nand UO_245 (O_245,N_12206,N_13681);
or UO_246 (O_246,N_14671,N_14515);
nand UO_247 (O_247,N_14243,N_12437);
nor UO_248 (O_248,N_12209,N_14915);
nand UO_249 (O_249,N_14813,N_14732);
and UO_250 (O_250,N_14444,N_13553);
and UO_251 (O_251,N_13798,N_12365);
nor UO_252 (O_252,N_12057,N_14340);
nor UO_253 (O_253,N_12088,N_14206);
and UO_254 (O_254,N_13370,N_13827);
and UO_255 (O_255,N_12132,N_12721);
nor UO_256 (O_256,N_14624,N_13480);
nor UO_257 (O_257,N_13799,N_14846);
nor UO_258 (O_258,N_13858,N_12387);
and UO_259 (O_259,N_12021,N_13819);
and UO_260 (O_260,N_13580,N_12499);
and UO_261 (O_261,N_12095,N_13772);
and UO_262 (O_262,N_14355,N_14144);
and UO_263 (O_263,N_14817,N_13387);
nand UO_264 (O_264,N_14465,N_13883);
and UO_265 (O_265,N_12287,N_13860);
or UO_266 (O_266,N_14576,N_12939);
or UO_267 (O_267,N_14746,N_13548);
nor UO_268 (O_268,N_13004,N_13210);
or UO_269 (O_269,N_12882,N_12228);
nor UO_270 (O_270,N_12417,N_13560);
and UO_271 (O_271,N_14263,N_14152);
and UO_272 (O_272,N_13209,N_13769);
nand UO_273 (O_273,N_13119,N_14053);
or UO_274 (O_274,N_13670,N_13092);
or UO_275 (O_275,N_12491,N_14114);
nand UO_276 (O_276,N_13402,N_14092);
and UO_277 (O_277,N_13737,N_13031);
nand UO_278 (O_278,N_12250,N_12385);
xor UO_279 (O_279,N_14333,N_13727);
xnor UO_280 (O_280,N_14427,N_14248);
and UO_281 (O_281,N_12703,N_12478);
or UO_282 (O_282,N_14010,N_12104);
nor UO_283 (O_283,N_12310,N_12647);
nor UO_284 (O_284,N_12755,N_12221);
nand UO_285 (O_285,N_13571,N_13849);
nand UO_286 (O_286,N_14605,N_13973);
nand UO_287 (O_287,N_14830,N_13633);
nor UO_288 (O_288,N_13189,N_13195);
nand UO_289 (O_289,N_12126,N_12576);
xor UO_290 (O_290,N_13590,N_14652);
nor UO_291 (O_291,N_14514,N_13982);
or UO_292 (O_292,N_13413,N_14245);
xor UO_293 (O_293,N_12130,N_13701);
and UO_294 (O_294,N_14699,N_14687);
nor UO_295 (O_295,N_13511,N_14541);
nor UO_296 (O_296,N_12886,N_13667);
or UO_297 (O_297,N_14507,N_14905);
and UO_298 (O_298,N_13637,N_12771);
nor UO_299 (O_299,N_12889,N_14731);
nor UO_300 (O_300,N_12037,N_12528);
nand UO_301 (O_301,N_14088,N_14653);
nor UO_302 (O_302,N_12293,N_14983);
or UO_303 (O_303,N_12615,N_13135);
nor UO_304 (O_304,N_12488,N_13933);
and UO_305 (O_305,N_14483,N_13631);
and UO_306 (O_306,N_13653,N_12972);
nor UO_307 (O_307,N_14319,N_14438);
nand UO_308 (O_308,N_14163,N_13743);
or UO_309 (O_309,N_13066,N_13703);
nand UO_310 (O_310,N_14161,N_13859);
or UO_311 (O_311,N_14393,N_12600);
or UO_312 (O_312,N_13197,N_12168);
nand UO_313 (O_313,N_13505,N_14870);
and UO_314 (O_314,N_12594,N_12416);
nand UO_315 (O_315,N_14406,N_13323);
nor UO_316 (O_316,N_14032,N_13522);
nor UO_317 (O_317,N_13786,N_13208);
and UO_318 (O_318,N_14184,N_12603);
nand UO_319 (O_319,N_13918,N_14225);
nand UO_320 (O_320,N_14043,N_13344);
nand UO_321 (O_321,N_12843,N_14691);
nand UO_322 (O_322,N_12698,N_13015);
or UO_323 (O_323,N_13996,N_14875);
or UO_324 (O_324,N_12896,N_12339);
nand UO_325 (O_325,N_14701,N_13729);
nor UO_326 (O_326,N_12866,N_12914);
nand UO_327 (O_327,N_12166,N_14745);
and UO_328 (O_328,N_14993,N_12974);
and UO_329 (O_329,N_13150,N_13125);
nand UO_330 (O_330,N_12342,N_14832);
or UO_331 (O_331,N_14679,N_14686);
nor UO_332 (O_332,N_14267,N_12957);
and UO_333 (O_333,N_13965,N_12808);
and UO_334 (O_334,N_13172,N_14840);
and UO_335 (O_335,N_14681,N_13305);
or UO_336 (O_336,N_13478,N_13175);
or UO_337 (O_337,N_14982,N_13717);
nor UO_338 (O_338,N_14430,N_13479);
nand UO_339 (O_339,N_12705,N_13532);
or UO_340 (O_340,N_13704,N_13026);
nand UO_341 (O_341,N_14105,N_12439);
nand UO_342 (O_342,N_13082,N_14611);
nand UO_343 (O_343,N_12734,N_14063);
nand UO_344 (O_344,N_13216,N_14005);
or UO_345 (O_345,N_12066,N_12536);
xor UO_346 (O_346,N_13830,N_12522);
nor UO_347 (O_347,N_13484,N_12542);
or UO_348 (O_348,N_14592,N_14867);
and UO_349 (O_349,N_14816,N_13147);
nand UO_350 (O_350,N_12640,N_14921);
nand UO_351 (O_351,N_12941,N_14853);
or UO_352 (O_352,N_14847,N_14591);
nand UO_353 (O_353,N_13447,N_12999);
xnor UO_354 (O_354,N_13855,N_14366);
nor UO_355 (O_355,N_14569,N_13124);
or UO_356 (O_356,N_13410,N_13512);
nor UO_357 (O_357,N_13003,N_12862);
nand UO_358 (O_358,N_13954,N_13991);
nand UO_359 (O_359,N_13614,N_12573);
nand UO_360 (O_360,N_13088,N_14392);
xor UO_361 (O_361,N_13776,N_12389);
or UO_362 (O_362,N_12509,N_12053);
and UO_363 (O_363,N_12813,N_13628);
xnor UO_364 (O_364,N_12276,N_13506);
or UO_365 (O_365,N_13389,N_14380);
nand UO_366 (O_366,N_13351,N_13876);
nor UO_367 (O_367,N_12159,N_12691);
or UO_368 (O_368,N_13474,N_13137);
nand UO_369 (O_369,N_13978,N_14097);
and UO_370 (O_370,N_13164,N_13441);
nand UO_371 (O_371,N_13043,N_12869);
nor UO_372 (O_372,N_12500,N_14590);
nand UO_373 (O_373,N_13747,N_14705);
nand UO_374 (O_374,N_14913,N_13375);
nand UO_375 (O_375,N_14607,N_12404);
and UO_376 (O_376,N_13029,N_12772);
nand UO_377 (O_377,N_13972,N_14046);
or UO_378 (O_378,N_14216,N_13350);
nand UO_379 (O_379,N_12811,N_13472);
and UO_380 (O_380,N_13090,N_12424);
nand UO_381 (O_381,N_13087,N_12282);
nor UO_382 (O_382,N_14492,N_12003);
and UO_383 (O_383,N_14302,N_14227);
nand UO_384 (O_384,N_14132,N_12392);
or UO_385 (O_385,N_14526,N_14889);
nor UO_386 (O_386,N_14399,N_13490);
and UO_387 (O_387,N_12020,N_14839);
and UO_388 (O_388,N_13010,N_12261);
or UO_389 (O_389,N_13764,N_14091);
nor UO_390 (O_390,N_13602,N_13230);
nand UO_391 (O_391,N_13741,N_14077);
nor UO_392 (O_392,N_12793,N_13736);
or UO_393 (O_393,N_13107,N_13549);
or UO_394 (O_394,N_14407,N_13591);
nand UO_395 (O_395,N_14597,N_14702);
xnor UO_396 (O_396,N_14595,N_12278);
nand UO_397 (O_397,N_13432,N_14955);
nor UO_398 (O_398,N_13673,N_13239);
and UO_399 (O_399,N_13863,N_12708);
nand UO_400 (O_400,N_14895,N_12857);
and UO_401 (O_401,N_13054,N_14615);
nor UO_402 (O_402,N_13028,N_14990);
nand UO_403 (O_403,N_13404,N_12163);
nor UO_404 (O_404,N_13049,N_14187);
or UO_405 (O_405,N_13438,N_13417);
or UO_406 (O_406,N_12047,N_14494);
and UO_407 (O_407,N_12015,N_12635);
nand UO_408 (O_408,N_14318,N_13770);
nand UO_409 (O_409,N_14622,N_12723);
and UO_410 (O_410,N_14898,N_12402);
and UO_411 (O_411,N_13577,N_14965);
nand UO_412 (O_412,N_12182,N_12661);
nand UO_413 (O_413,N_12883,N_12867);
or UO_414 (O_414,N_12133,N_13168);
or UO_415 (O_415,N_12900,N_13102);
and UO_416 (O_416,N_14610,N_13517);
and UO_417 (O_417,N_14644,N_12856);
or UO_418 (O_418,N_13609,N_14957);
nor UO_419 (O_419,N_13475,N_14706);
nand UO_420 (O_420,N_13042,N_13309);
nand UO_421 (O_421,N_13286,N_13738);
nand UO_422 (O_422,N_14946,N_13086);
nor UO_423 (O_423,N_12517,N_12617);
or UO_424 (O_424,N_14214,N_12038);
or UO_425 (O_425,N_14865,N_14800);
nor UO_426 (O_426,N_14327,N_14110);
xor UO_427 (O_427,N_12672,N_12359);
or UO_428 (O_428,N_13903,N_14274);
nand UO_429 (O_429,N_14819,N_12599);
or UO_430 (O_430,N_12158,N_12492);
and UO_431 (O_431,N_12111,N_12973);
and UO_432 (O_432,N_13191,N_12610);
nand UO_433 (O_433,N_12348,N_13321);
or UO_434 (O_434,N_14722,N_14101);
and UO_435 (O_435,N_12124,N_13570);
or UO_436 (O_436,N_13892,N_12052);
nor UO_437 (O_437,N_14704,N_13630);
or UO_438 (O_438,N_13064,N_13757);
or UO_439 (O_439,N_13452,N_14838);
nor UO_440 (O_440,N_14791,N_13061);
or UO_441 (O_441,N_12628,N_13154);
and UO_442 (O_442,N_13684,N_12039);
xnor UO_443 (O_443,N_12484,N_14372);
and UO_444 (O_444,N_13844,N_12006);
nand UO_445 (O_445,N_13381,N_13222);
or UO_446 (O_446,N_14467,N_12595);
nor UO_447 (O_447,N_12927,N_12906);
and UO_448 (O_448,N_14268,N_14435);
nor UO_449 (O_449,N_13039,N_13261);
nor UO_450 (O_450,N_12190,N_13977);
or UO_451 (O_451,N_13641,N_13235);
or UO_452 (O_452,N_14551,N_14943);
nor UO_453 (O_453,N_12490,N_14288);
or UO_454 (O_454,N_14798,N_14650);
or UO_455 (O_455,N_12236,N_12873);
and UO_456 (O_456,N_12720,N_12887);
nor UO_457 (O_457,N_13937,N_14818);
nor UO_458 (O_458,N_13144,N_13052);
nor UO_459 (O_459,N_14386,N_12493);
or UO_460 (O_460,N_13601,N_13750);
or UO_461 (O_461,N_13457,N_14096);
and UO_462 (O_462,N_14735,N_12780);
nand UO_463 (O_463,N_13500,N_14241);
or UO_464 (O_464,N_14630,N_13113);
nor UO_465 (O_465,N_13089,N_13588);
or UO_466 (O_466,N_14684,N_12920);
and UO_467 (O_467,N_14136,N_13995);
xnor UO_468 (O_468,N_14896,N_12636);
nor UO_469 (O_469,N_13584,N_12036);
nor UO_470 (O_470,N_12243,N_12259);
nand UO_471 (O_471,N_14255,N_12707);
or UO_472 (O_472,N_12639,N_13696);
or UO_473 (O_473,N_13740,N_13493);
or UO_474 (O_474,N_12966,N_12044);
nor UO_475 (O_475,N_13642,N_13820);
or UO_476 (O_476,N_13811,N_12382);
xnor UO_477 (O_477,N_14675,N_12529);
and UO_478 (O_478,N_14370,N_14296);
or UO_479 (O_479,N_14489,N_12467);
nand UO_480 (O_480,N_14747,N_14138);
and UO_481 (O_481,N_14720,N_14002);
and UO_482 (O_482,N_14412,N_12618);
and UO_483 (O_483,N_12891,N_14656);
and UO_484 (O_484,N_12198,N_13632);
and UO_485 (O_485,N_12477,N_12831);
or UO_486 (O_486,N_14540,N_14198);
nor UO_487 (O_487,N_12497,N_14127);
or UO_488 (O_488,N_13223,N_14356);
nand UO_489 (O_489,N_13034,N_12288);
or UO_490 (O_490,N_14281,N_14191);
or UO_491 (O_491,N_12400,N_12964);
nand UO_492 (O_492,N_13666,N_12260);
and UO_493 (O_493,N_12589,N_13554);
and UO_494 (O_494,N_12148,N_13659);
or UO_495 (O_495,N_12060,N_12289);
and UO_496 (O_496,N_12787,N_12346);
xnor UO_497 (O_497,N_12281,N_12955);
nor UO_498 (O_498,N_14293,N_12146);
nor UO_499 (O_499,N_14916,N_12061);
nand UO_500 (O_500,N_12344,N_12515);
nand UO_501 (O_501,N_12013,N_13782);
xor UO_502 (O_502,N_14261,N_14928);
nand UO_503 (O_503,N_13122,N_13136);
and UO_504 (O_504,N_14397,N_14244);
and UO_505 (O_505,N_14642,N_14040);
or UO_506 (O_506,N_13182,N_13562);
or UO_507 (O_507,N_13957,N_14716);
nand UO_508 (O_508,N_14822,N_14432);
nand UO_509 (O_509,N_14456,N_14775);
nand UO_510 (O_510,N_12009,N_13672);
and UO_511 (O_511,N_13145,N_14154);
and UO_512 (O_512,N_14060,N_14341);
or UO_513 (O_513,N_14550,N_14246);
or UO_514 (O_514,N_12568,N_13926);
nor UO_515 (O_515,N_14179,N_12455);
or UO_516 (O_516,N_12998,N_13048);
nand UO_517 (O_517,N_14282,N_13459);
nor UO_518 (O_518,N_13099,N_13299);
or UO_519 (O_519,N_13282,N_14606);
nor UO_520 (O_520,N_14911,N_14208);
or UO_521 (O_521,N_14219,N_12643);
nand UO_522 (O_522,N_14121,N_13678);
and UO_523 (O_523,N_13132,N_13170);
nor UO_524 (O_524,N_13536,N_14938);
or UO_525 (O_525,N_14103,N_14086);
or UO_526 (O_526,N_12627,N_13715);
and UO_527 (O_527,N_14475,N_13898);
and UO_528 (O_528,N_13330,N_12197);
and UO_529 (O_529,N_14850,N_13355);
nand UO_530 (O_530,N_12681,N_14977);
nor UO_531 (O_531,N_12987,N_13391);
nor UO_532 (O_532,N_14883,N_13595);
and UO_533 (O_533,N_13336,N_14554);
nor UO_534 (O_534,N_12853,N_13519);
nand UO_535 (O_535,N_14351,N_12408);
nand UO_536 (O_536,N_14070,N_13403);
nor UO_537 (O_537,N_13491,N_13271);
nand UO_538 (O_538,N_14771,N_14947);
and UO_539 (O_539,N_12561,N_14614);
and UO_540 (O_540,N_13963,N_12014);
nor UO_541 (O_541,N_13121,N_13932);
nor UO_542 (O_542,N_13340,N_12213);
nand UO_543 (O_543,N_13758,N_13839);
nand UO_544 (O_544,N_12504,N_14841);
and UO_545 (O_545,N_13018,N_12087);
nand UO_546 (O_546,N_13433,N_12527);
and UO_547 (O_547,N_13437,N_13509);
nand UO_548 (O_548,N_12651,N_14466);
nand UO_549 (O_549,N_14923,N_13748);
nand UO_550 (O_550,N_14417,N_13471);
nor UO_551 (O_551,N_12894,N_12711);
or UO_552 (O_552,N_12034,N_13497);
or UO_553 (O_553,N_14469,N_13427);
nor UO_554 (O_554,N_13458,N_12423);
nand UO_555 (O_555,N_12660,N_14968);
nor UO_556 (O_556,N_12930,N_13476);
or UO_557 (O_557,N_12171,N_14891);
or UO_558 (O_558,N_13944,N_14448);
and UO_559 (O_559,N_14885,N_13386);
nor UO_560 (O_560,N_14343,N_13702);
and UO_561 (O_561,N_12435,N_12608);
and UO_562 (O_562,N_12211,N_14068);
nor UO_563 (O_563,N_14286,N_13036);
or UO_564 (O_564,N_12376,N_14126);
nor UO_565 (O_565,N_13369,N_12065);
nand UO_566 (O_566,N_12237,N_12333);
nand UO_567 (O_567,N_14643,N_12495);
nor UO_568 (O_568,N_14153,N_14007);
nor UO_569 (O_569,N_14773,N_13600);
and UO_570 (O_570,N_12558,N_13565);
or UO_571 (O_571,N_12657,N_13032);
and UO_572 (O_572,N_14118,N_13339);
nor UO_573 (O_573,N_14056,N_14188);
nor UO_574 (O_574,N_14305,N_13211);
nand UO_575 (O_575,N_12471,N_12358);
and UO_576 (O_576,N_14689,N_14342);
nand UO_577 (O_577,N_14519,N_13940);
nand UO_578 (O_578,N_12899,N_13650);
and UO_579 (O_579,N_14420,N_12546);
nor UO_580 (O_580,N_14212,N_13989);
and UO_581 (O_581,N_13862,N_12350);
or UO_582 (O_582,N_13252,N_12238);
nand UO_583 (O_583,N_13074,N_14277);
nand UO_584 (O_584,N_14809,N_13907);
or UO_585 (O_585,N_13528,N_13011);
nor UO_586 (O_586,N_12580,N_13146);
nand UO_587 (O_587,N_12425,N_12170);
nor UO_588 (O_588,N_14416,N_12684);
and UO_589 (O_589,N_14347,N_12377);
nor UO_590 (O_590,N_12085,N_14980);
nor UO_591 (O_591,N_13573,N_12954);
and UO_592 (O_592,N_13735,N_13176);
and UO_593 (O_593,N_13364,N_14192);
nor UO_594 (O_594,N_14616,N_14396);
or UO_595 (O_595,N_12936,N_14141);
and UO_596 (O_596,N_12301,N_12353);
or UO_597 (O_597,N_13106,N_13686);
nand UO_598 (O_598,N_13334,N_12283);
nand UO_599 (O_599,N_13345,N_13935);
nand UO_600 (O_600,N_14304,N_14934);
and UO_601 (O_601,N_12195,N_14148);
and UO_602 (O_602,N_13171,N_12152);
nor UO_603 (O_603,N_14258,N_14067);
or UO_604 (O_604,N_12055,N_12028);
or UO_605 (O_605,N_12741,N_13643);
and UO_606 (O_606,N_14927,N_14139);
or UO_607 (O_607,N_13975,N_14019);
nand UO_608 (O_608,N_14662,N_13936);
nor UO_609 (O_609,N_13796,N_13605);
or UO_610 (O_610,N_14057,N_12801);
nor UO_611 (O_611,N_12176,N_13925);
nor UO_612 (O_612,N_12196,N_12943);
and UO_613 (O_613,N_13941,N_14522);
or UO_614 (O_614,N_14089,N_13473);
nor UO_615 (O_615,N_12481,N_13581);
nand UO_616 (O_616,N_14122,N_13422);
nand UO_617 (O_617,N_14029,N_14963);
nor UO_618 (O_618,N_13444,N_13275);
and UO_619 (O_619,N_14987,N_14612);
or UO_620 (O_620,N_13158,N_13138);
nor UO_621 (O_621,N_14012,N_13268);
and UO_622 (O_622,N_13535,N_12770);
xor UO_623 (O_623,N_14271,N_12928);
nor UO_624 (O_624,N_13376,N_13342);
nor UO_625 (O_625,N_14711,N_12436);
nand UO_626 (O_626,N_14690,N_13812);
nor UO_627 (O_627,N_12942,N_12128);
nor UO_628 (O_628,N_12655,N_12173);
nor UO_629 (O_629,N_14741,N_14786);
nor UO_630 (O_630,N_12090,N_13917);
and UO_631 (O_631,N_12751,N_14562);
and UO_632 (O_632,N_14834,N_14186);
nand UO_633 (O_633,N_12908,N_14868);
nor UO_634 (O_634,N_13674,N_12791);
or UO_635 (O_635,N_13994,N_12732);
and UO_636 (O_636,N_14753,N_12731);
nand UO_637 (O_637,N_13919,N_14641);
nor UO_638 (O_638,N_12798,N_13797);
nand UO_639 (O_639,N_13076,N_13555);
or UO_640 (O_640,N_12749,N_13183);
xnor UO_641 (O_641,N_14543,N_12979);
and UO_642 (O_642,N_12611,N_12859);
nor UO_643 (O_643,N_12706,N_13766);
nor UO_644 (O_644,N_13984,N_12918);
nor UO_645 (O_645,N_12165,N_12968);
and UO_646 (O_646,N_12907,N_12279);
or UO_647 (O_647,N_14301,N_12325);
and UO_648 (O_648,N_12685,N_14600);
and UO_649 (O_649,N_12563,N_13526);
or UO_650 (O_650,N_12406,N_12457);
or UO_651 (O_651,N_13636,N_13882);
nor UO_652 (O_652,N_12855,N_12924);
xor UO_653 (O_653,N_12877,N_12830);
nor UO_654 (O_654,N_13070,N_12909);
nor UO_655 (O_655,N_13360,N_12363);
or UO_656 (O_656,N_12833,N_12890);
nor UO_657 (O_657,N_13151,N_13062);
xor UO_658 (O_658,N_12337,N_13050);
nand UO_659 (O_659,N_12089,N_12696);
nand UO_660 (O_660,N_13448,N_12270);
or UO_661 (O_661,N_12520,N_14805);
nor UO_662 (O_662,N_13699,N_13658);
nand UO_663 (O_663,N_13871,N_14827);
xor UO_664 (O_664,N_12229,N_12072);
nand UO_665 (O_665,N_14539,N_12470);
and UO_666 (O_666,N_13081,N_13651);
and UO_667 (O_667,N_14888,N_12135);
and UO_668 (O_668,N_12432,N_14833);
nand UO_669 (O_669,N_12077,N_12161);
or UO_670 (O_670,N_12002,N_12442);
and UO_671 (O_671,N_13492,N_12981);
or UO_672 (O_672,N_14509,N_13806);
and UO_673 (O_673,N_14874,N_13325);
and UO_674 (O_674,N_13267,N_14365);
and UO_675 (O_675,N_13253,N_12338);
nand UO_676 (O_676,N_14434,N_13017);
and UO_677 (O_677,N_12485,N_13495);
or UO_678 (O_678,N_13468,N_13256);
or UO_679 (O_679,N_12683,N_14108);
nor UO_680 (O_680,N_13896,N_13691);
or UO_681 (O_681,N_13792,N_13270);
and UO_682 (O_682,N_12975,N_12572);
nand UO_683 (O_683,N_13787,N_12030);
nor UO_684 (O_684,N_13005,N_12824);
and UO_685 (O_685,N_12919,N_13359);
nand UO_686 (O_686,N_12024,N_14224);
nor UO_687 (O_687,N_14956,N_12290);
nor UO_688 (O_688,N_13349,N_14876);
nand UO_689 (O_689,N_12239,N_13971);
nor UO_690 (O_690,N_13529,N_13753);
nand UO_691 (O_691,N_12842,N_12368);
and UO_692 (O_692,N_13290,N_12666);
nor UO_693 (O_693,N_13213,N_13767);
nor UO_694 (O_694,N_12817,N_12145);
and UO_695 (O_695,N_13869,N_12727);
or UO_696 (O_696,N_13055,N_13022);
and UO_697 (O_697,N_12017,N_12421);
nor UO_698 (O_698,N_13450,N_12784);
nor UO_699 (O_699,N_13023,N_13778);
nor UO_700 (O_700,N_14408,N_14660);
and UO_701 (O_701,N_12123,N_12284);
or UO_702 (O_702,N_14897,N_12438);
nand UO_703 (O_703,N_14073,N_14473);
nand UO_704 (O_704,N_14081,N_13238);
nor UO_705 (O_705,N_12834,N_13730);
nand UO_706 (O_706,N_14454,N_14272);
or UO_707 (O_707,N_13890,N_14939);
nor UO_708 (O_708,N_13815,N_14453);
nand UO_709 (O_709,N_13915,N_14112);
nand UO_710 (O_710,N_13697,N_14193);
nor UO_711 (O_711,N_14440,N_12738);
nor UO_712 (O_712,N_12839,N_12729);
nor UO_713 (O_713,N_12067,N_13870);
or UO_714 (O_714,N_14632,N_13714);
nand UO_715 (O_715,N_12950,N_13131);
nor UO_716 (O_716,N_14782,N_14485);
nor UO_717 (O_717,N_14377,N_12386);
nor UO_718 (O_718,N_12965,N_12393);
nor UO_719 (O_719,N_12832,N_14949);
nand UO_720 (O_720,N_12483,N_12507);
or UO_721 (O_721,N_12776,N_12388);
nor UO_722 (O_722,N_13461,N_12895);
nand UO_723 (O_723,N_14729,N_13218);
nor UO_724 (O_724,N_14082,N_14215);
nand UO_725 (O_725,N_13754,N_13338);
nand UO_726 (O_726,N_13675,N_13117);
nor UO_727 (O_727,N_12686,N_14035);
nor UO_728 (O_728,N_12959,N_13308);
or UO_729 (O_729,N_13993,N_14678);
nor UO_730 (O_730,N_12414,N_14556);
and UO_731 (O_731,N_12326,N_13579);
nand UO_732 (O_732,N_14676,N_12321);
or UO_733 (O_733,N_12726,N_12556);
xor UO_734 (O_734,N_13431,N_13887);
and UO_735 (O_735,N_13514,N_14984);
nand UO_736 (O_736,N_13594,N_13421);
nor UO_737 (O_737,N_13303,N_13405);
and UO_738 (O_738,N_14147,N_12315);
nand UO_739 (O_739,N_13347,N_12825);
nand UO_740 (O_740,N_12335,N_13044);
and UO_741 (O_741,N_12687,N_13037);
or UO_742 (O_742,N_12000,N_14677);
xnor UO_743 (O_743,N_14265,N_13035);
nor UO_744 (O_744,N_14017,N_13206);
nand UO_745 (O_745,N_12523,N_13283);
nand UO_746 (O_746,N_13294,N_12786);
and UO_747 (O_747,N_12023,N_12136);
nand UO_748 (O_748,N_14221,N_13343);
xnor UO_749 (O_749,N_14009,N_14497);
or UO_750 (O_750,N_14229,N_14249);
or UO_751 (O_751,N_12223,N_14713);
nand UO_752 (O_752,N_14792,N_13606);
and UO_753 (O_753,N_12292,N_14508);
nand UO_754 (O_754,N_12383,N_12468);
and UO_755 (O_755,N_12027,N_12985);
nand UO_756 (O_756,N_14387,N_13518);
or UO_757 (O_757,N_12049,N_13014);
and UO_758 (O_758,N_14835,N_12554);
or UO_759 (O_759,N_12094,N_13566);
or UO_760 (O_760,N_14379,N_12074);
or UO_761 (O_761,N_13353,N_13306);
or UO_762 (O_762,N_12045,N_14001);
nor UO_763 (O_763,N_14969,N_14736);
nand UO_764 (O_764,N_12805,N_14168);
or UO_765 (O_765,N_12513,N_14436);
nand UO_766 (O_766,N_12220,N_14966);
or UO_767 (O_767,N_14223,N_12019);
and UO_768 (O_768,N_12252,N_13557);
and UO_769 (O_769,N_13482,N_12605);
nand UO_770 (O_770,N_14598,N_13615);
and UO_771 (O_771,N_12951,N_12754);
or UO_772 (O_772,N_14903,N_13962);
or UO_773 (O_773,N_13646,N_13719);
nor UO_774 (O_774,N_14772,N_14442);
nor UO_775 (O_775,N_14680,N_12836);
or UO_776 (O_776,N_12945,N_13310);
nand UO_777 (O_777,N_14447,N_14516);
or UO_778 (O_778,N_13012,N_13889);
and UO_779 (O_779,N_14649,N_14648);
nand UO_780 (O_780,N_13083,N_14176);
nand UO_781 (O_781,N_13731,N_14257);
nand UO_782 (O_782,N_12349,N_14395);
and UO_783 (O_783,N_12569,N_14696);
and UO_784 (O_784,N_13676,N_12648);
and UO_785 (O_785,N_12463,N_12792);
nor UO_786 (O_786,N_14177,N_14262);
nor UO_787 (O_787,N_13079,N_14628);
nor UO_788 (O_788,N_14918,N_14733);
nor UO_789 (O_789,N_13367,N_12783);
or UO_790 (O_790,N_13967,N_13992);
nor UO_791 (O_791,N_14880,N_12742);
nor UO_792 (O_792,N_12064,N_12418);
or UO_793 (O_793,N_14549,N_12240);
and UO_794 (O_794,N_14256,N_14031);
nand UO_795 (O_795,N_13755,N_14439);
and UO_796 (O_796,N_13530,N_14423);
or UO_797 (O_797,N_12487,N_14042);
or UO_798 (O_798,N_12125,N_12797);
and UO_799 (O_799,N_14345,N_13775);
and UO_800 (O_800,N_13412,N_14555);
and UO_801 (O_801,N_13466,N_14505);
nor UO_802 (O_802,N_14700,N_13295);
and UO_803 (O_803,N_12391,N_12818);
or UO_804 (O_804,N_12860,N_13593);
nand UO_805 (O_805,N_12079,N_12447);
or UO_806 (O_806,N_13563,N_13809);
and UO_807 (O_807,N_12804,N_12662);
nand UO_808 (O_808,N_12147,N_13943);
or UO_809 (O_809,N_13007,N_12412);
nand UO_810 (O_810,N_14728,N_14140);
nand UO_811 (O_811,N_12295,N_13728);
or UO_812 (O_812,N_12156,N_12384);
nand UO_813 (O_813,N_13828,N_13834);
nor UO_814 (O_814,N_14912,N_14368);
and UO_815 (O_815,N_13260,N_13552);
and UO_816 (O_816,N_12745,N_13589);
nor UO_817 (O_817,N_14329,N_12584);
nand UO_818 (O_818,N_14443,N_12526);
nand UO_819 (O_819,N_12314,N_13123);
or UO_820 (O_820,N_13583,N_14575);
or UO_821 (O_821,N_13332,N_13688);
xnor UO_822 (O_822,N_14848,N_14986);
nor UO_823 (O_823,N_14723,N_13399);
or UO_824 (O_824,N_12620,N_13826);
and UO_825 (O_825,N_12078,N_12369);
and UO_826 (O_826,N_12871,N_14052);
and UO_827 (O_827,N_12993,N_13374);
or UO_828 (O_828,N_14829,N_13435);
xor UO_829 (O_829,N_12118,N_12667);
nor UO_830 (O_830,N_12758,N_14945);
nor UO_831 (O_831,N_12007,N_12747);
or UO_832 (O_832,N_12407,N_14976);
and UO_833 (O_833,N_12352,N_14604);
or UO_834 (O_834,N_13156,N_12978);
or UO_835 (O_835,N_12989,N_12653);
nor UO_836 (O_836,N_14789,N_12854);
or UO_837 (O_837,N_13966,N_12829);
nand UO_838 (O_838,N_13534,N_14045);
nand UO_839 (O_839,N_13904,N_12311);
or UO_840 (O_840,N_13020,N_14190);
nand UO_841 (O_841,N_12779,N_13626);
nor UO_842 (O_842,N_13964,N_12498);
or UO_843 (O_843,N_12309,N_13439);
nor UO_844 (O_844,N_12560,N_12944);
nand UO_845 (O_845,N_14131,N_12875);
nor UO_846 (O_846,N_12616,N_14143);
nand UO_847 (O_847,N_12641,N_12453);
nand UO_848 (O_848,N_14317,N_14084);
nand UO_849 (O_849,N_13929,N_14533);
nor UO_850 (O_850,N_12139,N_12415);
nand UO_851 (O_851,N_13488,N_14173);
or UO_852 (O_852,N_13848,N_12650);
nand UO_853 (O_853,N_13075,N_12516);
and UO_854 (O_854,N_14535,N_13093);
or UO_855 (O_855,N_13853,N_12271);
nor UO_856 (O_856,N_13333,N_13385);
and UO_857 (O_857,N_13496,N_13568);
nand UO_858 (O_858,N_14083,N_13269);
and UO_859 (O_859,N_14159,N_12901);
nand UO_860 (O_860,N_12994,N_13931);
nor UO_861 (O_861,N_13902,N_14893);
or UO_862 (O_862,N_12489,N_12837);
or UO_863 (O_863,N_13856,N_14495);
nand UO_864 (O_864,N_14011,N_14226);
nand UO_865 (O_865,N_13999,N_14349);
or UO_866 (O_866,N_13802,N_12765);
or UO_867 (O_867,N_13501,N_13077);
nor UO_868 (O_868,N_13930,N_14536);
nand UO_869 (O_869,N_13187,N_12913);
and UO_870 (O_870,N_14586,N_14050);
nor UO_871 (O_871,N_14025,N_13361);
or UO_872 (O_872,N_13499,N_13095);
nand UO_873 (O_873,N_14080,N_13394);
or UO_874 (O_874,N_13813,N_13516);
nand UO_875 (O_875,N_13623,N_12056);
or UO_876 (O_876,N_14901,N_14768);
nor UO_877 (O_877,N_14703,N_14599);
nor UO_878 (O_878,N_14451,N_14557);
and UO_879 (O_879,N_12253,N_13841);
and UO_880 (O_880,N_14376,N_13446);
nor UO_881 (O_881,N_13720,N_12933);
xnor UO_882 (O_882,N_13297,N_13180);
nand UO_883 (O_883,N_14474,N_13250);
nor UO_884 (O_884,N_13315,N_14878);
or UO_885 (O_885,N_12462,N_14613);
and UO_886 (O_886,N_13224,N_13358);
or UO_887 (O_887,N_12555,N_14123);
or UO_888 (O_888,N_14646,N_14102);
nand UO_889 (O_889,N_14381,N_14359);
nor UO_890 (O_890,N_13793,N_12565);
nor UO_891 (O_891,N_12982,N_14790);
and UO_892 (O_892,N_14218,N_14250);
nor UO_893 (O_893,N_12469,N_12673);
nor UO_894 (O_894,N_14072,N_13440);
nand UO_895 (O_895,N_13454,N_14022);
nor UO_896 (O_896,N_12298,N_14117);
xor UO_897 (O_897,N_13521,N_14952);
nor UO_898 (O_898,N_14737,N_14740);
and UO_899 (O_899,N_13311,N_12736);
nor UO_900 (O_900,N_13744,N_13442);
and UO_901 (O_901,N_13610,N_13698);
nand UO_902 (O_902,N_13241,N_13033);
and UO_903 (O_903,N_12210,N_14275);
or UO_904 (O_904,N_14335,N_14437);
or UO_905 (O_905,N_12362,N_14207);
and UO_906 (O_906,N_13460,N_14185);
nand UO_907 (O_907,N_14338,N_12327);
or UO_908 (O_908,N_12948,N_12100);
nor UO_909 (O_909,N_14404,N_14326);
nand UO_910 (O_910,N_13976,N_14712);
nor UO_911 (O_911,N_12286,N_12598);
nor UO_912 (O_912,N_12644,N_14511);
or UO_913 (O_913,N_13335,N_12151);
or UO_914 (O_914,N_12121,N_14726);
nor UO_915 (O_915,N_13226,N_14048);
or UO_916 (O_916,N_13836,N_14942);
nor UO_917 (O_917,N_12807,N_14433);
and UO_918 (O_918,N_14115,N_12844);
nor UO_919 (O_919,N_13414,N_13221);
or UO_920 (O_920,N_13690,N_12961);
and UO_921 (O_921,N_13352,N_12709);
nand UO_922 (O_922,N_12430,N_14421);
or UO_923 (O_923,N_14672,N_14710);
nand UO_924 (O_924,N_13372,N_13833);
nor UO_925 (O_925,N_12422,N_13872);
nor UO_926 (O_926,N_12324,N_12319);
nand UO_927 (O_927,N_14358,N_14234);
or UO_928 (O_928,N_14666,N_14039);
or UO_929 (O_929,N_13185,N_12789);
nor UO_930 (O_930,N_14094,N_13464);
xnor UO_931 (O_931,N_14162,N_12847);
nor UO_932 (O_932,N_12852,N_14348);
and UO_933 (O_933,N_14402,N_12098);
nor UO_934 (O_934,N_14133,N_12070);
and UO_935 (O_935,N_14398,N_12935);
or UO_936 (O_936,N_13246,N_13363);
or UO_937 (O_937,N_12940,N_13520);
or UO_938 (O_938,N_14581,N_12604);
or UO_939 (O_939,N_13873,N_13789);
nor UO_940 (O_940,N_12172,N_12806);
and UO_941 (O_941,N_13027,N_12096);
nor UO_942 (O_942,N_14363,N_13316);
and UO_943 (O_943,N_12113,N_14354);
nor UO_944 (O_944,N_14504,N_14034);
nor UO_945 (O_945,N_13337,N_12677);
nor UO_946 (O_946,N_13314,N_14134);
or UO_947 (O_947,N_12233,N_12689);
nand UO_948 (O_948,N_12409,N_13946);
nor UO_949 (O_949,N_12244,N_14350);
nor UO_950 (O_950,N_13245,N_14626);
or UO_951 (O_951,N_14166,N_14307);
nor UO_952 (O_952,N_12275,N_12374);
and UO_953 (O_953,N_12320,N_14502);
and UO_954 (O_954,N_12531,N_12241);
nor UO_955 (O_955,N_13307,N_14814);
and UO_956 (O_956,N_13634,N_14770);
and UO_957 (O_957,N_13248,N_13773);
nor UO_958 (O_958,N_13808,N_13803);
nor UO_959 (O_959,N_12969,N_14744);
xnor UO_960 (O_960,N_13298,N_12562);
or UO_961 (O_961,N_13598,N_13829);
nand UO_962 (O_962,N_12186,N_13265);
nand UO_963 (O_963,N_14694,N_12266);
and UO_964 (O_964,N_12040,N_14196);
or UO_965 (O_965,N_12361,N_14914);
nor UO_966 (O_966,N_12632,N_13818);
nor UO_967 (O_967,N_13934,N_13293);
and UO_968 (O_968,N_13760,N_14006);
or UO_969 (O_969,N_14837,N_12845);
xnor UO_970 (O_970,N_14887,N_14128);
or UO_971 (O_971,N_14908,N_14950);
or UO_972 (O_972,N_12410,N_13722);
or UO_973 (O_973,N_12304,N_14018);
nand UO_974 (O_974,N_13569,N_14589);
nand UO_975 (O_975,N_14235,N_12486);
nand UO_976 (O_976,N_13207,N_13357);
and UO_977 (O_977,N_14044,N_12701);
xor UO_978 (O_978,N_13212,N_14692);
nor UO_979 (O_979,N_13742,N_12231);
or UO_980 (O_980,N_14546,N_12508);
nor UO_981 (O_981,N_13485,N_12149);
nand UO_982 (O_982,N_12946,N_14645);
nand UO_983 (O_983,N_14637,N_13761);
or UO_984 (O_984,N_12212,N_13411);
nand UO_985 (O_985,N_12760,N_12748);
or UO_986 (O_986,N_14124,N_13559);
nor UO_987 (O_987,N_14323,N_14099);
and UO_988 (O_988,N_12115,N_12858);
nand UO_989 (O_989,N_13785,N_13652);
nor UO_990 (O_990,N_14761,N_14530);
nand UO_991 (O_991,N_14663,N_13379);
nor UO_992 (O_992,N_12332,N_13244);
or UO_993 (O_993,N_14563,N_13831);
nand UO_994 (O_994,N_13451,N_12591);
nand UO_995 (O_995,N_13911,N_13377);
and UO_996 (O_996,N_12174,N_12140);
and UO_997 (O_997,N_13682,N_13768);
nor UO_998 (O_998,N_12291,N_12405);
and UO_999 (O_999,N_12506,N_14291);
nor UO_1000 (O_1000,N_12744,N_14222);
nand UO_1001 (O_1001,N_12285,N_12725);
and UO_1002 (O_1002,N_13914,N_14877);
and UO_1003 (O_1003,N_14970,N_13751);
or UO_1004 (O_1004,N_13163,N_14015);
nor UO_1005 (O_1005,N_14253,N_12502);
or UO_1006 (O_1006,N_12419,N_13979);
and UO_1007 (O_1007,N_13486,N_14884);
or UO_1008 (O_1008,N_14688,N_14797);
nor UO_1009 (O_1009,N_12850,N_12433);
nand UO_1010 (O_1010,N_13916,N_12790);
and UO_1011 (O_1011,N_12911,N_13469);
nor UO_1012 (O_1012,N_12581,N_12669);
nor UO_1013 (O_1013,N_12922,N_12395);
nor UO_1014 (O_1014,N_12693,N_12717);
or UO_1015 (O_1015,N_12923,N_13832);
nor UO_1016 (O_1016,N_12127,N_14113);
nand UO_1017 (O_1017,N_14640,N_12634);
and UO_1018 (O_1018,N_14499,N_14280);
nor UO_1019 (O_1019,N_12715,N_12879);
or UO_1020 (O_1020,N_12461,N_13327);
xor UO_1021 (O_1021,N_12567,N_14998);
or UO_1022 (O_1022,N_13958,N_12637);
nand UO_1023 (O_1023,N_14259,N_14383);
and UO_1024 (O_1024,N_14210,N_14183);
nand UO_1025 (O_1025,N_13780,N_14749);
nand UO_1026 (O_1026,N_12916,N_13852);
and UO_1027 (O_1027,N_12154,N_14585);
or UO_1028 (O_1028,N_14414,N_14778);
and UO_1029 (O_1029,N_12323,N_13551);
nor UO_1030 (O_1030,N_12328,N_13301);
or UO_1031 (O_1031,N_12305,N_12367);
nand UO_1032 (O_1032,N_12203,N_14202);
and UO_1033 (O_1033,N_14294,N_13974);
or UO_1034 (O_1034,N_14137,N_13913);
nor UO_1035 (O_1035,N_13531,N_13837);
nand UO_1036 (O_1036,N_13024,N_12401);
or UO_1037 (O_1037,N_13324,N_13312);
or UO_1038 (O_1038,N_14518,N_14106);
and UO_1039 (O_1039,N_14668,N_12718);
and UO_1040 (O_1040,N_13251,N_13019);
nand UO_1041 (O_1041,N_12884,N_14879);
and UO_1042 (O_1042,N_14796,N_14633);
nor UO_1043 (O_1043,N_12086,N_12659);
nor UO_1044 (O_1044,N_14405,N_13640);
and UO_1045 (O_1045,N_14284,N_13685);
nor UO_1046 (O_1046,N_13635,N_13822);
nor UO_1047 (O_1047,N_13354,N_13711);
nor UO_1048 (O_1048,N_14807,N_14821);
and UO_1049 (O_1049,N_12032,N_12494);
and UO_1050 (O_1050,N_12538,N_12814);
or UO_1051 (O_1051,N_14120,N_14567);
nand UO_1052 (O_1052,N_14559,N_14812);
nand UO_1053 (O_1053,N_13541,N_13879);
nand UO_1054 (O_1054,N_12630,N_14707);
or UO_1055 (O_1055,N_13341,N_14869);
nor UO_1056 (O_1056,N_13572,N_13864);
or UO_1057 (O_1057,N_14085,N_14743);
or UO_1058 (O_1058,N_13237,N_14156);
or UO_1059 (O_1059,N_13304,N_13779);
and UO_1060 (O_1060,N_14851,N_13655);
or UO_1061 (O_1061,N_14783,N_13502);
or UO_1062 (O_1062,N_13961,N_12256);
nor UO_1063 (O_1063,N_12885,N_14973);
nand UO_1064 (O_1064,N_14204,N_12626);
and UO_1065 (O_1065,N_12612,N_13880);
nor UO_1066 (O_1066,N_12980,N_14400);
nand UO_1067 (O_1067,N_14428,N_14787);
and UO_1068 (O_1068,N_14602,N_13430);
nor UO_1069 (O_1069,N_12588,N_13449);
or UO_1070 (O_1070,N_13453,N_14003);
and UO_1071 (O_1071,N_12264,N_12277);
nand UO_1072 (O_1072,N_14481,N_12861);
nor UO_1073 (O_1073,N_12336,N_14312);
and UO_1074 (O_1074,N_14971,N_13104);
and UO_1075 (O_1075,N_13204,N_14079);
nand UO_1076 (O_1076,N_13661,N_13788);
or UO_1077 (O_1077,N_13489,N_12129);
nand UO_1078 (O_1078,N_13540,N_14582);
or UO_1079 (O_1079,N_13233,N_12169);
nor UO_1080 (O_1080,N_12227,N_13264);
or UO_1081 (O_1081,N_12702,N_14788);
nor UO_1082 (O_1082,N_12881,N_14552);
nand UO_1083 (O_1083,N_13981,N_13429);
xor UO_1084 (O_1084,N_12018,N_14863);
nand UO_1085 (O_1085,N_14013,N_13618);
nand UO_1086 (O_1086,N_12674,N_14051);
and UO_1087 (O_1087,N_14512,N_12826);
nor UO_1088 (O_1088,N_14532,N_13947);
nand UO_1089 (O_1089,N_13127,N_14197);
nor UO_1090 (O_1090,N_13155,N_13679);
nand UO_1091 (O_1091,N_14194,N_14460);
nand UO_1092 (O_1092,N_13257,N_13586);
or UO_1093 (O_1093,N_12273,N_13851);
nor UO_1094 (O_1094,N_12815,N_14160);
or UO_1095 (O_1095,N_14175,N_13868);
and UO_1096 (O_1096,N_12730,N_12192);
and UO_1097 (O_1097,N_13952,N_14510);
or UO_1098 (O_1098,N_12440,N_14517);
nor UO_1099 (O_1099,N_14471,N_14715);
nand UO_1100 (O_1100,N_12267,N_13192);
or UO_1101 (O_1101,N_13203,N_13945);
or UO_1102 (O_1102,N_14266,N_13291);
nand UO_1103 (O_1103,N_13956,N_14996);
nand UO_1104 (O_1104,N_12537,N_14111);
nor UO_1105 (O_1105,N_12082,N_12378);
or UO_1106 (O_1106,N_12008,N_12904);
and UO_1107 (O_1107,N_14116,N_14426);
xor UO_1108 (O_1108,N_12593,N_13960);
or UO_1109 (O_1109,N_14506,N_14553);
nand UO_1110 (O_1110,N_14988,N_14388);
nor UO_1111 (O_1111,N_14337,N_12719);
nor UO_1112 (O_1112,N_14364,N_14228);
or UO_1113 (O_1113,N_14457,N_13924);
and UO_1114 (O_1114,N_13322,N_13725);
nor UO_1115 (O_1115,N_13821,N_13319);
or UO_1116 (O_1116,N_13202,N_12838);
nand UO_1117 (O_1117,N_13072,N_14298);
nand UO_1118 (O_1118,N_14375,N_14936);
and UO_1119 (O_1119,N_14578,N_13115);
nor UO_1120 (O_1120,N_14828,N_14793);
nand UO_1121 (O_1121,N_12583,N_12934);
xor UO_1122 (O_1122,N_13416,N_12343);
nor UO_1123 (O_1123,N_12602,N_12932);
nor UO_1124 (O_1124,N_12663,N_14468);
nor UO_1125 (O_1125,N_12514,N_12255);
or UO_1126 (O_1126,N_13348,N_12652);
nand UO_1127 (O_1127,N_13356,N_12216);
nand UO_1128 (O_1128,N_13968,N_13970);
nor UO_1129 (O_1129,N_12619,N_12541);
xnor UO_1130 (O_1130,N_13219,N_13141);
or UO_1131 (O_1131,N_13948,N_14858);
nor UO_1132 (O_1132,N_14297,N_13901);
or UO_1133 (O_1133,N_13752,N_13481);
nand UO_1134 (O_1134,N_13708,N_14760);
nand UO_1135 (O_1135,N_14933,N_13539);
nor UO_1136 (O_1136,N_13060,N_12411);
and UO_1137 (O_1137,N_14972,N_13927);
nor UO_1138 (O_1138,N_14654,N_14815);
and UO_1139 (O_1139,N_13987,N_12533);
or UO_1140 (O_1140,N_13395,N_13718);
xor UO_1141 (O_1141,N_12141,N_12763);
or UO_1142 (O_1142,N_12524,N_12670);
nand UO_1143 (O_1143,N_14779,N_14992);
and UO_1144 (O_1144,N_12519,N_12553);
nor UO_1145 (O_1145,N_14594,N_13118);
nand UO_1146 (O_1146,N_12688,N_13331);
nor UO_1147 (O_1147,N_14464,N_12782);
or UO_1148 (O_1148,N_12768,N_14674);
or UO_1149 (O_1149,N_14369,N_14844);
nand UO_1150 (O_1150,N_14529,N_14078);
and UO_1151 (O_1151,N_13647,N_14571);
or UO_1152 (O_1152,N_14037,N_12347);
and UO_1153 (O_1153,N_12794,N_13390);
or UO_1154 (O_1154,N_12396,N_14697);
and UO_1155 (O_1155,N_14295,N_14076);
or UO_1156 (O_1156,N_14411,N_13804);
and UO_1157 (O_1157,N_14930,N_14449);
nand UO_1158 (O_1158,N_13000,N_12114);
nand UO_1159 (O_1159,N_14561,N_14129);
nor UO_1160 (O_1160,N_12242,N_12570);
or UO_1161 (O_1161,N_12912,N_12312);
nand UO_1162 (O_1162,N_13951,N_13134);
nor UO_1163 (O_1163,N_14974,N_14021);
nand UO_1164 (O_1164,N_12629,N_12775);
nor UO_1165 (O_1165,N_13922,N_14413);
or UO_1166 (O_1166,N_13262,N_12201);
nand UO_1167 (O_1167,N_12394,N_13608);
or UO_1168 (O_1168,N_12191,N_13575);
nand UO_1169 (O_1169,N_13874,N_13120);
nor UO_1170 (O_1170,N_14478,N_12062);
nand UO_1171 (O_1171,N_12300,N_13525);
nor UO_1172 (O_1172,N_12112,N_14410);
or UO_1173 (O_1173,N_14785,N_12496);
or UO_1174 (O_1174,N_12822,N_12371);
or UO_1175 (O_1175,N_14059,N_12001);
nor UO_1176 (O_1176,N_12187,N_12441);
and UO_1177 (O_1177,N_14233,N_14458);
nand UO_1178 (O_1178,N_13313,N_12925);
and UO_1179 (O_1179,N_14954,N_12202);
or UO_1180 (O_1180,N_14727,N_13100);
or UO_1181 (O_1181,N_14020,N_13558);
or UO_1182 (O_1182,N_13425,N_14352);
or UO_1183 (O_1183,N_14994,N_12601);
nor UO_1184 (O_1184,N_13111,N_13545);
nor UO_1185 (O_1185,N_14252,N_13443);
nor UO_1186 (O_1186,N_13846,N_12597);
and UO_1187 (O_1187,N_13671,N_12799);
or UO_1188 (O_1188,N_12443,N_14608);
nor UO_1189 (O_1189,N_12063,N_13867);
or UO_1190 (O_1190,N_14574,N_12679);
and UO_1191 (O_1191,N_14278,N_14055);
and UO_1192 (O_1192,N_13498,N_12230);
and UO_1193 (O_1193,N_13420,N_13599);
and UO_1194 (O_1194,N_13533,N_14164);
nor UO_1195 (O_1195,N_14150,N_13217);
nand UO_1196 (O_1196,N_14493,N_13891);
or UO_1197 (O_1197,N_13668,N_13582);
and UO_1198 (O_1198,N_14172,N_12621);
and UO_1199 (O_1199,N_14065,N_14300);
nor UO_1200 (O_1200,N_14623,N_13317);
and UO_1201 (O_1201,N_12917,N_14618);
nand UO_1202 (O_1202,N_13847,N_13415);
or UO_1203 (O_1203,N_13051,N_12456);
nand UO_1204 (O_1204,N_12041,N_14534);
and UO_1205 (O_1205,N_14872,N_13510);
or UO_1206 (O_1206,N_12767,N_13909);
or UO_1207 (O_1207,N_13561,N_14008);
and UO_1208 (O_1208,N_13546,N_12571);
and UO_1209 (O_1209,N_12262,N_14316);
or UO_1210 (O_1210,N_13214,N_13694);
nand UO_1211 (O_1211,N_14367,N_14866);
nand UO_1212 (O_1212,N_14664,N_12160);
nor UO_1213 (O_1213,N_13408,N_12004);
nor UO_1214 (O_1214,N_12622,N_13162);
nand UO_1215 (O_1215,N_12245,N_13504);
nor UO_1216 (O_1216,N_12033,N_12762);
nor UO_1217 (O_1217,N_12888,N_13434);
and UO_1218 (O_1218,N_14418,N_12092);
and UO_1219 (O_1219,N_13097,N_14087);
nor UO_1220 (O_1220,N_12902,N_14978);
nor UO_1221 (O_1221,N_14766,N_12865);
and UO_1222 (O_1222,N_12025,N_12131);
nor UO_1223 (O_1223,N_12204,N_14047);
nor UO_1224 (O_1224,N_14548,N_13128);
nor UO_1225 (O_1225,N_14609,N_13897);
nand UO_1226 (O_1226,N_13835,N_14016);
or UO_1227 (O_1227,N_13777,N_12102);
nor UO_1228 (O_1228,N_13959,N_12093);
or UO_1229 (O_1229,N_14146,N_14997);
nor UO_1230 (O_1230,N_14477,N_13664);
nor UO_1231 (O_1231,N_12756,N_14631);
and UO_1232 (O_1232,N_14239,N_12992);
nor UO_1233 (O_1233,N_14095,N_12258);
and UO_1234 (O_1234,N_12960,N_12193);
nand UO_1235 (O_1235,N_13771,N_14238);
and UO_1236 (O_1236,N_12733,N_14292);
or UO_1237 (O_1237,N_12117,N_12614);
nor UO_1238 (O_1238,N_14498,N_13455);
nand UO_1239 (O_1239,N_13861,N_12466);
and UO_1240 (O_1240,N_13638,N_14171);
nand UO_1241 (O_1241,N_14487,N_13620);
nand UO_1242 (O_1242,N_14074,N_12097);
nand UO_1243 (O_1243,N_14287,N_12099);
nor UO_1244 (O_1244,N_12189,N_14100);
and UO_1245 (O_1245,N_13288,N_12949);
or UO_1246 (O_1246,N_12108,N_13428);
and UO_1247 (O_1247,N_14871,N_13456);
or UO_1248 (O_1248,N_13166,N_12680);
and UO_1249 (O_1249,N_13816,N_13200);
and UO_1250 (O_1250,N_14041,N_13939);
and UO_1251 (O_1251,N_14634,N_12690);
nand UO_1252 (O_1252,N_12042,N_14178);
and UO_1253 (O_1253,N_14864,N_14211);
nor UO_1254 (O_1254,N_14583,N_12307);
nand UO_1255 (O_1255,N_13071,N_13710);
nor UO_1256 (O_1256,N_14220,N_12851);
xor UO_1257 (O_1257,N_12543,N_14781);
nor UO_1258 (O_1258,N_14627,N_14558);
and UO_1259 (O_1259,N_13030,N_14026);
and UO_1260 (O_1260,N_12120,N_13038);
and UO_1261 (O_1261,N_12341,N_12272);
or UO_1262 (O_1262,N_12773,N_13053);
and UO_1263 (O_1263,N_13445,N_14360);
or UO_1264 (O_1264,N_13910,N_12953);
and UO_1265 (O_1265,N_13542,N_14777);
and UO_1266 (O_1266,N_13621,N_13949);
nor UO_1267 (O_1267,N_13477,N_13398);
nand UO_1268 (O_1268,N_12482,N_13380);
and UO_1269 (O_1269,N_14104,N_13056);
nand UO_1270 (O_1270,N_14346,N_12308);
nand UO_1271 (O_1271,N_12764,N_14836);
and UO_1272 (O_1272,N_12398,N_14521);
and UO_1273 (O_1273,N_13723,N_12306);
and UO_1274 (O_1274,N_12046,N_13739);
nand UO_1275 (O_1275,N_13726,N_13596);
or UO_1276 (O_1276,N_12316,N_13279);
nand UO_1277 (O_1277,N_13318,N_12205);
or UO_1278 (O_1278,N_14935,N_13800);
and UO_1279 (O_1279,N_14780,N_13188);
or UO_1280 (O_1280,N_12185,N_13205);
nand UO_1281 (O_1281,N_14170,N_12656);
nand UO_1282 (O_1282,N_12379,N_14289);
nand UO_1283 (O_1283,N_14708,N_13041);
nor UO_1284 (O_1284,N_14909,N_14669);
and UO_1285 (O_1285,N_12351,N_12215);
or UO_1286 (O_1286,N_14130,N_12633);
nand UO_1287 (O_1287,N_13436,N_13923);
and UO_1288 (O_1288,N_13148,N_12658);
nand UO_1289 (O_1289,N_14862,N_14230);
nand UO_1290 (O_1290,N_13660,N_14573);
or UO_1291 (O_1291,N_12150,N_13178);
xnor UO_1292 (O_1292,N_12257,N_13644);
nor UO_1293 (O_1293,N_12876,N_13705);
nor UO_1294 (O_1294,N_14823,N_14714);
xor UO_1295 (O_1295,N_12958,N_12265);
or UO_1296 (O_1296,N_12452,N_12340);
or UO_1297 (O_1297,N_12413,N_13801);
nor UO_1298 (O_1298,N_12578,N_14090);
nor UO_1299 (O_1299,N_13401,N_14378);
and UO_1300 (O_1300,N_14169,N_14803);
nand UO_1301 (O_1301,N_14765,N_12549);
or UO_1302 (O_1302,N_14401,N_12649);
nor UO_1303 (O_1303,N_14588,N_12446);
nor UO_1304 (O_1304,N_14685,N_13289);
nand UO_1305 (O_1305,N_12083,N_12381);
and UO_1306 (O_1306,N_13850,N_13167);
nor UO_1307 (O_1307,N_13096,N_14098);
nand UO_1308 (O_1308,N_13986,N_13990);
or UO_1309 (O_1309,N_14157,N_13840);
nand UO_1310 (O_1310,N_12054,N_12473);
or UO_1311 (O_1311,N_14625,N_12334);
and UO_1312 (O_1312,N_12313,N_13040);
nor UO_1313 (O_1313,N_12465,N_12586);
nor UO_1314 (O_1314,N_12750,N_14203);
nand UO_1315 (O_1315,N_14254,N_12510);
nand UO_1316 (O_1316,N_14719,N_13133);
nor UO_1317 (O_1317,N_14964,N_14362);
or UO_1318 (O_1318,N_12695,N_12540);
or UO_1319 (O_1319,N_14480,N_13928);
nand UO_1320 (O_1320,N_14756,N_14390);
and UO_1321 (O_1321,N_13462,N_13169);
nand UO_1322 (O_1322,N_12268,N_12592);
and UO_1323 (O_1323,N_12051,N_14181);
nor UO_1324 (O_1324,N_14036,N_13173);
nor UO_1325 (O_1325,N_12303,N_14991);
or UO_1326 (O_1326,N_14860,N_14501);
or UO_1327 (O_1327,N_12296,N_12728);
or UO_1328 (O_1328,N_14849,N_13073);
nand UO_1329 (O_1329,N_13893,N_14145);
nor UO_1330 (O_1330,N_12503,N_14661);
nor UO_1331 (O_1331,N_13920,N_14709);
xnor UO_1332 (O_1332,N_14810,N_12330);
nor UO_1333 (O_1333,N_12606,N_12996);
nand UO_1334 (O_1334,N_14769,N_13266);
and UO_1335 (O_1335,N_12809,N_12915);
xnor UO_1336 (O_1336,N_13255,N_13063);
or UO_1337 (O_1337,N_12587,N_14959);
or UO_1338 (O_1338,N_14167,N_13465);
and UO_1339 (O_1339,N_13085,N_13114);
or UO_1340 (O_1340,N_13196,N_12757);
nor UO_1341 (O_1341,N_12390,N_14251);
nand UO_1342 (O_1342,N_13988,N_14054);
or UO_1343 (O_1343,N_12397,N_14545);
or UO_1344 (O_1344,N_12138,N_13198);
nand UO_1345 (O_1345,N_13045,N_13105);
and UO_1346 (O_1346,N_13254,N_13578);
or UO_1347 (O_1347,N_13895,N_12480);
and UO_1348 (O_1348,N_12740,N_14962);
and UO_1349 (O_1349,N_12735,N_12898);
or UO_1350 (O_1350,N_13823,N_14484);
nand UO_1351 (O_1351,N_14373,N_13814);
or UO_1352 (O_1352,N_13383,N_14344);
nor UO_1353 (O_1353,N_14932,N_14064);
nand UO_1354 (O_1354,N_14855,N_13611);
nand UO_1355 (O_1355,N_13866,N_13400);
and UO_1356 (O_1356,N_14804,N_14236);
nand UO_1357 (O_1357,N_12753,N_14629);
and UO_1358 (O_1358,N_13878,N_14496);
nor UO_1359 (O_1359,N_14920,N_12109);
nand UO_1360 (O_1360,N_12076,N_14596);
or UO_1361 (O_1361,N_12525,N_13300);
or UO_1362 (O_1362,N_14856,N_14503);
nor UO_1363 (O_1363,N_12431,N_14182);
and UO_1364 (O_1364,N_13179,N_13378);
nand UO_1365 (O_1365,N_14886,N_14667);
and UO_1366 (O_1366,N_13649,N_13515);
and UO_1367 (O_1367,N_12048,N_12769);
or UO_1368 (O_1368,N_12427,N_12761);
and UO_1369 (O_1369,N_13174,N_12892);
and UO_1370 (O_1370,N_14665,N_12743);
or UO_1371 (O_1371,N_14038,N_14476);
nand UO_1372 (O_1372,N_14751,N_14180);
nor UO_1373 (O_1373,N_14314,N_13129);
or UO_1374 (O_1374,N_13296,N_14742);
nor UO_1375 (O_1375,N_14931,N_12354);
and UO_1376 (O_1376,N_13177,N_14568);
xnor UO_1377 (O_1377,N_12623,N_14999);
and UO_1378 (O_1378,N_12551,N_12137);
or UO_1379 (O_1379,N_14357,N_13662);
nor UO_1380 (O_1380,N_14873,N_13692);
nor UO_1381 (O_1381,N_13613,N_13843);
or UO_1382 (O_1382,N_14491,N_14904);
or UO_1383 (O_1383,N_13790,N_12429);
nand UO_1384 (O_1384,N_14000,N_13774);
or UO_1385 (O_1385,N_12613,N_13258);
nand UO_1386 (O_1386,N_12207,N_14639);
nor UO_1387 (O_1387,N_12778,N_13247);
nor UO_1388 (O_1388,N_13985,N_12370);
or UO_1389 (O_1389,N_14570,N_13547);
or UO_1390 (O_1390,N_14750,N_14232);
or UO_1391 (O_1391,N_13272,N_12474);
or UO_1392 (O_1392,N_14382,N_12878);
or UO_1393 (O_1393,N_12144,N_13397);
xnor UO_1394 (O_1394,N_12069,N_13021);
or UO_1395 (O_1395,N_13733,N_14482);
nor UO_1396 (O_1396,N_13854,N_13845);
or UO_1397 (O_1397,N_12511,N_12849);
nand UO_1398 (O_1398,N_14135,N_13877);
nand UO_1399 (O_1399,N_13229,N_14900);
and UO_1400 (O_1400,N_13487,N_14831);
nand UO_1401 (O_1401,N_12534,N_12366);
nand UO_1402 (O_1402,N_14361,N_12073);
and UO_1403 (O_1403,N_13276,N_13543);
or UO_1404 (O_1404,N_13160,N_13627);
nor UO_1405 (O_1405,N_14754,N_14826);
or UO_1406 (O_1406,N_12694,N_13184);
nor UO_1407 (O_1407,N_12043,N_12235);
nor UO_1408 (O_1408,N_14201,N_14845);
and UO_1409 (O_1409,N_13234,N_14033);
or UO_1410 (O_1410,N_13259,N_13194);
or UO_1411 (O_1411,N_14580,N_12143);
or UO_1412 (O_1412,N_13645,N_12746);
nand UO_1413 (O_1413,N_12142,N_12983);
nor UO_1414 (O_1414,N_12841,N_14237);
nand UO_1415 (O_1415,N_13424,N_14332);
nand UO_1416 (O_1416,N_12134,N_12819);
nor UO_1417 (O_1417,N_14757,N_12458);
and UO_1418 (O_1418,N_13908,N_14285);
or UO_1419 (O_1419,N_12091,N_12893);
or UO_1420 (O_1420,N_12986,N_13513);
and UO_1421 (O_1421,N_13508,N_14446);
nor UO_1422 (O_1422,N_13950,N_14062);
nor UO_1423 (O_1423,N_13756,N_12995);
and UO_1424 (O_1424,N_13058,N_12222);
nand UO_1425 (O_1425,N_13625,N_14693);
nor UO_1426 (O_1426,N_14441,N_13825);
and UO_1427 (O_1427,N_13112,N_14371);
and UO_1428 (O_1428,N_12226,N_13765);
or UO_1429 (O_1429,N_12544,N_14767);
and UO_1430 (O_1430,N_12249,N_12426);
nor UO_1431 (O_1431,N_13494,N_14071);
and UO_1432 (O_1432,N_14892,N_12607);
or UO_1433 (O_1433,N_12420,N_12234);
or UO_1434 (O_1434,N_13842,N_13152);
nand UO_1435 (O_1435,N_14385,N_13242);
nand UO_1436 (O_1436,N_12550,N_13240);
nand UO_1437 (O_1437,N_12926,N_13220);
and UO_1438 (O_1438,N_12646,N_14902);
and UO_1439 (O_1439,N_13225,N_14881);
nand UO_1440 (O_1440,N_12232,N_14852);
or UO_1441 (O_1441,N_12059,N_13228);
nor UO_1442 (O_1442,N_12194,N_13629);
nand UO_1443 (O_1443,N_13759,N_12164);
and UO_1444 (O_1444,N_13707,N_12977);
xnor UO_1445 (O_1445,N_13669,N_14231);
and UO_1446 (O_1446,N_13008,N_14882);
nand UO_1447 (O_1447,N_14279,N_14415);
nor UO_1448 (O_1448,N_13320,N_13236);
or UO_1449 (O_1449,N_14924,N_14303);
xor UO_1450 (O_1450,N_14264,N_14525);
nand UO_1451 (O_1451,N_13002,N_14520);
or UO_1452 (O_1452,N_13732,N_13745);
nor UO_1453 (O_1453,N_13709,N_14894);
and UO_1454 (O_1454,N_14854,N_14579);
nor UO_1455 (O_1455,N_13281,N_14620);
and UO_1456 (O_1456,N_14758,N_12217);
nand UO_1457 (O_1457,N_12828,N_13783);
nor UO_1458 (O_1458,N_12219,N_12821);
or UO_1459 (O_1459,N_14490,N_12910);
and UO_1460 (O_1460,N_12971,N_13159);
xor UO_1461 (O_1461,N_13161,N_14155);
and UO_1462 (O_1462,N_13544,N_13068);
and UO_1463 (O_1463,N_14213,N_13607);
nand UO_1464 (O_1464,N_14334,N_13139);
or UO_1465 (O_1465,N_13285,N_14799);
nor UO_1466 (O_1466,N_14209,N_13001);
nor UO_1467 (O_1467,N_13574,N_13537);
xor UO_1468 (O_1468,N_13881,N_14806);
nor UO_1469 (O_1469,N_12816,N_13109);
or UO_1470 (O_1470,N_14200,N_12795);
or UO_1471 (O_1471,N_14308,N_13292);
or UO_1472 (O_1472,N_13274,N_12963);
nor UO_1473 (O_1473,N_12179,N_12722);
nand UO_1474 (O_1474,N_14330,N_12434);
nand UO_1475 (O_1475,N_12785,N_12990);
or UO_1476 (O_1476,N_12155,N_12521);
nor UO_1477 (O_1477,N_13665,N_14313);
nor UO_1478 (O_1478,N_12110,N_12280);
or UO_1479 (O_1479,N_13622,N_12084);
or UO_1480 (O_1480,N_14734,N_13762);
nor UO_1481 (O_1481,N_14389,N_12823);
and UO_1482 (O_1482,N_13362,N_12181);
and UO_1483 (O_1483,N_13616,N_14695);
nand UO_1484 (O_1484,N_12372,N_14328);
and UO_1485 (O_1485,N_12512,N_14431);
xor UO_1486 (O_1486,N_12116,N_12574);
nand UO_1487 (O_1487,N_12774,N_14321);
or UO_1488 (O_1488,N_13838,N_13857);
nor UO_1489 (O_1489,N_12777,N_14486);
nand UO_1490 (O_1490,N_12263,N_13243);
nand UO_1491 (O_1491,N_14603,N_14403);
nand UO_1492 (O_1492,N_13227,N_14425);
nor UO_1493 (O_1493,N_14028,N_12464);
and UO_1494 (O_1494,N_14419,N_13418);
nand UO_1495 (O_1495,N_13149,N_14721);
and UO_1496 (O_1496,N_14027,N_13810);
and UO_1497 (O_1497,N_13683,N_13807);
nor UO_1498 (O_1498,N_13046,N_14890);
nand UO_1499 (O_1499,N_14651,N_12802);
nand UO_1500 (O_1500,N_12549,N_14151);
and UO_1501 (O_1501,N_12170,N_12987);
or UO_1502 (O_1502,N_13129,N_14940);
or UO_1503 (O_1503,N_14297,N_14475);
and UO_1504 (O_1504,N_14213,N_12896);
nand UO_1505 (O_1505,N_14030,N_12259);
nand UO_1506 (O_1506,N_12517,N_13526);
nor UO_1507 (O_1507,N_12496,N_12004);
nand UO_1508 (O_1508,N_14291,N_13659);
and UO_1509 (O_1509,N_14108,N_14695);
or UO_1510 (O_1510,N_12294,N_14381);
or UO_1511 (O_1511,N_13413,N_14766);
or UO_1512 (O_1512,N_12116,N_14878);
nor UO_1513 (O_1513,N_13808,N_12171);
and UO_1514 (O_1514,N_14723,N_13350);
nor UO_1515 (O_1515,N_13455,N_13842);
nor UO_1516 (O_1516,N_12032,N_14687);
or UO_1517 (O_1517,N_13139,N_12580);
and UO_1518 (O_1518,N_12825,N_14257);
nor UO_1519 (O_1519,N_12436,N_13180);
and UO_1520 (O_1520,N_12199,N_12642);
nand UO_1521 (O_1521,N_14773,N_13488);
xor UO_1522 (O_1522,N_12873,N_13189);
or UO_1523 (O_1523,N_13366,N_14401);
nand UO_1524 (O_1524,N_13787,N_12354);
nor UO_1525 (O_1525,N_12565,N_13090);
or UO_1526 (O_1526,N_12674,N_14251);
and UO_1527 (O_1527,N_13612,N_13756);
nor UO_1528 (O_1528,N_12792,N_13917);
or UO_1529 (O_1529,N_13113,N_14053);
and UO_1530 (O_1530,N_12733,N_14528);
nor UO_1531 (O_1531,N_12423,N_14858);
and UO_1532 (O_1532,N_13842,N_12940);
and UO_1533 (O_1533,N_14977,N_14740);
and UO_1534 (O_1534,N_14172,N_14895);
and UO_1535 (O_1535,N_13972,N_12247);
nor UO_1536 (O_1536,N_12189,N_14266);
or UO_1537 (O_1537,N_13247,N_14221);
and UO_1538 (O_1538,N_13188,N_13993);
xnor UO_1539 (O_1539,N_13292,N_14990);
xor UO_1540 (O_1540,N_13545,N_12008);
and UO_1541 (O_1541,N_14800,N_12970);
nand UO_1542 (O_1542,N_14093,N_12227);
or UO_1543 (O_1543,N_12337,N_14841);
and UO_1544 (O_1544,N_12454,N_14068);
and UO_1545 (O_1545,N_12746,N_13515);
and UO_1546 (O_1546,N_14262,N_14540);
nand UO_1547 (O_1547,N_14301,N_12120);
and UO_1548 (O_1548,N_12485,N_14443);
or UO_1549 (O_1549,N_12510,N_12381);
or UO_1550 (O_1550,N_12925,N_12068);
or UO_1551 (O_1551,N_12903,N_12849);
nor UO_1552 (O_1552,N_12274,N_14822);
and UO_1553 (O_1553,N_13697,N_14654);
nand UO_1554 (O_1554,N_12002,N_12834);
nand UO_1555 (O_1555,N_12051,N_12797);
nand UO_1556 (O_1556,N_13984,N_12070);
nand UO_1557 (O_1557,N_13984,N_13990);
or UO_1558 (O_1558,N_13113,N_13981);
nor UO_1559 (O_1559,N_14609,N_14117);
and UO_1560 (O_1560,N_12742,N_14478);
and UO_1561 (O_1561,N_13713,N_14422);
nor UO_1562 (O_1562,N_12710,N_14764);
nor UO_1563 (O_1563,N_12072,N_12028);
nor UO_1564 (O_1564,N_12533,N_12628);
or UO_1565 (O_1565,N_13533,N_12651);
nor UO_1566 (O_1566,N_13785,N_13129);
nor UO_1567 (O_1567,N_13688,N_13798);
nand UO_1568 (O_1568,N_14224,N_13369);
nor UO_1569 (O_1569,N_14984,N_13780);
nor UO_1570 (O_1570,N_14120,N_13459);
or UO_1571 (O_1571,N_12848,N_14099);
or UO_1572 (O_1572,N_12369,N_14081);
and UO_1573 (O_1573,N_13919,N_13945);
nand UO_1574 (O_1574,N_14717,N_14769);
nor UO_1575 (O_1575,N_13614,N_12444);
and UO_1576 (O_1576,N_13160,N_14819);
or UO_1577 (O_1577,N_12995,N_13149);
nor UO_1578 (O_1578,N_14872,N_13921);
or UO_1579 (O_1579,N_13823,N_12559);
nor UO_1580 (O_1580,N_12043,N_13646);
and UO_1581 (O_1581,N_14600,N_12374);
and UO_1582 (O_1582,N_13478,N_14934);
and UO_1583 (O_1583,N_14332,N_12129);
nor UO_1584 (O_1584,N_12465,N_12944);
or UO_1585 (O_1585,N_13053,N_13924);
nand UO_1586 (O_1586,N_14613,N_12652);
or UO_1587 (O_1587,N_14323,N_13088);
or UO_1588 (O_1588,N_13596,N_13715);
and UO_1589 (O_1589,N_14675,N_12986);
or UO_1590 (O_1590,N_14166,N_12533);
nand UO_1591 (O_1591,N_12118,N_14653);
nor UO_1592 (O_1592,N_13767,N_12854);
nand UO_1593 (O_1593,N_13679,N_14464);
or UO_1594 (O_1594,N_13479,N_12753);
nor UO_1595 (O_1595,N_14919,N_12455);
or UO_1596 (O_1596,N_13428,N_13619);
or UO_1597 (O_1597,N_13345,N_13429);
and UO_1598 (O_1598,N_14219,N_13764);
nor UO_1599 (O_1599,N_14652,N_14272);
or UO_1600 (O_1600,N_14244,N_14976);
nand UO_1601 (O_1601,N_12545,N_12961);
or UO_1602 (O_1602,N_14520,N_14113);
and UO_1603 (O_1603,N_14616,N_12493);
nand UO_1604 (O_1604,N_13866,N_12765);
and UO_1605 (O_1605,N_13769,N_13069);
and UO_1606 (O_1606,N_12798,N_12448);
or UO_1607 (O_1607,N_13996,N_13235);
and UO_1608 (O_1608,N_14218,N_13171);
or UO_1609 (O_1609,N_14915,N_14393);
nor UO_1610 (O_1610,N_13528,N_14263);
or UO_1611 (O_1611,N_12556,N_12209);
nor UO_1612 (O_1612,N_12877,N_13994);
and UO_1613 (O_1613,N_14922,N_12918);
xor UO_1614 (O_1614,N_14168,N_13172);
nor UO_1615 (O_1615,N_13776,N_13685);
and UO_1616 (O_1616,N_12513,N_12177);
nor UO_1617 (O_1617,N_13075,N_12208);
nor UO_1618 (O_1618,N_13734,N_13163);
and UO_1619 (O_1619,N_13725,N_12074);
and UO_1620 (O_1620,N_14943,N_12579);
or UO_1621 (O_1621,N_14670,N_13270);
or UO_1622 (O_1622,N_12141,N_14129);
and UO_1623 (O_1623,N_14676,N_13403);
nor UO_1624 (O_1624,N_13680,N_14106);
nor UO_1625 (O_1625,N_12022,N_14267);
xor UO_1626 (O_1626,N_14848,N_12062);
or UO_1627 (O_1627,N_14033,N_14532);
or UO_1628 (O_1628,N_14284,N_13986);
or UO_1629 (O_1629,N_14960,N_12295);
nand UO_1630 (O_1630,N_14655,N_12437);
and UO_1631 (O_1631,N_13390,N_13979);
nand UO_1632 (O_1632,N_13505,N_12407);
and UO_1633 (O_1633,N_12753,N_12011);
or UO_1634 (O_1634,N_12820,N_14688);
and UO_1635 (O_1635,N_13702,N_12685);
nand UO_1636 (O_1636,N_13022,N_14298);
nor UO_1637 (O_1637,N_12650,N_13917);
nand UO_1638 (O_1638,N_13547,N_13690);
and UO_1639 (O_1639,N_12707,N_13419);
nand UO_1640 (O_1640,N_12344,N_13067);
and UO_1641 (O_1641,N_13692,N_13395);
nand UO_1642 (O_1642,N_12583,N_14898);
nand UO_1643 (O_1643,N_12784,N_14057);
and UO_1644 (O_1644,N_14037,N_13984);
or UO_1645 (O_1645,N_14762,N_13872);
nand UO_1646 (O_1646,N_12203,N_12980);
nor UO_1647 (O_1647,N_14575,N_12692);
nand UO_1648 (O_1648,N_13038,N_12611);
nor UO_1649 (O_1649,N_14339,N_12294);
nor UO_1650 (O_1650,N_13307,N_13886);
nor UO_1651 (O_1651,N_13418,N_14177);
nor UO_1652 (O_1652,N_12329,N_13659);
and UO_1653 (O_1653,N_14997,N_14187);
nand UO_1654 (O_1654,N_13562,N_14294);
nor UO_1655 (O_1655,N_14226,N_14242);
nand UO_1656 (O_1656,N_14739,N_12694);
nand UO_1657 (O_1657,N_14942,N_14787);
or UO_1658 (O_1658,N_14188,N_12117);
or UO_1659 (O_1659,N_14972,N_14642);
or UO_1660 (O_1660,N_12962,N_14998);
or UO_1661 (O_1661,N_14933,N_12606);
nor UO_1662 (O_1662,N_12499,N_13272);
nand UO_1663 (O_1663,N_13406,N_13250);
nor UO_1664 (O_1664,N_13331,N_14650);
or UO_1665 (O_1665,N_12311,N_13413);
nand UO_1666 (O_1666,N_13300,N_14613);
or UO_1667 (O_1667,N_12379,N_14324);
nor UO_1668 (O_1668,N_14535,N_14729);
nor UO_1669 (O_1669,N_14636,N_14403);
and UO_1670 (O_1670,N_14391,N_13287);
nor UO_1671 (O_1671,N_14623,N_14974);
nand UO_1672 (O_1672,N_14948,N_14138);
nor UO_1673 (O_1673,N_13594,N_13493);
nor UO_1674 (O_1674,N_12192,N_12311);
and UO_1675 (O_1675,N_12643,N_14216);
or UO_1676 (O_1676,N_14797,N_13495);
and UO_1677 (O_1677,N_13898,N_12184);
nand UO_1678 (O_1678,N_14001,N_13136);
nand UO_1679 (O_1679,N_14887,N_13394);
xnor UO_1680 (O_1680,N_14240,N_14348);
or UO_1681 (O_1681,N_13915,N_13879);
xnor UO_1682 (O_1682,N_12273,N_13538);
or UO_1683 (O_1683,N_12611,N_12492);
nor UO_1684 (O_1684,N_12106,N_14746);
or UO_1685 (O_1685,N_14180,N_13331);
or UO_1686 (O_1686,N_13882,N_13036);
nand UO_1687 (O_1687,N_13295,N_14728);
nor UO_1688 (O_1688,N_14733,N_12012);
nor UO_1689 (O_1689,N_13162,N_13808);
nand UO_1690 (O_1690,N_12500,N_12986);
or UO_1691 (O_1691,N_14397,N_12705);
nor UO_1692 (O_1692,N_13934,N_12868);
nor UO_1693 (O_1693,N_14019,N_14676);
nor UO_1694 (O_1694,N_14228,N_14460);
and UO_1695 (O_1695,N_13313,N_13524);
nor UO_1696 (O_1696,N_12429,N_14857);
nor UO_1697 (O_1697,N_12617,N_12939);
nand UO_1698 (O_1698,N_13304,N_14973);
nand UO_1699 (O_1699,N_12345,N_13686);
or UO_1700 (O_1700,N_14436,N_13006);
and UO_1701 (O_1701,N_12318,N_14908);
or UO_1702 (O_1702,N_12380,N_14773);
and UO_1703 (O_1703,N_14201,N_13989);
and UO_1704 (O_1704,N_13487,N_12216);
and UO_1705 (O_1705,N_13638,N_14748);
or UO_1706 (O_1706,N_12334,N_14573);
and UO_1707 (O_1707,N_12972,N_14888);
nand UO_1708 (O_1708,N_13125,N_13616);
or UO_1709 (O_1709,N_12355,N_12757);
or UO_1710 (O_1710,N_13123,N_12288);
and UO_1711 (O_1711,N_14726,N_13938);
and UO_1712 (O_1712,N_12088,N_14090);
nor UO_1713 (O_1713,N_12563,N_14064);
nand UO_1714 (O_1714,N_14737,N_13767);
nand UO_1715 (O_1715,N_14523,N_14881);
nand UO_1716 (O_1716,N_12370,N_12807);
and UO_1717 (O_1717,N_14020,N_14953);
and UO_1718 (O_1718,N_13701,N_12923);
or UO_1719 (O_1719,N_12292,N_14548);
and UO_1720 (O_1720,N_12333,N_12486);
and UO_1721 (O_1721,N_13468,N_12315);
nand UO_1722 (O_1722,N_14789,N_14719);
nand UO_1723 (O_1723,N_12235,N_13161);
xnor UO_1724 (O_1724,N_12361,N_12159);
and UO_1725 (O_1725,N_12956,N_14723);
and UO_1726 (O_1726,N_14375,N_13697);
nand UO_1727 (O_1727,N_14213,N_14875);
and UO_1728 (O_1728,N_12076,N_13484);
nand UO_1729 (O_1729,N_12093,N_14206);
nand UO_1730 (O_1730,N_13255,N_14291);
nor UO_1731 (O_1731,N_14818,N_12644);
or UO_1732 (O_1732,N_12316,N_12182);
or UO_1733 (O_1733,N_13724,N_14433);
and UO_1734 (O_1734,N_12128,N_14224);
nor UO_1735 (O_1735,N_14778,N_13464);
nor UO_1736 (O_1736,N_12421,N_12922);
or UO_1737 (O_1737,N_13432,N_13214);
or UO_1738 (O_1738,N_13674,N_14973);
nor UO_1739 (O_1739,N_12480,N_14670);
xnor UO_1740 (O_1740,N_14715,N_13493);
nand UO_1741 (O_1741,N_12367,N_13694);
nand UO_1742 (O_1742,N_14936,N_12092);
nand UO_1743 (O_1743,N_12149,N_12956);
or UO_1744 (O_1744,N_14114,N_14077);
or UO_1745 (O_1745,N_13118,N_13318);
nor UO_1746 (O_1746,N_14943,N_12919);
or UO_1747 (O_1747,N_13944,N_13143);
nand UO_1748 (O_1748,N_14433,N_12081);
nand UO_1749 (O_1749,N_13718,N_13894);
nand UO_1750 (O_1750,N_12139,N_14866);
nand UO_1751 (O_1751,N_13491,N_14952);
nand UO_1752 (O_1752,N_12793,N_14542);
nand UO_1753 (O_1753,N_14863,N_14367);
nand UO_1754 (O_1754,N_12976,N_13557);
nor UO_1755 (O_1755,N_12697,N_14305);
and UO_1756 (O_1756,N_12147,N_14073);
and UO_1757 (O_1757,N_13738,N_13510);
or UO_1758 (O_1758,N_13153,N_13530);
or UO_1759 (O_1759,N_13034,N_14205);
nor UO_1760 (O_1760,N_12865,N_14753);
nor UO_1761 (O_1761,N_13738,N_12370);
or UO_1762 (O_1762,N_12766,N_14283);
and UO_1763 (O_1763,N_13580,N_12404);
or UO_1764 (O_1764,N_14140,N_13207);
or UO_1765 (O_1765,N_12977,N_14833);
or UO_1766 (O_1766,N_12196,N_13668);
or UO_1767 (O_1767,N_13231,N_13278);
and UO_1768 (O_1768,N_13705,N_14048);
and UO_1769 (O_1769,N_13379,N_14940);
and UO_1770 (O_1770,N_12814,N_12446);
nand UO_1771 (O_1771,N_14387,N_14393);
or UO_1772 (O_1772,N_14653,N_14917);
and UO_1773 (O_1773,N_12984,N_14721);
nand UO_1774 (O_1774,N_13695,N_13032);
and UO_1775 (O_1775,N_12170,N_14036);
nor UO_1776 (O_1776,N_13519,N_14779);
or UO_1777 (O_1777,N_14513,N_13447);
nand UO_1778 (O_1778,N_12672,N_12018);
or UO_1779 (O_1779,N_12754,N_14351);
xor UO_1780 (O_1780,N_14492,N_14318);
nand UO_1781 (O_1781,N_12581,N_13040);
and UO_1782 (O_1782,N_14887,N_13486);
nand UO_1783 (O_1783,N_14171,N_14198);
or UO_1784 (O_1784,N_13525,N_14875);
nor UO_1785 (O_1785,N_14734,N_12319);
nor UO_1786 (O_1786,N_13252,N_14813);
or UO_1787 (O_1787,N_14531,N_13872);
nor UO_1788 (O_1788,N_13925,N_14480);
and UO_1789 (O_1789,N_12400,N_12396);
nand UO_1790 (O_1790,N_14518,N_14322);
nor UO_1791 (O_1791,N_13782,N_12183);
or UO_1792 (O_1792,N_14521,N_12757);
or UO_1793 (O_1793,N_12845,N_12414);
nor UO_1794 (O_1794,N_13991,N_14540);
nand UO_1795 (O_1795,N_13809,N_14689);
and UO_1796 (O_1796,N_14299,N_12545);
nand UO_1797 (O_1797,N_13649,N_13722);
xor UO_1798 (O_1798,N_13007,N_13675);
nor UO_1799 (O_1799,N_13251,N_13201);
and UO_1800 (O_1800,N_14238,N_14012);
nand UO_1801 (O_1801,N_12896,N_13039);
and UO_1802 (O_1802,N_14006,N_12530);
and UO_1803 (O_1803,N_12272,N_13896);
xnor UO_1804 (O_1804,N_12289,N_14924);
or UO_1805 (O_1805,N_12708,N_12928);
nor UO_1806 (O_1806,N_12933,N_12493);
nor UO_1807 (O_1807,N_12522,N_14834);
or UO_1808 (O_1808,N_13442,N_14124);
xnor UO_1809 (O_1809,N_13300,N_12614);
or UO_1810 (O_1810,N_14850,N_14357);
nor UO_1811 (O_1811,N_13669,N_12365);
nor UO_1812 (O_1812,N_13890,N_13938);
nand UO_1813 (O_1813,N_13178,N_14733);
and UO_1814 (O_1814,N_12555,N_14260);
nor UO_1815 (O_1815,N_13222,N_13287);
nand UO_1816 (O_1816,N_14156,N_13363);
and UO_1817 (O_1817,N_12786,N_13835);
or UO_1818 (O_1818,N_12179,N_14978);
or UO_1819 (O_1819,N_14442,N_12219);
nand UO_1820 (O_1820,N_12043,N_13947);
nor UO_1821 (O_1821,N_13933,N_13758);
or UO_1822 (O_1822,N_14023,N_14584);
or UO_1823 (O_1823,N_13072,N_12942);
nand UO_1824 (O_1824,N_12583,N_14906);
nor UO_1825 (O_1825,N_14360,N_14562);
nand UO_1826 (O_1826,N_12443,N_13811);
nand UO_1827 (O_1827,N_14926,N_13409);
nor UO_1828 (O_1828,N_14569,N_14618);
nand UO_1829 (O_1829,N_12902,N_13008);
nor UO_1830 (O_1830,N_13446,N_13025);
nand UO_1831 (O_1831,N_12608,N_13710);
nand UO_1832 (O_1832,N_12958,N_13429);
nor UO_1833 (O_1833,N_13303,N_14704);
and UO_1834 (O_1834,N_12749,N_14697);
xnor UO_1835 (O_1835,N_12593,N_13178);
nand UO_1836 (O_1836,N_12396,N_13951);
xnor UO_1837 (O_1837,N_13902,N_14992);
and UO_1838 (O_1838,N_13085,N_12831);
nand UO_1839 (O_1839,N_13734,N_14807);
nor UO_1840 (O_1840,N_12577,N_13006);
nand UO_1841 (O_1841,N_14652,N_12371);
nand UO_1842 (O_1842,N_14074,N_14926);
and UO_1843 (O_1843,N_13550,N_13536);
nand UO_1844 (O_1844,N_13756,N_13259);
nand UO_1845 (O_1845,N_12232,N_14987);
or UO_1846 (O_1846,N_14867,N_12126);
nand UO_1847 (O_1847,N_13691,N_14263);
and UO_1848 (O_1848,N_12586,N_14314);
nand UO_1849 (O_1849,N_13305,N_14188);
nand UO_1850 (O_1850,N_12842,N_13642);
and UO_1851 (O_1851,N_12066,N_14713);
nor UO_1852 (O_1852,N_14989,N_14900);
or UO_1853 (O_1853,N_13601,N_12264);
or UO_1854 (O_1854,N_14255,N_13679);
or UO_1855 (O_1855,N_14869,N_14470);
or UO_1856 (O_1856,N_13237,N_12800);
nand UO_1857 (O_1857,N_12787,N_14002);
xnor UO_1858 (O_1858,N_12519,N_14828);
and UO_1859 (O_1859,N_14122,N_14143);
nor UO_1860 (O_1860,N_14967,N_12268);
and UO_1861 (O_1861,N_12376,N_13214);
nand UO_1862 (O_1862,N_14020,N_14677);
and UO_1863 (O_1863,N_14927,N_12623);
nor UO_1864 (O_1864,N_12416,N_13119);
nor UO_1865 (O_1865,N_14031,N_14167);
or UO_1866 (O_1866,N_13030,N_14609);
nand UO_1867 (O_1867,N_14226,N_14790);
nor UO_1868 (O_1868,N_13914,N_14421);
nand UO_1869 (O_1869,N_13762,N_12212);
or UO_1870 (O_1870,N_13985,N_13951);
nor UO_1871 (O_1871,N_13360,N_12224);
nor UO_1872 (O_1872,N_12795,N_13529);
nand UO_1873 (O_1873,N_14840,N_13708);
and UO_1874 (O_1874,N_14798,N_12695);
nor UO_1875 (O_1875,N_13127,N_13017);
and UO_1876 (O_1876,N_13769,N_12776);
or UO_1877 (O_1877,N_13399,N_12608);
and UO_1878 (O_1878,N_14387,N_12860);
nor UO_1879 (O_1879,N_13708,N_12972);
and UO_1880 (O_1880,N_14393,N_13484);
and UO_1881 (O_1881,N_13284,N_14498);
nor UO_1882 (O_1882,N_13788,N_13950);
nand UO_1883 (O_1883,N_13947,N_14021);
or UO_1884 (O_1884,N_12286,N_13255);
nand UO_1885 (O_1885,N_13108,N_14921);
nand UO_1886 (O_1886,N_12109,N_13758);
or UO_1887 (O_1887,N_12739,N_13557);
nor UO_1888 (O_1888,N_13125,N_14502);
or UO_1889 (O_1889,N_13414,N_14097);
and UO_1890 (O_1890,N_12761,N_12096);
nand UO_1891 (O_1891,N_13939,N_12266);
and UO_1892 (O_1892,N_14879,N_14806);
or UO_1893 (O_1893,N_14833,N_12141);
nand UO_1894 (O_1894,N_12945,N_13095);
nand UO_1895 (O_1895,N_13867,N_13777);
and UO_1896 (O_1896,N_14032,N_14204);
nand UO_1897 (O_1897,N_13738,N_12642);
nand UO_1898 (O_1898,N_14759,N_13537);
nand UO_1899 (O_1899,N_13624,N_12895);
nor UO_1900 (O_1900,N_14991,N_12075);
nor UO_1901 (O_1901,N_13636,N_12027);
nor UO_1902 (O_1902,N_14298,N_13421);
nor UO_1903 (O_1903,N_12004,N_14062);
or UO_1904 (O_1904,N_14695,N_13032);
and UO_1905 (O_1905,N_13203,N_12115);
and UO_1906 (O_1906,N_13894,N_12444);
nand UO_1907 (O_1907,N_14828,N_14856);
nand UO_1908 (O_1908,N_13781,N_12996);
and UO_1909 (O_1909,N_12984,N_13506);
nand UO_1910 (O_1910,N_14399,N_13401);
or UO_1911 (O_1911,N_13430,N_14605);
nor UO_1912 (O_1912,N_13741,N_14493);
and UO_1913 (O_1913,N_14103,N_13576);
or UO_1914 (O_1914,N_13533,N_12581);
nand UO_1915 (O_1915,N_14306,N_14566);
nor UO_1916 (O_1916,N_14482,N_13849);
or UO_1917 (O_1917,N_14219,N_14673);
nor UO_1918 (O_1918,N_13329,N_12639);
or UO_1919 (O_1919,N_12421,N_14881);
nor UO_1920 (O_1920,N_13103,N_12490);
and UO_1921 (O_1921,N_13800,N_12907);
nor UO_1922 (O_1922,N_14865,N_13459);
nand UO_1923 (O_1923,N_12682,N_13481);
nor UO_1924 (O_1924,N_13290,N_12230);
and UO_1925 (O_1925,N_13188,N_14179);
nor UO_1926 (O_1926,N_14095,N_14504);
nand UO_1927 (O_1927,N_12917,N_12118);
and UO_1928 (O_1928,N_13889,N_13626);
or UO_1929 (O_1929,N_12185,N_12906);
nand UO_1930 (O_1930,N_13996,N_13281);
nor UO_1931 (O_1931,N_14602,N_14740);
and UO_1932 (O_1932,N_14374,N_13262);
and UO_1933 (O_1933,N_14992,N_12100);
or UO_1934 (O_1934,N_14536,N_13430);
nor UO_1935 (O_1935,N_13872,N_13907);
and UO_1936 (O_1936,N_13948,N_13878);
or UO_1937 (O_1937,N_13539,N_12893);
nor UO_1938 (O_1938,N_12704,N_13128);
xor UO_1939 (O_1939,N_13741,N_12382);
or UO_1940 (O_1940,N_13236,N_14836);
and UO_1941 (O_1941,N_12709,N_14264);
or UO_1942 (O_1942,N_12524,N_14753);
nor UO_1943 (O_1943,N_12790,N_13636);
nand UO_1944 (O_1944,N_14709,N_14295);
nand UO_1945 (O_1945,N_13614,N_13965);
nand UO_1946 (O_1946,N_12229,N_13487);
nand UO_1947 (O_1947,N_14385,N_13419);
or UO_1948 (O_1948,N_12529,N_12832);
and UO_1949 (O_1949,N_12947,N_12691);
and UO_1950 (O_1950,N_12004,N_12029);
and UO_1951 (O_1951,N_14616,N_12017);
nor UO_1952 (O_1952,N_14104,N_12279);
or UO_1953 (O_1953,N_14561,N_14029);
nor UO_1954 (O_1954,N_13898,N_12438);
nand UO_1955 (O_1955,N_14440,N_14224);
and UO_1956 (O_1956,N_14811,N_14698);
and UO_1957 (O_1957,N_12723,N_12448);
nand UO_1958 (O_1958,N_13574,N_13441);
or UO_1959 (O_1959,N_12910,N_12627);
or UO_1960 (O_1960,N_14951,N_14833);
or UO_1961 (O_1961,N_12803,N_14319);
or UO_1962 (O_1962,N_13204,N_12464);
nand UO_1963 (O_1963,N_13320,N_13907);
nor UO_1964 (O_1964,N_13123,N_12718);
nand UO_1965 (O_1965,N_14174,N_13263);
and UO_1966 (O_1966,N_13055,N_14504);
nor UO_1967 (O_1967,N_14156,N_14899);
and UO_1968 (O_1968,N_13641,N_14344);
or UO_1969 (O_1969,N_13145,N_13752);
or UO_1970 (O_1970,N_12171,N_12354);
or UO_1971 (O_1971,N_12883,N_13321);
and UO_1972 (O_1972,N_14237,N_14817);
nand UO_1973 (O_1973,N_13752,N_13146);
and UO_1974 (O_1974,N_14919,N_12059);
or UO_1975 (O_1975,N_14320,N_13313);
or UO_1976 (O_1976,N_13131,N_14989);
nand UO_1977 (O_1977,N_14883,N_14790);
and UO_1978 (O_1978,N_14774,N_14852);
and UO_1979 (O_1979,N_12569,N_14761);
or UO_1980 (O_1980,N_14033,N_12436);
and UO_1981 (O_1981,N_13963,N_12463);
or UO_1982 (O_1982,N_13269,N_13251);
nand UO_1983 (O_1983,N_12693,N_14198);
nor UO_1984 (O_1984,N_13430,N_13852);
nor UO_1985 (O_1985,N_12676,N_14104);
and UO_1986 (O_1986,N_12594,N_14360);
and UO_1987 (O_1987,N_13072,N_12548);
or UO_1988 (O_1988,N_13589,N_12146);
nor UO_1989 (O_1989,N_13393,N_12373);
nor UO_1990 (O_1990,N_13084,N_13015);
and UO_1991 (O_1991,N_14654,N_12373);
nand UO_1992 (O_1992,N_12900,N_12395);
nand UO_1993 (O_1993,N_14536,N_12165);
nor UO_1994 (O_1994,N_13648,N_14120);
nor UO_1995 (O_1995,N_13179,N_13123);
or UO_1996 (O_1996,N_13981,N_12095);
nand UO_1997 (O_1997,N_14795,N_14306);
nand UO_1998 (O_1998,N_12656,N_14822);
nor UO_1999 (O_1999,N_13322,N_12509);
endmodule