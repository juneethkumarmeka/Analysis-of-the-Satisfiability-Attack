module basic_750_5000_1000_50_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_444,In_5);
or U1 (N_1,In_198,In_669);
nand U2 (N_2,In_357,In_633);
nand U3 (N_3,In_222,In_10);
nand U4 (N_4,In_91,In_156);
or U5 (N_5,In_187,In_8);
xnor U6 (N_6,In_558,In_711);
nand U7 (N_7,In_301,In_113);
and U8 (N_8,In_421,In_491);
and U9 (N_9,In_478,In_449);
nor U10 (N_10,In_404,In_583);
nor U11 (N_11,In_57,In_497);
or U12 (N_12,In_479,In_166);
nor U13 (N_13,In_721,In_487);
nand U14 (N_14,In_364,In_13);
nand U15 (N_15,In_739,In_111);
or U16 (N_16,In_33,In_426);
nand U17 (N_17,In_264,In_403);
nor U18 (N_18,In_297,In_385);
and U19 (N_19,In_212,In_471);
nand U20 (N_20,In_531,In_4);
nand U21 (N_21,In_326,In_717);
or U22 (N_22,In_622,In_293);
or U23 (N_23,In_363,In_578);
nand U24 (N_24,In_679,In_498);
xnor U25 (N_25,In_225,In_350);
and U26 (N_26,In_311,In_119);
or U27 (N_27,In_338,In_346);
nor U28 (N_28,In_96,In_109);
or U29 (N_29,In_232,In_697);
nor U30 (N_30,In_342,In_553);
and U31 (N_31,In_391,In_18);
xor U32 (N_32,In_83,In_539);
nor U33 (N_33,In_670,In_183);
or U34 (N_34,In_282,In_202);
and U35 (N_35,In_229,In_6);
or U36 (N_36,In_104,In_447);
or U37 (N_37,In_211,In_2);
or U38 (N_38,In_50,In_593);
or U39 (N_39,In_394,In_501);
or U40 (N_40,In_432,In_496);
xor U41 (N_41,In_580,In_59);
xnor U42 (N_42,In_67,In_660);
nand U43 (N_43,In_210,In_436);
or U44 (N_44,In_149,In_464);
xor U45 (N_45,In_681,In_123);
or U46 (N_46,In_528,In_493);
nor U47 (N_47,In_567,In_712);
nor U48 (N_48,In_223,In_359);
nor U49 (N_49,In_179,In_292);
xnor U50 (N_50,In_351,In_625);
or U51 (N_51,In_136,In_416);
or U52 (N_52,In_352,In_79);
nor U53 (N_53,In_549,In_554);
or U54 (N_54,In_538,In_72);
nor U55 (N_55,In_16,In_68);
nor U56 (N_56,In_275,In_741);
nand U57 (N_57,In_263,In_635);
nand U58 (N_58,In_564,In_167);
and U59 (N_59,In_683,In_269);
or U60 (N_60,In_172,In_325);
and U61 (N_61,In_298,In_81);
nand U62 (N_62,In_598,In_77);
nand U63 (N_63,In_286,In_565);
or U64 (N_64,In_268,In_406);
and U65 (N_65,In_253,In_243);
and U66 (N_66,In_695,In_398);
nand U67 (N_67,In_709,In_312);
nand U68 (N_68,In_692,In_315);
and U69 (N_69,In_361,In_500);
nor U70 (N_70,In_430,In_360);
xor U71 (N_71,In_427,In_586);
nor U72 (N_72,In_170,In_90);
and U73 (N_73,In_685,In_65);
nand U74 (N_74,In_550,In_749);
or U75 (N_75,In_551,In_373);
and U76 (N_76,In_61,In_313);
and U77 (N_77,In_3,In_488);
nand U78 (N_78,In_372,In_483);
xnor U79 (N_79,In_610,In_654);
or U80 (N_80,In_621,In_217);
xnor U81 (N_81,In_196,In_646);
and U82 (N_82,In_370,In_450);
nand U83 (N_83,In_157,In_706);
xor U84 (N_84,In_525,In_437);
nand U85 (N_85,In_134,In_45);
and U86 (N_86,In_380,In_145);
and U87 (N_87,In_469,In_51);
nand U88 (N_88,In_19,In_715);
or U89 (N_89,In_105,In_204);
and U90 (N_90,In_112,In_675);
nand U91 (N_91,In_98,In_600);
nand U92 (N_92,In_601,In_340);
nand U93 (N_93,In_589,In_146);
nor U94 (N_94,In_270,In_141);
nand U95 (N_95,In_547,In_147);
or U96 (N_96,In_566,In_285);
nand U97 (N_97,In_283,In_193);
and U98 (N_98,In_82,In_748);
nor U99 (N_99,In_429,In_594);
nor U100 (N_100,In_186,N_90);
or U101 (N_101,In_516,In_630);
or U102 (N_102,In_664,In_203);
or U103 (N_103,In_671,In_431);
or U104 (N_104,In_335,In_476);
nand U105 (N_105,In_228,In_349);
nand U106 (N_106,In_742,In_348);
and U107 (N_107,In_414,In_233);
or U108 (N_108,In_678,In_384);
xnor U109 (N_109,N_4,N_71);
or U110 (N_110,In_176,In_732);
or U111 (N_111,In_453,In_546);
xnor U112 (N_112,In_354,In_40);
and U113 (N_113,In_674,In_88);
xor U114 (N_114,In_184,In_323);
nand U115 (N_115,N_14,In_744);
nand U116 (N_116,In_468,In_728);
nor U117 (N_117,In_522,In_133);
or U118 (N_118,In_631,N_20);
and U119 (N_119,In_737,In_611);
or U120 (N_120,In_629,In_219);
nor U121 (N_121,N_64,In_543);
and U122 (N_122,In_597,In_616);
and U123 (N_123,In_255,In_462);
nor U124 (N_124,In_482,In_571);
and U125 (N_125,In_336,N_78);
xor U126 (N_126,In_129,In_287);
nor U127 (N_127,In_314,N_79);
or U128 (N_128,In_396,N_66);
nor U129 (N_129,In_53,In_648);
and U130 (N_130,In_624,In_517);
nor U131 (N_131,In_560,In_194);
nand U132 (N_132,In_209,In_238);
nor U133 (N_133,In_461,N_50);
and U134 (N_134,In_316,In_256);
and U135 (N_135,In_559,In_356);
nor U136 (N_136,In_295,N_44);
and U137 (N_137,In_262,In_634);
or U138 (N_138,In_224,In_688);
or U139 (N_139,N_3,In_389);
nor U140 (N_140,In_510,In_495);
or U141 (N_141,In_237,In_35);
nand U142 (N_142,In_87,In_169);
or U143 (N_143,In_103,In_707);
xor U144 (N_144,In_708,In_377);
nor U145 (N_145,In_653,In_513);
and U146 (N_146,N_49,In_250);
nor U147 (N_147,In_657,In_173);
and U148 (N_148,In_480,In_523);
and U149 (N_149,N_13,In_667);
and U150 (N_150,In_647,In_192);
nand U151 (N_151,In_661,N_33);
xnor U152 (N_152,In_317,N_40);
or U153 (N_153,N_21,In_216);
or U154 (N_154,In_613,In_278);
xnor U155 (N_155,In_30,N_23);
nor U156 (N_156,In_602,N_38);
nor U157 (N_157,In_620,In_175);
nor U158 (N_158,In_46,In_490);
and U159 (N_159,In_177,In_422);
nor U160 (N_160,In_591,In_445);
nor U161 (N_161,In_642,In_365);
xor U162 (N_162,In_376,N_89);
or U163 (N_163,In_249,N_87);
nand U164 (N_164,In_727,In_582);
xor U165 (N_165,In_595,In_443);
or U166 (N_166,In_254,N_12);
nor U167 (N_167,In_636,In_439);
nor U168 (N_168,In_321,In_623);
nor U169 (N_169,In_509,In_64);
nand U170 (N_170,In_698,In_310);
nand U171 (N_171,N_94,In_322);
and U172 (N_172,In_617,In_502);
nand U173 (N_173,In_694,In_180);
or U174 (N_174,In_526,In_411);
and U175 (N_175,In_608,In_44);
nor U176 (N_176,In_399,In_56);
and U177 (N_177,In_66,In_54);
or U178 (N_178,In_682,In_85);
xnor U179 (N_179,In_368,In_58);
xnor U180 (N_180,N_68,In_279);
nor U181 (N_181,In_171,In_723);
nor U182 (N_182,In_542,In_457);
nor U183 (N_183,In_652,In_734);
or U184 (N_184,In_703,N_6);
nor U185 (N_185,N_0,In_402);
nand U186 (N_186,In_120,In_719);
nand U187 (N_187,In_208,In_21);
nor U188 (N_188,In_131,In_231);
xor U189 (N_189,In_484,In_252);
and U190 (N_190,In_168,In_151);
nor U191 (N_191,In_726,N_41);
nor U192 (N_192,In_75,In_668);
nor U193 (N_193,In_590,In_691);
nor U194 (N_194,In_561,In_390);
nor U195 (N_195,N_55,In_11);
nand U196 (N_196,In_334,N_70);
or U197 (N_197,In_158,N_39);
nor U198 (N_198,In_215,In_304);
and U199 (N_199,In_410,In_693);
nand U200 (N_200,In_29,In_424);
nand U201 (N_201,In_672,N_74);
xor U202 (N_202,In_115,In_62);
nand U203 (N_203,In_596,N_176);
nor U204 (N_204,In_435,N_84);
nand U205 (N_205,N_166,In_200);
or U206 (N_206,N_24,In_201);
xor U207 (N_207,In_433,In_506);
nor U208 (N_208,In_143,In_26);
nor U209 (N_209,In_614,N_143);
and U210 (N_210,In_25,N_54);
nor U211 (N_211,In_94,N_125);
xor U212 (N_212,In_665,In_277);
or U213 (N_213,In_1,In_419);
and U214 (N_214,In_508,In_230);
xnor U215 (N_215,In_533,In_154);
and U216 (N_216,N_30,In_440);
or U217 (N_217,N_159,N_7);
or U218 (N_218,In_673,In_24);
nor U219 (N_219,In_52,In_745);
nand U220 (N_220,In_632,In_327);
or U221 (N_221,In_540,In_442);
xor U222 (N_222,N_93,In_366);
xnor U223 (N_223,In_274,In_100);
or U224 (N_224,N_174,In_235);
nand U225 (N_225,N_56,In_165);
nor U226 (N_226,In_246,In_704);
nor U227 (N_227,N_27,N_8);
and U228 (N_228,In_102,In_213);
or U229 (N_229,N_152,In_343);
nand U230 (N_230,N_173,In_272);
nand U231 (N_231,N_17,N_10);
nand U232 (N_232,In_574,N_63);
xnor U233 (N_233,N_182,In_556);
and U234 (N_234,N_58,N_164);
or U235 (N_235,In_418,In_248);
or U236 (N_236,In_353,In_573);
nor U237 (N_237,N_113,N_116);
or U238 (N_238,N_198,In_530);
and U239 (N_239,In_375,In_126);
or U240 (N_240,In_150,N_161);
nand U241 (N_241,In_36,In_226);
nor U242 (N_242,In_73,N_60);
nor U243 (N_243,In_362,In_687);
nand U244 (N_244,In_161,N_150);
and U245 (N_245,N_83,N_65);
and U246 (N_246,In_740,N_193);
or U247 (N_247,N_148,In_266);
nor U248 (N_248,In_512,N_28);
nand U249 (N_249,In_409,N_121);
and U250 (N_250,N_1,In_320);
nand U251 (N_251,N_137,In_515);
and U252 (N_252,N_130,In_618);
and U253 (N_253,N_31,In_722);
nor U254 (N_254,In_662,In_541);
nand U255 (N_255,In_460,In_345);
xnor U256 (N_256,In_641,In_358);
and U257 (N_257,In_446,N_175);
nand U258 (N_258,In_412,In_178);
or U259 (N_259,N_99,In_23);
xor U260 (N_260,In_155,In_197);
nand U261 (N_261,In_643,In_650);
nor U262 (N_262,In_452,In_288);
nor U263 (N_263,In_455,N_73);
nand U264 (N_264,N_168,In_257);
nand U265 (N_265,In_78,In_122);
or U266 (N_266,In_273,In_428);
xnor U267 (N_267,N_188,In_140);
or U268 (N_268,N_46,N_131);
or U269 (N_269,N_67,In_536);
xnor U270 (N_270,N_62,In_441);
and U271 (N_271,N_189,In_381);
and U272 (N_272,In_684,In_729);
or U273 (N_273,In_276,In_645);
nand U274 (N_274,In_63,N_172);
nand U275 (N_275,In_388,In_92);
or U276 (N_276,N_11,N_104);
xor U277 (N_277,In_110,In_520);
or U278 (N_278,N_157,N_163);
and U279 (N_279,N_158,In_333);
and U280 (N_280,In_9,N_140);
nor U281 (N_281,In_392,N_147);
nor U282 (N_282,In_400,In_413);
xor U283 (N_283,In_537,In_12);
or U284 (N_284,In_107,N_97);
nor U285 (N_285,In_655,In_47);
and U286 (N_286,In_332,In_330);
nor U287 (N_287,N_43,In_505);
or U288 (N_288,In_355,In_236);
nor U289 (N_289,In_367,In_55);
and U290 (N_290,N_98,In_474);
nor U291 (N_291,N_77,In_481);
nand U292 (N_292,N_88,In_639);
nand U293 (N_293,In_477,In_463);
nand U294 (N_294,N_96,In_651);
nand U295 (N_295,N_91,In_20);
nor U296 (N_296,In_747,In_746);
or U297 (N_297,In_579,In_182);
or U298 (N_298,In_534,In_41);
nor U299 (N_299,In_383,N_105);
nor U300 (N_300,In_341,In_604);
and U301 (N_301,N_254,In_736);
and U302 (N_302,In_369,In_318);
and U303 (N_303,In_307,In_291);
nand U304 (N_304,In_148,In_80);
nor U305 (N_305,In_659,In_244);
nor U306 (N_306,In_290,In_206);
nor U307 (N_307,N_128,In_569);
and U308 (N_308,In_101,N_32);
nand U309 (N_309,In_118,N_253);
or U310 (N_310,N_76,N_248);
nand U311 (N_311,N_236,N_120);
or U312 (N_312,In_117,N_34);
or U313 (N_313,N_103,N_151);
nor U314 (N_314,In_267,N_149);
nand U315 (N_315,In_308,In_174);
xnor U316 (N_316,In_329,N_235);
xor U317 (N_317,N_255,In_397);
nand U318 (N_318,N_246,In_240);
and U319 (N_319,In_34,In_401);
and U320 (N_320,In_227,N_153);
or U321 (N_321,In_371,In_135);
nor U322 (N_322,In_185,N_106);
and U323 (N_323,N_252,N_115);
nor U324 (N_324,In_420,N_299);
xnor U325 (N_325,N_244,N_112);
nand U326 (N_326,In_640,N_256);
and U327 (N_327,N_271,In_296);
nor U328 (N_328,In_378,N_234);
and U329 (N_329,In_699,N_129);
nor U330 (N_330,In_705,In_710);
and U331 (N_331,In_76,N_126);
nor U332 (N_332,N_281,In_572);
nand U333 (N_333,N_192,N_75);
nor U334 (N_334,N_197,N_25);
nand U335 (N_335,In_504,In_486);
and U336 (N_336,In_241,In_162);
nor U337 (N_337,In_666,In_22);
nand U338 (N_338,N_211,N_225);
or U339 (N_339,N_177,In_163);
nor U340 (N_340,N_293,In_423);
and U341 (N_341,In_407,In_570);
and U342 (N_342,N_82,In_69);
and U343 (N_343,In_199,In_557);
nor U344 (N_344,In_607,In_568);
nand U345 (N_345,In_294,N_218);
nor U346 (N_346,In_448,N_204);
nor U347 (N_347,In_507,N_290);
nand U348 (N_348,In_37,N_134);
nor U349 (N_349,In_221,In_575);
nor U350 (N_350,N_260,In_686);
nor U351 (N_351,In_511,N_107);
nor U352 (N_352,In_27,In_124);
nor U353 (N_353,In_139,In_408);
nand U354 (N_354,In_218,N_238);
nor U355 (N_355,In_289,N_187);
nor U356 (N_356,In_615,N_51);
nor U357 (N_357,N_224,N_35);
nand U358 (N_358,In_48,N_216);
or U359 (N_359,N_250,N_274);
or U360 (N_360,N_29,N_111);
and U361 (N_361,In_544,In_458);
or U362 (N_362,In_95,In_470);
or U363 (N_363,N_266,N_279);
and U364 (N_364,In_106,N_286);
and U365 (N_365,In_456,In_114);
xnor U366 (N_366,In_271,In_130);
nor U367 (N_367,In_676,N_285);
nand U368 (N_368,In_555,N_57);
and U369 (N_369,In_585,In_663);
nand U370 (N_370,In_499,In_328);
or U371 (N_371,In_245,In_205);
nand U372 (N_372,In_160,In_720);
nor U373 (N_373,In_121,In_306);
and U374 (N_374,N_95,In_612);
nor U375 (N_375,N_206,N_242);
xor U376 (N_376,N_270,N_102);
or U377 (N_377,In_14,N_208);
or U378 (N_378,In_84,In_303);
nor U379 (N_379,N_142,N_9);
nor U380 (N_380,In_39,N_85);
nand U381 (N_381,In_716,In_638);
nor U382 (N_382,N_280,N_283);
nand U383 (N_383,N_296,N_222);
or U384 (N_384,In_284,N_139);
or U385 (N_385,In_626,In_300);
nor U386 (N_386,N_146,In_637);
nor U387 (N_387,N_2,N_212);
nor U388 (N_388,N_47,In_552);
or U389 (N_389,In_535,N_196);
xnor U390 (N_390,N_22,N_184);
nor U391 (N_391,In_195,N_213);
nor U392 (N_392,In_337,N_291);
and U393 (N_393,N_264,N_243);
or U394 (N_394,In_563,N_167);
and U395 (N_395,N_36,In_714);
nor U396 (N_396,In_592,In_503);
nor U397 (N_397,In_309,N_179);
and U398 (N_398,In_207,In_31);
nor U399 (N_399,In_239,In_189);
xor U400 (N_400,N_165,N_289);
or U401 (N_401,In_319,N_295);
or U402 (N_402,N_326,In_93);
xor U403 (N_403,In_628,In_127);
and U404 (N_404,In_188,N_101);
and U405 (N_405,In_649,N_292);
nand U406 (N_406,N_348,N_277);
and U407 (N_407,N_346,N_298);
or U408 (N_408,N_186,In_32);
or U409 (N_409,N_203,N_393);
or U410 (N_410,In_475,N_169);
and U411 (N_411,N_114,In_17);
xnor U412 (N_412,N_180,In_302);
and U413 (N_413,N_259,N_19);
nand U414 (N_414,N_261,N_344);
or U415 (N_415,In_28,N_132);
or U416 (N_416,N_275,N_338);
or U417 (N_417,N_162,N_265);
and U418 (N_418,N_219,In_42);
nor U419 (N_419,In_609,N_372);
nor U420 (N_420,In_344,N_92);
or U421 (N_421,In_339,N_358);
nor U422 (N_422,N_200,In_576);
and U423 (N_423,N_118,N_145);
and U424 (N_424,N_233,N_315);
nor U425 (N_425,N_217,N_313);
or U426 (N_426,N_267,In_153);
or U427 (N_427,N_359,N_321);
or U428 (N_428,N_319,N_377);
or U429 (N_429,N_170,N_389);
nor U430 (N_430,N_122,N_127);
or U431 (N_431,N_154,N_310);
nor U432 (N_432,N_136,N_317);
and U433 (N_433,In_724,N_61);
and U434 (N_434,N_302,N_343);
or U435 (N_435,In_718,N_201);
and U436 (N_436,N_397,In_467);
or U437 (N_437,In_191,In_374);
or U438 (N_438,In_690,N_347);
nand U439 (N_439,N_386,In_472);
nor U440 (N_440,N_373,N_272);
nor U441 (N_441,N_303,N_245);
and U442 (N_442,N_330,In_379);
nor U443 (N_443,In_459,In_70);
or U444 (N_444,N_383,N_144);
nor U445 (N_445,N_396,N_350);
or U446 (N_446,In_425,N_325);
or U447 (N_447,N_374,In_138);
nand U448 (N_448,In_7,In_548);
xnor U449 (N_449,In_545,N_138);
nand U450 (N_450,N_185,N_297);
nor U451 (N_451,N_220,In_730);
nand U452 (N_452,N_191,N_288);
nand U453 (N_453,N_205,N_306);
and U454 (N_454,In_214,In_128);
nor U455 (N_455,N_356,N_160);
nor U456 (N_456,N_229,N_376);
nand U457 (N_457,In_524,N_353);
and U458 (N_458,N_382,N_391);
or U459 (N_459,N_141,N_327);
nand U460 (N_460,N_135,N_183);
nor U461 (N_461,N_388,N_309);
or U462 (N_462,N_379,N_156);
nand U463 (N_463,In_700,In_387);
or U464 (N_464,N_332,N_215);
nand U465 (N_465,N_394,In_599);
nand U466 (N_466,In_696,N_133);
or U467 (N_467,In_605,In_242);
and U468 (N_468,N_333,In_99);
or U469 (N_469,N_80,N_199);
nand U470 (N_470,In_680,N_37);
or U471 (N_471,N_392,N_155);
or U472 (N_472,In_466,N_53);
nor U473 (N_473,N_278,In_281);
or U474 (N_474,N_282,In_247);
nand U475 (N_475,In_71,N_69);
nand U476 (N_476,In_725,N_375);
or U477 (N_477,In_393,In_331);
xnor U478 (N_478,N_45,N_378);
and U479 (N_479,In_116,N_307);
and U480 (N_480,In_587,N_354);
or U481 (N_481,N_247,N_171);
xor U482 (N_482,In_43,In_518);
or U483 (N_483,N_119,In_164);
and U484 (N_484,In_438,N_249);
nand U485 (N_485,In_485,In_382);
nor U486 (N_486,N_294,In_689);
nor U487 (N_487,N_380,N_370);
or U488 (N_488,In_415,N_258);
nor U489 (N_489,In_86,In_190);
or U490 (N_490,In_713,In_644);
nor U491 (N_491,In_743,N_381);
or U492 (N_492,N_52,In_261);
and U493 (N_493,In_137,In_454);
or U494 (N_494,N_322,N_334);
or U495 (N_495,N_305,In_144);
or U496 (N_496,In_280,N_231);
xnor U497 (N_497,N_124,N_385);
and U498 (N_498,In_562,N_340);
or U499 (N_499,In_529,N_110);
nand U500 (N_500,N_194,N_18);
and U501 (N_501,N_455,N_329);
or U502 (N_502,In_142,N_427);
or U503 (N_503,N_485,N_335);
and U504 (N_504,N_223,In_265);
nand U505 (N_505,N_365,N_403);
nand U506 (N_506,In_152,N_357);
and U507 (N_507,N_390,In_619);
nor U508 (N_508,In_132,N_466);
nand U509 (N_509,N_437,In_606);
nor U510 (N_510,N_367,In_627);
nor U511 (N_511,In_489,In_514);
nand U512 (N_512,In_0,N_411);
nor U513 (N_513,N_262,N_445);
or U514 (N_514,N_237,In_581);
and U515 (N_515,N_489,N_472);
and U516 (N_516,In_656,In_735);
or U517 (N_517,In_738,N_263);
nor U518 (N_518,N_227,N_457);
or U519 (N_519,N_123,In_519);
or U520 (N_520,In_60,N_408);
and U521 (N_521,N_498,In_434);
nor U522 (N_522,In_49,N_331);
or U523 (N_523,N_434,N_463);
and U524 (N_524,N_412,N_371);
nor U525 (N_525,N_473,In_473);
nor U526 (N_526,N_304,N_475);
nor U527 (N_527,N_5,In_658);
nand U528 (N_528,N_478,N_456);
and U529 (N_529,N_482,N_465);
xor U530 (N_530,N_349,In_305);
or U531 (N_531,N_207,In_38);
nand U532 (N_532,N_494,In_299);
xnor U533 (N_533,N_496,N_178);
and U534 (N_534,N_487,N_405);
or U535 (N_535,N_251,N_492);
nand U536 (N_536,In_74,N_341);
nand U537 (N_537,In_15,N_469);
nor U538 (N_538,In_733,N_461);
or U539 (N_539,N_479,N_312);
and U540 (N_540,N_195,N_490);
and U541 (N_541,N_301,N_459);
nand U542 (N_542,N_352,In_577);
or U543 (N_543,N_424,N_241);
nand U544 (N_544,N_59,N_410);
and U545 (N_545,In_677,N_439);
nand U546 (N_546,N_477,N_48);
nand U547 (N_547,N_276,N_15);
nor U548 (N_548,N_433,N_407);
and U549 (N_549,N_499,N_230);
and U550 (N_550,N_426,N_273);
nand U551 (N_551,In_731,N_399);
xor U552 (N_552,N_351,N_423);
and U553 (N_553,N_484,N_414);
nand U554 (N_554,N_474,N_429);
nor U555 (N_555,N_226,N_368);
xor U556 (N_556,N_460,N_324);
nor U557 (N_557,N_109,N_404);
nor U558 (N_558,In_260,In_258);
nor U559 (N_559,N_384,N_453);
and U560 (N_560,N_395,In_386);
and U561 (N_561,N_181,N_432);
or U562 (N_562,N_117,N_240);
and U563 (N_563,N_428,N_257);
nand U564 (N_564,N_311,N_467);
or U565 (N_565,N_318,N_476);
or U566 (N_566,N_214,N_443);
and U567 (N_567,N_269,N_361);
nand U568 (N_568,In_347,N_232);
nand U569 (N_569,In_395,N_430);
nand U570 (N_570,In_220,In_465);
xor U571 (N_571,N_398,In_527);
or U572 (N_572,N_416,In_417);
nand U573 (N_573,In_125,N_316);
nand U574 (N_574,N_300,N_406);
nand U575 (N_575,N_284,N_421);
nand U576 (N_576,N_464,N_336);
or U577 (N_577,N_450,N_228);
nand U578 (N_578,In_159,In_108);
xnor U579 (N_579,N_314,N_337);
and U580 (N_580,N_417,In_701);
nor U581 (N_581,In_494,N_100);
nand U582 (N_582,N_442,N_42);
or U583 (N_583,N_449,In_234);
nor U584 (N_584,N_420,N_446);
and U585 (N_585,N_328,N_355);
nand U586 (N_586,In_251,N_454);
and U587 (N_587,N_422,N_468);
nor U588 (N_588,N_108,N_483);
or U589 (N_589,N_413,N_491);
or U590 (N_590,In_521,N_221);
xnor U591 (N_591,N_497,N_441);
nand U592 (N_592,N_488,N_480);
or U593 (N_593,N_308,N_409);
nor U594 (N_594,N_440,N_447);
nand U595 (N_595,N_425,N_209);
nor U596 (N_596,N_400,N_26);
nor U597 (N_597,In_603,N_452);
or U598 (N_598,N_345,N_495);
nand U599 (N_599,N_239,N_486);
and U600 (N_600,N_540,N_320);
nand U601 (N_601,N_503,N_16);
nor U602 (N_602,N_431,N_593);
or U603 (N_603,N_598,N_526);
nand U604 (N_604,N_587,N_507);
nor U605 (N_605,In_324,N_462);
xnor U606 (N_606,N_86,N_592);
or U607 (N_607,In_492,N_551);
or U608 (N_608,N_547,N_501);
or U609 (N_609,N_578,N_550);
or U610 (N_610,N_518,In_181);
or U611 (N_611,In_584,N_202);
and U612 (N_612,N_590,N_585);
or U613 (N_613,N_504,N_596);
and U614 (N_614,N_435,In_588);
nor U615 (N_615,N_506,N_519);
nand U616 (N_616,N_562,N_567);
nand U617 (N_617,N_402,N_584);
and U618 (N_618,N_510,N_438);
xor U619 (N_619,N_522,N_529);
nor U620 (N_620,N_493,N_500);
or U621 (N_621,N_508,N_287);
nor U622 (N_622,N_401,N_520);
nand U623 (N_623,N_533,N_339);
nand U624 (N_624,N_555,In_405);
nor U625 (N_625,N_514,N_444);
and U626 (N_626,N_458,N_538);
nor U627 (N_627,N_512,N_470);
nor U628 (N_628,N_419,N_72);
or U629 (N_629,N_471,N_536);
and U630 (N_630,N_436,N_570);
nor U631 (N_631,N_481,N_505);
or U632 (N_632,N_268,N_556);
and U633 (N_633,N_366,N_535);
xor U634 (N_634,N_586,In_532);
nand U635 (N_635,N_559,N_582);
nand U636 (N_636,N_580,N_594);
or U637 (N_637,N_565,N_581);
nor U638 (N_638,N_560,N_577);
and U639 (N_639,N_553,N_528);
nor U640 (N_640,N_568,N_525);
nor U641 (N_641,In_259,N_588);
or U642 (N_642,N_571,In_702);
nor U643 (N_643,N_546,In_97);
or U644 (N_644,N_564,N_210);
xor U645 (N_645,N_591,N_574);
xor U646 (N_646,N_524,N_502);
nor U647 (N_647,N_563,N_599);
or U648 (N_648,N_342,N_575);
nand U649 (N_649,N_369,N_539);
nand U650 (N_650,N_589,N_448);
nand U651 (N_651,N_521,N_418);
or U652 (N_652,N_573,N_572);
nor U653 (N_653,N_415,N_323);
and U654 (N_654,N_541,In_451);
nor U655 (N_655,In_89,N_523);
and U656 (N_656,N_579,N_549);
and U657 (N_657,N_576,N_558);
or U658 (N_658,N_360,N_561);
xor U659 (N_659,N_517,N_516);
nand U660 (N_660,N_544,N_534);
nor U661 (N_661,N_511,N_552);
nor U662 (N_662,N_513,N_509);
or U663 (N_663,N_81,N_543);
or U664 (N_664,N_569,N_515);
and U665 (N_665,N_530,N_537);
nor U666 (N_666,N_542,N_364);
nor U667 (N_667,N_362,N_595);
and U668 (N_668,N_554,N_387);
and U669 (N_669,N_597,N_566);
xor U670 (N_670,N_583,N_190);
or U671 (N_671,N_531,N_363);
or U672 (N_672,N_557,N_451);
or U673 (N_673,N_532,N_548);
nor U674 (N_674,N_527,N_545);
or U675 (N_675,N_532,N_573);
and U676 (N_676,N_521,N_520);
nand U677 (N_677,N_500,N_517);
xnor U678 (N_678,N_552,N_16);
and U679 (N_679,N_571,In_181);
xor U680 (N_680,N_536,In_181);
nand U681 (N_681,N_500,N_588);
nor U682 (N_682,N_529,N_16);
nand U683 (N_683,N_493,N_530);
nand U684 (N_684,In_451,N_505);
nand U685 (N_685,N_557,N_401);
nand U686 (N_686,In_702,N_547);
or U687 (N_687,N_190,N_562);
and U688 (N_688,N_542,N_401);
nor U689 (N_689,N_578,N_544);
nor U690 (N_690,N_558,In_588);
and U691 (N_691,N_591,N_514);
or U692 (N_692,N_543,N_549);
nand U693 (N_693,N_521,N_545);
nand U694 (N_694,N_481,N_526);
or U695 (N_695,N_586,N_585);
nand U696 (N_696,N_567,N_580);
nor U697 (N_697,N_584,N_543);
nand U698 (N_698,N_514,N_508);
nand U699 (N_699,N_548,N_567);
or U700 (N_700,N_688,N_697);
xor U701 (N_701,N_689,N_676);
nand U702 (N_702,N_687,N_629);
xnor U703 (N_703,N_699,N_661);
and U704 (N_704,N_628,N_655);
or U705 (N_705,N_694,N_634);
nand U706 (N_706,N_601,N_645);
and U707 (N_707,N_671,N_633);
nor U708 (N_708,N_632,N_622);
nor U709 (N_709,N_635,N_624);
nor U710 (N_710,N_693,N_620);
nor U711 (N_711,N_643,N_684);
nor U712 (N_712,N_658,N_659);
and U713 (N_713,N_617,N_642);
and U714 (N_714,N_611,N_641);
and U715 (N_715,N_683,N_623);
and U716 (N_716,N_606,N_652);
and U717 (N_717,N_660,N_657);
or U718 (N_718,N_662,N_626);
nand U719 (N_719,N_609,N_682);
nand U720 (N_720,N_648,N_610);
nand U721 (N_721,N_672,N_696);
nand U722 (N_722,N_603,N_667);
or U723 (N_723,N_680,N_690);
nor U724 (N_724,N_686,N_646);
or U725 (N_725,N_668,N_612);
or U726 (N_726,N_621,N_625);
nor U727 (N_727,N_638,N_637);
nand U728 (N_728,N_644,N_630);
and U729 (N_729,N_651,N_607);
or U730 (N_730,N_631,N_669);
nor U731 (N_731,N_677,N_679);
xor U732 (N_732,N_600,N_608);
nand U733 (N_733,N_692,N_698);
or U734 (N_734,N_618,N_616);
nor U735 (N_735,N_604,N_670);
nor U736 (N_736,N_614,N_605);
xnor U737 (N_737,N_673,N_678);
and U738 (N_738,N_639,N_619);
and U739 (N_739,N_649,N_650);
nand U740 (N_740,N_654,N_685);
and U741 (N_741,N_656,N_681);
nor U742 (N_742,N_627,N_695);
xor U743 (N_743,N_602,N_675);
and U744 (N_744,N_653,N_665);
and U745 (N_745,N_640,N_691);
nand U746 (N_746,N_613,N_663);
and U747 (N_747,N_666,N_674);
nand U748 (N_748,N_636,N_664);
or U749 (N_749,N_647,N_615);
nand U750 (N_750,N_651,N_660);
nand U751 (N_751,N_611,N_668);
nor U752 (N_752,N_697,N_660);
xor U753 (N_753,N_653,N_641);
xor U754 (N_754,N_600,N_643);
or U755 (N_755,N_692,N_632);
and U756 (N_756,N_692,N_676);
nor U757 (N_757,N_690,N_642);
or U758 (N_758,N_661,N_682);
or U759 (N_759,N_693,N_616);
nand U760 (N_760,N_621,N_672);
nor U761 (N_761,N_634,N_628);
and U762 (N_762,N_653,N_602);
and U763 (N_763,N_692,N_685);
nor U764 (N_764,N_610,N_625);
nand U765 (N_765,N_605,N_672);
and U766 (N_766,N_694,N_652);
or U767 (N_767,N_634,N_667);
or U768 (N_768,N_673,N_666);
and U769 (N_769,N_682,N_611);
nor U770 (N_770,N_603,N_635);
and U771 (N_771,N_649,N_640);
nor U772 (N_772,N_668,N_633);
nor U773 (N_773,N_601,N_659);
nor U774 (N_774,N_621,N_612);
xor U775 (N_775,N_668,N_665);
nor U776 (N_776,N_639,N_686);
and U777 (N_777,N_665,N_618);
or U778 (N_778,N_643,N_697);
xor U779 (N_779,N_674,N_617);
nand U780 (N_780,N_633,N_693);
or U781 (N_781,N_608,N_650);
nor U782 (N_782,N_625,N_605);
nand U783 (N_783,N_630,N_609);
and U784 (N_784,N_603,N_600);
and U785 (N_785,N_661,N_678);
nand U786 (N_786,N_698,N_664);
and U787 (N_787,N_696,N_637);
or U788 (N_788,N_644,N_639);
nor U789 (N_789,N_629,N_685);
xnor U790 (N_790,N_671,N_626);
nand U791 (N_791,N_600,N_627);
or U792 (N_792,N_629,N_611);
nor U793 (N_793,N_673,N_604);
nand U794 (N_794,N_671,N_690);
nand U795 (N_795,N_614,N_688);
xnor U796 (N_796,N_673,N_647);
nor U797 (N_797,N_683,N_639);
nand U798 (N_798,N_698,N_616);
and U799 (N_799,N_670,N_600);
nor U800 (N_800,N_767,N_770);
nor U801 (N_801,N_753,N_702);
and U802 (N_802,N_748,N_766);
or U803 (N_803,N_788,N_785);
or U804 (N_804,N_738,N_731);
nand U805 (N_805,N_722,N_745);
nor U806 (N_806,N_713,N_741);
or U807 (N_807,N_782,N_790);
and U808 (N_808,N_720,N_740);
or U809 (N_809,N_726,N_776);
nor U810 (N_810,N_715,N_794);
and U811 (N_811,N_708,N_796);
and U812 (N_812,N_727,N_742);
or U813 (N_813,N_771,N_709);
and U814 (N_814,N_746,N_732);
or U815 (N_815,N_778,N_755);
or U816 (N_816,N_749,N_779);
and U817 (N_817,N_798,N_700);
nand U818 (N_818,N_735,N_799);
or U819 (N_819,N_780,N_758);
nor U820 (N_820,N_723,N_712);
and U821 (N_821,N_764,N_774);
nor U822 (N_822,N_724,N_772);
and U823 (N_823,N_707,N_734);
nand U824 (N_824,N_759,N_705);
nand U825 (N_825,N_730,N_791);
nand U826 (N_826,N_717,N_714);
nand U827 (N_827,N_718,N_769);
or U828 (N_828,N_793,N_789);
xnor U829 (N_829,N_721,N_737);
nand U830 (N_830,N_761,N_773);
or U831 (N_831,N_752,N_728);
nand U832 (N_832,N_765,N_725);
and U833 (N_833,N_750,N_763);
and U834 (N_834,N_795,N_775);
or U835 (N_835,N_736,N_797);
or U836 (N_836,N_751,N_703);
nor U837 (N_837,N_760,N_792);
or U838 (N_838,N_747,N_756);
nand U839 (N_839,N_719,N_743);
nor U840 (N_840,N_710,N_706);
nor U841 (N_841,N_744,N_757);
or U842 (N_842,N_786,N_781);
nor U843 (N_843,N_704,N_783);
and U844 (N_844,N_701,N_768);
nor U845 (N_845,N_762,N_739);
and U846 (N_846,N_777,N_729);
xnor U847 (N_847,N_787,N_733);
nand U848 (N_848,N_784,N_716);
nor U849 (N_849,N_711,N_754);
or U850 (N_850,N_740,N_753);
or U851 (N_851,N_799,N_781);
and U852 (N_852,N_704,N_745);
nor U853 (N_853,N_701,N_762);
xnor U854 (N_854,N_790,N_747);
and U855 (N_855,N_729,N_753);
nand U856 (N_856,N_707,N_709);
or U857 (N_857,N_753,N_723);
or U858 (N_858,N_767,N_766);
nand U859 (N_859,N_770,N_772);
nor U860 (N_860,N_709,N_780);
or U861 (N_861,N_719,N_773);
and U862 (N_862,N_710,N_753);
nor U863 (N_863,N_751,N_720);
and U864 (N_864,N_700,N_727);
and U865 (N_865,N_736,N_786);
and U866 (N_866,N_709,N_708);
nor U867 (N_867,N_703,N_706);
nand U868 (N_868,N_705,N_764);
nor U869 (N_869,N_708,N_731);
or U870 (N_870,N_747,N_788);
and U871 (N_871,N_760,N_708);
and U872 (N_872,N_773,N_727);
and U873 (N_873,N_707,N_745);
and U874 (N_874,N_709,N_785);
nor U875 (N_875,N_702,N_782);
nor U876 (N_876,N_777,N_792);
xnor U877 (N_877,N_793,N_770);
nor U878 (N_878,N_767,N_704);
and U879 (N_879,N_758,N_713);
nor U880 (N_880,N_750,N_701);
or U881 (N_881,N_761,N_784);
nand U882 (N_882,N_776,N_717);
and U883 (N_883,N_746,N_762);
nand U884 (N_884,N_781,N_710);
or U885 (N_885,N_721,N_770);
nor U886 (N_886,N_791,N_760);
nand U887 (N_887,N_758,N_741);
or U888 (N_888,N_766,N_712);
nand U889 (N_889,N_743,N_705);
xnor U890 (N_890,N_715,N_726);
nor U891 (N_891,N_756,N_719);
nor U892 (N_892,N_741,N_772);
nor U893 (N_893,N_707,N_712);
and U894 (N_894,N_758,N_717);
and U895 (N_895,N_786,N_767);
and U896 (N_896,N_716,N_770);
nor U897 (N_897,N_731,N_786);
xnor U898 (N_898,N_720,N_744);
nor U899 (N_899,N_719,N_738);
or U900 (N_900,N_893,N_812);
nand U901 (N_901,N_890,N_881);
and U902 (N_902,N_800,N_838);
and U903 (N_903,N_877,N_804);
or U904 (N_904,N_841,N_847);
or U905 (N_905,N_818,N_823);
and U906 (N_906,N_851,N_832);
xnor U907 (N_907,N_822,N_856);
nor U908 (N_908,N_892,N_882);
xnor U909 (N_909,N_839,N_858);
or U910 (N_910,N_867,N_855);
nor U911 (N_911,N_869,N_883);
and U912 (N_912,N_844,N_816);
and U913 (N_913,N_854,N_828);
or U914 (N_914,N_850,N_891);
nand U915 (N_915,N_808,N_888);
nor U916 (N_916,N_885,N_821);
or U917 (N_917,N_860,N_861);
nor U918 (N_918,N_807,N_866);
or U919 (N_919,N_842,N_899);
nor U920 (N_920,N_889,N_837);
nand U921 (N_921,N_805,N_825);
nand U922 (N_922,N_829,N_873);
and U923 (N_923,N_886,N_814);
or U924 (N_924,N_896,N_843);
nor U925 (N_925,N_874,N_879);
nand U926 (N_926,N_831,N_806);
or U927 (N_927,N_863,N_817);
or U928 (N_928,N_826,N_801);
nand U929 (N_929,N_864,N_849);
or U930 (N_930,N_834,N_853);
or U931 (N_931,N_884,N_833);
nor U932 (N_932,N_809,N_830);
xnor U933 (N_933,N_845,N_871);
or U934 (N_934,N_875,N_887);
or U935 (N_935,N_811,N_870);
and U936 (N_936,N_824,N_848);
xor U937 (N_937,N_803,N_880);
and U938 (N_938,N_810,N_813);
nor U939 (N_939,N_857,N_868);
nor U940 (N_940,N_872,N_876);
xnor U941 (N_941,N_835,N_897);
nand U942 (N_942,N_878,N_836);
and U943 (N_943,N_859,N_840);
or U944 (N_944,N_895,N_894);
and U945 (N_945,N_819,N_846);
nor U946 (N_946,N_898,N_865);
xnor U947 (N_947,N_820,N_827);
nand U948 (N_948,N_862,N_815);
nand U949 (N_949,N_852,N_802);
nand U950 (N_950,N_850,N_861);
and U951 (N_951,N_801,N_844);
or U952 (N_952,N_832,N_896);
nor U953 (N_953,N_814,N_807);
or U954 (N_954,N_899,N_817);
and U955 (N_955,N_804,N_808);
nand U956 (N_956,N_835,N_855);
nor U957 (N_957,N_804,N_820);
xnor U958 (N_958,N_866,N_881);
xnor U959 (N_959,N_860,N_826);
and U960 (N_960,N_816,N_866);
nand U961 (N_961,N_802,N_849);
xor U962 (N_962,N_850,N_875);
or U963 (N_963,N_867,N_841);
nand U964 (N_964,N_828,N_837);
nand U965 (N_965,N_818,N_805);
nand U966 (N_966,N_814,N_834);
and U967 (N_967,N_851,N_810);
or U968 (N_968,N_890,N_800);
or U969 (N_969,N_820,N_825);
nand U970 (N_970,N_824,N_853);
nor U971 (N_971,N_827,N_886);
nor U972 (N_972,N_819,N_886);
or U973 (N_973,N_874,N_831);
nand U974 (N_974,N_884,N_816);
and U975 (N_975,N_869,N_836);
and U976 (N_976,N_850,N_800);
xnor U977 (N_977,N_893,N_898);
xnor U978 (N_978,N_860,N_802);
and U979 (N_979,N_875,N_855);
or U980 (N_980,N_892,N_858);
or U981 (N_981,N_863,N_839);
and U982 (N_982,N_873,N_850);
or U983 (N_983,N_813,N_856);
nand U984 (N_984,N_838,N_896);
and U985 (N_985,N_819,N_884);
nor U986 (N_986,N_819,N_812);
and U987 (N_987,N_823,N_822);
nor U988 (N_988,N_820,N_810);
nor U989 (N_989,N_802,N_815);
xnor U990 (N_990,N_815,N_812);
or U991 (N_991,N_844,N_810);
and U992 (N_992,N_849,N_806);
xor U993 (N_993,N_820,N_883);
nor U994 (N_994,N_876,N_887);
or U995 (N_995,N_899,N_857);
or U996 (N_996,N_832,N_877);
nand U997 (N_997,N_825,N_855);
nor U998 (N_998,N_856,N_850);
xor U999 (N_999,N_832,N_874);
nand U1000 (N_1000,N_981,N_948);
or U1001 (N_1001,N_900,N_908);
or U1002 (N_1002,N_935,N_924);
or U1003 (N_1003,N_950,N_914);
and U1004 (N_1004,N_956,N_959);
and U1005 (N_1005,N_953,N_931);
nor U1006 (N_1006,N_954,N_927);
and U1007 (N_1007,N_955,N_973);
or U1008 (N_1008,N_910,N_961);
xnor U1009 (N_1009,N_934,N_975);
nor U1010 (N_1010,N_998,N_974);
or U1011 (N_1011,N_964,N_905);
and U1012 (N_1012,N_904,N_971);
nor U1013 (N_1013,N_937,N_962);
nand U1014 (N_1014,N_940,N_915);
and U1015 (N_1015,N_988,N_939);
nor U1016 (N_1016,N_976,N_923);
nand U1017 (N_1017,N_979,N_930);
and U1018 (N_1018,N_968,N_949);
and U1019 (N_1019,N_989,N_938);
or U1020 (N_1020,N_967,N_991);
nor U1021 (N_1021,N_926,N_946);
or U1022 (N_1022,N_902,N_996);
nor U1023 (N_1023,N_994,N_960);
or U1024 (N_1024,N_990,N_941);
nand U1025 (N_1025,N_997,N_918);
nand U1026 (N_1026,N_909,N_912);
xor U1027 (N_1027,N_983,N_925);
xnor U1028 (N_1028,N_957,N_928);
nor U1029 (N_1029,N_917,N_932);
nor U1030 (N_1030,N_958,N_995);
and U1031 (N_1031,N_906,N_943);
nand U1032 (N_1032,N_977,N_993);
nor U1033 (N_1033,N_985,N_969);
and U1034 (N_1034,N_933,N_978);
or U1035 (N_1035,N_916,N_929);
xnor U1036 (N_1036,N_901,N_984);
or U1037 (N_1037,N_945,N_944);
or U1038 (N_1038,N_963,N_922);
nand U1039 (N_1039,N_999,N_952);
or U1040 (N_1040,N_965,N_947);
nand U1041 (N_1041,N_992,N_970);
and U1042 (N_1042,N_920,N_982);
nand U1043 (N_1043,N_986,N_987);
and U1044 (N_1044,N_942,N_911);
or U1045 (N_1045,N_980,N_921);
and U1046 (N_1046,N_919,N_907);
and U1047 (N_1047,N_936,N_966);
and U1048 (N_1048,N_913,N_972);
or U1049 (N_1049,N_903,N_951);
nand U1050 (N_1050,N_930,N_931);
or U1051 (N_1051,N_952,N_989);
nand U1052 (N_1052,N_904,N_994);
and U1053 (N_1053,N_902,N_946);
and U1054 (N_1054,N_964,N_952);
nor U1055 (N_1055,N_956,N_979);
or U1056 (N_1056,N_960,N_921);
and U1057 (N_1057,N_997,N_978);
and U1058 (N_1058,N_988,N_932);
nand U1059 (N_1059,N_963,N_936);
xnor U1060 (N_1060,N_987,N_914);
nor U1061 (N_1061,N_914,N_974);
xor U1062 (N_1062,N_950,N_958);
and U1063 (N_1063,N_920,N_987);
nor U1064 (N_1064,N_980,N_929);
nor U1065 (N_1065,N_940,N_969);
xor U1066 (N_1066,N_956,N_936);
and U1067 (N_1067,N_915,N_942);
and U1068 (N_1068,N_958,N_935);
and U1069 (N_1069,N_981,N_946);
and U1070 (N_1070,N_995,N_908);
nand U1071 (N_1071,N_926,N_917);
xor U1072 (N_1072,N_935,N_944);
nand U1073 (N_1073,N_927,N_935);
nand U1074 (N_1074,N_988,N_964);
or U1075 (N_1075,N_943,N_932);
and U1076 (N_1076,N_990,N_944);
nand U1077 (N_1077,N_924,N_919);
nand U1078 (N_1078,N_971,N_965);
or U1079 (N_1079,N_974,N_919);
xor U1080 (N_1080,N_967,N_927);
xnor U1081 (N_1081,N_945,N_963);
or U1082 (N_1082,N_968,N_977);
and U1083 (N_1083,N_947,N_949);
nor U1084 (N_1084,N_940,N_971);
and U1085 (N_1085,N_952,N_974);
nor U1086 (N_1086,N_934,N_915);
nor U1087 (N_1087,N_947,N_993);
nor U1088 (N_1088,N_919,N_956);
nor U1089 (N_1089,N_958,N_941);
xor U1090 (N_1090,N_905,N_995);
nand U1091 (N_1091,N_934,N_940);
nand U1092 (N_1092,N_999,N_982);
nand U1093 (N_1093,N_923,N_975);
xnor U1094 (N_1094,N_973,N_954);
and U1095 (N_1095,N_930,N_955);
and U1096 (N_1096,N_918,N_930);
nor U1097 (N_1097,N_902,N_965);
nor U1098 (N_1098,N_962,N_940);
and U1099 (N_1099,N_977,N_989);
xor U1100 (N_1100,N_1046,N_1059);
nand U1101 (N_1101,N_1010,N_1056);
and U1102 (N_1102,N_1015,N_1044);
or U1103 (N_1103,N_1035,N_1011);
nand U1104 (N_1104,N_1084,N_1073);
nand U1105 (N_1105,N_1045,N_1094);
xor U1106 (N_1106,N_1022,N_1013);
and U1107 (N_1107,N_1079,N_1017);
nor U1108 (N_1108,N_1086,N_1019);
and U1109 (N_1109,N_1002,N_1003);
nor U1110 (N_1110,N_1052,N_1066);
and U1111 (N_1111,N_1006,N_1061);
and U1112 (N_1112,N_1053,N_1036);
nor U1113 (N_1113,N_1091,N_1055);
or U1114 (N_1114,N_1038,N_1042);
nor U1115 (N_1115,N_1093,N_1025);
nor U1116 (N_1116,N_1007,N_1050);
and U1117 (N_1117,N_1040,N_1085);
nor U1118 (N_1118,N_1001,N_1037);
nor U1119 (N_1119,N_1058,N_1074);
nor U1120 (N_1120,N_1078,N_1057);
or U1121 (N_1121,N_1027,N_1092);
and U1122 (N_1122,N_1099,N_1071);
or U1123 (N_1123,N_1004,N_1032);
nand U1124 (N_1124,N_1067,N_1062);
nand U1125 (N_1125,N_1014,N_1068);
xnor U1126 (N_1126,N_1020,N_1008);
or U1127 (N_1127,N_1077,N_1060);
xnor U1128 (N_1128,N_1081,N_1049);
and U1129 (N_1129,N_1088,N_1031);
nand U1130 (N_1130,N_1030,N_1070);
xor U1131 (N_1131,N_1087,N_1048);
or U1132 (N_1132,N_1064,N_1029);
and U1133 (N_1133,N_1016,N_1023);
nand U1134 (N_1134,N_1076,N_1026);
nor U1135 (N_1135,N_1034,N_1018);
and U1136 (N_1136,N_1028,N_1075);
and U1137 (N_1137,N_1069,N_1098);
nor U1138 (N_1138,N_1005,N_1012);
or U1139 (N_1139,N_1072,N_1080);
nor U1140 (N_1140,N_1065,N_1054);
or U1141 (N_1141,N_1082,N_1009);
or U1142 (N_1142,N_1041,N_1097);
or U1143 (N_1143,N_1047,N_1051);
or U1144 (N_1144,N_1090,N_1096);
and U1145 (N_1145,N_1039,N_1089);
or U1146 (N_1146,N_1000,N_1033);
nand U1147 (N_1147,N_1063,N_1021);
xor U1148 (N_1148,N_1083,N_1043);
nor U1149 (N_1149,N_1095,N_1024);
nor U1150 (N_1150,N_1048,N_1085);
nand U1151 (N_1151,N_1043,N_1001);
nor U1152 (N_1152,N_1023,N_1053);
nand U1153 (N_1153,N_1083,N_1072);
nand U1154 (N_1154,N_1078,N_1065);
xor U1155 (N_1155,N_1074,N_1098);
or U1156 (N_1156,N_1039,N_1020);
and U1157 (N_1157,N_1017,N_1050);
nand U1158 (N_1158,N_1024,N_1011);
nor U1159 (N_1159,N_1072,N_1099);
nor U1160 (N_1160,N_1006,N_1039);
or U1161 (N_1161,N_1020,N_1031);
nor U1162 (N_1162,N_1016,N_1021);
nand U1163 (N_1163,N_1065,N_1063);
or U1164 (N_1164,N_1012,N_1094);
or U1165 (N_1165,N_1089,N_1014);
or U1166 (N_1166,N_1046,N_1009);
and U1167 (N_1167,N_1039,N_1085);
xor U1168 (N_1168,N_1023,N_1034);
nor U1169 (N_1169,N_1062,N_1005);
nor U1170 (N_1170,N_1007,N_1046);
xnor U1171 (N_1171,N_1099,N_1050);
xor U1172 (N_1172,N_1056,N_1087);
and U1173 (N_1173,N_1044,N_1099);
and U1174 (N_1174,N_1086,N_1024);
nand U1175 (N_1175,N_1071,N_1045);
or U1176 (N_1176,N_1028,N_1080);
or U1177 (N_1177,N_1048,N_1089);
and U1178 (N_1178,N_1014,N_1029);
nor U1179 (N_1179,N_1024,N_1074);
nand U1180 (N_1180,N_1065,N_1093);
or U1181 (N_1181,N_1022,N_1058);
and U1182 (N_1182,N_1056,N_1096);
and U1183 (N_1183,N_1049,N_1032);
nor U1184 (N_1184,N_1044,N_1025);
nor U1185 (N_1185,N_1080,N_1063);
and U1186 (N_1186,N_1053,N_1065);
nor U1187 (N_1187,N_1052,N_1048);
nand U1188 (N_1188,N_1069,N_1027);
and U1189 (N_1189,N_1033,N_1054);
nand U1190 (N_1190,N_1020,N_1005);
xnor U1191 (N_1191,N_1089,N_1067);
nor U1192 (N_1192,N_1055,N_1082);
nor U1193 (N_1193,N_1027,N_1053);
xnor U1194 (N_1194,N_1004,N_1092);
nor U1195 (N_1195,N_1076,N_1065);
and U1196 (N_1196,N_1082,N_1028);
or U1197 (N_1197,N_1008,N_1003);
and U1198 (N_1198,N_1003,N_1052);
nor U1199 (N_1199,N_1092,N_1093);
nor U1200 (N_1200,N_1193,N_1186);
and U1201 (N_1201,N_1101,N_1120);
and U1202 (N_1202,N_1122,N_1109);
and U1203 (N_1203,N_1124,N_1105);
or U1204 (N_1204,N_1151,N_1164);
xor U1205 (N_1205,N_1155,N_1141);
nor U1206 (N_1206,N_1102,N_1167);
nand U1207 (N_1207,N_1196,N_1183);
nor U1208 (N_1208,N_1146,N_1156);
nor U1209 (N_1209,N_1180,N_1154);
nand U1210 (N_1210,N_1168,N_1199);
or U1211 (N_1211,N_1138,N_1169);
nand U1212 (N_1212,N_1106,N_1136);
and U1213 (N_1213,N_1135,N_1103);
or U1214 (N_1214,N_1191,N_1182);
and U1215 (N_1215,N_1192,N_1187);
xnor U1216 (N_1216,N_1179,N_1118);
xnor U1217 (N_1217,N_1134,N_1127);
or U1218 (N_1218,N_1119,N_1140);
nand U1219 (N_1219,N_1112,N_1113);
xnor U1220 (N_1220,N_1137,N_1129);
nor U1221 (N_1221,N_1130,N_1117);
or U1222 (N_1222,N_1100,N_1115);
or U1223 (N_1223,N_1176,N_1152);
nand U1224 (N_1224,N_1178,N_1147);
or U1225 (N_1225,N_1184,N_1165);
and U1226 (N_1226,N_1139,N_1158);
nand U1227 (N_1227,N_1174,N_1116);
nand U1228 (N_1228,N_1150,N_1143);
or U1229 (N_1229,N_1161,N_1110);
nand U1230 (N_1230,N_1173,N_1121);
and U1231 (N_1231,N_1195,N_1107);
and U1232 (N_1232,N_1170,N_1125);
nand U1233 (N_1233,N_1145,N_1142);
nor U1234 (N_1234,N_1126,N_1194);
xor U1235 (N_1235,N_1163,N_1190);
and U1236 (N_1236,N_1132,N_1189);
nor U1237 (N_1237,N_1198,N_1144);
and U1238 (N_1238,N_1148,N_1133);
nor U1239 (N_1239,N_1111,N_1175);
nor U1240 (N_1240,N_1108,N_1157);
nand U1241 (N_1241,N_1177,N_1128);
nand U1242 (N_1242,N_1185,N_1153);
and U1243 (N_1243,N_1114,N_1149);
or U1244 (N_1244,N_1123,N_1197);
nand U1245 (N_1245,N_1188,N_1162);
nand U1246 (N_1246,N_1171,N_1159);
or U1247 (N_1247,N_1104,N_1181);
xnor U1248 (N_1248,N_1172,N_1160);
xor U1249 (N_1249,N_1166,N_1131);
or U1250 (N_1250,N_1103,N_1174);
or U1251 (N_1251,N_1131,N_1133);
or U1252 (N_1252,N_1115,N_1196);
or U1253 (N_1253,N_1166,N_1141);
nand U1254 (N_1254,N_1164,N_1153);
or U1255 (N_1255,N_1184,N_1109);
nor U1256 (N_1256,N_1148,N_1143);
nor U1257 (N_1257,N_1186,N_1112);
nand U1258 (N_1258,N_1178,N_1165);
nand U1259 (N_1259,N_1135,N_1177);
or U1260 (N_1260,N_1180,N_1177);
nand U1261 (N_1261,N_1195,N_1140);
nand U1262 (N_1262,N_1161,N_1189);
nor U1263 (N_1263,N_1138,N_1168);
and U1264 (N_1264,N_1152,N_1192);
nand U1265 (N_1265,N_1174,N_1167);
or U1266 (N_1266,N_1145,N_1123);
xnor U1267 (N_1267,N_1140,N_1104);
or U1268 (N_1268,N_1120,N_1106);
nand U1269 (N_1269,N_1166,N_1151);
xnor U1270 (N_1270,N_1153,N_1154);
nand U1271 (N_1271,N_1158,N_1116);
nand U1272 (N_1272,N_1157,N_1167);
or U1273 (N_1273,N_1171,N_1180);
and U1274 (N_1274,N_1185,N_1186);
or U1275 (N_1275,N_1170,N_1158);
and U1276 (N_1276,N_1132,N_1140);
xor U1277 (N_1277,N_1171,N_1134);
nand U1278 (N_1278,N_1147,N_1161);
or U1279 (N_1279,N_1193,N_1131);
nor U1280 (N_1280,N_1115,N_1180);
nor U1281 (N_1281,N_1113,N_1126);
nand U1282 (N_1282,N_1182,N_1197);
nor U1283 (N_1283,N_1177,N_1119);
nor U1284 (N_1284,N_1117,N_1192);
nor U1285 (N_1285,N_1182,N_1196);
or U1286 (N_1286,N_1175,N_1105);
and U1287 (N_1287,N_1197,N_1186);
xor U1288 (N_1288,N_1110,N_1139);
nand U1289 (N_1289,N_1120,N_1189);
or U1290 (N_1290,N_1104,N_1107);
xnor U1291 (N_1291,N_1188,N_1102);
and U1292 (N_1292,N_1176,N_1100);
nor U1293 (N_1293,N_1116,N_1149);
or U1294 (N_1294,N_1170,N_1199);
nor U1295 (N_1295,N_1128,N_1114);
or U1296 (N_1296,N_1165,N_1135);
and U1297 (N_1297,N_1118,N_1144);
and U1298 (N_1298,N_1170,N_1149);
or U1299 (N_1299,N_1156,N_1180);
or U1300 (N_1300,N_1203,N_1241);
nand U1301 (N_1301,N_1298,N_1213);
nand U1302 (N_1302,N_1222,N_1242);
or U1303 (N_1303,N_1209,N_1223);
nand U1304 (N_1304,N_1225,N_1239);
and U1305 (N_1305,N_1257,N_1252);
nor U1306 (N_1306,N_1260,N_1210);
or U1307 (N_1307,N_1285,N_1294);
nand U1308 (N_1308,N_1277,N_1289);
or U1309 (N_1309,N_1279,N_1275);
nor U1310 (N_1310,N_1270,N_1268);
nand U1311 (N_1311,N_1282,N_1218);
and U1312 (N_1312,N_1284,N_1206);
and U1313 (N_1313,N_1271,N_1297);
nor U1314 (N_1314,N_1296,N_1202);
nor U1315 (N_1315,N_1287,N_1233);
nand U1316 (N_1316,N_1246,N_1272);
or U1317 (N_1317,N_1278,N_1232);
or U1318 (N_1318,N_1240,N_1236);
or U1319 (N_1319,N_1288,N_1243);
nand U1320 (N_1320,N_1256,N_1208);
or U1321 (N_1321,N_1248,N_1249);
and U1322 (N_1322,N_1212,N_1221);
nand U1323 (N_1323,N_1259,N_1238);
xor U1324 (N_1324,N_1231,N_1253);
or U1325 (N_1325,N_1280,N_1214);
nand U1326 (N_1326,N_1200,N_1292);
nand U1327 (N_1327,N_1269,N_1299);
nand U1328 (N_1328,N_1227,N_1215);
nor U1329 (N_1329,N_1211,N_1258);
nor U1330 (N_1330,N_1266,N_1245);
nor U1331 (N_1331,N_1220,N_1228);
nor U1332 (N_1332,N_1273,N_1274);
or U1333 (N_1333,N_1290,N_1235);
and U1334 (N_1334,N_1250,N_1291);
or U1335 (N_1335,N_1207,N_1286);
xor U1336 (N_1336,N_1237,N_1281);
or U1337 (N_1337,N_1247,N_1265);
and U1338 (N_1338,N_1267,N_1204);
nand U1339 (N_1339,N_1251,N_1217);
xor U1340 (N_1340,N_1261,N_1293);
and U1341 (N_1341,N_1216,N_1234);
or U1342 (N_1342,N_1283,N_1295);
or U1343 (N_1343,N_1201,N_1230);
and U1344 (N_1344,N_1276,N_1262);
nor U1345 (N_1345,N_1244,N_1264);
nand U1346 (N_1346,N_1255,N_1254);
and U1347 (N_1347,N_1229,N_1226);
or U1348 (N_1348,N_1219,N_1224);
or U1349 (N_1349,N_1263,N_1205);
and U1350 (N_1350,N_1296,N_1261);
nand U1351 (N_1351,N_1247,N_1291);
nand U1352 (N_1352,N_1298,N_1249);
xor U1353 (N_1353,N_1268,N_1247);
nand U1354 (N_1354,N_1216,N_1284);
nand U1355 (N_1355,N_1218,N_1285);
nor U1356 (N_1356,N_1226,N_1223);
nand U1357 (N_1357,N_1265,N_1242);
or U1358 (N_1358,N_1226,N_1266);
and U1359 (N_1359,N_1229,N_1295);
and U1360 (N_1360,N_1241,N_1259);
nand U1361 (N_1361,N_1263,N_1238);
or U1362 (N_1362,N_1255,N_1213);
nor U1363 (N_1363,N_1268,N_1216);
and U1364 (N_1364,N_1247,N_1234);
and U1365 (N_1365,N_1226,N_1221);
and U1366 (N_1366,N_1291,N_1207);
or U1367 (N_1367,N_1218,N_1276);
nand U1368 (N_1368,N_1253,N_1227);
nand U1369 (N_1369,N_1212,N_1238);
or U1370 (N_1370,N_1222,N_1281);
nand U1371 (N_1371,N_1274,N_1209);
or U1372 (N_1372,N_1239,N_1223);
xnor U1373 (N_1373,N_1222,N_1288);
and U1374 (N_1374,N_1297,N_1259);
nand U1375 (N_1375,N_1207,N_1240);
nand U1376 (N_1376,N_1268,N_1223);
and U1377 (N_1377,N_1202,N_1243);
and U1378 (N_1378,N_1296,N_1266);
nand U1379 (N_1379,N_1257,N_1280);
and U1380 (N_1380,N_1281,N_1223);
nand U1381 (N_1381,N_1269,N_1209);
nand U1382 (N_1382,N_1202,N_1258);
and U1383 (N_1383,N_1204,N_1230);
and U1384 (N_1384,N_1217,N_1262);
nor U1385 (N_1385,N_1275,N_1274);
nand U1386 (N_1386,N_1295,N_1218);
xnor U1387 (N_1387,N_1265,N_1220);
and U1388 (N_1388,N_1241,N_1298);
nand U1389 (N_1389,N_1259,N_1249);
or U1390 (N_1390,N_1215,N_1255);
or U1391 (N_1391,N_1209,N_1228);
xnor U1392 (N_1392,N_1262,N_1280);
nor U1393 (N_1393,N_1291,N_1256);
and U1394 (N_1394,N_1287,N_1203);
or U1395 (N_1395,N_1248,N_1226);
or U1396 (N_1396,N_1262,N_1203);
nand U1397 (N_1397,N_1242,N_1298);
or U1398 (N_1398,N_1277,N_1266);
or U1399 (N_1399,N_1222,N_1298);
and U1400 (N_1400,N_1373,N_1354);
nor U1401 (N_1401,N_1335,N_1374);
nand U1402 (N_1402,N_1364,N_1350);
and U1403 (N_1403,N_1329,N_1312);
nor U1404 (N_1404,N_1399,N_1383);
xnor U1405 (N_1405,N_1310,N_1358);
or U1406 (N_1406,N_1382,N_1369);
nand U1407 (N_1407,N_1365,N_1352);
nand U1408 (N_1408,N_1362,N_1315);
and U1409 (N_1409,N_1349,N_1305);
nand U1410 (N_1410,N_1341,N_1301);
nor U1411 (N_1411,N_1351,N_1300);
nor U1412 (N_1412,N_1334,N_1342);
nand U1413 (N_1413,N_1359,N_1353);
nand U1414 (N_1414,N_1327,N_1337);
nand U1415 (N_1415,N_1308,N_1360);
or U1416 (N_1416,N_1378,N_1381);
and U1417 (N_1417,N_1309,N_1338);
and U1418 (N_1418,N_1393,N_1321);
nand U1419 (N_1419,N_1398,N_1303);
and U1420 (N_1420,N_1372,N_1385);
nand U1421 (N_1421,N_1376,N_1397);
nor U1422 (N_1422,N_1357,N_1366);
or U1423 (N_1423,N_1361,N_1380);
or U1424 (N_1424,N_1306,N_1304);
and U1425 (N_1425,N_1339,N_1384);
xor U1426 (N_1426,N_1348,N_1392);
and U1427 (N_1427,N_1316,N_1394);
nor U1428 (N_1428,N_1313,N_1318);
nand U1429 (N_1429,N_1368,N_1379);
nand U1430 (N_1430,N_1346,N_1320);
and U1431 (N_1431,N_1311,N_1336);
nand U1432 (N_1432,N_1317,N_1340);
xnor U1433 (N_1433,N_1375,N_1367);
or U1434 (N_1434,N_1388,N_1319);
nor U1435 (N_1435,N_1395,N_1332);
nor U1436 (N_1436,N_1314,N_1347);
or U1437 (N_1437,N_1363,N_1356);
nand U1438 (N_1438,N_1386,N_1396);
nor U1439 (N_1439,N_1370,N_1307);
nand U1440 (N_1440,N_1323,N_1371);
nand U1441 (N_1441,N_1326,N_1377);
xor U1442 (N_1442,N_1390,N_1328);
nand U1443 (N_1443,N_1343,N_1389);
or U1444 (N_1444,N_1387,N_1355);
nor U1445 (N_1445,N_1331,N_1325);
nor U1446 (N_1446,N_1302,N_1333);
xor U1447 (N_1447,N_1330,N_1324);
nand U1448 (N_1448,N_1344,N_1345);
nor U1449 (N_1449,N_1322,N_1391);
nor U1450 (N_1450,N_1311,N_1322);
nor U1451 (N_1451,N_1364,N_1366);
or U1452 (N_1452,N_1308,N_1375);
or U1453 (N_1453,N_1373,N_1324);
and U1454 (N_1454,N_1393,N_1305);
xnor U1455 (N_1455,N_1364,N_1385);
nand U1456 (N_1456,N_1304,N_1317);
or U1457 (N_1457,N_1353,N_1369);
nor U1458 (N_1458,N_1314,N_1356);
and U1459 (N_1459,N_1300,N_1397);
xor U1460 (N_1460,N_1339,N_1374);
nand U1461 (N_1461,N_1311,N_1334);
and U1462 (N_1462,N_1355,N_1395);
nor U1463 (N_1463,N_1350,N_1336);
xor U1464 (N_1464,N_1362,N_1329);
or U1465 (N_1465,N_1325,N_1367);
xor U1466 (N_1466,N_1394,N_1352);
or U1467 (N_1467,N_1395,N_1391);
or U1468 (N_1468,N_1319,N_1347);
nor U1469 (N_1469,N_1395,N_1334);
nand U1470 (N_1470,N_1369,N_1367);
nand U1471 (N_1471,N_1326,N_1352);
or U1472 (N_1472,N_1333,N_1329);
or U1473 (N_1473,N_1345,N_1383);
nand U1474 (N_1474,N_1398,N_1308);
xor U1475 (N_1475,N_1328,N_1345);
xor U1476 (N_1476,N_1335,N_1372);
or U1477 (N_1477,N_1398,N_1364);
and U1478 (N_1478,N_1352,N_1334);
nand U1479 (N_1479,N_1352,N_1316);
xnor U1480 (N_1480,N_1332,N_1331);
and U1481 (N_1481,N_1365,N_1304);
or U1482 (N_1482,N_1376,N_1309);
and U1483 (N_1483,N_1307,N_1316);
nand U1484 (N_1484,N_1307,N_1329);
nand U1485 (N_1485,N_1392,N_1366);
or U1486 (N_1486,N_1339,N_1376);
nor U1487 (N_1487,N_1305,N_1351);
or U1488 (N_1488,N_1376,N_1392);
nand U1489 (N_1489,N_1371,N_1329);
and U1490 (N_1490,N_1363,N_1315);
nor U1491 (N_1491,N_1349,N_1366);
or U1492 (N_1492,N_1397,N_1389);
nor U1493 (N_1493,N_1376,N_1383);
nor U1494 (N_1494,N_1364,N_1306);
nand U1495 (N_1495,N_1313,N_1388);
xnor U1496 (N_1496,N_1319,N_1350);
and U1497 (N_1497,N_1311,N_1302);
and U1498 (N_1498,N_1349,N_1322);
and U1499 (N_1499,N_1324,N_1382);
nor U1500 (N_1500,N_1473,N_1402);
nand U1501 (N_1501,N_1465,N_1410);
and U1502 (N_1502,N_1449,N_1495);
nand U1503 (N_1503,N_1426,N_1434);
or U1504 (N_1504,N_1423,N_1442);
or U1505 (N_1505,N_1413,N_1448);
nor U1506 (N_1506,N_1421,N_1427);
or U1507 (N_1507,N_1403,N_1429);
nand U1508 (N_1508,N_1460,N_1405);
and U1509 (N_1509,N_1425,N_1428);
and U1510 (N_1510,N_1494,N_1499);
nor U1511 (N_1511,N_1455,N_1487);
or U1512 (N_1512,N_1468,N_1407);
nand U1513 (N_1513,N_1488,N_1489);
nor U1514 (N_1514,N_1415,N_1486);
nor U1515 (N_1515,N_1461,N_1471);
nor U1516 (N_1516,N_1457,N_1422);
nor U1517 (N_1517,N_1464,N_1463);
xnor U1518 (N_1518,N_1445,N_1469);
or U1519 (N_1519,N_1485,N_1479);
nor U1520 (N_1520,N_1491,N_1454);
and U1521 (N_1521,N_1431,N_1476);
nor U1522 (N_1522,N_1443,N_1437);
nor U1523 (N_1523,N_1424,N_1412);
nor U1524 (N_1524,N_1408,N_1466);
nand U1525 (N_1525,N_1452,N_1409);
nor U1526 (N_1526,N_1417,N_1404);
nor U1527 (N_1527,N_1444,N_1496);
or U1528 (N_1528,N_1492,N_1498);
or U1529 (N_1529,N_1414,N_1477);
and U1530 (N_1530,N_1436,N_1480);
nor U1531 (N_1531,N_1416,N_1472);
nor U1532 (N_1532,N_1475,N_1440);
nor U1533 (N_1533,N_1484,N_1411);
nand U1534 (N_1534,N_1432,N_1451);
and U1535 (N_1535,N_1481,N_1474);
nand U1536 (N_1536,N_1497,N_1482);
or U1537 (N_1537,N_1418,N_1478);
or U1538 (N_1538,N_1441,N_1456);
xnor U1539 (N_1539,N_1470,N_1493);
nand U1540 (N_1540,N_1453,N_1430);
nor U1541 (N_1541,N_1406,N_1433);
and U1542 (N_1542,N_1462,N_1420);
and U1543 (N_1543,N_1459,N_1447);
nand U1544 (N_1544,N_1490,N_1439);
or U1545 (N_1545,N_1438,N_1400);
and U1546 (N_1546,N_1446,N_1401);
and U1547 (N_1547,N_1435,N_1458);
nor U1548 (N_1548,N_1483,N_1419);
nand U1549 (N_1549,N_1450,N_1467);
nand U1550 (N_1550,N_1482,N_1425);
nor U1551 (N_1551,N_1469,N_1439);
nand U1552 (N_1552,N_1447,N_1426);
or U1553 (N_1553,N_1489,N_1413);
nand U1554 (N_1554,N_1473,N_1492);
and U1555 (N_1555,N_1484,N_1437);
nand U1556 (N_1556,N_1486,N_1438);
nand U1557 (N_1557,N_1467,N_1413);
xnor U1558 (N_1558,N_1457,N_1414);
nand U1559 (N_1559,N_1434,N_1437);
nand U1560 (N_1560,N_1458,N_1445);
nand U1561 (N_1561,N_1424,N_1472);
or U1562 (N_1562,N_1418,N_1437);
nor U1563 (N_1563,N_1440,N_1411);
or U1564 (N_1564,N_1482,N_1410);
or U1565 (N_1565,N_1428,N_1478);
and U1566 (N_1566,N_1495,N_1494);
and U1567 (N_1567,N_1476,N_1493);
and U1568 (N_1568,N_1408,N_1458);
nor U1569 (N_1569,N_1421,N_1433);
nand U1570 (N_1570,N_1477,N_1411);
nor U1571 (N_1571,N_1489,N_1438);
nor U1572 (N_1572,N_1474,N_1442);
or U1573 (N_1573,N_1483,N_1417);
nor U1574 (N_1574,N_1484,N_1402);
nor U1575 (N_1575,N_1455,N_1450);
or U1576 (N_1576,N_1478,N_1417);
and U1577 (N_1577,N_1413,N_1455);
nor U1578 (N_1578,N_1403,N_1476);
nand U1579 (N_1579,N_1448,N_1420);
xnor U1580 (N_1580,N_1450,N_1462);
nand U1581 (N_1581,N_1413,N_1462);
xnor U1582 (N_1582,N_1475,N_1425);
nand U1583 (N_1583,N_1455,N_1498);
nand U1584 (N_1584,N_1485,N_1432);
nor U1585 (N_1585,N_1472,N_1420);
nand U1586 (N_1586,N_1448,N_1406);
xnor U1587 (N_1587,N_1461,N_1420);
nor U1588 (N_1588,N_1473,N_1452);
nor U1589 (N_1589,N_1494,N_1433);
and U1590 (N_1590,N_1428,N_1411);
nand U1591 (N_1591,N_1483,N_1405);
or U1592 (N_1592,N_1400,N_1410);
and U1593 (N_1593,N_1434,N_1443);
nor U1594 (N_1594,N_1432,N_1401);
nor U1595 (N_1595,N_1461,N_1453);
nor U1596 (N_1596,N_1406,N_1425);
xor U1597 (N_1597,N_1412,N_1440);
nand U1598 (N_1598,N_1428,N_1488);
xor U1599 (N_1599,N_1463,N_1441);
nor U1600 (N_1600,N_1533,N_1532);
nand U1601 (N_1601,N_1521,N_1569);
nand U1602 (N_1602,N_1582,N_1544);
nand U1603 (N_1603,N_1509,N_1540);
nor U1604 (N_1604,N_1546,N_1551);
nand U1605 (N_1605,N_1539,N_1513);
and U1606 (N_1606,N_1585,N_1592);
and U1607 (N_1607,N_1514,N_1531);
and U1608 (N_1608,N_1568,N_1570);
or U1609 (N_1609,N_1571,N_1552);
nor U1610 (N_1610,N_1512,N_1529);
and U1611 (N_1611,N_1555,N_1541);
or U1612 (N_1612,N_1516,N_1588);
nand U1613 (N_1613,N_1524,N_1523);
nor U1614 (N_1614,N_1564,N_1504);
and U1615 (N_1615,N_1511,N_1554);
or U1616 (N_1616,N_1591,N_1538);
nor U1617 (N_1617,N_1589,N_1596);
or U1618 (N_1618,N_1553,N_1518);
nor U1619 (N_1619,N_1599,N_1549);
nor U1620 (N_1620,N_1594,N_1583);
or U1621 (N_1621,N_1561,N_1595);
and U1622 (N_1622,N_1575,N_1580);
or U1623 (N_1623,N_1515,N_1528);
nand U1624 (N_1624,N_1572,N_1530);
nor U1625 (N_1625,N_1502,N_1556);
and U1626 (N_1626,N_1506,N_1507);
nand U1627 (N_1627,N_1503,N_1573);
or U1628 (N_1628,N_1598,N_1565);
nor U1629 (N_1629,N_1584,N_1587);
and U1630 (N_1630,N_1574,N_1567);
and U1631 (N_1631,N_1577,N_1517);
nor U1632 (N_1632,N_1576,N_1526);
or U1633 (N_1633,N_1597,N_1548);
nor U1634 (N_1634,N_1519,N_1578);
nand U1635 (N_1635,N_1545,N_1508);
xor U1636 (N_1636,N_1563,N_1557);
nand U1637 (N_1637,N_1559,N_1558);
nand U1638 (N_1638,N_1522,N_1500);
and U1639 (N_1639,N_1505,N_1581);
nand U1640 (N_1640,N_1535,N_1536);
nand U1641 (N_1641,N_1593,N_1527);
or U1642 (N_1642,N_1590,N_1501);
nor U1643 (N_1643,N_1566,N_1579);
or U1644 (N_1644,N_1550,N_1525);
nor U1645 (N_1645,N_1542,N_1510);
or U1646 (N_1646,N_1537,N_1560);
xor U1647 (N_1647,N_1547,N_1534);
nand U1648 (N_1648,N_1562,N_1543);
nand U1649 (N_1649,N_1520,N_1586);
nand U1650 (N_1650,N_1520,N_1523);
or U1651 (N_1651,N_1575,N_1532);
nand U1652 (N_1652,N_1510,N_1561);
or U1653 (N_1653,N_1556,N_1585);
nor U1654 (N_1654,N_1536,N_1583);
nand U1655 (N_1655,N_1552,N_1589);
xnor U1656 (N_1656,N_1597,N_1505);
nor U1657 (N_1657,N_1594,N_1593);
nor U1658 (N_1658,N_1520,N_1585);
xor U1659 (N_1659,N_1567,N_1583);
nor U1660 (N_1660,N_1590,N_1543);
or U1661 (N_1661,N_1580,N_1544);
and U1662 (N_1662,N_1589,N_1572);
nor U1663 (N_1663,N_1585,N_1586);
nor U1664 (N_1664,N_1527,N_1564);
nor U1665 (N_1665,N_1554,N_1588);
and U1666 (N_1666,N_1500,N_1507);
or U1667 (N_1667,N_1505,N_1571);
nand U1668 (N_1668,N_1502,N_1512);
xor U1669 (N_1669,N_1565,N_1586);
nand U1670 (N_1670,N_1571,N_1576);
xnor U1671 (N_1671,N_1578,N_1568);
or U1672 (N_1672,N_1557,N_1554);
nor U1673 (N_1673,N_1591,N_1554);
and U1674 (N_1674,N_1533,N_1581);
nor U1675 (N_1675,N_1572,N_1503);
and U1676 (N_1676,N_1507,N_1550);
nor U1677 (N_1677,N_1526,N_1535);
or U1678 (N_1678,N_1526,N_1541);
nor U1679 (N_1679,N_1566,N_1552);
and U1680 (N_1680,N_1559,N_1544);
or U1681 (N_1681,N_1521,N_1537);
nand U1682 (N_1682,N_1523,N_1539);
nor U1683 (N_1683,N_1565,N_1532);
nor U1684 (N_1684,N_1546,N_1562);
nor U1685 (N_1685,N_1561,N_1557);
and U1686 (N_1686,N_1549,N_1575);
nor U1687 (N_1687,N_1524,N_1566);
nand U1688 (N_1688,N_1588,N_1560);
nor U1689 (N_1689,N_1508,N_1588);
and U1690 (N_1690,N_1547,N_1542);
nand U1691 (N_1691,N_1561,N_1555);
and U1692 (N_1692,N_1541,N_1581);
and U1693 (N_1693,N_1529,N_1520);
nor U1694 (N_1694,N_1555,N_1558);
or U1695 (N_1695,N_1539,N_1542);
or U1696 (N_1696,N_1557,N_1530);
xor U1697 (N_1697,N_1584,N_1511);
and U1698 (N_1698,N_1534,N_1503);
nor U1699 (N_1699,N_1570,N_1557);
or U1700 (N_1700,N_1631,N_1608);
or U1701 (N_1701,N_1640,N_1653);
nor U1702 (N_1702,N_1638,N_1622);
nor U1703 (N_1703,N_1679,N_1615);
and U1704 (N_1704,N_1656,N_1683);
or U1705 (N_1705,N_1630,N_1614);
or U1706 (N_1706,N_1674,N_1691);
nor U1707 (N_1707,N_1625,N_1658);
nand U1708 (N_1708,N_1610,N_1619);
nand U1709 (N_1709,N_1606,N_1600);
and U1710 (N_1710,N_1621,N_1633);
nor U1711 (N_1711,N_1675,N_1666);
nand U1712 (N_1712,N_1686,N_1670);
nand U1713 (N_1713,N_1612,N_1644);
nand U1714 (N_1714,N_1671,N_1663);
nor U1715 (N_1715,N_1669,N_1696);
nor U1716 (N_1716,N_1618,N_1639);
nand U1717 (N_1717,N_1678,N_1613);
and U1718 (N_1718,N_1657,N_1697);
nand U1719 (N_1719,N_1623,N_1667);
nor U1720 (N_1720,N_1655,N_1665);
nand U1721 (N_1721,N_1641,N_1607);
nand U1722 (N_1722,N_1647,N_1634);
or U1723 (N_1723,N_1668,N_1681);
nor U1724 (N_1724,N_1680,N_1673);
nor U1725 (N_1725,N_1603,N_1651);
nor U1726 (N_1726,N_1661,N_1616);
nor U1727 (N_1727,N_1649,N_1617);
nor U1728 (N_1728,N_1602,N_1684);
and U1729 (N_1729,N_1635,N_1699);
xor U1730 (N_1730,N_1629,N_1605);
xnor U1731 (N_1731,N_1664,N_1685);
or U1732 (N_1732,N_1652,N_1643);
or U1733 (N_1733,N_1693,N_1628);
nand U1734 (N_1734,N_1660,N_1604);
xnor U1735 (N_1735,N_1688,N_1662);
nor U1736 (N_1736,N_1645,N_1689);
and U1737 (N_1737,N_1677,N_1632);
and U1738 (N_1738,N_1601,N_1687);
and U1739 (N_1739,N_1672,N_1659);
or U1740 (N_1740,N_1654,N_1627);
or U1741 (N_1741,N_1682,N_1646);
and U1742 (N_1742,N_1694,N_1650);
xor U1743 (N_1743,N_1648,N_1624);
or U1744 (N_1744,N_1626,N_1636);
nor U1745 (N_1745,N_1692,N_1637);
and U1746 (N_1746,N_1695,N_1609);
nand U1747 (N_1747,N_1611,N_1676);
and U1748 (N_1748,N_1690,N_1620);
nor U1749 (N_1749,N_1642,N_1698);
nor U1750 (N_1750,N_1652,N_1664);
and U1751 (N_1751,N_1605,N_1681);
or U1752 (N_1752,N_1616,N_1605);
and U1753 (N_1753,N_1696,N_1682);
nor U1754 (N_1754,N_1664,N_1621);
nand U1755 (N_1755,N_1698,N_1674);
and U1756 (N_1756,N_1623,N_1620);
nor U1757 (N_1757,N_1635,N_1600);
and U1758 (N_1758,N_1664,N_1600);
and U1759 (N_1759,N_1611,N_1631);
or U1760 (N_1760,N_1686,N_1640);
nand U1761 (N_1761,N_1606,N_1694);
nor U1762 (N_1762,N_1647,N_1643);
and U1763 (N_1763,N_1612,N_1648);
nand U1764 (N_1764,N_1606,N_1666);
or U1765 (N_1765,N_1652,N_1613);
nand U1766 (N_1766,N_1600,N_1610);
nand U1767 (N_1767,N_1639,N_1607);
nor U1768 (N_1768,N_1652,N_1641);
nor U1769 (N_1769,N_1604,N_1628);
xnor U1770 (N_1770,N_1652,N_1688);
nor U1771 (N_1771,N_1621,N_1671);
nor U1772 (N_1772,N_1689,N_1663);
or U1773 (N_1773,N_1670,N_1637);
and U1774 (N_1774,N_1683,N_1691);
nor U1775 (N_1775,N_1677,N_1614);
nor U1776 (N_1776,N_1663,N_1605);
or U1777 (N_1777,N_1647,N_1651);
or U1778 (N_1778,N_1689,N_1658);
nand U1779 (N_1779,N_1636,N_1620);
or U1780 (N_1780,N_1606,N_1644);
nor U1781 (N_1781,N_1671,N_1680);
and U1782 (N_1782,N_1622,N_1612);
and U1783 (N_1783,N_1653,N_1630);
nor U1784 (N_1784,N_1690,N_1614);
nand U1785 (N_1785,N_1632,N_1671);
nor U1786 (N_1786,N_1678,N_1667);
and U1787 (N_1787,N_1635,N_1651);
or U1788 (N_1788,N_1669,N_1666);
nand U1789 (N_1789,N_1688,N_1694);
nand U1790 (N_1790,N_1666,N_1603);
or U1791 (N_1791,N_1631,N_1686);
xnor U1792 (N_1792,N_1608,N_1681);
nor U1793 (N_1793,N_1613,N_1698);
nand U1794 (N_1794,N_1653,N_1683);
nor U1795 (N_1795,N_1614,N_1649);
nor U1796 (N_1796,N_1645,N_1665);
and U1797 (N_1797,N_1692,N_1621);
or U1798 (N_1798,N_1639,N_1687);
nand U1799 (N_1799,N_1618,N_1690);
or U1800 (N_1800,N_1733,N_1760);
and U1801 (N_1801,N_1781,N_1770);
nor U1802 (N_1802,N_1771,N_1721);
nand U1803 (N_1803,N_1709,N_1798);
nor U1804 (N_1804,N_1725,N_1785);
and U1805 (N_1805,N_1739,N_1766);
or U1806 (N_1806,N_1753,N_1743);
nor U1807 (N_1807,N_1796,N_1735);
nor U1808 (N_1808,N_1740,N_1789);
and U1809 (N_1809,N_1754,N_1723);
nor U1810 (N_1810,N_1722,N_1706);
and U1811 (N_1811,N_1727,N_1710);
or U1812 (N_1812,N_1745,N_1729);
and U1813 (N_1813,N_1780,N_1757);
nand U1814 (N_1814,N_1700,N_1799);
and U1815 (N_1815,N_1704,N_1715);
or U1816 (N_1816,N_1788,N_1756);
or U1817 (N_1817,N_1732,N_1765);
nand U1818 (N_1818,N_1777,N_1741);
or U1819 (N_1819,N_1751,N_1784);
and U1820 (N_1820,N_1748,N_1791);
or U1821 (N_1821,N_1786,N_1714);
xnor U1822 (N_1822,N_1737,N_1779);
and U1823 (N_1823,N_1763,N_1731);
or U1824 (N_1824,N_1762,N_1761);
and U1825 (N_1825,N_1794,N_1712);
nor U1826 (N_1826,N_1720,N_1705);
and U1827 (N_1827,N_1768,N_1797);
nor U1828 (N_1828,N_1767,N_1759);
and U1829 (N_1829,N_1730,N_1782);
or U1830 (N_1830,N_1764,N_1776);
or U1831 (N_1831,N_1728,N_1773);
or U1832 (N_1832,N_1758,N_1718);
and U1833 (N_1833,N_1746,N_1702);
nor U1834 (N_1834,N_1747,N_1736);
or U1835 (N_1835,N_1738,N_1708);
nor U1836 (N_1836,N_1774,N_1775);
xnor U1837 (N_1837,N_1792,N_1716);
nor U1838 (N_1838,N_1711,N_1713);
nand U1839 (N_1839,N_1755,N_1793);
nand U1840 (N_1840,N_1707,N_1724);
nand U1841 (N_1841,N_1778,N_1742);
or U1842 (N_1842,N_1795,N_1717);
nor U1843 (N_1843,N_1726,N_1701);
or U1844 (N_1844,N_1744,N_1719);
nand U1845 (N_1845,N_1750,N_1769);
nor U1846 (N_1846,N_1783,N_1734);
or U1847 (N_1847,N_1703,N_1752);
xnor U1848 (N_1848,N_1749,N_1790);
and U1849 (N_1849,N_1787,N_1772);
or U1850 (N_1850,N_1755,N_1766);
nor U1851 (N_1851,N_1788,N_1775);
nor U1852 (N_1852,N_1765,N_1745);
xor U1853 (N_1853,N_1718,N_1774);
or U1854 (N_1854,N_1765,N_1778);
or U1855 (N_1855,N_1719,N_1706);
xnor U1856 (N_1856,N_1762,N_1758);
or U1857 (N_1857,N_1761,N_1713);
and U1858 (N_1858,N_1746,N_1773);
nor U1859 (N_1859,N_1708,N_1755);
or U1860 (N_1860,N_1745,N_1762);
and U1861 (N_1861,N_1736,N_1739);
nand U1862 (N_1862,N_1702,N_1744);
nand U1863 (N_1863,N_1730,N_1776);
or U1864 (N_1864,N_1710,N_1737);
or U1865 (N_1865,N_1772,N_1755);
xnor U1866 (N_1866,N_1761,N_1730);
and U1867 (N_1867,N_1763,N_1726);
nand U1868 (N_1868,N_1782,N_1715);
nor U1869 (N_1869,N_1737,N_1788);
or U1870 (N_1870,N_1731,N_1762);
or U1871 (N_1871,N_1722,N_1703);
nand U1872 (N_1872,N_1723,N_1762);
or U1873 (N_1873,N_1766,N_1733);
and U1874 (N_1874,N_1787,N_1728);
nor U1875 (N_1875,N_1744,N_1785);
and U1876 (N_1876,N_1711,N_1763);
or U1877 (N_1877,N_1753,N_1711);
and U1878 (N_1878,N_1762,N_1765);
or U1879 (N_1879,N_1734,N_1747);
nand U1880 (N_1880,N_1712,N_1711);
nand U1881 (N_1881,N_1740,N_1752);
or U1882 (N_1882,N_1783,N_1760);
or U1883 (N_1883,N_1718,N_1795);
or U1884 (N_1884,N_1731,N_1708);
nor U1885 (N_1885,N_1749,N_1735);
and U1886 (N_1886,N_1792,N_1723);
nand U1887 (N_1887,N_1792,N_1790);
nor U1888 (N_1888,N_1746,N_1701);
or U1889 (N_1889,N_1722,N_1738);
or U1890 (N_1890,N_1769,N_1796);
nor U1891 (N_1891,N_1755,N_1794);
nand U1892 (N_1892,N_1738,N_1728);
nor U1893 (N_1893,N_1765,N_1727);
and U1894 (N_1894,N_1775,N_1782);
or U1895 (N_1895,N_1781,N_1745);
xnor U1896 (N_1896,N_1780,N_1750);
or U1897 (N_1897,N_1720,N_1730);
nand U1898 (N_1898,N_1793,N_1714);
nor U1899 (N_1899,N_1760,N_1797);
xor U1900 (N_1900,N_1894,N_1823);
or U1901 (N_1901,N_1862,N_1825);
or U1902 (N_1902,N_1831,N_1834);
and U1903 (N_1903,N_1824,N_1801);
nor U1904 (N_1904,N_1870,N_1813);
nand U1905 (N_1905,N_1858,N_1871);
nand U1906 (N_1906,N_1890,N_1852);
nor U1907 (N_1907,N_1878,N_1895);
nor U1908 (N_1908,N_1836,N_1844);
nor U1909 (N_1909,N_1865,N_1807);
and U1910 (N_1910,N_1875,N_1816);
nor U1911 (N_1911,N_1872,N_1851);
nand U1912 (N_1912,N_1857,N_1841);
or U1913 (N_1913,N_1863,N_1887);
nor U1914 (N_1914,N_1873,N_1879);
and U1915 (N_1915,N_1883,N_1859);
or U1916 (N_1916,N_1888,N_1835);
nor U1917 (N_1917,N_1898,N_1810);
or U1918 (N_1918,N_1892,N_1820);
or U1919 (N_1919,N_1854,N_1848);
nand U1920 (N_1920,N_1847,N_1819);
nor U1921 (N_1921,N_1837,N_1866);
and U1922 (N_1922,N_1882,N_1803);
and U1923 (N_1923,N_1853,N_1849);
nor U1924 (N_1924,N_1829,N_1830);
nor U1925 (N_1925,N_1889,N_1864);
nor U1926 (N_1926,N_1869,N_1808);
and U1927 (N_1927,N_1891,N_1897);
or U1928 (N_1928,N_1884,N_1893);
or U1929 (N_1929,N_1868,N_1867);
or U1930 (N_1930,N_1881,N_1896);
xor U1931 (N_1931,N_1826,N_1809);
nand U1932 (N_1932,N_1805,N_1840);
xor U1933 (N_1933,N_1850,N_1806);
or U1934 (N_1934,N_1877,N_1885);
nand U1935 (N_1935,N_1839,N_1800);
and U1936 (N_1936,N_1833,N_1811);
nand U1937 (N_1937,N_1874,N_1802);
xnor U1938 (N_1938,N_1817,N_1818);
nand U1939 (N_1939,N_1832,N_1804);
and U1940 (N_1940,N_1822,N_1838);
or U1941 (N_1941,N_1876,N_1880);
nor U1942 (N_1942,N_1845,N_1842);
and U1943 (N_1943,N_1814,N_1827);
and U1944 (N_1944,N_1846,N_1821);
and U1945 (N_1945,N_1815,N_1860);
and U1946 (N_1946,N_1856,N_1828);
nand U1947 (N_1947,N_1886,N_1861);
and U1948 (N_1948,N_1899,N_1843);
nor U1949 (N_1949,N_1855,N_1812);
nor U1950 (N_1950,N_1810,N_1805);
or U1951 (N_1951,N_1800,N_1821);
nand U1952 (N_1952,N_1869,N_1812);
and U1953 (N_1953,N_1837,N_1895);
xnor U1954 (N_1954,N_1872,N_1808);
nor U1955 (N_1955,N_1884,N_1836);
xnor U1956 (N_1956,N_1827,N_1805);
or U1957 (N_1957,N_1886,N_1859);
nor U1958 (N_1958,N_1801,N_1854);
nand U1959 (N_1959,N_1856,N_1874);
or U1960 (N_1960,N_1805,N_1874);
nor U1961 (N_1961,N_1846,N_1849);
nand U1962 (N_1962,N_1864,N_1808);
xnor U1963 (N_1963,N_1877,N_1821);
or U1964 (N_1964,N_1855,N_1810);
or U1965 (N_1965,N_1863,N_1843);
nand U1966 (N_1966,N_1844,N_1826);
nor U1967 (N_1967,N_1895,N_1888);
xnor U1968 (N_1968,N_1805,N_1835);
and U1969 (N_1969,N_1884,N_1847);
nand U1970 (N_1970,N_1884,N_1883);
nand U1971 (N_1971,N_1880,N_1883);
nand U1972 (N_1972,N_1872,N_1870);
xnor U1973 (N_1973,N_1810,N_1834);
and U1974 (N_1974,N_1891,N_1863);
nand U1975 (N_1975,N_1858,N_1870);
or U1976 (N_1976,N_1836,N_1883);
nor U1977 (N_1977,N_1815,N_1847);
or U1978 (N_1978,N_1809,N_1843);
xnor U1979 (N_1979,N_1885,N_1863);
and U1980 (N_1980,N_1882,N_1861);
nor U1981 (N_1981,N_1871,N_1894);
nor U1982 (N_1982,N_1818,N_1866);
xor U1983 (N_1983,N_1814,N_1877);
or U1984 (N_1984,N_1886,N_1885);
nand U1985 (N_1985,N_1846,N_1890);
nor U1986 (N_1986,N_1888,N_1894);
or U1987 (N_1987,N_1806,N_1821);
or U1988 (N_1988,N_1847,N_1832);
and U1989 (N_1989,N_1885,N_1842);
nand U1990 (N_1990,N_1894,N_1840);
and U1991 (N_1991,N_1811,N_1835);
nand U1992 (N_1992,N_1859,N_1837);
nor U1993 (N_1993,N_1829,N_1843);
or U1994 (N_1994,N_1868,N_1846);
and U1995 (N_1995,N_1805,N_1889);
or U1996 (N_1996,N_1863,N_1803);
and U1997 (N_1997,N_1898,N_1812);
and U1998 (N_1998,N_1833,N_1887);
xnor U1999 (N_1999,N_1819,N_1808);
xnor U2000 (N_2000,N_1905,N_1980);
nor U2001 (N_2001,N_1940,N_1935);
and U2002 (N_2002,N_1941,N_1928);
nor U2003 (N_2003,N_1932,N_1904);
xnor U2004 (N_2004,N_1990,N_1957);
nor U2005 (N_2005,N_1988,N_1908);
nand U2006 (N_2006,N_1995,N_1927);
nor U2007 (N_2007,N_1969,N_1993);
nor U2008 (N_2008,N_1983,N_1944);
nor U2009 (N_2009,N_1966,N_1910);
and U2010 (N_2010,N_1919,N_1925);
nor U2011 (N_2011,N_1933,N_1909);
nor U2012 (N_2012,N_1970,N_1985);
and U2013 (N_2013,N_1955,N_1911);
and U2014 (N_2014,N_1939,N_1920);
nand U2015 (N_2015,N_1953,N_1916);
nor U2016 (N_2016,N_1930,N_1934);
nand U2017 (N_2017,N_1931,N_1949);
or U2018 (N_2018,N_1954,N_1947);
nand U2019 (N_2019,N_1915,N_1923);
and U2020 (N_2020,N_1964,N_1929);
nand U2021 (N_2021,N_1971,N_1978);
nand U2022 (N_2022,N_1981,N_1938);
nor U2023 (N_2023,N_1912,N_1979);
and U2024 (N_2024,N_1942,N_1976);
nor U2025 (N_2025,N_1913,N_1906);
nor U2026 (N_2026,N_1986,N_1921);
or U2027 (N_2027,N_1999,N_1907);
nand U2028 (N_2028,N_1922,N_1958);
nor U2029 (N_2029,N_1902,N_1950);
nor U2030 (N_2030,N_1997,N_1961);
nand U2031 (N_2031,N_1963,N_1984);
xnor U2032 (N_2032,N_1926,N_1977);
nor U2033 (N_2033,N_1918,N_1974);
nor U2034 (N_2034,N_1924,N_1914);
or U2035 (N_2035,N_1968,N_1967);
or U2036 (N_2036,N_1989,N_1901);
nand U2037 (N_2037,N_1998,N_1945);
nor U2038 (N_2038,N_1946,N_1917);
or U2039 (N_2039,N_1975,N_1972);
nand U2040 (N_2040,N_1965,N_1943);
or U2041 (N_2041,N_1937,N_1996);
nand U2042 (N_2042,N_1982,N_1903);
nor U2043 (N_2043,N_1973,N_1987);
nand U2044 (N_2044,N_1952,N_1956);
and U2045 (N_2045,N_1948,N_1994);
or U2046 (N_2046,N_1960,N_1959);
and U2047 (N_2047,N_1936,N_1992);
xnor U2048 (N_2048,N_1900,N_1962);
nor U2049 (N_2049,N_1951,N_1991);
nand U2050 (N_2050,N_1934,N_1923);
and U2051 (N_2051,N_1993,N_1990);
and U2052 (N_2052,N_1911,N_1994);
or U2053 (N_2053,N_1906,N_1927);
xor U2054 (N_2054,N_1937,N_1913);
or U2055 (N_2055,N_1963,N_1962);
and U2056 (N_2056,N_1926,N_1921);
xor U2057 (N_2057,N_1935,N_1961);
xnor U2058 (N_2058,N_1993,N_1903);
and U2059 (N_2059,N_1948,N_1901);
or U2060 (N_2060,N_1908,N_1914);
xor U2061 (N_2061,N_1911,N_1962);
and U2062 (N_2062,N_1922,N_1949);
nor U2063 (N_2063,N_1975,N_1950);
nand U2064 (N_2064,N_1928,N_1931);
nand U2065 (N_2065,N_1927,N_1973);
or U2066 (N_2066,N_1987,N_1929);
and U2067 (N_2067,N_1977,N_1956);
and U2068 (N_2068,N_1941,N_1965);
and U2069 (N_2069,N_1968,N_1991);
and U2070 (N_2070,N_1982,N_1950);
nand U2071 (N_2071,N_1958,N_1901);
and U2072 (N_2072,N_1901,N_1943);
nor U2073 (N_2073,N_1997,N_1996);
or U2074 (N_2074,N_1934,N_1945);
and U2075 (N_2075,N_1951,N_1963);
nand U2076 (N_2076,N_1944,N_1916);
and U2077 (N_2077,N_1998,N_1926);
nand U2078 (N_2078,N_1938,N_1952);
and U2079 (N_2079,N_1904,N_1974);
nor U2080 (N_2080,N_1976,N_1968);
and U2081 (N_2081,N_1981,N_1908);
nand U2082 (N_2082,N_1917,N_1919);
and U2083 (N_2083,N_1936,N_1987);
or U2084 (N_2084,N_1993,N_1922);
and U2085 (N_2085,N_1976,N_1982);
and U2086 (N_2086,N_1954,N_1958);
nand U2087 (N_2087,N_1975,N_1981);
xnor U2088 (N_2088,N_1958,N_1920);
or U2089 (N_2089,N_1960,N_1907);
nor U2090 (N_2090,N_1991,N_1942);
xor U2091 (N_2091,N_1948,N_1900);
xor U2092 (N_2092,N_1962,N_1959);
xnor U2093 (N_2093,N_1982,N_1925);
nand U2094 (N_2094,N_1982,N_1927);
nand U2095 (N_2095,N_1922,N_1956);
or U2096 (N_2096,N_1913,N_1953);
and U2097 (N_2097,N_1977,N_1949);
and U2098 (N_2098,N_1958,N_1933);
or U2099 (N_2099,N_1925,N_1936);
nand U2100 (N_2100,N_2006,N_2077);
and U2101 (N_2101,N_2016,N_2010);
nor U2102 (N_2102,N_2002,N_2045);
or U2103 (N_2103,N_2086,N_2065);
or U2104 (N_2104,N_2051,N_2081);
nor U2105 (N_2105,N_2091,N_2030);
nor U2106 (N_2106,N_2056,N_2035);
and U2107 (N_2107,N_2079,N_2022);
xnor U2108 (N_2108,N_2037,N_2026);
xnor U2109 (N_2109,N_2089,N_2067);
nor U2110 (N_2110,N_2025,N_2049);
nand U2111 (N_2111,N_2044,N_2012);
and U2112 (N_2112,N_2092,N_2073);
and U2113 (N_2113,N_2011,N_2083);
xor U2114 (N_2114,N_2075,N_2059);
nor U2115 (N_2115,N_2034,N_2048);
nand U2116 (N_2116,N_2043,N_2036);
nand U2117 (N_2117,N_2095,N_2096);
xor U2118 (N_2118,N_2020,N_2098);
or U2119 (N_2119,N_2021,N_2064);
nor U2120 (N_2120,N_2009,N_2015);
and U2121 (N_2121,N_2018,N_2046);
or U2122 (N_2122,N_2099,N_2023);
and U2123 (N_2123,N_2008,N_2066);
nor U2124 (N_2124,N_2052,N_2063);
or U2125 (N_2125,N_2074,N_2014);
and U2126 (N_2126,N_2071,N_2004);
nand U2127 (N_2127,N_2039,N_2076);
nand U2128 (N_2128,N_2017,N_2001);
and U2129 (N_2129,N_2060,N_2032);
nand U2130 (N_2130,N_2024,N_2055);
xnor U2131 (N_2131,N_2061,N_2078);
nor U2132 (N_2132,N_2028,N_2003);
or U2133 (N_2133,N_2072,N_2038);
or U2134 (N_2134,N_2040,N_2084);
or U2135 (N_2135,N_2062,N_2013);
xor U2136 (N_2136,N_2093,N_2042);
nor U2137 (N_2137,N_2094,N_2031);
or U2138 (N_2138,N_2090,N_2033);
xnor U2139 (N_2139,N_2050,N_2082);
xnor U2140 (N_2140,N_2097,N_2041);
nor U2141 (N_2141,N_2088,N_2047);
nor U2142 (N_2142,N_2053,N_2027);
nor U2143 (N_2143,N_2080,N_2058);
nor U2144 (N_2144,N_2085,N_2029);
and U2145 (N_2145,N_2054,N_2068);
nand U2146 (N_2146,N_2087,N_2057);
nor U2147 (N_2147,N_2000,N_2019);
and U2148 (N_2148,N_2070,N_2007);
and U2149 (N_2149,N_2069,N_2005);
or U2150 (N_2150,N_2016,N_2074);
and U2151 (N_2151,N_2057,N_2007);
nor U2152 (N_2152,N_2052,N_2003);
and U2153 (N_2153,N_2047,N_2003);
nor U2154 (N_2154,N_2080,N_2022);
nor U2155 (N_2155,N_2071,N_2000);
nor U2156 (N_2156,N_2087,N_2074);
nand U2157 (N_2157,N_2034,N_2043);
nand U2158 (N_2158,N_2060,N_2093);
nor U2159 (N_2159,N_2009,N_2094);
and U2160 (N_2160,N_2013,N_2026);
nor U2161 (N_2161,N_2088,N_2024);
and U2162 (N_2162,N_2092,N_2052);
nand U2163 (N_2163,N_2001,N_2090);
or U2164 (N_2164,N_2037,N_2002);
and U2165 (N_2165,N_2002,N_2010);
or U2166 (N_2166,N_2003,N_2066);
and U2167 (N_2167,N_2002,N_2042);
or U2168 (N_2168,N_2036,N_2087);
and U2169 (N_2169,N_2080,N_2024);
nor U2170 (N_2170,N_2029,N_2055);
and U2171 (N_2171,N_2077,N_2031);
nand U2172 (N_2172,N_2082,N_2045);
and U2173 (N_2173,N_2068,N_2058);
nand U2174 (N_2174,N_2057,N_2097);
xor U2175 (N_2175,N_2089,N_2021);
nor U2176 (N_2176,N_2036,N_2062);
nand U2177 (N_2177,N_2095,N_2099);
nand U2178 (N_2178,N_2044,N_2091);
nand U2179 (N_2179,N_2093,N_2032);
nor U2180 (N_2180,N_2068,N_2031);
xnor U2181 (N_2181,N_2088,N_2015);
nand U2182 (N_2182,N_2000,N_2045);
nor U2183 (N_2183,N_2088,N_2032);
or U2184 (N_2184,N_2058,N_2046);
or U2185 (N_2185,N_2023,N_2051);
and U2186 (N_2186,N_2081,N_2096);
nand U2187 (N_2187,N_2038,N_2046);
and U2188 (N_2188,N_2067,N_2001);
and U2189 (N_2189,N_2073,N_2058);
and U2190 (N_2190,N_2011,N_2004);
nor U2191 (N_2191,N_2070,N_2050);
xnor U2192 (N_2192,N_2050,N_2048);
nand U2193 (N_2193,N_2013,N_2006);
or U2194 (N_2194,N_2088,N_2073);
nor U2195 (N_2195,N_2063,N_2027);
and U2196 (N_2196,N_2004,N_2017);
nand U2197 (N_2197,N_2024,N_2062);
or U2198 (N_2198,N_2008,N_2007);
nand U2199 (N_2199,N_2021,N_2006);
or U2200 (N_2200,N_2185,N_2163);
or U2201 (N_2201,N_2195,N_2194);
nand U2202 (N_2202,N_2177,N_2132);
nand U2203 (N_2203,N_2102,N_2196);
nand U2204 (N_2204,N_2174,N_2123);
and U2205 (N_2205,N_2161,N_2158);
nand U2206 (N_2206,N_2188,N_2138);
nand U2207 (N_2207,N_2153,N_2110);
nor U2208 (N_2208,N_2159,N_2179);
nor U2209 (N_2209,N_2128,N_2108);
xnor U2210 (N_2210,N_2180,N_2100);
and U2211 (N_2211,N_2183,N_2125);
nor U2212 (N_2212,N_2109,N_2107);
nand U2213 (N_2213,N_2145,N_2127);
and U2214 (N_2214,N_2117,N_2149);
nand U2215 (N_2215,N_2137,N_2119);
nor U2216 (N_2216,N_2199,N_2198);
and U2217 (N_2217,N_2131,N_2167);
xor U2218 (N_2218,N_2178,N_2171);
and U2219 (N_2219,N_2134,N_2186);
nand U2220 (N_2220,N_2106,N_2111);
and U2221 (N_2221,N_2120,N_2165);
or U2222 (N_2222,N_2187,N_2126);
xor U2223 (N_2223,N_2113,N_2172);
and U2224 (N_2224,N_2193,N_2160);
or U2225 (N_2225,N_2155,N_2115);
or U2226 (N_2226,N_2118,N_2147);
and U2227 (N_2227,N_2122,N_2129);
nand U2228 (N_2228,N_2103,N_2169);
or U2229 (N_2229,N_2150,N_2139);
or U2230 (N_2230,N_2173,N_2144);
and U2231 (N_2231,N_2175,N_2116);
and U2232 (N_2232,N_2192,N_2141);
nor U2233 (N_2233,N_2176,N_2162);
or U2234 (N_2234,N_2136,N_2140);
or U2235 (N_2235,N_2189,N_2143);
or U2236 (N_2236,N_2154,N_2182);
or U2237 (N_2237,N_2114,N_2121);
or U2238 (N_2238,N_2124,N_2148);
nand U2239 (N_2239,N_2184,N_2152);
nor U2240 (N_2240,N_2104,N_2166);
and U2241 (N_2241,N_2105,N_2170);
nor U2242 (N_2242,N_2157,N_2101);
or U2243 (N_2243,N_2197,N_2164);
nor U2244 (N_2244,N_2135,N_2133);
nand U2245 (N_2245,N_2142,N_2190);
or U2246 (N_2246,N_2151,N_2191);
nor U2247 (N_2247,N_2181,N_2130);
and U2248 (N_2248,N_2146,N_2112);
nand U2249 (N_2249,N_2156,N_2168);
and U2250 (N_2250,N_2177,N_2113);
nand U2251 (N_2251,N_2109,N_2144);
or U2252 (N_2252,N_2113,N_2160);
or U2253 (N_2253,N_2147,N_2122);
nor U2254 (N_2254,N_2110,N_2128);
or U2255 (N_2255,N_2199,N_2183);
or U2256 (N_2256,N_2156,N_2141);
nand U2257 (N_2257,N_2174,N_2109);
nor U2258 (N_2258,N_2197,N_2177);
and U2259 (N_2259,N_2143,N_2190);
nor U2260 (N_2260,N_2135,N_2175);
nor U2261 (N_2261,N_2187,N_2160);
xnor U2262 (N_2262,N_2158,N_2180);
or U2263 (N_2263,N_2141,N_2105);
or U2264 (N_2264,N_2107,N_2121);
and U2265 (N_2265,N_2110,N_2147);
nor U2266 (N_2266,N_2119,N_2199);
and U2267 (N_2267,N_2117,N_2163);
or U2268 (N_2268,N_2186,N_2135);
or U2269 (N_2269,N_2101,N_2107);
nand U2270 (N_2270,N_2154,N_2189);
nand U2271 (N_2271,N_2131,N_2136);
and U2272 (N_2272,N_2199,N_2112);
nor U2273 (N_2273,N_2165,N_2176);
nor U2274 (N_2274,N_2121,N_2148);
nor U2275 (N_2275,N_2113,N_2123);
or U2276 (N_2276,N_2183,N_2177);
or U2277 (N_2277,N_2123,N_2117);
or U2278 (N_2278,N_2104,N_2119);
or U2279 (N_2279,N_2139,N_2125);
nor U2280 (N_2280,N_2116,N_2168);
xor U2281 (N_2281,N_2124,N_2133);
and U2282 (N_2282,N_2110,N_2181);
nor U2283 (N_2283,N_2177,N_2164);
or U2284 (N_2284,N_2185,N_2186);
or U2285 (N_2285,N_2112,N_2190);
nand U2286 (N_2286,N_2128,N_2180);
and U2287 (N_2287,N_2120,N_2138);
or U2288 (N_2288,N_2125,N_2188);
or U2289 (N_2289,N_2105,N_2190);
nor U2290 (N_2290,N_2148,N_2157);
nor U2291 (N_2291,N_2116,N_2152);
nand U2292 (N_2292,N_2157,N_2166);
xor U2293 (N_2293,N_2188,N_2126);
nor U2294 (N_2294,N_2137,N_2123);
nand U2295 (N_2295,N_2137,N_2145);
xnor U2296 (N_2296,N_2146,N_2158);
nand U2297 (N_2297,N_2128,N_2193);
and U2298 (N_2298,N_2152,N_2155);
or U2299 (N_2299,N_2108,N_2164);
or U2300 (N_2300,N_2245,N_2284);
nand U2301 (N_2301,N_2252,N_2225);
nand U2302 (N_2302,N_2261,N_2213);
or U2303 (N_2303,N_2275,N_2292);
nor U2304 (N_2304,N_2204,N_2203);
or U2305 (N_2305,N_2217,N_2264);
nand U2306 (N_2306,N_2297,N_2212);
and U2307 (N_2307,N_2250,N_2243);
xor U2308 (N_2308,N_2242,N_2223);
and U2309 (N_2309,N_2287,N_2262);
nand U2310 (N_2310,N_2282,N_2201);
or U2311 (N_2311,N_2230,N_2236);
nand U2312 (N_2312,N_2229,N_2226);
nor U2313 (N_2313,N_2258,N_2294);
nand U2314 (N_2314,N_2221,N_2268);
xnor U2315 (N_2315,N_2231,N_2214);
or U2316 (N_2316,N_2205,N_2234);
or U2317 (N_2317,N_2259,N_2291);
nor U2318 (N_2318,N_2215,N_2202);
xor U2319 (N_2319,N_2219,N_2273);
nand U2320 (N_2320,N_2255,N_2286);
xnor U2321 (N_2321,N_2228,N_2299);
nand U2322 (N_2322,N_2295,N_2239);
nor U2323 (N_2323,N_2241,N_2269);
and U2324 (N_2324,N_2224,N_2220);
xnor U2325 (N_2325,N_2267,N_2288);
nor U2326 (N_2326,N_2266,N_2251);
or U2327 (N_2327,N_2209,N_2263);
nor U2328 (N_2328,N_2277,N_2208);
or U2329 (N_2329,N_2207,N_2274);
or U2330 (N_2330,N_2281,N_2270);
nor U2331 (N_2331,N_2237,N_2246);
nand U2332 (N_2332,N_2260,N_2227);
xnor U2333 (N_2333,N_2222,N_2200);
xor U2334 (N_2334,N_2265,N_2211);
or U2335 (N_2335,N_2232,N_2279);
and U2336 (N_2336,N_2283,N_2210);
nand U2337 (N_2337,N_2233,N_2248);
nor U2338 (N_2338,N_2296,N_2280);
xnor U2339 (N_2339,N_2249,N_2216);
nor U2340 (N_2340,N_2240,N_2285);
xnor U2341 (N_2341,N_2278,N_2254);
nor U2342 (N_2342,N_2298,N_2276);
or U2343 (N_2343,N_2206,N_2290);
and U2344 (N_2344,N_2244,N_2272);
and U2345 (N_2345,N_2256,N_2247);
and U2346 (N_2346,N_2218,N_2289);
and U2347 (N_2347,N_2271,N_2257);
nand U2348 (N_2348,N_2238,N_2293);
xnor U2349 (N_2349,N_2253,N_2235);
nand U2350 (N_2350,N_2260,N_2271);
or U2351 (N_2351,N_2285,N_2283);
nor U2352 (N_2352,N_2249,N_2204);
nor U2353 (N_2353,N_2205,N_2213);
or U2354 (N_2354,N_2251,N_2203);
or U2355 (N_2355,N_2259,N_2241);
or U2356 (N_2356,N_2258,N_2212);
nand U2357 (N_2357,N_2262,N_2293);
nand U2358 (N_2358,N_2245,N_2250);
and U2359 (N_2359,N_2245,N_2287);
or U2360 (N_2360,N_2205,N_2235);
nand U2361 (N_2361,N_2290,N_2201);
nand U2362 (N_2362,N_2247,N_2214);
and U2363 (N_2363,N_2283,N_2270);
and U2364 (N_2364,N_2274,N_2267);
nor U2365 (N_2365,N_2224,N_2274);
nor U2366 (N_2366,N_2216,N_2280);
and U2367 (N_2367,N_2281,N_2283);
nor U2368 (N_2368,N_2224,N_2233);
nand U2369 (N_2369,N_2299,N_2234);
and U2370 (N_2370,N_2201,N_2297);
or U2371 (N_2371,N_2271,N_2217);
and U2372 (N_2372,N_2256,N_2252);
nand U2373 (N_2373,N_2273,N_2298);
nor U2374 (N_2374,N_2249,N_2271);
nand U2375 (N_2375,N_2258,N_2291);
and U2376 (N_2376,N_2255,N_2260);
and U2377 (N_2377,N_2272,N_2263);
xor U2378 (N_2378,N_2216,N_2299);
and U2379 (N_2379,N_2252,N_2205);
xnor U2380 (N_2380,N_2291,N_2265);
or U2381 (N_2381,N_2294,N_2281);
xnor U2382 (N_2382,N_2266,N_2230);
nand U2383 (N_2383,N_2224,N_2211);
nand U2384 (N_2384,N_2240,N_2292);
or U2385 (N_2385,N_2298,N_2210);
nor U2386 (N_2386,N_2244,N_2270);
xor U2387 (N_2387,N_2231,N_2295);
xor U2388 (N_2388,N_2217,N_2230);
or U2389 (N_2389,N_2230,N_2222);
and U2390 (N_2390,N_2277,N_2283);
and U2391 (N_2391,N_2263,N_2253);
or U2392 (N_2392,N_2251,N_2243);
nor U2393 (N_2393,N_2253,N_2225);
nor U2394 (N_2394,N_2216,N_2206);
or U2395 (N_2395,N_2227,N_2217);
nand U2396 (N_2396,N_2223,N_2239);
nand U2397 (N_2397,N_2240,N_2260);
nor U2398 (N_2398,N_2223,N_2200);
or U2399 (N_2399,N_2216,N_2236);
or U2400 (N_2400,N_2367,N_2384);
or U2401 (N_2401,N_2358,N_2330);
or U2402 (N_2402,N_2347,N_2332);
nand U2403 (N_2403,N_2397,N_2307);
xor U2404 (N_2404,N_2351,N_2343);
or U2405 (N_2405,N_2385,N_2338);
and U2406 (N_2406,N_2304,N_2339);
or U2407 (N_2407,N_2378,N_2300);
or U2408 (N_2408,N_2366,N_2323);
nor U2409 (N_2409,N_2383,N_2348);
and U2410 (N_2410,N_2342,N_2381);
xnor U2411 (N_2411,N_2318,N_2377);
nand U2412 (N_2412,N_2370,N_2329);
or U2413 (N_2413,N_2368,N_2324);
nor U2414 (N_2414,N_2306,N_2305);
xnor U2415 (N_2415,N_2387,N_2311);
nor U2416 (N_2416,N_2372,N_2398);
nor U2417 (N_2417,N_2389,N_2321);
nor U2418 (N_2418,N_2317,N_2341);
and U2419 (N_2419,N_2392,N_2325);
and U2420 (N_2420,N_2380,N_2308);
nor U2421 (N_2421,N_2312,N_2359);
nor U2422 (N_2422,N_2388,N_2399);
nor U2423 (N_2423,N_2369,N_2357);
and U2424 (N_2424,N_2350,N_2393);
nor U2425 (N_2425,N_2360,N_2349);
nand U2426 (N_2426,N_2365,N_2379);
xnor U2427 (N_2427,N_2303,N_2382);
nand U2428 (N_2428,N_2395,N_2322);
and U2429 (N_2429,N_2344,N_2313);
nor U2430 (N_2430,N_2354,N_2327);
or U2431 (N_2431,N_2364,N_2375);
and U2432 (N_2432,N_2374,N_2386);
or U2433 (N_2433,N_2319,N_2363);
and U2434 (N_2434,N_2335,N_2328);
and U2435 (N_2435,N_2326,N_2315);
and U2436 (N_2436,N_2391,N_2356);
and U2437 (N_2437,N_2352,N_2346);
nand U2438 (N_2438,N_2336,N_2310);
and U2439 (N_2439,N_2345,N_2337);
or U2440 (N_2440,N_2316,N_2334);
xor U2441 (N_2441,N_2373,N_2390);
or U2442 (N_2442,N_2394,N_2340);
nor U2443 (N_2443,N_2302,N_2361);
or U2444 (N_2444,N_2314,N_2355);
nor U2445 (N_2445,N_2309,N_2353);
nand U2446 (N_2446,N_2371,N_2331);
nor U2447 (N_2447,N_2362,N_2320);
nor U2448 (N_2448,N_2376,N_2396);
xnor U2449 (N_2449,N_2301,N_2333);
or U2450 (N_2450,N_2348,N_2301);
nand U2451 (N_2451,N_2300,N_2306);
nor U2452 (N_2452,N_2309,N_2368);
xor U2453 (N_2453,N_2319,N_2338);
xor U2454 (N_2454,N_2356,N_2390);
or U2455 (N_2455,N_2330,N_2393);
nand U2456 (N_2456,N_2308,N_2393);
nor U2457 (N_2457,N_2310,N_2300);
xor U2458 (N_2458,N_2387,N_2310);
and U2459 (N_2459,N_2324,N_2389);
xnor U2460 (N_2460,N_2391,N_2304);
nor U2461 (N_2461,N_2326,N_2316);
and U2462 (N_2462,N_2362,N_2391);
and U2463 (N_2463,N_2318,N_2365);
nand U2464 (N_2464,N_2399,N_2347);
nand U2465 (N_2465,N_2334,N_2331);
nor U2466 (N_2466,N_2368,N_2375);
or U2467 (N_2467,N_2359,N_2344);
and U2468 (N_2468,N_2348,N_2382);
nand U2469 (N_2469,N_2348,N_2381);
and U2470 (N_2470,N_2330,N_2327);
nand U2471 (N_2471,N_2386,N_2354);
nand U2472 (N_2472,N_2383,N_2341);
or U2473 (N_2473,N_2308,N_2365);
nand U2474 (N_2474,N_2390,N_2352);
nand U2475 (N_2475,N_2320,N_2359);
nand U2476 (N_2476,N_2320,N_2318);
xnor U2477 (N_2477,N_2300,N_2374);
nand U2478 (N_2478,N_2340,N_2381);
and U2479 (N_2479,N_2355,N_2388);
or U2480 (N_2480,N_2344,N_2354);
nand U2481 (N_2481,N_2335,N_2318);
and U2482 (N_2482,N_2365,N_2315);
and U2483 (N_2483,N_2310,N_2368);
and U2484 (N_2484,N_2307,N_2391);
nand U2485 (N_2485,N_2309,N_2330);
or U2486 (N_2486,N_2395,N_2367);
nor U2487 (N_2487,N_2327,N_2335);
nor U2488 (N_2488,N_2353,N_2369);
and U2489 (N_2489,N_2332,N_2325);
and U2490 (N_2490,N_2361,N_2307);
or U2491 (N_2491,N_2353,N_2333);
and U2492 (N_2492,N_2393,N_2366);
or U2493 (N_2493,N_2396,N_2344);
and U2494 (N_2494,N_2336,N_2314);
nor U2495 (N_2495,N_2348,N_2358);
nor U2496 (N_2496,N_2362,N_2313);
nand U2497 (N_2497,N_2365,N_2321);
and U2498 (N_2498,N_2330,N_2336);
xnor U2499 (N_2499,N_2367,N_2325);
and U2500 (N_2500,N_2411,N_2417);
and U2501 (N_2501,N_2459,N_2471);
and U2502 (N_2502,N_2447,N_2463);
nand U2503 (N_2503,N_2437,N_2433);
nor U2504 (N_2504,N_2413,N_2421);
or U2505 (N_2505,N_2431,N_2462);
xnor U2506 (N_2506,N_2434,N_2448);
nand U2507 (N_2507,N_2493,N_2477);
and U2508 (N_2508,N_2481,N_2478);
nor U2509 (N_2509,N_2440,N_2479);
and U2510 (N_2510,N_2427,N_2465);
and U2511 (N_2511,N_2484,N_2457);
nand U2512 (N_2512,N_2424,N_2451);
or U2513 (N_2513,N_2470,N_2419);
or U2514 (N_2514,N_2499,N_2405);
nand U2515 (N_2515,N_2444,N_2497);
xnor U2516 (N_2516,N_2488,N_2400);
nor U2517 (N_2517,N_2487,N_2414);
nor U2518 (N_2518,N_2408,N_2452);
xnor U2519 (N_2519,N_2468,N_2423);
or U2520 (N_2520,N_2415,N_2435);
nand U2521 (N_2521,N_2456,N_2475);
nor U2522 (N_2522,N_2403,N_2445);
and U2523 (N_2523,N_2474,N_2443);
and U2524 (N_2524,N_2401,N_2428);
or U2525 (N_2525,N_2438,N_2409);
nand U2526 (N_2526,N_2422,N_2496);
nor U2527 (N_2527,N_2402,N_2426);
nor U2528 (N_2528,N_2432,N_2489);
xor U2529 (N_2529,N_2454,N_2467);
xnor U2530 (N_2530,N_2450,N_2461);
and U2531 (N_2531,N_2404,N_2472);
xor U2532 (N_2532,N_2483,N_2486);
nand U2533 (N_2533,N_2416,N_2498);
nand U2534 (N_2534,N_2418,N_2466);
or U2535 (N_2535,N_2407,N_2410);
nand U2536 (N_2536,N_2491,N_2485);
nor U2537 (N_2537,N_2420,N_2436);
nand U2538 (N_2538,N_2425,N_2476);
nand U2539 (N_2539,N_2406,N_2469);
nor U2540 (N_2540,N_2429,N_2439);
and U2541 (N_2541,N_2460,N_2482);
nor U2542 (N_2542,N_2453,N_2441);
nor U2543 (N_2543,N_2412,N_2455);
or U2544 (N_2544,N_2446,N_2449);
nand U2545 (N_2545,N_2480,N_2464);
nand U2546 (N_2546,N_2430,N_2458);
nor U2547 (N_2547,N_2490,N_2495);
nand U2548 (N_2548,N_2442,N_2494);
and U2549 (N_2549,N_2492,N_2473);
nand U2550 (N_2550,N_2461,N_2414);
or U2551 (N_2551,N_2478,N_2461);
xor U2552 (N_2552,N_2453,N_2486);
xnor U2553 (N_2553,N_2433,N_2492);
and U2554 (N_2554,N_2407,N_2472);
and U2555 (N_2555,N_2450,N_2483);
nor U2556 (N_2556,N_2402,N_2478);
or U2557 (N_2557,N_2414,N_2416);
nand U2558 (N_2558,N_2466,N_2414);
xor U2559 (N_2559,N_2495,N_2411);
or U2560 (N_2560,N_2431,N_2427);
and U2561 (N_2561,N_2415,N_2472);
nand U2562 (N_2562,N_2452,N_2419);
nor U2563 (N_2563,N_2447,N_2466);
nor U2564 (N_2564,N_2403,N_2488);
nor U2565 (N_2565,N_2452,N_2435);
or U2566 (N_2566,N_2460,N_2487);
nor U2567 (N_2567,N_2460,N_2434);
nand U2568 (N_2568,N_2414,N_2425);
or U2569 (N_2569,N_2497,N_2455);
and U2570 (N_2570,N_2407,N_2420);
nand U2571 (N_2571,N_2400,N_2481);
nor U2572 (N_2572,N_2427,N_2437);
nand U2573 (N_2573,N_2443,N_2459);
and U2574 (N_2574,N_2479,N_2468);
and U2575 (N_2575,N_2433,N_2420);
nand U2576 (N_2576,N_2416,N_2456);
xor U2577 (N_2577,N_2463,N_2458);
xnor U2578 (N_2578,N_2464,N_2434);
nand U2579 (N_2579,N_2445,N_2428);
nor U2580 (N_2580,N_2452,N_2418);
xnor U2581 (N_2581,N_2406,N_2482);
nand U2582 (N_2582,N_2471,N_2498);
or U2583 (N_2583,N_2409,N_2450);
nand U2584 (N_2584,N_2460,N_2426);
and U2585 (N_2585,N_2415,N_2448);
nor U2586 (N_2586,N_2417,N_2479);
nor U2587 (N_2587,N_2484,N_2495);
nor U2588 (N_2588,N_2402,N_2484);
and U2589 (N_2589,N_2498,N_2460);
or U2590 (N_2590,N_2445,N_2488);
nand U2591 (N_2591,N_2447,N_2443);
nor U2592 (N_2592,N_2406,N_2497);
or U2593 (N_2593,N_2423,N_2410);
xnor U2594 (N_2594,N_2487,N_2453);
xor U2595 (N_2595,N_2459,N_2479);
nor U2596 (N_2596,N_2480,N_2430);
and U2597 (N_2597,N_2468,N_2431);
nand U2598 (N_2598,N_2401,N_2494);
nand U2599 (N_2599,N_2477,N_2424);
and U2600 (N_2600,N_2594,N_2574);
nand U2601 (N_2601,N_2581,N_2569);
xor U2602 (N_2602,N_2590,N_2500);
nor U2603 (N_2603,N_2522,N_2504);
nor U2604 (N_2604,N_2591,N_2538);
xnor U2605 (N_2605,N_2584,N_2518);
nand U2606 (N_2606,N_2524,N_2544);
nand U2607 (N_2607,N_2552,N_2516);
or U2608 (N_2608,N_2567,N_2558);
nand U2609 (N_2609,N_2572,N_2585);
and U2610 (N_2610,N_2543,N_2551);
nand U2611 (N_2611,N_2555,N_2531);
and U2612 (N_2612,N_2545,N_2530);
or U2613 (N_2613,N_2534,N_2562);
and U2614 (N_2614,N_2507,N_2539);
nand U2615 (N_2615,N_2592,N_2570);
or U2616 (N_2616,N_2580,N_2533);
nand U2617 (N_2617,N_2532,N_2564);
or U2618 (N_2618,N_2514,N_2525);
or U2619 (N_2619,N_2557,N_2578);
and U2620 (N_2620,N_2583,N_2573);
nand U2621 (N_2621,N_2517,N_2576);
nor U2622 (N_2622,N_2535,N_2561);
or U2623 (N_2623,N_2589,N_2515);
nor U2624 (N_2624,N_2527,N_2502);
or U2625 (N_2625,N_2537,N_2529);
or U2626 (N_2626,N_2521,N_2560);
nor U2627 (N_2627,N_2526,N_2553);
xnor U2628 (N_2628,N_2501,N_2520);
and U2629 (N_2629,N_2565,N_2509);
nand U2630 (N_2630,N_2566,N_2575);
nor U2631 (N_2631,N_2512,N_2579);
or U2632 (N_2632,N_2546,N_2554);
nand U2633 (N_2633,N_2528,N_2547);
nor U2634 (N_2634,N_2568,N_2548);
nand U2635 (N_2635,N_2536,N_2556);
nor U2636 (N_2636,N_2540,N_2588);
or U2637 (N_2637,N_2519,N_2511);
or U2638 (N_2638,N_2593,N_2510);
or U2639 (N_2639,N_2563,N_2596);
nor U2640 (N_2640,N_2599,N_2503);
nand U2641 (N_2641,N_2542,N_2577);
or U2642 (N_2642,N_2550,N_2541);
or U2643 (N_2643,N_2587,N_2549);
nor U2644 (N_2644,N_2597,N_2571);
or U2645 (N_2645,N_2523,N_2595);
nand U2646 (N_2646,N_2559,N_2513);
or U2647 (N_2647,N_2582,N_2508);
nor U2648 (N_2648,N_2505,N_2506);
or U2649 (N_2649,N_2586,N_2598);
or U2650 (N_2650,N_2594,N_2504);
nand U2651 (N_2651,N_2526,N_2516);
or U2652 (N_2652,N_2500,N_2532);
nor U2653 (N_2653,N_2544,N_2558);
and U2654 (N_2654,N_2547,N_2592);
nand U2655 (N_2655,N_2560,N_2551);
nand U2656 (N_2656,N_2544,N_2557);
nor U2657 (N_2657,N_2507,N_2592);
nor U2658 (N_2658,N_2555,N_2512);
nand U2659 (N_2659,N_2596,N_2568);
and U2660 (N_2660,N_2529,N_2575);
nand U2661 (N_2661,N_2536,N_2537);
nand U2662 (N_2662,N_2509,N_2555);
nand U2663 (N_2663,N_2549,N_2527);
or U2664 (N_2664,N_2584,N_2529);
nand U2665 (N_2665,N_2544,N_2563);
nand U2666 (N_2666,N_2527,N_2510);
or U2667 (N_2667,N_2591,N_2571);
nand U2668 (N_2668,N_2550,N_2543);
nor U2669 (N_2669,N_2547,N_2549);
or U2670 (N_2670,N_2570,N_2565);
or U2671 (N_2671,N_2575,N_2500);
and U2672 (N_2672,N_2508,N_2549);
or U2673 (N_2673,N_2528,N_2538);
nand U2674 (N_2674,N_2567,N_2535);
and U2675 (N_2675,N_2507,N_2594);
or U2676 (N_2676,N_2515,N_2523);
and U2677 (N_2677,N_2585,N_2584);
nand U2678 (N_2678,N_2566,N_2501);
nand U2679 (N_2679,N_2568,N_2555);
nand U2680 (N_2680,N_2535,N_2541);
nand U2681 (N_2681,N_2543,N_2576);
nor U2682 (N_2682,N_2598,N_2574);
nand U2683 (N_2683,N_2568,N_2517);
nor U2684 (N_2684,N_2544,N_2571);
or U2685 (N_2685,N_2556,N_2542);
xnor U2686 (N_2686,N_2530,N_2592);
or U2687 (N_2687,N_2516,N_2542);
or U2688 (N_2688,N_2547,N_2598);
or U2689 (N_2689,N_2567,N_2501);
or U2690 (N_2690,N_2538,N_2587);
or U2691 (N_2691,N_2537,N_2570);
nand U2692 (N_2692,N_2552,N_2595);
nor U2693 (N_2693,N_2522,N_2512);
nand U2694 (N_2694,N_2505,N_2527);
nor U2695 (N_2695,N_2589,N_2559);
nor U2696 (N_2696,N_2508,N_2551);
nand U2697 (N_2697,N_2583,N_2562);
and U2698 (N_2698,N_2593,N_2526);
and U2699 (N_2699,N_2570,N_2529);
and U2700 (N_2700,N_2641,N_2652);
and U2701 (N_2701,N_2677,N_2624);
or U2702 (N_2702,N_2671,N_2696);
or U2703 (N_2703,N_2619,N_2655);
or U2704 (N_2704,N_2664,N_2683);
xor U2705 (N_2705,N_2634,N_2632);
and U2706 (N_2706,N_2629,N_2697);
or U2707 (N_2707,N_2657,N_2605);
nand U2708 (N_2708,N_2653,N_2666);
and U2709 (N_2709,N_2693,N_2637);
or U2710 (N_2710,N_2680,N_2648);
nor U2711 (N_2711,N_2681,N_2670);
nor U2712 (N_2712,N_2631,N_2695);
nand U2713 (N_2713,N_2626,N_2674);
and U2714 (N_2714,N_2610,N_2668);
and U2715 (N_2715,N_2673,N_2614);
xnor U2716 (N_2716,N_2644,N_2620);
nand U2717 (N_2717,N_2609,N_2643);
and U2718 (N_2718,N_2690,N_2679);
or U2719 (N_2719,N_2633,N_2659);
nor U2720 (N_2720,N_2662,N_2667);
or U2721 (N_2721,N_2640,N_2685);
xor U2722 (N_2722,N_2694,N_2654);
or U2723 (N_2723,N_2621,N_2611);
or U2724 (N_2724,N_2617,N_2661);
xnor U2725 (N_2725,N_2636,N_2678);
and U2726 (N_2726,N_2630,N_2602);
nand U2727 (N_2727,N_2658,N_2608);
nand U2728 (N_2728,N_2606,N_2647);
or U2729 (N_2729,N_2600,N_2625);
and U2730 (N_2730,N_2687,N_2651);
and U2731 (N_2731,N_2627,N_2622);
nor U2732 (N_2732,N_2618,N_2688);
or U2733 (N_2733,N_2691,N_2639);
nand U2734 (N_2734,N_2603,N_2613);
nand U2735 (N_2735,N_2684,N_2689);
and U2736 (N_2736,N_2635,N_2604);
nand U2737 (N_2737,N_2645,N_2675);
and U2738 (N_2738,N_2616,N_2649);
and U2739 (N_2739,N_2665,N_2642);
xnor U2740 (N_2740,N_2628,N_2601);
nand U2741 (N_2741,N_2669,N_2686);
and U2742 (N_2742,N_2672,N_2650);
nor U2743 (N_2743,N_2682,N_2698);
nor U2744 (N_2744,N_2615,N_2692);
or U2745 (N_2745,N_2612,N_2660);
or U2746 (N_2746,N_2646,N_2699);
and U2747 (N_2747,N_2656,N_2607);
and U2748 (N_2748,N_2676,N_2623);
or U2749 (N_2749,N_2638,N_2663);
or U2750 (N_2750,N_2682,N_2686);
nand U2751 (N_2751,N_2648,N_2624);
nand U2752 (N_2752,N_2696,N_2609);
nand U2753 (N_2753,N_2612,N_2621);
and U2754 (N_2754,N_2603,N_2645);
or U2755 (N_2755,N_2613,N_2643);
xor U2756 (N_2756,N_2631,N_2654);
nor U2757 (N_2757,N_2654,N_2638);
nand U2758 (N_2758,N_2626,N_2678);
nand U2759 (N_2759,N_2666,N_2644);
nor U2760 (N_2760,N_2620,N_2693);
nor U2761 (N_2761,N_2630,N_2614);
nor U2762 (N_2762,N_2624,N_2689);
nor U2763 (N_2763,N_2607,N_2672);
nand U2764 (N_2764,N_2689,N_2670);
nand U2765 (N_2765,N_2697,N_2694);
nand U2766 (N_2766,N_2643,N_2631);
nor U2767 (N_2767,N_2664,N_2605);
and U2768 (N_2768,N_2600,N_2619);
or U2769 (N_2769,N_2652,N_2633);
and U2770 (N_2770,N_2692,N_2671);
and U2771 (N_2771,N_2680,N_2635);
and U2772 (N_2772,N_2626,N_2603);
or U2773 (N_2773,N_2630,N_2654);
or U2774 (N_2774,N_2691,N_2670);
or U2775 (N_2775,N_2657,N_2622);
or U2776 (N_2776,N_2600,N_2641);
nand U2777 (N_2777,N_2651,N_2674);
nand U2778 (N_2778,N_2621,N_2638);
or U2779 (N_2779,N_2687,N_2621);
nor U2780 (N_2780,N_2675,N_2609);
nand U2781 (N_2781,N_2602,N_2637);
nor U2782 (N_2782,N_2648,N_2679);
xnor U2783 (N_2783,N_2679,N_2617);
xnor U2784 (N_2784,N_2671,N_2661);
nor U2785 (N_2785,N_2682,N_2618);
and U2786 (N_2786,N_2666,N_2681);
and U2787 (N_2787,N_2604,N_2608);
or U2788 (N_2788,N_2693,N_2685);
nand U2789 (N_2789,N_2691,N_2692);
or U2790 (N_2790,N_2648,N_2654);
nor U2791 (N_2791,N_2651,N_2689);
nor U2792 (N_2792,N_2668,N_2639);
nor U2793 (N_2793,N_2683,N_2632);
nand U2794 (N_2794,N_2671,N_2609);
nor U2795 (N_2795,N_2618,N_2652);
nand U2796 (N_2796,N_2691,N_2611);
or U2797 (N_2797,N_2662,N_2697);
nand U2798 (N_2798,N_2674,N_2610);
nor U2799 (N_2799,N_2600,N_2662);
nor U2800 (N_2800,N_2798,N_2755);
nand U2801 (N_2801,N_2751,N_2780);
or U2802 (N_2802,N_2736,N_2759);
xnor U2803 (N_2803,N_2792,N_2797);
or U2804 (N_2804,N_2761,N_2764);
or U2805 (N_2805,N_2730,N_2776);
nor U2806 (N_2806,N_2735,N_2795);
or U2807 (N_2807,N_2744,N_2734);
or U2808 (N_2808,N_2785,N_2756);
or U2809 (N_2809,N_2724,N_2763);
or U2810 (N_2810,N_2741,N_2773);
nand U2811 (N_2811,N_2758,N_2746);
nand U2812 (N_2812,N_2700,N_2719);
nand U2813 (N_2813,N_2778,N_2771);
and U2814 (N_2814,N_2767,N_2768);
xor U2815 (N_2815,N_2718,N_2733);
nand U2816 (N_2816,N_2747,N_2743);
or U2817 (N_2817,N_2714,N_2715);
or U2818 (N_2818,N_2777,N_2721);
and U2819 (N_2819,N_2701,N_2799);
and U2820 (N_2820,N_2775,N_2706);
nor U2821 (N_2821,N_2765,N_2749);
nor U2822 (N_2822,N_2731,N_2716);
nor U2823 (N_2823,N_2791,N_2740);
or U2824 (N_2824,N_2769,N_2707);
nand U2825 (N_2825,N_2711,N_2781);
nand U2826 (N_2826,N_2748,N_2766);
or U2827 (N_2827,N_2722,N_2705);
and U2828 (N_2828,N_2782,N_2720);
nand U2829 (N_2829,N_2750,N_2774);
and U2830 (N_2830,N_2702,N_2784);
nor U2831 (N_2831,N_2772,N_2738);
nor U2832 (N_2832,N_2710,N_2796);
nor U2833 (N_2833,N_2723,N_2728);
nand U2834 (N_2834,N_2712,N_2783);
nand U2835 (N_2835,N_2788,N_2708);
nand U2836 (N_2836,N_2794,N_2745);
or U2837 (N_2837,N_2729,N_2704);
nor U2838 (N_2838,N_2760,N_2726);
nand U2839 (N_2839,N_2739,N_2770);
nand U2840 (N_2840,N_2779,N_2787);
xnor U2841 (N_2841,N_2757,N_2793);
nand U2842 (N_2842,N_2790,N_2742);
nor U2843 (N_2843,N_2789,N_2727);
nand U2844 (N_2844,N_2737,N_2709);
nor U2845 (N_2845,N_2713,N_2754);
nand U2846 (N_2846,N_2752,N_2732);
and U2847 (N_2847,N_2725,N_2762);
nand U2848 (N_2848,N_2703,N_2786);
or U2849 (N_2849,N_2717,N_2753);
nor U2850 (N_2850,N_2713,N_2742);
or U2851 (N_2851,N_2718,N_2737);
or U2852 (N_2852,N_2726,N_2705);
xor U2853 (N_2853,N_2700,N_2765);
or U2854 (N_2854,N_2793,N_2704);
and U2855 (N_2855,N_2792,N_2718);
or U2856 (N_2856,N_2711,N_2747);
nand U2857 (N_2857,N_2724,N_2717);
nor U2858 (N_2858,N_2773,N_2737);
or U2859 (N_2859,N_2704,N_2712);
nor U2860 (N_2860,N_2750,N_2773);
and U2861 (N_2861,N_2730,N_2784);
nand U2862 (N_2862,N_2737,N_2751);
nand U2863 (N_2863,N_2762,N_2711);
or U2864 (N_2864,N_2715,N_2798);
or U2865 (N_2865,N_2777,N_2764);
nor U2866 (N_2866,N_2769,N_2702);
xor U2867 (N_2867,N_2735,N_2758);
and U2868 (N_2868,N_2762,N_2759);
or U2869 (N_2869,N_2770,N_2757);
xnor U2870 (N_2870,N_2785,N_2781);
xnor U2871 (N_2871,N_2730,N_2734);
or U2872 (N_2872,N_2719,N_2785);
and U2873 (N_2873,N_2788,N_2725);
and U2874 (N_2874,N_2789,N_2765);
or U2875 (N_2875,N_2796,N_2752);
nand U2876 (N_2876,N_2795,N_2747);
nor U2877 (N_2877,N_2700,N_2749);
or U2878 (N_2878,N_2754,N_2703);
or U2879 (N_2879,N_2724,N_2721);
nand U2880 (N_2880,N_2778,N_2718);
and U2881 (N_2881,N_2708,N_2707);
nor U2882 (N_2882,N_2739,N_2748);
and U2883 (N_2883,N_2713,N_2722);
nor U2884 (N_2884,N_2734,N_2792);
and U2885 (N_2885,N_2738,N_2764);
xor U2886 (N_2886,N_2711,N_2797);
nand U2887 (N_2887,N_2735,N_2752);
and U2888 (N_2888,N_2791,N_2729);
nor U2889 (N_2889,N_2775,N_2789);
and U2890 (N_2890,N_2731,N_2717);
and U2891 (N_2891,N_2751,N_2791);
nor U2892 (N_2892,N_2764,N_2796);
and U2893 (N_2893,N_2734,N_2778);
nand U2894 (N_2894,N_2759,N_2763);
nor U2895 (N_2895,N_2776,N_2738);
or U2896 (N_2896,N_2737,N_2763);
and U2897 (N_2897,N_2767,N_2746);
and U2898 (N_2898,N_2724,N_2707);
or U2899 (N_2899,N_2745,N_2702);
nand U2900 (N_2900,N_2872,N_2827);
nand U2901 (N_2901,N_2886,N_2859);
nor U2902 (N_2902,N_2821,N_2894);
nor U2903 (N_2903,N_2858,N_2812);
nor U2904 (N_2904,N_2882,N_2829);
and U2905 (N_2905,N_2860,N_2855);
and U2906 (N_2906,N_2875,N_2834);
nor U2907 (N_2907,N_2801,N_2879);
or U2908 (N_2908,N_2848,N_2856);
nor U2909 (N_2909,N_2853,N_2805);
or U2910 (N_2910,N_2868,N_2840);
xor U2911 (N_2911,N_2892,N_2846);
or U2912 (N_2912,N_2863,N_2841);
nor U2913 (N_2913,N_2803,N_2830);
or U2914 (N_2914,N_2865,N_2874);
xor U2915 (N_2915,N_2824,N_2850);
and U2916 (N_2916,N_2836,N_2826);
nor U2917 (N_2917,N_2822,N_2896);
xor U2918 (N_2918,N_2873,N_2823);
and U2919 (N_2919,N_2897,N_2809);
nand U2920 (N_2920,N_2889,N_2808);
or U2921 (N_2921,N_2814,N_2844);
or U2922 (N_2922,N_2837,N_2828);
nand U2923 (N_2923,N_2866,N_2891);
nand U2924 (N_2924,N_2815,N_2849);
nand U2925 (N_2925,N_2835,N_2867);
or U2926 (N_2926,N_2878,N_2816);
nor U2927 (N_2927,N_2876,N_2869);
nand U2928 (N_2928,N_2883,N_2843);
and U2929 (N_2929,N_2832,N_2806);
nor U2930 (N_2930,N_2813,N_2831);
nand U2931 (N_2931,N_2802,N_2864);
or U2932 (N_2932,N_2851,N_2811);
or U2933 (N_2933,N_2893,N_2888);
xnor U2934 (N_2934,N_2820,N_2862);
nor U2935 (N_2935,N_2838,N_2895);
and U2936 (N_2936,N_2857,N_2845);
and U2937 (N_2937,N_2861,N_2817);
nand U2938 (N_2938,N_2852,N_2810);
nand U2939 (N_2939,N_2885,N_2884);
or U2940 (N_2940,N_2847,N_2825);
nor U2941 (N_2941,N_2899,N_2818);
or U2942 (N_2942,N_2880,N_2800);
nor U2943 (N_2943,N_2881,N_2807);
nand U2944 (N_2944,N_2819,N_2898);
nor U2945 (N_2945,N_2854,N_2842);
nor U2946 (N_2946,N_2890,N_2804);
or U2947 (N_2947,N_2887,N_2870);
and U2948 (N_2948,N_2871,N_2839);
or U2949 (N_2949,N_2833,N_2877);
nor U2950 (N_2950,N_2892,N_2811);
or U2951 (N_2951,N_2857,N_2882);
nand U2952 (N_2952,N_2827,N_2812);
and U2953 (N_2953,N_2892,N_2803);
nor U2954 (N_2954,N_2812,N_2850);
nor U2955 (N_2955,N_2829,N_2810);
and U2956 (N_2956,N_2893,N_2868);
xnor U2957 (N_2957,N_2809,N_2866);
nor U2958 (N_2958,N_2849,N_2846);
and U2959 (N_2959,N_2856,N_2804);
and U2960 (N_2960,N_2845,N_2812);
or U2961 (N_2961,N_2827,N_2854);
or U2962 (N_2962,N_2824,N_2842);
and U2963 (N_2963,N_2815,N_2857);
nand U2964 (N_2964,N_2830,N_2899);
and U2965 (N_2965,N_2896,N_2869);
and U2966 (N_2966,N_2887,N_2849);
and U2967 (N_2967,N_2892,N_2881);
nand U2968 (N_2968,N_2873,N_2826);
and U2969 (N_2969,N_2886,N_2858);
and U2970 (N_2970,N_2874,N_2860);
or U2971 (N_2971,N_2849,N_2862);
nor U2972 (N_2972,N_2837,N_2827);
nor U2973 (N_2973,N_2814,N_2891);
and U2974 (N_2974,N_2851,N_2889);
nand U2975 (N_2975,N_2840,N_2812);
nor U2976 (N_2976,N_2829,N_2824);
or U2977 (N_2977,N_2827,N_2808);
and U2978 (N_2978,N_2808,N_2892);
and U2979 (N_2979,N_2881,N_2827);
nand U2980 (N_2980,N_2834,N_2802);
nand U2981 (N_2981,N_2859,N_2838);
xor U2982 (N_2982,N_2862,N_2824);
and U2983 (N_2983,N_2888,N_2813);
and U2984 (N_2984,N_2860,N_2825);
nand U2985 (N_2985,N_2820,N_2832);
and U2986 (N_2986,N_2801,N_2854);
and U2987 (N_2987,N_2806,N_2887);
or U2988 (N_2988,N_2865,N_2863);
nand U2989 (N_2989,N_2899,N_2866);
and U2990 (N_2990,N_2859,N_2814);
and U2991 (N_2991,N_2873,N_2812);
and U2992 (N_2992,N_2870,N_2839);
and U2993 (N_2993,N_2873,N_2895);
nand U2994 (N_2994,N_2838,N_2819);
nand U2995 (N_2995,N_2807,N_2875);
nor U2996 (N_2996,N_2830,N_2868);
or U2997 (N_2997,N_2867,N_2813);
or U2998 (N_2998,N_2845,N_2827);
and U2999 (N_2999,N_2825,N_2889);
and U3000 (N_3000,N_2972,N_2975);
nand U3001 (N_3001,N_2996,N_2903);
and U3002 (N_3002,N_2931,N_2928);
or U3003 (N_3003,N_2902,N_2942);
xor U3004 (N_3004,N_2933,N_2943);
and U3005 (N_3005,N_2939,N_2971);
and U3006 (N_3006,N_2987,N_2995);
nand U3007 (N_3007,N_2945,N_2934);
nand U3008 (N_3008,N_2980,N_2908);
and U3009 (N_3009,N_2957,N_2953);
nor U3010 (N_3010,N_2966,N_2914);
xnor U3011 (N_3011,N_2923,N_2994);
nand U3012 (N_3012,N_2924,N_2958);
nand U3013 (N_3013,N_2973,N_2990);
nand U3014 (N_3014,N_2962,N_2913);
or U3015 (N_3015,N_2984,N_2985);
nand U3016 (N_3016,N_2950,N_2999);
and U3017 (N_3017,N_2956,N_2946);
nor U3018 (N_3018,N_2926,N_2978);
or U3019 (N_3019,N_2977,N_2963);
or U3020 (N_3020,N_2965,N_2920);
and U3021 (N_3021,N_2900,N_2982);
and U3022 (N_3022,N_2918,N_2915);
or U3023 (N_3023,N_2930,N_2979);
nand U3024 (N_3024,N_2925,N_2974);
nor U3025 (N_3025,N_2992,N_2906);
nand U3026 (N_3026,N_2969,N_2935);
or U3027 (N_3027,N_2949,N_2961);
nand U3028 (N_3028,N_2952,N_2964);
nand U3029 (N_3029,N_2940,N_2941);
nand U3030 (N_3030,N_2986,N_2932);
xnor U3031 (N_3031,N_2922,N_2968);
and U3032 (N_3032,N_2905,N_2948);
xnor U3033 (N_3033,N_2921,N_2976);
or U3034 (N_3034,N_2947,N_2988);
nand U3035 (N_3035,N_2997,N_2910);
or U3036 (N_3036,N_2938,N_2954);
nor U3037 (N_3037,N_2951,N_2907);
nand U3038 (N_3038,N_2901,N_2967);
and U3039 (N_3039,N_2937,N_2983);
or U3040 (N_3040,N_2989,N_2991);
nor U3041 (N_3041,N_2944,N_2904);
or U3042 (N_3042,N_2960,N_2909);
nand U3043 (N_3043,N_2927,N_2981);
nor U3044 (N_3044,N_2919,N_2916);
and U3045 (N_3045,N_2959,N_2912);
nand U3046 (N_3046,N_2911,N_2970);
xnor U3047 (N_3047,N_2917,N_2929);
and U3048 (N_3048,N_2998,N_2955);
and U3049 (N_3049,N_2936,N_2993);
nand U3050 (N_3050,N_2962,N_2925);
or U3051 (N_3051,N_2991,N_2914);
and U3052 (N_3052,N_2963,N_2950);
nor U3053 (N_3053,N_2917,N_2912);
or U3054 (N_3054,N_2956,N_2983);
nand U3055 (N_3055,N_2974,N_2982);
or U3056 (N_3056,N_2910,N_2959);
and U3057 (N_3057,N_2919,N_2966);
xnor U3058 (N_3058,N_2930,N_2952);
or U3059 (N_3059,N_2943,N_2902);
nand U3060 (N_3060,N_2973,N_2985);
nor U3061 (N_3061,N_2967,N_2903);
nand U3062 (N_3062,N_2905,N_2937);
nor U3063 (N_3063,N_2904,N_2902);
nor U3064 (N_3064,N_2957,N_2950);
xnor U3065 (N_3065,N_2931,N_2922);
nor U3066 (N_3066,N_2966,N_2954);
and U3067 (N_3067,N_2900,N_2964);
nand U3068 (N_3068,N_2966,N_2944);
nor U3069 (N_3069,N_2927,N_2951);
nor U3070 (N_3070,N_2933,N_2948);
or U3071 (N_3071,N_2928,N_2952);
xor U3072 (N_3072,N_2990,N_2993);
and U3073 (N_3073,N_2999,N_2980);
xor U3074 (N_3074,N_2907,N_2953);
or U3075 (N_3075,N_2943,N_2910);
and U3076 (N_3076,N_2957,N_2948);
or U3077 (N_3077,N_2962,N_2970);
nand U3078 (N_3078,N_2968,N_2943);
or U3079 (N_3079,N_2951,N_2937);
and U3080 (N_3080,N_2932,N_2969);
nor U3081 (N_3081,N_2916,N_2927);
nand U3082 (N_3082,N_2983,N_2944);
nor U3083 (N_3083,N_2903,N_2915);
nand U3084 (N_3084,N_2922,N_2928);
and U3085 (N_3085,N_2925,N_2985);
and U3086 (N_3086,N_2903,N_2930);
nand U3087 (N_3087,N_2912,N_2979);
or U3088 (N_3088,N_2943,N_2989);
xor U3089 (N_3089,N_2928,N_2941);
nor U3090 (N_3090,N_2901,N_2937);
xnor U3091 (N_3091,N_2946,N_2943);
and U3092 (N_3092,N_2927,N_2933);
nor U3093 (N_3093,N_2995,N_2955);
nor U3094 (N_3094,N_2946,N_2963);
and U3095 (N_3095,N_2954,N_2923);
and U3096 (N_3096,N_2903,N_2964);
nand U3097 (N_3097,N_2930,N_2920);
and U3098 (N_3098,N_2965,N_2955);
nand U3099 (N_3099,N_2950,N_2990);
or U3100 (N_3100,N_3097,N_3004);
xor U3101 (N_3101,N_3057,N_3040);
nand U3102 (N_3102,N_3081,N_3034);
and U3103 (N_3103,N_3010,N_3079);
nor U3104 (N_3104,N_3023,N_3095);
xnor U3105 (N_3105,N_3007,N_3009);
or U3106 (N_3106,N_3094,N_3016);
nor U3107 (N_3107,N_3027,N_3042);
and U3108 (N_3108,N_3087,N_3065);
or U3109 (N_3109,N_3026,N_3037);
and U3110 (N_3110,N_3088,N_3035);
or U3111 (N_3111,N_3025,N_3078);
and U3112 (N_3112,N_3062,N_3055);
nor U3113 (N_3113,N_3031,N_3092);
or U3114 (N_3114,N_3072,N_3093);
and U3115 (N_3115,N_3067,N_3038);
nand U3116 (N_3116,N_3083,N_3061);
or U3117 (N_3117,N_3086,N_3032);
or U3118 (N_3118,N_3099,N_3068);
and U3119 (N_3119,N_3054,N_3080);
and U3120 (N_3120,N_3096,N_3012);
nor U3121 (N_3121,N_3013,N_3029);
or U3122 (N_3122,N_3058,N_3020);
and U3123 (N_3123,N_3033,N_3085);
and U3124 (N_3124,N_3048,N_3008);
nor U3125 (N_3125,N_3077,N_3074);
or U3126 (N_3126,N_3030,N_3071);
or U3127 (N_3127,N_3051,N_3041);
and U3128 (N_3128,N_3091,N_3064);
or U3129 (N_3129,N_3098,N_3043);
nor U3130 (N_3130,N_3053,N_3017);
xnor U3131 (N_3131,N_3014,N_3002);
or U3132 (N_3132,N_3001,N_3006);
or U3133 (N_3133,N_3021,N_3005);
and U3134 (N_3134,N_3039,N_3070);
and U3135 (N_3135,N_3089,N_3018);
and U3136 (N_3136,N_3063,N_3028);
and U3137 (N_3137,N_3052,N_3044);
nor U3138 (N_3138,N_3075,N_3090);
nor U3139 (N_3139,N_3015,N_3047);
nor U3140 (N_3140,N_3036,N_3076);
and U3141 (N_3141,N_3046,N_3069);
or U3142 (N_3142,N_3084,N_3066);
and U3143 (N_3143,N_3000,N_3003);
nor U3144 (N_3144,N_3082,N_3073);
nand U3145 (N_3145,N_3024,N_3060);
and U3146 (N_3146,N_3011,N_3059);
and U3147 (N_3147,N_3056,N_3049);
and U3148 (N_3148,N_3019,N_3045);
or U3149 (N_3149,N_3050,N_3022);
nor U3150 (N_3150,N_3082,N_3089);
or U3151 (N_3151,N_3046,N_3022);
and U3152 (N_3152,N_3017,N_3024);
and U3153 (N_3153,N_3072,N_3054);
nor U3154 (N_3154,N_3061,N_3079);
nand U3155 (N_3155,N_3007,N_3010);
nor U3156 (N_3156,N_3095,N_3078);
and U3157 (N_3157,N_3076,N_3038);
nand U3158 (N_3158,N_3052,N_3037);
nor U3159 (N_3159,N_3031,N_3069);
nor U3160 (N_3160,N_3024,N_3082);
and U3161 (N_3161,N_3054,N_3070);
nor U3162 (N_3162,N_3075,N_3012);
nand U3163 (N_3163,N_3086,N_3047);
or U3164 (N_3164,N_3089,N_3054);
nand U3165 (N_3165,N_3022,N_3064);
or U3166 (N_3166,N_3089,N_3006);
nand U3167 (N_3167,N_3090,N_3050);
or U3168 (N_3168,N_3072,N_3045);
xnor U3169 (N_3169,N_3047,N_3026);
nor U3170 (N_3170,N_3085,N_3025);
nand U3171 (N_3171,N_3013,N_3062);
nand U3172 (N_3172,N_3033,N_3074);
nor U3173 (N_3173,N_3091,N_3081);
or U3174 (N_3174,N_3024,N_3077);
and U3175 (N_3175,N_3056,N_3064);
xor U3176 (N_3176,N_3083,N_3035);
nor U3177 (N_3177,N_3081,N_3014);
nor U3178 (N_3178,N_3005,N_3096);
nor U3179 (N_3179,N_3027,N_3069);
or U3180 (N_3180,N_3039,N_3092);
and U3181 (N_3181,N_3063,N_3061);
xor U3182 (N_3182,N_3040,N_3073);
and U3183 (N_3183,N_3006,N_3036);
or U3184 (N_3184,N_3014,N_3097);
nand U3185 (N_3185,N_3044,N_3084);
or U3186 (N_3186,N_3067,N_3008);
and U3187 (N_3187,N_3002,N_3032);
or U3188 (N_3188,N_3027,N_3060);
or U3189 (N_3189,N_3063,N_3070);
nand U3190 (N_3190,N_3002,N_3060);
and U3191 (N_3191,N_3012,N_3069);
or U3192 (N_3192,N_3003,N_3068);
nor U3193 (N_3193,N_3003,N_3080);
nand U3194 (N_3194,N_3094,N_3063);
and U3195 (N_3195,N_3055,N_3053);
or U3196 (N_3196,N_3070,N_3037);
and U3197 (N_3197,N_3067,N_3021);
and U3198 (N_3198,N_3084,N_3095);
and U3199 (N_3199,N_3088,N_3042);
nor U3200 (N_3200,N_3114,N_3186);
nand U3201 (N_3201,N_3134,N_3145);
or U3202 (N_3202,N_3171,N_3144);
and U3203 (N_3203,N_3160,N_3198);
xnor U3204 (N_3204,N_3156,N_3169);
or U3205 (N_3205,N_3112,N_3115);
nor U3206 (N_3206,N_3182,N_3157);
xnor U3207 (N_3207,N_3128,N_3141);
xor U3208 (N_3208,N_3123,N_3151);
or U3209 (N_3209,N_3172,N_3127);
nand U3210 (N_3210,N_3106,N_3150);
nand U3211 (N_3211,N_3100,N_3138);
nor U3212 (N_3212,N_3164,N_3113);
xor U3213 (N_3213,N_3193,N_3111);
or U3214 (N_3214,N_3168,N_3140);
or U3215 (N_3215,N_3129,N_3136);
nand U3216 (N_3216,N_3149,N_3126);
nand U3217 (N_3217,N_3105,N_3154);
nand U3218 (N_3218,N_3125,N_3142);
or U3219 (N_3219,N_3122,N_3101);
nand U3220 (N_3220,N_3147,N_3159);
nand U3221 (N_3221,N_3189,N_3180);
or U3222 (N_3222,N_3132,N_3137);
or U3223 (N_3223,N_3148,N_3192);
nor U3224 (N_3224,N_3158,N_3161);
nor U3225 (N_3225,N_3191,N_3185);
xor U3226 (N_3226,N_3110,N_3121);
or U3227 (N_3227,N_3116,N_3162);
nand U3228 (N_3228,N_3102,N_3118);
nor U3229 (N_3229,N_3181,N_3176);
nor U3230 (N_3230,N_3143,N_3124);
nor U3231 (N_3231,N_3199,N_3152);
or U3232 (N_3232,N_3139,N_3195);
nor U3233 (N_3233,N_3103,N_3174);
nor U3234 (N_3234,N_3196,N_3175);
nand U3235 (N_3235,N_3177,N_3163);
nor U3236 (N_3236,N_3190,N_3131);
and U3237 (N_3237,N_3109,N_3153);
nor U3238 (N_3238,N_3173,N_3117);
nand U3239 (N_3239,N_3167,N_3107);
or U3240 (N_3240,N_3188,N_3197);
xor U3241 (N_3241,N_3183,N_3146);
and U3242 (N_3242,N_3194,N_3165);
and U3243 (N_3243,N_3184,N_3130);
nand U3244 (N_3244,N_3135,N_3120);
nor U3245 (N_3245,N_3179,N_3155);
nand U3246 (N_3246,N_3178,N_3133);
nor U3247 (N_3247,N_3187,N_3104);
nand U3248 (N_3248,N_3108,N_3119);
nor U3249 (N_3249,N_3166,N_3170);
nor U3250 (N_3250,N_3124,N_3179);
and U3251 (N_3251,N_3161,N_3135);
nand U3252 (N_3252,N_3153,N_3192);
nor U3253 (N_3253,N_3199,N_3139);
nor U3254 (N_3254,N_3115,N_3152);
nor U3255 (N_3255,N_3167,N_3189);
xor U3256 (N_3256,N_3107,N_3188);
nor U3257 (N_3257,N_3154,N_3153);
and U3258 (N_3258,N_3168,N_3153);
nand U3259 (N_3259,N_3169,N_3176);
nand U3260 (N_3260,N_3136,N_3177);
or U3261 (N_3261,N_3171,N_3198);
and U3262 (N_3262,N_3165,N_3187);
and U3263 (N_3263,N_3178,N_3193);
nor U3264 (N_3264,N_3101,N_3134);
or U3265 (N_3265,N_3136,N_3117);
and U3266 (N_3266,N_3135,N_3160);
nand U3267 (N_3267,N_3178,N_3125);
and U3268 (N_3268,N_3125,N_3139);
or U3269 (N_3269,N_3175,N_3100);
nand U3270 (N_3270,N_3188,N_3196);
or U3271 (N_3271,N_3167,N_3113);
or U3272 (N_3272,N_3198,N_3181);
nor U3273 (N_3273,N_3182,N_3138);
nand U3274 (N_3274,N_3128,N_3110);
and U3275 (N_3275,N_3128,N_3170);
nand U3276 (N_3276,N_3139,N_3144);
nor U3277 (N_3277,N_3160,N_3168);
nor U3278 (N_3278,N_3153,N_3121);
nor U3279 (N_3279,N_3150,N_3103);
nor U3280 (N_3280,N_3141,N_3131);
or U3281 (N_3281,N_3178,N_3155);
nand U3282 (N_3282,N_3126,N_3116);
or U3283 (N_3283,N_3145,N_3161);
and U3284 (N_3284,N_3121,N_3157);
xor U3285 (N_3285,N_3120,N_3110);
and U3286 (N_3286,N_3116,N_3165);
and U3287 (N_3287,N_3123,N_3102);
or U3288 (N_3288,N_3127,N_3112);
nand U3289 (N_3289,N_3199,N_3140);
nor U3290 (N_3290,N_3114,N_3128);
nor U3291 (N_3291,N_3114,N_3124);
or U3292 (N_3292,N_3169,N_3108);
nor U3293 (N_3293,N_3122,N_3163);
or U3294 (N_3294,N_3133,N_3139);
or U3295 (N_3295,N_3181,N_3127);
nand U3296 (N_3296,N_3108,N_3192);
nand U3297 (N_3297,N_3169,N_3123);
xnor U3298 (N_3298,N_3189,N_3149);
or U3299 (N_3299,N_3183,N_3152);
or U3300 (N_3300,N_3238,N_3263);
xor U3301 (N_3301,N_3216,N_3251);
or U3302 (N_3302,N_3250,N_3243);
and U3303 (N_3303,N_3269,N_3212);
nand U3304 (N_3304,N_3276,N_3252);
nand U3305 (N_3305,N_3268,N_3266);
nor U3306 (N_3306,N_3297,N_3298);
nand U3307 (N_3307,N_3200,N_3292);
and U3308 (N_3308,N_3271,N_3291);
or U3309 (N_3309,N_3246,N_3229);
nand U3310 (N_3310,N_3247,N_3217);
nor U3311 (N_3311,N_3281,N_3272);
nor U3312 (N_3312,N_3213,N_3259);
nand U3313 (N_3313,N_3218,N_3262);
nand U3314 (N_3314,N_3285,N_3226);
xor U3315 (N_3315,N_3235,N_3234);
and U3316 (N_3316,N_3240,N_3278);
and U3317 (N_3317,N_3214,N_3237);
xnor U3318 (N_3318,N_3248,N_3279);
xnor U3319 (N_3319,N_3293,N_3230);
nand U3320 (N_3320,N_3258,N_3242);
nor U3321 (N_3321,N_3254,N_3224);
nand U3322 (N_3322,N_3255,N_3288);
nand U3323 (N_3323,N_3232,N_3205);
and U3324 (N_3324,N_3256,N_3239);
or U3325 (N_3325,N_3209,N_3245);
nand U3326 (N_3326,N_3260,N_3233);
and U3327 (N_3327,N_3215,N_3284);
nor U3328 (N_3328,N_3227,N_3253);
nand U3329 (N_3329,N_3208,N_3287);
nand U3330 (N_3330,N_3204,N_3295);
nor U3331 (N_3331,N_3280,N_3202);
nor U3332 (N_3332,N_3277,N_3231);
and U3333 (N_3333,N_3236,N_3228);
nor U3334 (N_3334,N_3283,N_3296);
or U3335 (N_3335,N_3201,N_3274);
xor U3336 (N_3336,N_3211,N_3207);
nand U3337 (N_3337,N_3261,N_3210);
xnor U3338 (N_3338,N_3203,N_3264);
nor U3339 (N_3339,N_3282,N_3225);
nand U3340 (N_3340,N_3294,N_3249);
xnor U3341 (N_3341,N_3241,N_3275);
nand U3342 (N_3342,N_3244,N_3289);
nor U3343 (N_3343,N_3286,N_3273);
and U3344 (N_3344,N_3206,N_3219);
nor U3345 (N_3345,N_3290,N_3220);
or U3346 (N_3346,N_3299,N_3223);
nand U3347 (N_3347,N_3222,N_3221);
or U3348 (N_3348,N_3267,N_3265);
and U3349 (N_3349,N_3257,N_3270);
and U3350 (N_3350,N_3284,N_3233);
nor U3351 (N_3351,N_3294,N_3200);
xnor U3352 (N_3352,N_3248,N_3287);
and U3353 (N_3353,N_3225,N_3265);
nand U3354 (N_3354,N_3299,N_3284);
nor U3355 (N_3355,N_3281,N_3214);
xnor U3356 (N_3356,N_3267,N_3283);
nor U3357 (N_3357,N_3269,N_3271);
xor U3358 (N_3358,N_3236,N_3284);
and U3359 (N_3359,N_3282,N_3283);
nor U3360 (N_3360,N_3243,N_3245);
nand U3361 (N_3361,N_3203,N_3266);
or U3362 (N_3362,N_3266,N_3279);
nor U3363 (N_3363,N_3273,N_3266);
or U3364 (N_3364,N_3218,N_3233);
nand U3365 (N_3365,N_3264,N_3224);
nand U3366 (N_3366,N_3278,N_3207);
and U3367 (N_3367,N_3269,N_3211);
and U3368 (N_3368,N_3272,N_3226);
or U3369 (N_3369,N_3204,N_3211);
xnor U3370 (N_3370,N_3291,N_3287);
or U3371 (N_3371,N_3256,N_3241);
nor U3372 (N_3372,N_3281,N_3292);
nor U3373 (N_3373,N_3293,N_3212);
and U3374 (N_3374,N_3241,N_3208);
nand U3375 (N_3375,N_3203,N_3238);
or U3376 (N_3376,N_3287,N_3295);
and U3377 (N_3377,N_3237,N_3265);
xor U3378 (N_3378,N_3225,N_3288);
or U3379 (N_3379,N_3254,N_3260);
and U3380 (N_3380,N_3280,N_3263);
and U3381 (N_3381,N_3280,N_3279);
and U3382 (N_3382,N_3200,N_3215);
or U3383 (N_3383,N_3274,N_3208);
nor U3384 (N_3384,N_3280,N_3293);
nor U3385 (N_3385,N_3257,N_3288);
and U3386 (N_3386,N_3298,N_3230);
nor U3387 (N_3387,N_3234,N_3214);
or U3388 (N_3388,N_3220,N_3256);
nand U3389 (N_3389,N_3249,N_3202);
nand U3390 (N_3390,N_3274,N_3299);
or U3391 (N_3391,N_3217,N_3269);
and U3392 (N_3392,N_3263,N_3274);
or U3393 (N_3393,N_3265,N_3234);
and U3394 (N_3394,N_3213,N_3230);
or U3395 (N_3395,N_3239,N_3252);
nand U3396 (N_3396,N_3298,N_3272);
nand U3397 (N_3397,N_3233,N_3225);
nand U3398 (N_3398,N_3247,N_3200);
nand U3399 (N_3399,N_3254,N_3250);
nor U3400 (N_3400,N_3334,N_3305);
and U3401 (N_3401,N_3382,N_3322);
xor U3402 (N_3402,N_3323,N_3335);
nor U3403 (N_3403,N_3393,N_3337);
nor U3404 (N_3404,N_3354,N_3391);
or U3405 (N_3405,N_3341,N_3326);
nand U3406 (N_3406,N_3388,N_3313);
or U3407 (N_3407,N_3333,N_3359);
and U3408 (N_3408,N_3349,N_3357);
xor U3409 (N_3409,N_3376,N_3332);
and U3410 (N_3410,N_3336,N_3330);
xor U3411 (N_3411,N_3386,N_3364);
nor U3412 (N_3412,N_3345,N_3340);
nand U3413 (N_3413,N_3346,N_3302);
and U3414 (N_3414,N_3320,N_3312);
nand U3415 (N_3415,N_3347,N_3316);
and U3416 (N_3416,N_3343,N_3324);
nand U3417 (N_3417,N_3383,N_3315);
or U3418 (N_3418,N_3377,N_3314);
or U3419 (N_3419,N_3344,N_3342);
nor U3420 (N_3420,N_3389,N_3353);
or U3421 (N_3421,N_3367,N_3307);
nor U3422 (N_3422,N_3321,N_3375);
and U3423 (N_3423,N_3309,N_3300);
or U3424 (N_3424,N_3331,N_3390);
and U3425 (N_3425,N_3394,N_3370);
and U3426 (N_3426,N_3311,N_3361);
nor U3427 (N_3427,N_3366,N_3396);
nor U3428 (N_3428,N_3356,N_3387);
nor U3429 (N_3429,N_3350,N_3372);
nand U3430 (N_3430,N_3327,N_3365);
and U3431 (N_3431,N_3368,N_3318);
or U3432 (N_3432,N_3355,N_3329);
or U3433 (N_3433,N_3358,N_3303);
and U3434 (N_3434,N_3317,N_3371);
nor U3435 (N_3435,N_3384,N_3362);
nand U3436 (N_3436,N_3399,N_3325);
nand U3437 (N_3437,N_3306,N_3374);
xor U3438 (N_3438,N_3319,N_3308);
nand U3439 (N_3439,N_3395,N_3397);
xor U3440 (N_3440,N_3352,N_3360);
nor U3441 (N_3441,N_3301,N_3398);
or U3442 (N_3442,N_3385,N_3348);
xnor U3443 (N_3443,N_3381,N_3380);
and U3444 (N_3444,N_3363,N_3392);
nor U3445 (N_3445,N_3339,N_3378);
and U3446 (N_3446,N_3328,N_3338);
and U3447 (N_3447,N_3304,N_3379);
nand U3448 (N_3448,N_3369,N_3373);
nand U3449 (N_3449,N_3310,N_3351);
xor U3450 (N_3450,N_3344,N_3363);
and U3451 (N_3451,N_3352,N_3351);
or U3452 (N_3452,N_3335,N_3360);
nand U3453 (N_3453,N_3370,N_3374);
and U3454 (N_3454,N_3327,N_3394);
or U3455 (N_3455,N_3331,N_3343);
and U3456 (N_3456,N_3384,N_3300);
nor U3457 (N_3457,N_3317,N_3382);
nand U3458 (N_3458,N_3366,N_3331);
nand U3459 (N_3459,N_3383,N_3352);
xor U3460 (N_3460,N_3311,N_3386);
nor U3461 (N_3461,N_3304,N_3327);
nand U3462 (N_3462,N_3328,N_3333);
and U3463 (N_3463,N_3357,N_3384);
nor U3464 (N_3464,N_3385,N_3333);
or U3465 (N_3465,N_3386,N_3376);
nand U3466 (N_3466,N_3365,N_3346);
nand U3467 (N_3467,N_3330,N_3380);
nor U3468 (N_3468,N_3359,N_3302);
and U3469 (N_3469,N_3306,N_3389);
and U3470 (N_3470,N_3399,N_3362);
or U3471 (N_3471,N_3327,N_3358);
or U3472 (N_3472,N_3305,N_3386);
nand U3473 (N_3473,N_3361,N_3396);
nand U3474 (N_3474,N_3383,N_3376);
or U3475 (N_3475,N_3358,N_3325);
and U3476 (N_3476,N_3385,N_3389);
and U3477 (N_3477,N_3339,N_3307);
nand U3478 (N_3478,N_3378,N_3393);
nor U3479 (N_3479,N_3314,N_3356);
nand U3480 (N_3480,N_3398,N_3312);
and U3481 (N_3481,N_3368,N_3361);
or U3482 (N_3482,N_3323,N_3391);
nor U3483 (N_3483,N_3336,N_3381);
nand U3484 (N_3484,N_3340,N_3301);
nor U3485 (N_3485,N_3332,N_3314);
nand U3486 (N_3486,N_3380,N_3366);
or U3487 (N_3487,N_3371,N_3370);
and U3488 (N_3488,N_3376,N_3389);
and U3489 (N_3489,N_3347,N_3381);
nand U3490 (N_3490,N_3315,N_3343);
or U3491 (N_3491,N_3322,N_3336);
nand U3492 (N_3492,N_3332,N_3309);
nor U3493 (N_3493,N_3349,N_3390);
nor U3494 (N_3494,N_3392,N_3376);
or U3495 (N_3495,N_3364,N_3369);
or U3496 (N_3496,N_3357,N_3338);
or U3497 (N_3497,N_3339,N_3324);
or U3498 (N_3498,N_3350,N_3339);
nor U3499 (N_3499,N_3368,N_3308);
nor U3500 (N_3500,N_3445,N_3458);
nand U3501 (N_3501,N_3452,N_3470);
nand U3502 (N_3502,N_3495,N_3417);
and U3503 (N_3503,N_3483,N_3469);
nor U3504 (N_3504,N_3498,N_3466);
nand U3505 (N_3505,N_3436,N_3457);
nor U3506 (N_3506,N_3403,N_3428);
nand U3507 (N_3507,N_3492,N_3488);
and U3508 (N_3508,N_3494,N_3491);
xnor U3509 (N_3509,N_3499,N_3450);
nand U3510 (N_3510,N_3468,N_3474);
or U3511 (N_3511,N_3459,N_3462);
nand U3512 (N_3512,N_3496,N_3454);
nor U3513 (N_3513,N_3490,N_3430);
and U3514 (N_3514,N_3406,N_3441);
or U3515 (N_3515,N_3472,N_3429);
nor U3516 (N_3516,N_3414,N_3421);
nor U3517 (N_3517,N_3410,N_3487);
and U3518 (N_3518,N_3415,N_3440);
nor U3519 (N_3519,N_3477,N_3427);
nor U3520 (N_3520,N_3416,N_3432);
and U3521 (N_3521,N_3456,N_3408);
and U3522 (N_3522,N_3476,N_3442);
nor U3523 (N_3523,N_3418,N_3401);
or U3524 (N_3524,N_3419,N_3460);
nor U3525 (N_3525,N_3438,N_3426);
or U3526 (N_3526,N_3431,N_3409);
and U3527 (N_3527,N_3402,N_3451);
or U3528 (N_3528,N_3475,N_3425);
and U3529 (N_3529,N_3461,N_3449);
nor U3530 (N_3530,N_3420,N_3412);
nor U3531 (N_3531,N_3448,N_3400);
nand U3532 (N_3532,N_3422,N_3482);
xnor U3533 (N_3533,N_3486,N_3405);
or U3534 (N_3534,N_3437,N_3424);
and U3535 (N_3535,N_3489,N_3444);
or U3536 (N_3536,N_3446,N_3485);
nand U3537 (N_3537,N_3435,N_3404);
and U3538 (N_3538,N_3465,N_3413);
nor U3539 (N_3539,N_3481,N_3480);
nand U3540 (N_3540,N_3447,N_3471);
xor U3541 (N_3541,N_3463,N_3493);
or U3542 (N_3542,N_3478,N_3434);
and U3543 (N_3543,N_3433,N_3411);
xnor U3544 (N_3544,N_3473,N_3407);
nand U3545 (N_3545,N_3455,N_3467);
and U3546 (N_3546,N_3497,N_3464);
xnor U3547 (N_3547,N_3479,N_3439);
xor U3548 (N_3548,N_3423,N_3453);
or U3549 (N_3549,N_3443,N_3484);
or U3550 (N_3550,N_3428,N_3437);
nor U3551 (N_3551,N_3437,N_3498);
nor U3552 (N_3552,N_3460,N_3492);
or U3553 (N_3553,N_3458,N_3478);
nor U3554 (N_3554,N_3421,N_3474);
nor U3555 (N_3555,N_3440,N_3499);
xor U3556 (N_3556,N_3417,N_3461);
nand U3557 (N_3557,N_3460,N_3407);
nor U3558 (N_3558,N_3481,N_3423);
or U3559 (N_3559,N_3481,N_3464);
nor U3560 (N_3560,N_3434,N_3447);
or U3561 (N_3561,N_3488,N_3431);
or U3562 (N_3562,N_3402,N_3430);
nor U3563 (N_3563,N_3441,N_3494);
xor U3564 (N_3564,N_3464,N_3460);
and U3565 (N_3565,N_3430,N_3455);
or U3566 (N_3566,N_3428,N_3449);
nand U3567 (N_3567,N_3472,N_3490);
or U3568 (N_3568,N_3430,N_3479);
or U3569 (N_3569,N_3431,N_3469);
nand U3570 (N_3570,N_3436,N_3469);
or U3571 (N_3571,N_3417,N_3407);
and U3572 (N_3572,N_3412,N_3473);
nand U3573 (N_3573,N_3439,N_3495);
nand U3574 (N_3574,N_3482,N_3465);
xnor U3575 (N_3575,N_3447,N_3478);
nand U3576 (N_3576,N_3407,N_3459);
and U3577 (N_3577,N_3486,N_3412);
and U3578 (N_3578,N_3445,N_3470);
xnor U3579 (N_3579,N_3487,N_3479);
nor U3580 (N_3580,N_3401,N_3424);
and U3581 (N_3581,N_3478,N_3401);
nor U3582 (N_3582,N_3462,N_3486);
nand U3583 (N_3583,N_3486,N_3483);
nand U3584 (N_3584,N_3485,N_3473);
and U3585 (N_3585,N_3464,N_3434);
or U3586 (N_3586,N_3424,N_3464);
xor U3587 (N_3587,N_3476,N_3420);
nand U3588 (N_3588,N_3427,N_3450);
and U3589 (N_3589,N_3477,N_3483);
nand U3590 (N_3590,N_3465,N_3429);
and U3591 (N_3591,N_3416,N_3434);
or U3592 (N_3592,N_3483,N_3424);
or U3593 (N_3593,N_3426,N_3491);
xnor U3594 (N_3594,N_3416,N_3453);
or U3595 (N_3595,N_3453,N_3419);
or U3596 (N_3596,N_3496,N_3476);
nand U3597 (N_3597,N_3415,N_3483);
and U3598 (N_3598,N_3470,N_3409);
xor U3599 (N_3599,N_3417,N_3475);
xnor U3600 (N_3600,N_3589,N_3502);
and U3601 (N_3601,N_3556,N_3508);
or U3602 (N_3602,N_3585,N_3594);
or U3603 (N_3603,N_3595,N_3535);
or U3604 (N_3604,N_3530,N_3504);
and U3605 (N_3605,N_3536,N_3563);
xor U3606 (N_3606,N_3529,N_3518);
nand U3607 (N_3607,N_3571,N_3579);
nor U3608 (N_3608,N_3546,N_3576);
and U3609 (N_3609,N_3531,N_3543);
nor U3610 (N_3610,N_3548,N_3510);
xnor U3611 (N_3611,N_3588,N_3586);
and U3612 (N_3612,N_3509,N_3575);
nor U3613 (N_3613,N_3517,N_3568);
or U3614 (N_3614,N_3538,N_3567);
or U3615 (N_3615,N_3514,N_3569);
and U3616 (N_3616,N_3525,N_3507);
nand U3617 (N_3617,N_3553,N_3512);
xnor U3618 (N_3618,N_3524,N_3534);
nor U3619 (N_3619,N_3513,N_3582);
or U3620 (N_3620,N_3501,N_3540);
or U3621 (N_3621,N_3599,N_3597);
or U3622 (N_3622,N_3584,N_3506);
nand U3623 (N_3623,N_3572,N_3528);
nor U3624 (N_3624,N_3592,N_3596);
nand U3625 (N_3625,N_3578,N_3573);
nor U3626 (N_3626,N_3558,N_3551);
nor U3627 (N_3627,N_3574,N_3537);
nor U3628 (N_3628,N_3523,N_3552);
nand U3629 (N_3629,N_3541,N_3516);
or U3630 (N_3630,N_3593,N_3519);
and U3631 (N_3631,N_3522,N_3561);
nand U3632 (N_3632,N_3565,N_3555);
and U3633 (N_3633,N_3559,N_3526);
nand U3634 (N_3634,N_3577,N_3580);
and U3635 (N_3635,N_3542,N_3562);
or U3636 (N_3636,N_3527,N_3505);
nor U3637 (N_3637,N_3511,N_3557);
and U3638 (N_3638,N_3539,N_3547);
nor U3639 (N_3639,N_3503,N_3500);
nand U3640 (N_3640,N_3554,N_3566);
or U3641 (N_3641,N_3544,N_3520);
nor U3642 (N_3642,N_3591,N_3550);
xnor U3643 (N_3643,N_3533,N_3521);
and U3644 (N_3644,N_3564,N_3598);
xor U3645 (N_3645,N_3532,N_3545);
xor U3646 (N_3646,N_3583,N_3570);
or U3647 (N_3647,N_3581,N_3549);
xnor U3648 (N_3648,N_3515,N_3587);
nand U3649 (N_3649,N_3590,N_3560);
nand U3650 (N_3650,N_3565,N_3558);
nor U3651 (N_3651,N_3572,N_3542);
xor U3652 (N_3652,N_3542,N_3589);
nor U3653 (N_3653,N_3535,N_3533);
xnor U3654 (N_3654,N_3591,N_3513);
and U3655 (N_3655,N_3564,N_3503);
and U3656 (N_3656,N_3508,N_3566);
and U3657 (N_3657,N_3561,N_3510);
or U3658 (N_3658,N_3583,N_3532);
and U3659 (N_3659,N_3570,N_3519);
nand U3660 (N_3660,N_3516,N_3584);
or U3661 (N_3661,N_3597,N_3522);
or U3662 (N_3662,N_3519,N_3514);
and U3663 (N_3663,N_3526,N_3546);
xor U3664 (N_3664,N_3500,N_3582);
nor U3665 (N_3665,N_3518,N_3566);
or U3666 (N_3666,N_3534,N_3577);
nor U3667 (N_3667,N_3570,N_3520);
nor U3668 (N_3668,N_3562,N_3533);
nor U3669 (N_3669,N_3587,N_3539);
nand U3670 (N_3670,N_3543,N_3552);
nor U3671 (N_3671,N_3532,N_3550);
nand U3672 (N_3672,N_3561,N_3589);
or U3673 (N_3673,N_3590,N_3547);
nor U3674 (N_3674,N_3562,N_3503);
nor U3675 (N_3675,N_3580,N_3541);
nor U3676 (N_3676,N_3578,N_3542);
xnor U3677 (N_3677,N_3542,N_3584);
and U3678 (N_3678,N_3517,N_3596);
and U3679 (N_3679,N_3546,N_3550);
or U3680 (N_3680,N_3502,N_3517);
nor U3681 (N_3681,N_3541,N_3513);
nand U3682 (N_3682,N_3593,N_3598);
or U3683 (N_3683,N_3563,N_3511);
nor U3684 (N_3684,N_3593,N_3538);
or U3685 (N_3685,N_3525,N_3591);
or U3686 (N_3686,N_3587,N_3576);
nand U3687 (N_3687,N_3569,N_3583);
or U3688 (N_3688,N_3591,N_3586);
or U3689 (N_3689,N_3575,N_3564);
nor U3690 (N_3690,N_3594,N_3543);
and U3691 (N_3691,N_3582,N_3565);
and U3692 (N_3692,N_3524,N_3593);
nand U3693 (N_3693,N_3506,N_3541);
nand U3694 (N_3694,N_3575,N_3572);
nor U3695 (N_3695,N_3577,N_3582);
or U3696 (N_3696,N_3518,N_3515);
nor U3697 (N_3697,N_3550,N_3505);
or U3698 (N_3698,N_3593,N_3553);
nand U3699 (N_3699,N_3539,N_3515);
or U3700 (N_3700,N_3635,N_3685);
nand U3701 (N_3701,N_3619,N_3636);
nand U3702 (N_3702,N_3649,N_3609);
and U3703 (N_3703,N_3675,N_3628);
nand U3704 (N_3704,N_3600,N_3645);
and U3705 (N_3705,N_3604,N_3625);
xnor U3706 (N_3706,N_3655,N_3690);
nand U3707 (N_3707,N_3669,N_3681);
nor U3708 (N_3708,N_3616,N_3667);
nand U3709 (N_3709,N_3664,N_3634);
or U3710 (N_3710,N_3605,N_3684);
nor U3711 (N_3711,N_3683,N_3601);
or U3712 (N_3712,N_3657,N_3697);
or U3713 (N_3713,N_3631,N_3644);
xnor U3714 (N_3714,N_3696,N_3629);
and U3715 (N_3715,N_3647,N_3654);
and U3716 (N_3716,N_3671,N_3615);
xor U3717 (N_3717,N_3620,N_3672);
and U3718 (N_3718,N_3668,N_3682);
or U3719 (N_3719,N_3648,N_3680);
nor U3720 (N_3720,N_3624,N_3689);
and U3721 (N_3721,N_3676,N_3618);
nor U3722 (N_3722,N_3606,N_3695);
nand U3723 (N_3723,N_3674,N_3699);
and U3724 (N_3724,N_3607,N_3639);
xnor U3725 (N_3725,N_3623,N_3622);
nand U3726 (N_3726,N_3692,N_3640);
nand U3727 (N_3727,N_3613,N_3656);
nor U3728 (N_3728,N_3603,N_3650);
nor U3729 (N_3729,N_3663,N_3611);
or U3730 (N_3730,N_3679,N_3677);
xnor U3731 (N_3731,N_3670,N_3627);
nor U3732 (N_3732,N_3617,N_3614);
or U3733 (N_3733,N_3691,N_3608);
xor U3734 (N_3734,N_3687,N_3632);
and U3735 (N_3735,N_3694,N_3651);
nand U3736 (N_3736,N_3638,N_3661);
or U3737 (N_3737,N_3686,N_3658);
and U3738 (N_3738,N_3637,N_3646);
and U3739 (N_3739,N_3641,N_3693);
and U3740 (N_3740,N_3652,N_3642);
nor U3741 (N_3741,N_3666,N_3626);
nand U3742 (N_3742,N_3659,N_3665);
nor U3743 (N_3743,N_3643,N_3602);
nor U3744 (N_3744,N_3612,N_3698);
nor U3745 (N_3745,N_3678,N_3633);
and U3746 (N_3746,N_3621,N_3610);
or U3747 (N_3747,N_3688,N_3630);
nand U3748 (N_3748,N_3673,N_3660);
nor U3749 (N_3749,N_3662,N_3653);
nand U3750 (N_3750,N_3638,N_3695);
nor U3751 (N_3751,N_3649,N_3619);
or U3752 (N_3752,N_3639,N_3614);
nor U3753 (N_3753,N_3636,N_3657);
or U3754 (N_3754,N_3612,N_3695);
nor U3755 (N_3755,N_3656,N_3626);
nor U3756 (N_3756,N_3676,N_3608);
nor U3757 (N_3757,N_3688,N_3619);
and U3758 (N_3758,N_3673,N_3629);
and U3759 (N_3759,N_3658,N_3661);
or U3760 (N_3760,N_3696,N_3681);
and U3761 (N_3761,N_3606,N_3658);
or U3762 (N_3762,N_3607,N_3658);
or U3763 (N_3763,N_3641,N_3671);
nand U3764 (N_3764,N_3676,N_3684);
nand U3765 (N_3765,N_3680,N_3687);
or U3766 (N_3766,N_3627,N_3616);
or U3767 (N_3767,N_3671,N_3657);
nor U3768 (N_3768,N_3669,N_3617);
or U3769 (N_3769,N_3668,N_3638);
and U3770 (N_3770,N_3611,N_3636);
nor U3771 (N_3771,N_3651,N_3621);
and U3772 (N_3772,N_3636,N_3656);
xnor U3773 (N_3773,N_3667,N_3606);
nor U3774 (N_3774,N_3602,N_3658);
nand U3775 (N_3775,N_3633,N_3695);
or U3776 (N_3776,N_3634,N_3636);
nor U3777 (N_3777,N_3683,N_3612);
nor U3778 (N_3778,N_3661,N_3616);
and U3779 (N_3779,N_3653,N_3601);
nand U3780 (N_3780,N_3648,N_3693);
and U3781 (N_3781,N_3656,N_3676);
nand U3782 (N_3782,N_3684,N_3649);
and U3783 (N_3783,N_3633,N_3623);
and U3784 (N_3784,N_3637,N_3689);
nand U3785 (N_3785,N_3659,N_3663);
and U3786 (N_3786,N_3616,N_3695);
or U3787 (N_3787,N_3624,N_3661);
xnor U3788 (N_3788,N_3638,N_3674);
xor U3789 (N_3789,N_3664,N_3658);
nor U3790 (N_3790,N_3638,N_3611);
or U3791 (N_3791,N_3682,N_3637);
or U3792 (N_3792,N_3666,N_3605);
xnor U3793 (N_3793,N_3626,N_3611);
nor U3794 (N_3794,N_3696,N_3619);
nand U3795 (N_3795,N_3641,N_3686);
xnor U3796 (N_3796,N_3632,N_3652);
nand U3797 (N_3797,N_3679,N_3624);
and U3798 (N_3798,N_3639,N_3646);
and U3799 (N_3799,N_3602,N_3661);
or U3800 (N_3800,N_3717,N_3730);
nor U3801 (N_3801,N_3705,N_3761);
nor U3802 (N_3802,N_3722,N_3767);
nor U3803 (N_3803,N_3798,N_3729);
or U3804 (N_3804,N_3736,N_3728);
and U3805 (N_3805,N_3768,N_3707);
xor U3806 (N_3806,N_3737,N_3796);
and U3807 (N_3807,N_3791,N_3762);
or U3808 (N_3808,N_3799,N_3734);
xnor U3809 (N_3809,N_3740,N_3756);
nand U3810 (N_3810,N_3714,N_3718);
or U3811 (N_3811,N_3792,N_3778);
xnor U3812 (N_3812,N_3702,N_3758);
nand U3813 (N_3813,N_3742,N_3727);
nand U3814 (N_3814,N_3738,N_3724);
nor U3815 (N_3815,N_3704,N_3754);
nor U3816 (N_3816,N_3732,N_3711);
or U3817 (N_3817,N_3710,N_3771);
xor U3818 (N_3818,N_3735,N_3706);
xor U3819 (N_3819,N_3721,N_3769);
nor U3820 (N_3820,N_3760,N_3783);
nor U3821 (N_3821,N_3700,N_3753);
nor U3822 (N_3822,N_3716,N_3752);
and U3823 (N_3823,N_3773,N_3770);
and U3824 (N_3824,N_3741,N_3794);
or U3825 (N_3825,N_3723,N_3720);
and U3826 (N_3826,N_3788,N_3797);
or U3827 (N_3827,N_3763,N_3712);
nor U3828 (N_3828,N_3787,N_3708);
xor U3829 (N_3829,N_3782,N_3726);
or U3830 (N_3830,N_3759,N_3765);
nor U3831 (N_3831,N_3785,N_3795);
and U3832 (N_3832,N_3779,N_3755);
nand U3833 (N_3833,N_3749,N_3703);
nand U3834 (N_3834,N_3790,N_3789);
or U3835 (N_3835,N_3772,N_3709);
and U3836 (N_3836,N_3748,N_3780);
nor U3837 (N_3837,N_3775,N_3786);
nor U3838 (N_3838,N_3777,N_3715);
nor U3839 (N_3839,N_3781,N_3743);
nand U3840 (N_3840,N_3751,N_3744);
and U3841 (N_3841,N_3739,N_3766);
or U3842 (N_3842,N_3719,N_3733);
nand U3843 (N_3843,N_3764,N_3776);
nand U3844 (N_3844,N_3713,N_3731);
nand U3845 (N_3845,N_3757,N_3774);
nand U3846 (N_3846,N_3750,N_3793);
or U3847 (N_3847,N_3701,N_3725);
nand U3848 (N_3848,N_3746,N_3784);
and U3849 (N_3849,N_3747,N_3745);
nand U3850 (N_3850,N_3704,N_3710);
and U3851 (N_3851,N_3724,N_3791);
nand U3852 (N_3852,N_3738,N_3739);
or U3853 (N_3853,N_3708,N_3707);
and U3854 (N_3854,N_3752,N_3789);
or U3855 (N_3855,N_3761,N_3765);
or U3856 (N_3856,N_3761,N_3786);
or U3857 (N_3857,N_3762,N_3703);
and U3858 (N_3858,N_3777,N_3738);
and U3859 (N_3859,N_3732,N_3772);
nor U3860 (N_3860,N_3731,N_3777);
nand U3861 (N_3861,N_3746,N_3721);
nand U3862 (N_3862,N_3723,N_3787);
nor U3863 (N_3863,N_3734,N_3764);
or U3864 (N_3864,N_3786,N_3708);
or U3865 (N_3865,N_3756,N_3789);
nor U3866 (N_3866,N_3704,N_3712);
xnor U3867 (N_3867,N_3742,N_3745);
nor U3868 (N_3868,N_3795,N_3758);
nand U3869 (N_3869,N_3776,N_3729);
nand U3870 (N_3870,N_3767,N_3769);
and U3871 (N_3871,N_3769,N_3714);
nand U3872 (N_3872,N_3786,N_3772);
xor U3873 (N_3873,N_3791,N_3795);
and U3874 (N_3874,N_3747,N_3755);
or U3875 (N_3875,N_3745,N_3755);
and U3876 (N_3876,N_3787,N_3724);
or U3877 (N_3877,N_3719,N_3765);
nor U3878 (N_3878,N_3756,N_3716);
or U3879 (N_3879,N_3714,N_3705);
nand U3880 (N_3880,N_3768,N_3710);
xor U3881 (N_3881,N_3796,N_3722);
xor U3882 (N_3882,N_3736,N_3722);
or U3883 (N_3883,N_3790,N_3700);
nor U3884 (N_3884,N_3779,N_3791);
or U3885 (N_3885,N_3704,N_3715);
nand U3886 (N_3886,N_3713,N_3775);
nor U3887 (N_3887,N_3769,N_3793);
and U3888 (N_3888,N_3717,N_3748);
or U3889 (N_3889,N_3700,N_3730);
nand U3890 (N_3890,N_3778,N_3752);
xnor U3891 (N_3891,N_3780,N_3726);
nor U3892 (N_3892,N_3728,N_3727);
nor U3893 (N_3893,N_3744,N_3733);
nand U3894 (N_3894,N_3770,N_3720);
or U3895 (N_3895,N_3725,N_3753);
or U3896 (N_3896,N_3749,N_3706);
nand U3897 (N_3897,N_3727,N_3730);
and U3898 (N_3898,N_3720,N_3782);
or U3899 (N_3899,N_3708,N_3701);
nor U3900 (N_3900,N_3852,N_3880);
nor U3901 (N_3901,N_3859,N_3897);
or U3902 (N_3902,N_3837,N_3824);
xnor U3903 (N_3903,N_3866,N_3844);
nor U3904 (N_3904,N_3876,N_3847);
xor U3905 (N_3905,N_3865,N_3812);
nor U3906 (N_3906,N_3839,N_3860);
nor U3907 (N_3907,N_3826,N_3815);
xnor U3908 (N_3908,N_3863,N_3885);
nand U3909 (N_3909,N_3810,N_3807);
and U3910 (N_3910,N_3804,N_3870);
nor U3911 (N_3911,N_3864,N_3823);
nor U3912 (N_3912,N_3838,N_3855);
nor U3913 (N_3913,N_3825,N_3883);
or U3914 (N_3914,N_3875,N_3829);
or U3915 (N_3915,N_3878,N_3830);
nand U3916 (N_3916,N_3813,N_3888);
nor U3917 (N_3917,N_3884,N_3898);
nand U3918 (N_3918,N_3803,N_3842);
or U3919 (N_3919,N_3854,N_3801);
and U3920 (N_3920,N_3821,N_3892);
xnor U3921 (N_3921,N_3820,N_3879);
nand U3922 (N_3922,N_3840,N_3836);
xor U3923 (N_3923,N_3881,N_3887);
or U3924 (N_3924,N_3845,N_3886);
nor U3925 (N_3925,N_3873,N_3872);
xnor U3926 (N_3926,N_3871,N_3861);
and U3927 (N_3927,N_3802,N_3805);
and U3928 (N_3928,N_3808,N_3819);
nand U3929 (N_3929,N_3869,N_3858);
nand U3930 (N_3930,N_3833,N_3814);
xor U3931 (N_3931,N_3868,N_3895);
or U3932 (N_3932,N_3827,N_3857);
xnor U3933 (N_3933,N_3843,N_3882);
or U3934 (N_3934,N_3806,N_3818);
or U3935 (N_3935,N_3856,N_3832);
or U3936 (N_3936,N_3817,N_3874);
nand U3937 (N_3937,N_3890,N_3867);
or U3938 (N_3938,N_3851,N_3862);
and U3939 (N_3939,N_3877,N_3846);
or U3940 (N_3940,N_3894,N_3809);
nand U3941 (N_3941,N_3899,N_3831);
nand U3942 (N_3942,N_3816,N_3889);
or U3943 (N_3943,N_3835,N_3828);
or U3944 (N_3944,N_3893,N_3896);
and U3945 (N_3945,N_3848,N_3811);
nor U3946 (N_3946,N_3853,N_3849);
xnor U3947 (N_3947,N_3822,N_3834);
xor U3948 (N_3948,N_3800,N_3891);
and U3949 (N_3949,N_3841,N_3850);
nand U3950 (N_3950,N_3872,N_3868);
nor U3951 (N_3951,N_3889,N_3811);
nor U3952 (N_3952,N_3812,N_3888);
or U3953 (N_3953,N_3817,N_3870);
nand U3954 (N_3954,N_3887,N_3879);
nand U3955 (N_3955,N_3801,N_3857);
and U3956 (N_3956,N_3867,N_3842);
and U3957 (N_3957,N_3889,N_3827);
nor U3958 (N_3958,N_3824,N_3882);
nor U3959 (N_3959,N_3828,N_3892);
or U3960 (N_3960,N_3862,N_3845);
xor U3961 (N_3961,N_3828,N_3856);
and U3962 (N_3962,N_3832,N_3893);
nor U3963 (N_3963,N_3800,N_3817);
nand U3964 (N_3964,N_3819,N_3860);
nor U3965 (N_3965,N_3824,N_3821);
and U3966 (N_3966,N_3841,N_3863);
nor U3967 (N_3967,N_3864,N_3814);
nor U3968 (N_3968,N_3839,N_3861);
nand U3969 (N_3969,N_3839,N_3803);
nand U3970 (N_3970,N_3833,N_3895);
nor U3971 (N_3971,N_3830,N_3829);
or U3972 (N_3972,N_3882,N_3855);
nor U3973 (N_3973,N_3826,N_3888);
or U3974 (N_3974,N_3847,N_3878);
or U3975 (N_3975,N_3869,N_3820);
and U3976 (N_3976,N_3885,N_3889);
and U3977 (N_3977,N_3835,N_3870);
xor U3978 (N_3978,N_3880,N_3895);
and U3979 (N_3979,N_3896,N_3872);
nor U3980 (N_3980,N_3847,N_3807);
nor U3981 (N_3981,N_3881,N_3859);
or U3982 (N_3982,N_3828,N_3810);
nor U3983 (N_3983,N_3866,N_3856);
nor U3984 (N_3984,N_3814,N_3840);
and U3985 (N_3985,N_3887,N_3822);
nor U3986 (N_3986,N_3849,N_3846);
and U3987 (N_3987,N_3882,N_3823);
nand U3988 (N_3988,N_3832,N_3837);
or U3989 (N_3989,N_3851,N_3881);
and U3990 (N_3990,N_3849,N_3888);
and U3991 (N_3991,N_3808,N_3874);
nand U3992 (N_3992,N_3871,N_3822);
nand U3993 (N_3993,N_3818,N_3873);
and U3994 (N_3994,N_3872,N_3898);
and U3995 (N_3995,N_3813,N_3844);
nor U3996 (N_3996,N_3876,N_3820);
nor U3997 (N_3997,N_3801,N_3811);
xnor U3998 (N_3998,N_3831,N_3862);
nor U3999 (N_3999,N_3887,N_3892);
nor U4000 (N_4000,N_3917,N_3930);
nand U4001 (N_4001,N_3936,N_3939);
nor U4002 (N_4002,N_3942,N_3967);
nand U4003 (N_4003,N_3998,N_3937);
and U4004 (N_4004,N_3924,N_3990);
nand U4005 (N_4005,N_3950,N_3916);
nand U4006 (N_4006,N_3904,N_3919);
or U4007 (N_4007,N_3925,N_3977);
nand U4008 (N_4008,N_3915,N_3932);
or U4009 (N_4009,N_3953,N_3928);
and U4010 (N_4010,N_3945,N_3906);
xnor U4011 (N_4011,N_3933,N_3980);
nand U4012 (N_4012,N_3991,N_3934);
or U4013 (N_4013,N_3970,N_3905);
nor U4014 (N_4014,N_3901,N_3976);
xor U4015 (N_4015,N_3927,N_3997);
and U4016 (N_4016,N_3903,N_3994);
or U4017 (N_4017,N_3913,N_3983);
and U4018 (N_4018,N_3964,N_3922);
nor U4019 (N_4019,N_3992,N_3959);
xor U4020 (N_4020,N_3918,N_3956);
xor U4021 (N_4021,N_3962,N_3946);
and U4022 (N_4022,N_3975,N_3902);
or U4023 (N_4023,N_3951,N_3944);
nand U4024 (N_4024,N_3973,N_3931);
xor U4025 (N_4025,N_3968,N_3971);
nand U4026 (N_4026,N_3978,N_3958);
nand U4027 (N_4027,N_3909,N_3940);
nor U4028 (N_4028,N_3974,N_3947);
and U4029 (N_4029,N_3943,N_3969);
and U4030 (N_4030,N_3979,N_3987);
nor U4031 (N_4031,N_3965,N_3955);
nor U4032 (N_4032,N_3938,N_3995);
nand U4033 (N_4033,N_3984,N_3985);
and U4034 (N_4034,N_3960,N_3993);
nor U4035 (N_4035,N_3966,N_3989);
nor U4036 (N_4036,N_3911,N_3941);
or U4037 (N_4037,N_3996,N_3986);
and U4038 (N_4038,N_3972,N_3999);
xnor U4039 (N_4039,N_3954,N_3957);
xnor U4040 (N_4040,N_3961,N_3921);
and U4041 (N_4041,N_3912,N_3920);
or U4042 (N_4042,N_3952,N_3929);
nor U4043 (N_4043,N_3935,N_3900);
and U4044 (N_4044,N_3926,N_3923);
nand U4045 (N_4045,N_3982,N_3981);
or U4046 (N_4046,N_3948,N_3907);
and U4047 (N_4047,N_3914,N_3988);
and U4048 (N_4048,N_3908,N_3949);
nor U4049 (N_4049,N_3910,N_3963);
nor U4050 (N_4050,N_3944,N_3969);
nand U4051 (N_4051,N_3919,N_3923);
nand U4052 (N_4052,N_3980,N_3913);
and U4053 (N_4053,N_3957,N_3923);
nand U4054 (N_4054,N_3906,N_3995);
nor U4055 (N_4055,N_3965,N_3990);
and U4056 (N_4056,N_3957,N_3900);
nor U4057 (N_4057,N_3933,N_3955);
and U4058 (N_4058,N_3982,N_3971);
or U4059 (N_4059,N_3967,N_3995);
or U4060 (N_4060,N_3938,N_3929);
nand U4061 (N_4061,N_3968,N_3980);
or U4062 (N_4062,N_3933,N_3994);
nor U4063 (N_4063,N_3979,N_3998);
and U4064 (N_4064,N_3941,N_3931);
nor U4065 (N_4065,N_3910,N_3978);
nor U4066 (N_4066,N_3947,N_3986);
or U4067 (N_4067,N_3932,N_3973);
nor U4068 (N_4068,N_3980,N_3962);
nor U4069 (N_4069,N_3986,N_3917);
nand U4070 (N_4070,N_3959,N_3921);
nand U4071 (N_4071,N_3999,N_3948);
nor U4072 (N_4072,N_3907,N_3931);
or U4073 (N_4073,N_3955,N_3945);
or U4074 (N_4074,N_3946,N_3992);
xnor U4075 (N_4075,N_3927,N_3978);
and U4076 (N_4076,N_3965,N_3944);
xnor U4077 (N_4077,N_3978,N_3962);
and U4078 (N_4078,N_3948,N_3954);
nor U4079 (N_4079,N_3983,N_3998);
or U4080 (N_4080,N_3913,N_3998);
xor U4081 (N_4081,N_3918,N_3978);
and U4082 (N_4082,N_3925,N_3948);
or U4083 (N_4083,N_3978,N_3948);
and U4084 (N_4084,N_3957,N_3912);
nor U4085 (N_4085,N_3994,N_3943);
nand U4086 (N_4086,N_3995,N_3952);
nor U4087 (N_4087,N_3964,N_3902);
and U4088 (N_4088,N_3985,N_3916);
nand U4089 (N_4089,N_3925,N_3931);
or U4090 (N_4090,N_3901,N_3939);
nor U4091 (N_4091,N_3924,N_3989);
or U4092 (N_4092,N_3953,N_3972);
nand U4093 (N_4093,N_3996,N_3917);
xor U4094 (N_4094,N_3918,N_3909);
and U4095 (N_4095,N_3975,N_3986);
nor U4096 (N_4096,N_3990,N_3926);
nor U4097 (N_4097,N_3968,N_3975);
nand U4098 (N_4098,N_3993,N_3954);
and U4099 (N_4099,N_3941,N_3980);
nand U4100 (N_4100,N_4032,N_4021);
nand U4101 (N_4101,N_4041,N_4099);
nor U4102 (N_4102,N_4045,N_4089);
nand U4103 (N_4103,N_4007,N_4027);
and U4104 (N_4104,N_4048,N_4012);
nand U4105 (N_4105,N_4001,N_4075);
xor U4106 (N_4106,N_4073,N_4005);
nor U4107 (N_4107,N_4093,N_4056);
xor U4108 (N_4108,N_4008,N_4016);
xnor U4109 (N_4109,N_4057,N_4025);
or U4110 (N_4110,N_4014,N_4072);
nor U4111 (N_4111,N_4039,N_4063);
nor U4112 (N_4112,N_4026,N_4061);
nor U4113 (N_4113,N_4029,N_4082);
or U4114 (N_4114,N_4004,N_4055);
nor U4115 (N_4115,N_4080,N_4047);
or U4116 (N_4116,N_4002,N_4023);
or U4117 (N_4117,N_4046,N_4017);
nand U4118 (N_4118,N_4062,N_4069);
nor U4119 (N_4119,N_4050,N_4053);
and U4120 (N_4120,N_4013,N_4003);
nor U4121 (N_4121,N_4054,N_4084);
and U4122 (N_4122,N_4051,N_4019);
or U4123 (N_4123,N_4030,N_4074);
or U4124 (N_4124,N_4092,N_4096);
and U4125 (N_4125,N_4037,N_4036);
nand U4126 (N_4126,N_4083,N_4000);
xnor U4127 (N_4127,N_4091,N_4024);
and U4128 (N_4128,N_4079,N_4040);
nand U4129 (N_4129,N_4087,N_4076);
nand U4130 (N_4130,N_4071,N_4035);
nor U4131 (N_4131,N_4067,N_4094);
and U4132 (N_4132,N_4011,N_4033);
nand U4133 (N_4133,N_4006,N_4085);
nand U4134 (N_4134,N_4086,N_4049);
nor U4135 (N_4135,N_4010,N_4031);
nor U4136 (N_4136,N_4044,N_4060);
nand U4137 (N_4137,N_4042,N_4090);
nand U4138 (N_4138,N_4043,N_4098);
nand U4139 (N_4139,N_4088,N_4034);
or U4140 (N_4140,N_4052,N_4077);
or U4141 (N_4141,N_4009,N_4058);
nor U4142 (N_4142,N_4066,N_4081);
and U4143 (N_4143,N_4020,N_4097);
nand U4144 (N_4144,N_4028,N_4064);
and U4145 (N_4145,N_4078,N_4068);
nor U4146 (N_4146,N_4070,N_4065);
nand U4147 (N_4147,N_4022,N_4059);
nand U4148 (N_4148,N_4018,N_4038);
or U4149 (N_4149,N_4015,N_4095);
nand U4150 (N_4150,N_4089,N_4059);
xor U4151 (N_4151,N_4069,N_4091);
nand U4152 (N_4152,N_4064,N_4026);
nor U4153 (N_4153,N_4073,N_4014);
nand U4154 (N_4154,N_4026,N_4050);
nand U4155 (N_4155,N_4034,N_4024);
nor U4156 (N_4156,N_4056,N_4022);
nand U4157 (N_4157,N_4038,N_4098);
or U4158 (N_4158,N_4059,N_4072);
xor U4159 (N_4159,N_4059,N_4051);
or U4160 (N_4160,N_4008,N_4038);
xnor U4161 (N_4161,N_4050,N_4025);
nand U4162 (N_4162,N_4044,N_4063);
nor U4163 (N_4163,N_4080,N_4032);
nor U4164 (N_4164,N_4015,N_4000);
or U4165 (N_4165,N_4081,N_4097);
nand U4166 (N_4166,N_4095,N_4012);
nor U4167 (N_4167,N_4026,N_4098);
nand U4168 (N_4168,N_4041,N_4048);
and U4169 (N_4169,N_4022,N_4096);
and U4170 (N_4170,N_4084,N_4077);
nor U4171 (N_4171,N_4029,N_4020);
or U4172 (N_4172,N_4082,N_4005);
nor U4173 (N_4173,N_4020,N_4064);
and U4174 (N_4174,N_4066,N_4009);
nand U4175 (N_4175,N_4034,N_4082);
nor U4176 (N_4176,N_4076,N_4030);
or U4177 (N_4177,N_4052,N_4072);
nor U4178 (N_4178,N_4027,N_4025);
xnor U4179 (N_4179,N_4014,N_4092);
or U4180 (N_4180,N_4090,N_4064);
nand U4181 (N_4181,N_4019,N_4049);
xnor U4182 (N_4182,N_4040,N_4023);
and U4183 (N_4183,N_4012,N_4056);
or U4184 (N_4184,N_4057,N_4029);
xor U4185 (N_4185,N_4093,N_4041);
nor U4186 (N_4186,N_4043,N_4096);
nor U4187 (N_4187,N_4040,N_4074);
and U4188 (N_4188,N_4015,N_4058);
nand U4189 (N_4189,N_4068,N_4033);
and U4190 (N_4190,N_4026,N_4046);
nand U4191 (N_4191,N_4061,N_4049);
xor U4192 (N_4192,N_4057,N_4081);
nand U4193 (N_4193,N_4070,N_4002);
nor U4194 (N_4194,N_4005,N_4034);
nand U4195 (N_4195,N_4018,N_4025);
and U4196 (N_4196,N_4035,N_4099);
and U4197 (N_4197,N_4087,N_4071);
nand U4198 (N_4198,N_4005,N_4051);
nor U4199 (N_4199,N_4068,N_4036);
nor U4200 (N_4200,N_4130,N_4104);
nand U4201 (N_4201,N_4101,N_4193);
nor U4202 (N_4202,N_4105,N_4143);
nor U4203 (N_4203,N_4138,N_4163);
or U4204 (N_4204,N_4103,N_4128);
and U4205 (N_4205,N_4183,N_4179);
nor U4206 (N_4206,N_4181,N_4172);
nand U4207 (N_4207,N_4127,N_4135);
and U4208 (N_4208,N_4190,N_4159);
or U4209 (N_4209,N_4165,N_4182);
and U4210 (N_4210,N_4116,N_4114);
nand U4211 (N_4211,N_4160,N_4144);
nor U4212 (N_4212,N_4155,N_4170);
nor U4213 (N_4213,N_4198,N_4121);
and U4214 (N_4214,N_4152,N_4123);
and U4215 (N_4215,N_4187,N_4147);
nand U4216 (N_4216,N_4186,N_4175);
xor U4217 (N_4217,N_4100,N_4176);
nand U4218 (N_4218,N_4197,N_4189);
or U4219 (N_4219,N_4196,N_4195);
nor U4220 (N_4220,N_4111,N_4120);
nand U4221 (N_4221,N_4137,N_4108);
or U4222 (N_4222,N_4199,N_4122);
and U4223 (N_4223,N_4157,N_4180);
and U4224 (N_4224,N_4113,N_4148);
nand U4225 (N_4225,N_4115,N_4149);
or U4226 (N_4226,N_4166,N_4188);
nand U4227 (N_4227,N_4129,N_4136);
and U4228 (N_4228,N_4146,N_4132);
or U4229 (N_4229,N_4185,N_4161);
and U4230 (N_4230,N_4178,N_4153);
nand U4231 (N_4231,N_4168,N_4133);
xor U4232 (N_4232,N_4194,N_4192);
nor U4233 (N_4233,N_4158,N_4124);
and U4234 (N_4234,N_4139,N_4164);
xor U4235 (N_4235,N_4167,N_4191);
xor U4236 (N_4236,N_4140,N_4162);
nor U4237 (N_4237,N_4106,N_4131);
nand U4238 (N_4238,N_4118,N_4171);
and U4239 (N_4239,N_4102,N_4177);
or U4240 (N_4240,N_4109,N_4184);
nor U4241 (N_4241,N_4150,N_4151);
nand U4242 (N_4242,N_4110,N_4145);
and U4243 (N_4243,N_4126,N_4134);
xor U4244 (N_4244,N_4156,N_4173);
nand U4245 (N_4245,N_4141,N_4169);
nand U4246 (N_4246,N_4117,N_4107);
nand U4247 (N_4247,N_4119,N_4142);
or U4248 (N_4248,N_4174,N_4154);
nor U4249 (N_4249,N_4125,N_4112);
and U4250 (N_4250,N_4143,N_4146);
or U4251 (N_4251,N_4193,N_4149);
nand U4252 (N_4252,N_4142,N_4156);
nand U4253 (N_4253,N_4187,N_4186);
nor U4254 (N_4254,N_4139,N_4173);
and U4255 (N_4255,N_4128,N_4155);
nand U4256 (N_4256,N_4193,N_4198);
and U4257 (N_4257,N_4112,N_4183);
nor U4258 (N_4258,N_4146,N_4153);
nand U4259 (N_4259,N_4138,N_4177);
and U4260 (N_4260,N_4164,N_4111);
nand U4261 (N_4261,N_4127,N_4177);
xnor U4262 (N_4262,N_4190,N_4191);
nor U4263 (N_4263,N_4125,N_4173);
nand U4264 (N_4264,N_4190,N_4132);
and U4265 (N_4265,N_4130,N_4152);
xor U4266 (N_4266,N_4148,N_4170);
nand U4267 (N_4267,N_4173,N_4140);
and U4268 (N_4268,N_4186,N_4100);
nor U4269 (N_4269,N_4193,N_4144);
nand U4270 (N_4270,N_4150,N_4183);
nand U4271 (N_4271,N_4144,N_4174);
or U4272 (N_4272,N_4154,N_4110);
nand U4273 (N_4273,N_4117,N_4110);
or U4274 (N_4274,N_4182,N_4177);
and U4275 (N_4275,N_4119,N_4160);
and U4276 (N_4276,N_4181,N_4129);
and U4277 (N_4277,N_4172,N_4152);
and U4278 (N_4278,N_4155,N_4138);
or U4279 (N_4279,N_4149,N_4120);
nand U4280 (N_4280,N_4112,N_4114);
and U4281 (N_4281,N_4170,N_4105);
nand U4282 (N_4282,N_4169,N_4132);
or U4283 (N_4283,N_4130,N_4103);
nor U4284 (N_4284,N_4163,N_4154);
nand U4285 (N_4285,N_4184,N_4195);
or U4286 (N_4286,N_4144,N_4139);
or U4287 (N_4287,N_4150,N_4145);
or U4288 (N_4288,N_4154,N_4129);
or U4289 (N_4289,N_4156,N_4165);
or U4290 (N_4290,N_4178,N_4154);
and U4291 (N_4291,N_4104,N_4157);
and U4292 (N_4292,N_4137,N_4144);
or U4293 (N_4293,N_4138,N_4181);
nor U4294 (N_4294,N_4141,N_4167);
nor U4295 (N_4295,N_4119,N_4125);
xnor U4296 (N_4296,N_4137,N_4135);
xor U4297 (N_4297,N_4172,N_4113);
or U4298 (N_4298,N_4181,N_4182);
nand U4299 (N_4299,N_4115,N_4192);
nor U4300 (N_4300,N_4273,N_4293);
nor U4301 (N_4301,N_4286,N_4299);
nor U4302 (N_4302,N_4265,N_4296);
nor U4303 (N_4303,N_4292,N_4242);
or U4304 (N_4304,N_4274,N_4221);
xor U4305 (N_4305,N_4263,N_4230);
nand U4306 (N_4306,N_4211,N_4257);
or U4307 (N_4307,N_4244,N_4264);
and U4308 (N_4308,N_4222,N_4297);
nand U4309 (N_4309,N_4258,N_4232);
nor U4310 (N_4310,N_4216,N_4250);
and U4311 (N_4311,N_4248,N_4226);
or U4312 (N_4312,N_4231,N_4288);
or U4313 (N_4313,N_4215,N_4236);
and U4314 (N_4314,N_4253,N_4219);
and U4315 (N_4315,N_4285,N_4278);
or U4316 (N_4316,N_4251,N_4280);
nor U4317 (N_4317,N_4256,N_4246);
nor U4318 (N_4318,N_4213,N_4233);
or U4319 (N_4319,N_4247,N_4268);
nand U4320 (N_4320,N_4243,N_4209);
and U4321 (N_4321,N_4212,N_4239);
or U4322 (N_4322,N_4262,N_4270);
nand U4323 (N_4323,N_4291,N_4290);
nor U4324 (N_4324,N_4240,N_4217);
and U4325 (N_4325,N_4252,N_4295);
nor U4326 (N_4326,N_4284,N_4279);
nor U4327 (N_4327,N_4261,N_4289);
nand U4328 (N_4328,N_4224,N_4218);
nor U4329 (N_4329,N_4241,N_4237);
or U4330 (N_4330,N_4249,N_4201);
nand U4331 (N_4331,N_4260,N_4254);
and U4332 (N_4332,N_4234,N_4275);
nand U4333 (N_4333,N_4229,N_4210);
and U4334 (N_4334,N_4294,N_4205);
nor U4335 (N_4335,N_4266,N_4225);
or U4336 (N_4336,N_4204,N_4206);
nor U4337 (N_4337,N_4283,N_4271);
nor U4338 (N_4338,N_4277,N_4207);
or U4339 (N_4339,N_4202,N_4220);
nand U4340 (N_4340,N_4267,N_4298);
and U4341 (N_4341,N_4259,N_4228);
and U4342 (N_4342,N_4203,N_4272);
or U4343 (N_4343,N_4281,N_4223);
or U4344 (N_4344,N_4287,N_4200);
and U4345 (N_4345,N_4276,N_4255);
and U4346 (N_4346,N_4245,N_4227);
or U4347 (N_4347,N_4235,N_4238);
and U4348 (N_4348,N_4282,N_4208);
xor U4349 (N_4349,N_4269,N_4214);
nor U4350 (N_4350,N_4288,N_4258);
nor U4351 (N_4351,N_4264,N_4294);
nor U4352 (N_4352,N_4271,N_4255);
or U4353 (N_4353,N_4212,N_4242);
or U4354 (N_4354,N_4295,N_4218);
nor U4355 (N_4355,N_4244,N_4206);
nor U4356 (N_4356,N_4211,N_4217);
nor U4357 (N_4357,N_4252,N_4294);
nand U4358 (N_4358,N_4293,N_4223);
or U4359 (N_4359,N_4226,N_4243);
nand U4360 (N_4360,N_4236,N_4204);
nor U4361 (N_4361,N_4244,N_4288);
nor U4362 (N_4362,N_4244,N_4260);
nand U4363 (N_4363,N_4280,N_4243);
nand U4364 (N_4364,N_4288,N_4282);
nor U4365 (N_4365,N_4261,N_4275);
or U4366 (N_4366,N_4207,N_4210);
and U4367 (N_4367,N_4227,N_4207);
or U4368 (N_4368,N_4267,N_4296);
nand U4369 (N_4369,N_4215,N_4257);
nor U4370 (N_4370,N_4212,N_4250);
nor U4371 (N_4371,N_4273,N_4255);
nor U4372 (N_4372,N_4231,N_4272);
or U4373 (N_4373,N_4246,N_4290);
nand U4374 (N_4374,N_4203,N_4278);
nor U4375 (N_4375,N_4275,N_4245);
nand U4376 (N_4376,N_4245,N_4290);
and U4377 (N_4377,N_4237,N_4220);
nand U4378 (N_4378,N_4258,N_4265);
or U4379 (N_4379,N_4209,N_4233);
and U4380 (N_4380,N_4236,N_4299);
or U4381 (N_4381,N_4263,N_4213);
and U4382 (N_4382,N_4274,N_4250);
xor U4383 (N_4383,N_4259,N_4286);
or U4384 (N_4384,N_4265,N_4241);
and U4385 (N_4385,N_4264,N_4254);
or U4386 (N_4386,N_4277,N_4213);
or U4387 (N_4387,N_4230,N_4209);
and U4388 (N_4388,N_4291,N_4203);
nor U4389 (N_4389,N_4237,N_4277);
nor U4390 (N_4390,N_4210,N_4271);
or U4391 (N_4391,N_4268,N_4222);
or U4392 (N_4392,N_4287,N_4235);
nor U4393 (N_4393,N_4294,N_4280);
and U4394 (N_4394,N_4205,N_4209);
or U4395 (N_4395,N_4223,N_4276);
or U4396 (N_4396,N_4240,N_4205);
nor U4397 (N_4397,N_4269,N_4237);
nand U4398 (N_4398,N_4245,N_4288);
nand U4399 (N_4399,N_4269,N_4210);
and U4400 (N_4400,N_4367,N_4375);
and U4401 (N_4401,N_4384,N_4352);
or U4402 (N_4402,N_4338,N_4381);
or U4403 (N_4403,N_4368,N_4306);
or U4404 (N_4404,N_4399,N_4359);
and U4405 (N_4405,N_4353,N_4309);
nor U4406 (N_4406,N_4350,N_4330);
xor U4407 (N_4407,N_4337,N_4312);
nor U4408 (N_4408,N_4383,N_4374);
nor U4409 (N_4409,N_4328,N_4391);
nand U4410 (N_4410,N_4394,N_4346);
nand U4411 (N_4411,N_4378,N_4348);
nand U4412 (N_4412,N_4322,N_4372);
or U4413 (N_4413,N_4389,N_4339);
or U4414 (N_4414,N_4379,N_4371);
and U4415 (N_4415,N_4377,N_4315);
or U4416 (N_4416,N_4363,N_4304);
or U4417 (N_4417,N_4398,N_4369);
and U4418 (N_4418,N_4347,N_4303);
nand U4419 (N_4419,N_4390,N_4329);
nand U4420 (N_4420,N_4321,N_4333);
and U4421 (N_4421,N_4385,N_4317);
or U4422 (N_4422,N_4326,N_4319);
or U4423 (N_4423,N_4366,N_4331);
and U4424 (N_4424,N_4356,N_4358);
nand U4425 (N_4425,N_4313,N_4364);
nor U4426 (N_4426,N_4365,N_4361);
nand U4427 (N_4427,N_4314,N_4362);
nand U4428 (N_4428,N_4327,N_4334);
nand U4429 (N_4429,N_4336,N_4341);
and U4430 (N_4430,N_4395,N_4344);
nand U4431 (N_4431,N_4380,N_4354);
nand U4432 (N_4432,N_4397,N_4387);
nand U4433 (N_4433,N_4355,N_4396);
xnor U4434 (N_4434,N_4301,N_4382);
xor U4435 (N_4435,N_4386,N_4345);
or U4436 (N_4436,N_4335,N_4370);
or U4437 (N_4437,N_4324,N_4308);
nand U4438 (N_4438,N_4342,N_4318);
nor U4439 (N_4439,N_4302,N_4357);
and U4440 (N_4440,N_4392,N_4325);
nor U4441 (N_4441,N_4311,N_4373);
nand U4442 (N_4442,N_4310,N_4340);
xnor U4443 (N_4443,N_4343,N_4360);
nand U4444 (N_4444,N_4349,N_4316);
xnor U4445 (N_4445,N_4376,N_4323);
xor U4446 (N_4446,N_4393,N_4300);
and U4447 (N_4447,N_4305,N_4351);
nor U4448 (N_4448,N_4307,N_4388);
or U4449 (N_4449,N_4320,N_4332);
and U4450 (N_4450,N_4373,N_4357);
and U4451 (N_4451,N_4378,N_4324);
nand U4452 (N_4452,N_4310,N_4386);
nand U4453 (N_4453,N_4391,N_4377);
or U4454 (N_4454,N_4332,N_4330);
or U4455 (N_4455,N_4381,N_4321);
nor U4456 (N_4456,N_4389,N_4374);
or U4457 (N_4457,N_4336,N_4374);
or U4458 (N_4458,N_4334,N_4302);
and U4459 (N_4459,N_4322,N_4351);
xor U4460 (N_4460,N_4361,N_4308);
and U4461 (N_4461,N_4384,N_4333);
or U4462 (N_4462,N_4303,N_4364);
nand U4463 (N_4463,N_4333,N_4361);
and U4464 (N_4464,N_4385,N_4354);
and U4465 (N_4465,N_4355,N_4347);
or U4466 (N_4466,N_4332,N_4390);
and U4467 (N_4467,N_4308,N_4388);
or U4468 (N_4468,N_4366,N_4318);
or U4469 (N_4469,N_4394,N_4328);
xnor U4470 (N_4470,N_4326,N_4347);
and U4471 (N_4471,N_4356,N_4322);
and U4472 (N_4472,N_4375,N_4363);
or U4473 (N_4473,N_4347,N_4357);
and U4474 (N_4474,N_4361,N_4332);
and U4475 (N_4475,N_4385,N_4324);
nor U4476 (N_4476,N_4357,N_4324);
nor U4477 (N_4477,N_4324,N_4300);
or U4478 (N_4478,N_4355,N_4358);
nor U4479 (N_4479,N_4349,N_4342);
or U4480 (N_4480,N_4304,N_4361);
nand U4481 (N_4481,N_4341,N_4381);
xor U4482 (N_4482,N_4387,N_4331);
or U4483 (N_4483,N_4352,N_4360);
nor U4484 (N_4484,N_4347,N_4319);
nand U4485 (N_4485,N_4322,N_4332);
xnor U4486 (N_4486,N_4351,N_4381);
and U4487 (N_4487,N_4305,N_4387);
xor U4488 (N_4488,N_4392,N_4381);
nand U4489 (N_4489,N_4319,N_4353);
or U4490 (N_4490,N_4354,N_4335);
or U4491 (N_4491,N_4331,N_4305);
or U4492 (N_4492,N_4361,N_4395);
nor U4493 (N_4493,N_4378,N_4304);
xnor U4494 (N_4494,N_4314,N_4312);
nand U4495 (N_4495,N_4390,N_4353);
nand U4496 (N_4496,N_4350,N_4333);
xor U4497 (N_4497,N_4307,N_4321);
xor U4498 (N_4498,N_4396,N_4337);
nand U4499 (N_4499,N_4376,N_4314);
and U4500 (N_4500,N_4408,N_4420);
and U4501 (N_4501,N_4496,N_4424);
nand U4502 (N_4502,N_4449,N_4441);
nor U4503 (N_4503,N_4416,N_4461);
xnor U4504 (N_4504,N_4433,N_4409);
and U4505 (N_4505,N_4467,N_4415);
nor U4506 (N_4506,N_4469,N_4491);
nand U4507 (N_4507,N_4498,N_4473);
or U4508 (N_4508,N_4426,N_4410);
or U4509 (N_4509,N_4471,N_4456);
nor U4510 (N_4510,N_4445,N_4484);
or U4511 (N_4511,N_4482,N_4468);
nor U4512 (N_4512,N_4497,N_4428);
xor U4513 (N_4513,N_4417,N_4460);
or U4514 (N_4514,N_4413,N_4439);
xnor U4515 (N_4515,N_4442,N_4404);
or U4516 (N_4516,N_4485,N_4400);
nor U4517 (N_4517,N_4458,N_4477);
nand U4518 (N_4518,N_4405,N_4444);
nand U4519 (N_4519,N_4488,N_4462);
nor U4520 (N_4520,N_4494,N_4483);
or U4521 (N_4521,N_4435,N_4479);
and U4522 (N_4522,N_4440,N_4411);
nand U4523 (N_4523,N_4447,N_4443);
and U4524 (N_4524,N_4475,N_4434);
and U4525 (N_4525,N_4455,N_4407);
and U4526 (N_4526,N_4478,N_4402);
and U4527 (N_4527,N_4463,N_4425);
and U4528 (N_4528,N_4486,N_4421);
nor U4529 (N_4529,N_4457,N_4436);
or U4530 (N_4530,N_4437,N_4430);
nor U4531 (N_4531,N_4452,N_4472);
nand U4532 (N_4532,N_4451,N_4470);
nor U4533 (N_4533,N_4490,N_4466);
nand U4534 (N_4534,N_4474,N_4489);
or U4535 (N_4535,N_4480,N_4414);
nand U4536 (N_4536,N_4459,N_4481);
nor U4537 (N_4537,N_4499,N_4454);
and U4538 (N_4538,N_4401,N_4487);
nor U4539 (N_4539,N_4432,N_4495);
or U4540 (N_4540,N_4423,N_4492);
and U4541 (N_4541,N_4412,N_4464);
nor U4542 (N_4542,N_4429,N_4431);
nand U4543 (N_4543,N_4406,N_4418);
nor U4544 (N_4544,N_4438,N_4453);
and U4545 (N_4545,N_4493,N_4419);
nand U4546 (N_4546,N_4476,N_4446);
and U4547 (N_4547,N_4465,N_4427);
nand U4548 (N_4548,N_4448,N_4450);
nand U4549 (N_4549,N_4422,N_4403);
and U4550 (N_4550,N_4400,N_4414);
nor U4551 (N_4551,N_4484,N_4499);
and U4552 (N_4552,N_4477,N_4424);
nor U4553 (N_4553,N_4420,N_4467);
nand U4554 (N_4554,N_4468,N_4490);
and U4555 (N_4555,N_4415,N_4447);
or U4556 (N_4556,N_4494,N_4476);
or U4557 (N_4557,N_4443,N_4427);
nor U4558 (N_4558,N_4411,N_4456);
or U4559 (N_4559,N_4403,N_4429);
xnor U4560 (N_4560,N_4452,N_4464);
or U4561 (N_4561,N_4495,N_4441);
nor U4562 (N_4562,N_4427,N_4488);
and U4563 (N_4563,N_4432,N_4438);
or U4564 (N_4564,N_4499,N_4485);
and U4565 (N_4565,N_4401,N_4494);
xor U4566 (N_4566,N_4463,N_4441);
or U4567 (N_4567,N_4428,N_4429);
or U4568 (N_4568,N_4497,N_4488);
or U4569 (N_4569,N_4454,N_4451);
nor U4570 (N_4570,N_4437,N_4457);
xnor U4571 (N_4571,N_4464,N_4486);
nand U4572 (N_4572,N_4493,N_4436);
or U4573 (N_4573,N_4475,N_4478);
and U4574 (N_4574,N_4439,N_4463);
nor U4575 (N_4575,N_4418,N_4430);
xnor U4576 (N_4576,N_4453,N_4487);
and U4577 (N_4577,N_4489,N_4482);
or U4578 (N_4578,N_4437,N_4409);
nor U4579 (N_4579,N_4415,N_4464);
nand U4580 (N_4580,N_4429,N_4495);
or U4581 (N_4581,N_4443,N_4435);
or U4582 (N_4582,N_4418,N_4411);
and U4583 (N_4583,N_4464,N_4408);
or U4584 (N_4584,N_4426,N_4452);
nor U4585 (N_4585,N_4428,N_4443);
nor U4586 (N_4586,N_4469,N_4475);
or U4587 (N_4587,N_4463,N_4466);
nor U4588 (N_4588,N_4441,N_4411);
and U4589 (N_4589,N_4492,N_4420);
nor U4590 (N_4590,N_4476,N_4495);
or U4591 (N_4591,N_4477,N_4426);
nand U4592 (N_4592,N_4405,N_4404);
xnor U4593 (N_4593,N_4405,N_4411);
and U4594 (N_4594,N_4431,N_4450);
or U4595 (N_4595,N_4445,N_4473);
and U4596 (N_4596,N_4473,N_4482);
xor U4597 (N_4597,N_4485,N_4458);
nor U4598 (N_4598,N_4454,N_4449);
or U4599 (N_4599,N_4446,N_4407);
nand U4600 (N_4600,N_4553,N_4596);
or U4601 (N_4601,N_4526,N_4599);
and U4602 (N_4602,N_4581,N_4559);
nor U4603 (N_4603,N_4584,N_4514);
or U4604 (N_4604,N_4594,N_4527);
xnor U4605 (N_4605,N_4576,N_4525);
nand U4606 (N_4606,N_4564,N_4516);
nand U4607 (N_4607,N_4565,N_4580);
nor U4608 (N_4608,N_4546,N_4552);
nand U4609 (N_4609,N_4508,N_4515);
and U4610 (N_4610,N_4535,N_4517);
nor U4611 (N_4611,N_4561,N_4536);
nor U4612 (N_4612,N_4533,N_4543);
nand U4613 (N_4613,N_4502,N_4542);
or U4614 (N_4614,N_4569,N_4540);
and U4615 (N_4615,N_4597,N_4510);
nand U4616 (N_4616,N_4504,N_4587);
and U4617 (N_4617,N_4529,N_4549);
and U4618 (N_4618,N_4560,N_4550);
nor U4619 (N_4619,N_4588,N_4520);
or U4620 (N_4620,N_4562,N_4573);
nor U4621 (N_4621,N_4575,N_4500);
nor U4622 (N_4622,N_4501,N_4590);
or U4623 (N_4623,N_4571,N_4589);
xnor U4624 (N_4624,N_4503,N_4505);
or U4625 (N_4625,N_4556,N_4583);
and U4626 (N_4626,N_4577,N_4544);
nand U4627 (N_4627,N_4528,N_4523);
or U4628 (N_4628,N_4511,N_4585);
and U4629 (N_4629,N_4545,N_4551);
nand U4630 (N_4630,N_4579,N_4595);
and U4631 (N_4631,N_4530,N_4563);
nand U4632 (N_4632,N_4537,N_4572);
xnor U4633 (N_4633,N_4507,N_4586);
nor U4634 (N_4634,N_4538,N_4519);
nor U4635 (N_4635,N_4518,N_4591);
nor U4636 (N_4636,N_4592,N_4532);
nand U4637 (N_4637,N_4541,N_4568);
or U4638 (N_4638,N_4554,N_4522);
or U4639 (N_4639,N_4598,N_4555);
nand U4640 (N_4640,N_4512,N_4582);
nor U4641 (N_4641,N_4570,N_4548);
nand U4642 (N_4642,N_4558,N_4534);
nor U4643 (N_4643,N_4557,N_4578);
xor U4644 (N_4644,N_4513,N_4509);
and U4645 (N_4645,N_4566,N_4539);
xor U4646 (N_4646,N_4567,N_4547);
nand U4647 (N_4647,N_4574,N_4531);
nand U4648 (N_4648,N_4521,N_4506);
nor U4649 (N_4649,N_4593,N_4524);
and U4650 (N_4650,N_4514,N_4537);
and U4651 (N_4651,N_4560,N_4582);
and U4652 (N_4652,N_4547,N_4587);
nor U4653 (N_4653,N_4517,N_4558);
or U4654 (N_4654,N_4596,N_4562);
xnor U4655 (N_4655,N_4569,N_4506);
or U4656 (N_4656,N_4552,N_4567);
and U4657 (N_4657,N_4531,N_4576);
or U4658 (N_4658,N_4534,N_4516);
and U4659 (N_4659,N_4528,N_4550);
nand U4660 (N_4660,N_4554,N_4520);
nand U4661 (N_4661,N_4560,N_4528);
xor U4662 (N_4662,N_4526,N_4569);
or U4663 (N_4663,N_4594,N_4570);
nand U4664 (N_4664,N_4595,N_4585);
or U4665 (N_4665,N_4568,N_4504);
nand U4666 (N_4666,N_4573,N_4539);
nand U4667 (N_4667,N_4520,N_4536);
and U4668 (N_4668,N_4548,N_4590);
nand U4669 (N_4669,N_4573,N_4508);
nor U4670 (N_4670,N_4560,N_4531);
or U4671 (N_4671,N_4578,N_4549);
nand U4672 (N_4672,N_4503,N_4593);
and U4673 (N_4673,N_4550,N_4577);
or U4674 (N_4674,N_4590,N_4504);
xor U4675 (N_4675,N_4520,N_4543);
nand U4676 (N_4676,N_4521,N_4545);
or U4677 (N_4677,N_4540,N_4507);
and U4678 (N_4678,N_4503,N_4566);
nor U4679 (N_4679,N_4510,N_4512);
nand U4680 (N_4680,N_4524,N_4500);
or U4681 (N_4681,N_4596,N_4558);
nor U4682 (N_4682,N_4542,N_4531);
or U4683 (N_4683,N_4543,N_4567);
or U4684 (N_4684,N_4543,N_4505);
and U4685 (N_4685,N_4573,N_4507);
or U4686 (N_4686,N_4551,N_4544);
and U4687 (N_4687,N_4544,N_4534);
and U4688 (N_4688,N_4503,N_4510);
xor U4689 (N_4689,N_4566,N_4596);
and U4690 (N_4690,N_4519,N_4501);
xnor U4691 (N_4691,N_4598,N_4581);
or U4692 (N_4692,N_4500,N_4565);
and U4693 (N_4693,N_4592,N_4573);
or U4694 (N_4694,N_4517,N_4508);
or U4695 (N_4695,N_4501,N_4582);
or U4696 (N_4696,N_4579,N_4533);
xnor U4697 (N_4697,N_4579,N_4530);
and U4698 (N_4698,N_4501,N_4579);
or U4699 (N_4699,N_4560,N_4557);
nor U4700 (N_4700,N_4659,N_4666);
xor U4701 (N_4701,N_4671,N_4670);
xnor U4702 (N_4702,N_4635,N_4678);
and U4703 (N_4703,N_4665,N_4660);
or U4704 (N_4704,N_4610,N_4656);
nand U4705 (N_4705,N_4694,N_4650);
or U4706 (N_4706,N_4686,N_4624);
nand U4707 (N_4707,N_4693,N_4631);
nand U4708 (N_4708,N_4628,N_4661);
or U4709 (N_4709,N_4695,N_4629);
or U4710 (N_4710,N_4618,N_4684);
or U4711 (N_4711,N_4607,N_4603);
and U4712 (N_4712,N_4625,N_4675);
and U4713 (N_4713,N_4609,N_4657);
nor U4714 (N_4714,N_4680,N_4622);
nor U4715 (N_4715,N_4600,N_4667);
nor U4716 (N_4716,N_4692,N_4652);
or U4717 (N_4717,N_4651,N_4687);
and U4718 (N_4718,N_4617,N_4672);
nor U4719 (N_4719,N_4654,N_4682);
or U4720 (N_4720,N_4679,N_4698);
nand U4721 (N_4721,N_4606,N_4604);
nor U4722 (N_4722,N_4602,N_4611);
nor U4723 (N_4723,N_4608,N_4674);
nand U4724 (N_4724,N_4627,N_4649);
or U4725 (N_4725,N_4653,N_4676);
nand U4726 (N_4726,N_4688,N_4668);
nor U4727 (N_4727,N_4612,N_4632);
nand U4728 (N_4728,N_4646,N_4699);
or U4729 (N_4729,N_4639,N_4615);
nand U4730 (N_4730,N_4658,N_4633);
nand U4731 (N_4731,N_4636,N_4643);
nand U4732 (N_4732,N_4689,N_4638);
and U4733 (N_4733,N_4662,N_4621);
or U4734 (N_4734,N_4681,N_4620);
nand U4735 (N_4735,N_4644,N_4630);
and U4736 (N_4736,N_4616,N_4634);
nand U4737 (N_4737,N_4673,N_4685);
nand U4738 (N_4738,N_4683,N_4623);
nand U4739 (N_4739,N_4663,N_4664);
nor U4740 (N_4740,N_4696,N_4613);
and U4741 (N_4741,N_4626,N_4605);
xor U4742 (N_4742,N_4691,N_4614);
nand U4743 (N_4743,N_4641,N_4645);
xor U4744 (N_4744,N_4669,N_4647);
and U4745 (N_4745,N_4655,N_4619);
nand U4746 (N_4746,N_4642,N_4677);
nand U4747 (N_4747,N_4637,N_4640);
or U4748 (N_4748,N_4690,N_4697);
and U4749 (N_4749,N_4601,N_4648);
and U4750 (N_4750,N_4646,N_4661);
or U4751 (N_4751,N_4635,N_4611);
nor U4752 (N_4752,N_4600,N_4619);
and U4753 (N_4753,N_4673,N_4614);
nand U4754 (N_4754,N_4607,N_4672);
or U4755 (N_4755,N_4688,N_4606);
nor U4756 (N_4756,N_4615,N_4637);
nor U4757 (N_4757,N_4654,N_4680);
nand U4758 (N_4758,N_4651,N_4600);
nand U4759 (N_4759,N_4659,N_4647);
xor U4760 (N_4760,N_4657,N_4641);
nand U4761 (N_4761,N_4631,N_4664);
and U4762 (N_4762,N_4619,N_4654);
and U4763 (N_4763,N_4692,N_4607);
or U4764 (N_4764,N_4664,N_4680);
or U4765 (N_4765,N_4666,N_4603);
nand U4766 (N_4766,N_4642,N_4665);
nand U4767 (N_4767,N_4683,N_4650);
nor U4768 (N_4768,N_4647,N_4625);
nand U4769 (N_4769,N_4604,N_4643);
nor U4770 (N_4770,N_4664,N_4628);
nor U4771 (N_4771,N_4609,N_4623);
and U4772 (N_4772,N_4649,N_4677);
or U4773 (N_4773,N_4620,N_4669);
nor U4774 (N_4774,N_4680,N_4647);
or U4775 (N_4775,N_4606,N_4645);
or U4776 (N_4776,N_4634,N_4694);
nand U4777 (N_4777,N_4697,N_4691);
or U4778 (N_4778,N_4670,N_4642);
nor U4779 (N_4779,N_4641,N_4626);
nor U4780 (N_4780,N_4672,N_4692);
nand U4781 (N_4781,N_4688,N_4634);
nand U4782 (N_4782,N_4647,N_4672);
nor U4783 (N_4783,N_4678,N_4692);
nand U4784 (N_4784,N_4626,N_4646);
nor U4785 (N_4785,N_4638,N_4666);
xor U4786 (N_4786,N_4679,N_4674);
nand U4787 (N_4787,N_4680,N_4623);
or U4788 (N_4788,N_4600,N_4649);
nor U4789 (N_4789,N_4694,N_4659);
nor U4790 (N_4790,N_4686,N_4618);
nand U4791 (N_4791,N_4618,N_4641);
xnor U4792 (N_4792,N_4632,N_4660);
or U4793 (N_4793,N_4637,N_4627);
nor U4794 (N_4794,N_4681,N_4619);
or U4795 (N_4795,N_4650,N_4647);
nand U4796 (N_4796,N_4620,N_4699);
or U4797 (N_4797,N_4634,N_4627);
xor U4798 (N_4798,N_4680,N_4661);
or U4799 (N_4799,N_4680,N_4652);
nand U4800 (N_4800,N_4799,N_4766);
nor U4801 (N_4801,N_4747,N_4763);
nand U4802 (N_4802,N_4717,N_4791);
and U4803 (N_4803,N_4740,N_4708);
nor U4804 (N_4804,N_4758,N_4737);
and U4805 (N_4805,N_4782,N_4769);
nand U4806 (N_4806,N_4785,N_4728);
nor U4807 (N_4807,N_4727,N_4724);
nand U4808 (N_4808,N_4706,N_4729);
and U4809 (N_4809,N_4722,N_4721);
nand U4810 (N_4810,N_4783,N_4751);
xnor U4811 (N_4811,N_4762,N_4732);
and U4812 (N_4812,N_4794,N_4773);
or U4813 (N_4813,N_4718,N_4771);
and U4814 (N_4814,N_4746,N_4749);
xor U4815 (N_4815,N_4712,N_4784);
nand U4816 (N_4816,N_4792,N_4700);
or U4817 (N_4817,N_4754,N_4701);
and U4818 (N_4818,N_4767,N_4704);
nor U4819 (N_4819,N_4743,N_4755);
nand U4820 (N_4820,N_4715,N_4714);
nor U4821 (N_4821,N_4793,N_4770);
or U4822 (N_4822,N_4707,N_4703);
or U4823 (N_4823,N_4781,N_4786);
nand U4824 (N_4824,N_4705,N_4735);
xnor U4825 (N_4825,N_4716,N_4789);
nor U4826 (N_4826,N_4733,N_4726);
and U4827 (N_4827,N_4730,N_4795);
or U4828 (N_4828,N_4738,N_4702);
nand U4829 (N_4829,N_4752,N_4760);
nand U4830 (N_4830,N_4768,N_4797);
xnor U4831 (N_4831,N_4796,N_4775);
nor U4832 (N_4832,N_4761,N_4779);
and U4833 (N_4833,N_4776,N_4753);
nand U4834 (N_4834,N_4759,N_4744);
nor U4835 (N_4835,N_4765,N_4720);
nor U4836 (N_4836,N_4788,N_4772);
or U4837 (N_4837,N_4790,N_4780);
nand U4838 (N_4838,N_4745,N_4757);
and U4839 (N_4839,N_4709,N_4723);
nor U4840 (N_4840,N_4774,N_4739);
nand U4841 (N_4841,N_4756,N_4798);
nor U4842 (N_4842,N_4719,N_4710);
or U4843 (N_4843,N_4731,N_4713);
nor U4844 (N_4844,N_4777,N_4711);
and U4845 (N_4845,N_4750,N_4748);
nor U4846 (N_4846,N_4736,N_4741);
or U4847 (N_4847,N_4734,N_4725);
xnor U4848 (N_4848,N_4778,N_4787);
and U4849 (N_4849,N_4742,N_4764);
and U4850 (N_4850,N_4758,N_4734);
or U4851 (N_4851,N_4769,N_4756);
and U4852 (N_4852,N_4786,N_4751);
and U4853 (N_4853,N_4798,N_4783);
nand U4854 (N_4854,N_4754,N_4769);
and U4855 (N_4855,N_4701,N_4772);
or U4856 (N_4856,N_4746,N_4794);
nand U4857 (N_4857,N_4772,N_4746);
nand U4858 (N_4858,N_4705,N_4791);
nand U4859 (N_4859,N_4756,N_4797);
or U4860 (N_4860,N_4749,N_4721);
and U4861 (N_4861,N_4704,N_4724);
nand U4862 (N_4862,N_4708,N_4747);
nor U4863 (N_4863,N_4797,N_4705);
xor U4864 (N_4864,N_4706,N_4745);
nand U4865 (N_4865,N_4741,N_4747);
nor U4866 (N_4866,N_4770,N_4749);
nor U4867 (N_4867,N_4706,N_4791);
and U4868 (N_4868,N_4757,N_4706);
nand U4869 (N_4869,N_4705,N_4734);
nor U4870 (N_4870,N_4714,N_4725);
or U4871 (N_4871,N_4744,N_4733);
nand U4872 (N_4872,N_4788,N_4728);
and U4873 (N_4873,N_4756,N_4781);
nor U4874 (N_4874,N_4771,N_4716);
nor U4875 (N_4875,N_4790,N_4788);
nor U4876 (N_4876,N_4722,N_4701);
or U4877 (N_4877,N_4756,N_4729);
nor U4878 (N_4878,N_4784,N_4730);
and U4879 (N_4879,N_4712,N_4796);
nand U4880 (N_4880,N_4729,N_4750);
nor U4881 (N_4881,N_4745,N_4755);
or U4882 (N_4882,N_4715,N_4739);
and U4883 (N_4883,N_4768,N_4721);
or U4884 (N_4884,N_4745,N_4797);
or U4885 (N_4885,N_4737,N_4721);
nand U4886 (N_4886,N_4754,N_4732);
nand U4887 (N_4887,N_4700,N_4769);
and U4888 (N_4888,N_4766,N_4756);
nor U4889 (N_4889,N_4769,N_4757);
nor U4890 (N_4890,N_4765,N_4781);
nor U4891 (N_4891,N_4743,N_4739);
nand U4892 (N_4892,N_4757,N_4753);
nand U4893 (N_4893,N_4777,N_4778);
nand U4894 (N_4894,N_4775,N_4745);
and U4895 (N_4895,N_4714,N_4735);
and U4896 (N_4896,N_4731,N_4754);
or U4897 (N_4897,N_4798,N_4728);
nor U4898 (N_4898,N_4772,N_4700);
and U4899 (N_4899,N_4712,N_4720);
nor U4900 (N_4900,N_4835,N_4867);
or U4901 (N_4901,N_4880,N_4877);
and U4902 (N_4902,N_4853,N_4852);
nor U4903 (N_4903,N_4895,N_4823);
nor U4904 (N_4904,N_4854,N_4818);
and U4905 (N_4905,N_4817,N_4862);
or U4906 (N_4906,N_4861,N_4879);
nand U4907 (N_4907,N_4856,N_4884);
nor U4908 (N_4908,N_4891,N_4869);
nor U4909 (N_4909,N_4808,N_4810);
and U4910 (N_4910,N_4830,N_4829);
or U4911 (N_4911,N_4868,N_4834);
or U4912 (N_4912,N_4894,N_4863);
nor U4913 (N_4913,N_4885,N_4836);
and U4914 (N_4914,N_4832,N_4848);
nor U4915 (N_4915,N_4888,N_4815);
nand U4916 (N_4916,N_4842,N_4871);
xor U4917 (N_4917,N_4831,N_4865);
or U4918 (N_4918,N_4846,N_4813);
or U4919 (N_4919,N_4821,N_4866);
nor U4920 (N_4920,N_4857,N_4827);
or U4921 (N_4921,N_4822,N_4825);
nor U4922 (N_4922,N_4893,N_4841);
or U4923 (N_4923,N_4859,N_4864);
nand U4924 (N_4924,N_4839,N_4883);
nor U4925 (N_4925,N_4896,N_4803);
or U4926 (N_4926,N_4897,N_4845);
nand U4927 (N_4927,N_4824,N_4881);
nor U4928 (N_4928,N_4840,N_4882);
and U4929 (N_4929,N_4814,N_4860);
nand U4930 (N_4930,N_4875,N_4802);
xnor U4931 (N_4931,N_4849,N_4892);
and U4932 (N_4932,N_4843,N_4801);
and U4933 (N_4933,N_4826,N_4858);
and U4934 (N_4934,N_4819,N_4889);
nor U4935 (N_4935,N_4872,N_4873);
nor U4936 (N_4936,N_4812,N_4820);
and U4937 (N_4937,N_4828,N_4838);
xnor U4938 (N_4938,N_4850,N_4809);
or U4939 (N_4939,N_4816,N_4887);
nor U4940 (N_4940,N_4804,N_4844);
or U4941 (N_4941,N_4805,N_4886);
and U4942 (N_4942,N_4890,N_4851);
and U4943 (N_4943,N_4800,N_4837);
nand U4944 (N_4944,N_4807,N_4855);
nand U4945 (N_4945,N_4874,N_4806);
or U4946 (N_4946,N_4898,N_4878);
nand U4947 (N_4947,N_4899,N_4870);
nor U4948 (N_4948,N_4876,N_4811);
and U4949 (N_4949,N_4833,N_4847);
nor U4950 (N_4950,N_4872,N_4843);
or U4951 (N_4951,N_4892,N_4887);
nor U4952 (N_4952,N_4897,N_4805);
or U4953 (N_4953,N_4840,N_4852);
or U4954 (N_4954,N_4800,N_4818);
and U4955 (N_4955,N_4823,N_4804);
or U4956 (N_4956,N_4899,N_4821);
and U4957 (N_4957,N_4829,N_4844);
and U4958 (N_4958,N_4891,N_4845);
nor U4959 (N_4959,N_4855,N_4888);
nor U4960 (N_4960,N_4839,N_4880);
nand U4961 (N_4961,N_4868,N_4848);
or U4962 (N_4962,N_4804,N_4880);
and U4963 (N_4963,N_4855,N_4872);
or U4964 (N_4964,N_4827,N_4825);
nor U4965 (N_4965,N_4838,N_4890);
nor U4966 (N_4966,N_4824,N_4800);
and U4967 (N_4967,N_4879,N_4881);
or U4968 (N_4968,N_4826,N_4883);
nor U4969 (N_4969,N_4836,N_4809);
nor U4970 (N_4970,N_4807,N_4880);
and U4971 (N_4971,N_4845,N_4813);
and U4972 (N_4972,N_4879,N_4849);
nor U4973 (N_4973,N_4899,N_4887);
and U4974 (N_4974,N_4892,N_4881);
or U4975 (N_4975,N_4818,N_4881);
nand U4976 (N_4976,N_4811,N_4837);
or U4977 (N_4977,N_4898,N_4804);
xor U4978 (N_4978,N_4872,N_4875);
and U4979 (N_4979,N_4822,N_4838);
or U4980 (N_4980,N_4869,N_4870);
or U4981 (N_4981,N_4837,N_4832);
nand U4982 (N_4982,N_4857,N_4819);
or U4983 (N_4983,N_4820,N_4893);
xor U4984 (N_4984,N_4884,N_4873);
nor U4985 (N_4985,N_4802,N_4878);
and U4986 (N_4986,N_4883,N_4838);
nand U4987 (N_4987,N_4880,N_4895);
nand U4988 (N_4988,N_4812,N_4821);
nor U4989 (N_4989,N_4860,N_4895);
xor U4990 (N_4990,N_4859,N_4855);
or U4991 (N_4991,N_4847,N_4880);
nand U4992 (N_4992,N_4869,N_4856);
nor U4993 (N_4993,N_4848,N_4802);
nand U4994 (N_4994,N_4890,N_4868);
xor U4995 (N_4995,N_4858,N_4875);
xnor U4996 (N_4996,N_4801,N_4866);
nor U4997 (N_4997,N_4887,N_4894);
or U4998 (N_4998,N_4886,N_4884);
and U4999 (N_4999,N_4883,N_4802);
nor UO_0 (O_0,N_4949,N_4921);
nor UO_1 (O_1,N_4999,N_4908);
and UO_2 (O_2,N_4922,N_4986);
or UO_3 (O_3,N_4974,N_4948);
nand UO_4 (O_4,N_4951,N_4987);
and UO_5 (O_5,N_4932,N_4997);
nand UO_6 (O_6,N_4919,N_4998);
and UO_7 (O_7,N_4980,N_4952);
and UO_8 (O_8,N_4916,N_4931);
nor UO_9 (O_9,N_4903,N_4970);
and UO_10 (O_10,N_4992,N_4902);
xor UO_11 (O_11,N_4937,N_4901);
and UO_12 (O_12,N_4979,N_4946);
and UO_13 (O_13,N_4945,N_4959);
nand UO_14 (O_14,N_4944,N_4984);
and UO_15 (O_15,N_4918,N_4973);
and UO_16 (O_16,N_4964,N_4925);
nand UO_17 (O_17,N_4912,N_4909);
nand UO_18 (O_18,N_4954,N_4996);
and UO_19 (O_19,N_4960,N_4978);
or UO_20 (O_20,N_4920,N_4928);
or UO_21 (O_21,N_4989,N_4965);
or UO_22 (O_22,N_4913,N_4933);
xor UO_23 (O_23,N_4968,N_4915);
xnor UO_24 (O_24,N_4962,N_4956);
nand UO_25 (O_25,N_4907,N_4966);
or UO_26 (O_26,N_4938,N_4977);
nand UO_27 (O_27,N_4953,N_4982);
nor UO_28 (O_28,N_4900,N_4994);
nand UO_29 (O_29,N_4905,N_4957);
nand UO_30 (O_30,N_4929,N_4939);
nor UO_31 (O_31,N_4969,N_4975);
nand UO_32 (O_32,N_4940,N_4950);
or UO_33 (O_33,N_4917,N_4963);
xnor UO_34 (O_34,N_4967,N_4930);
nor UO_35 (O_35,N_4910,N_4935);
nor UO_36 (O_36,N_4983,N_4942);
xor UO_37 (O_37,N_4926,N_4961);
nand UO_38 (O_38,N_4971,N_4941);
and UO_39 (O_39,N_4972,N_4985);
nand UO_40 (O_40,N_4927,N_4988);
and UO_41 (O_41,N_4943,N_4991);
xor UO_42 (O_42,N_4904,N_4981);
nor UO_43 (O_43,N_4936,N_4955);
nand UO_44 (O_44,N_4906,N_4923);
nor UO_45 (O_45,N_4958,N_4947);
xnor UO_46 (O_46,N_4976,N_4934);
and UO_47 (O_47,N_4990,N_4914);
or UO_48 (O_48,N_4995,N_4924);
or UO_49 (O_49,N_4993,N_4911);
xor UO_50 (O_50,N_4950,N_4916);
or UO_51 (O_51,N_4990,N_4906);
nor UO_52 (O_52,N_4968,N_4922);
nor UO_53 (O_53,N_4980,N_4956);
nor UO_54 (O_54,N_4957,N_4996);
nand UO_55 (O_55,N_4991,N_4918);
and UO_56 (O_56,N_4983,N_4931);
or UO_57 (O_57,N_4983,N_4978);
xnor UO_58 (O_58,N_4936,N_4942);
and UO_59 (O_59,N_4921,N_4905);
or UO_60 (O_60,N_4954,N_4915);
and UO_61 (O_61,N_4971,N_4911);
or UO_62 (O_62,N_4991,N_4972);
and UO_63 (O_63,N_4944,N_4938);
nand UO_64 (O_64,N_4902,N_4943);
nand UO_65 (O_65,N_4905,N_4968);
and UO_66 (O_66,N_4921,N_4935);
and UO_67 (O_67,N_4917,N_4927);
nor UO_68 (O_68,N_4992,N_4940);
xnor UO_69 (O_69,N_4986,N_4997);
nor UO_70 (O_70,N_4913,N_4917);
nand UO_71 (O_71,N_4931,N_4960);
nand UO_72 (O_72,N_4989,N_4960);
nor UO_73 (O_73,N_4908,N_4929);
and UO_74 (O_74,N_4997,N_4925);
nor UO_75 (O_75,N_4940,N_4901);
and UO_76 (O_76,N_4917,N_4971);
nand UO_77 (O_77,N_4966,N_4927);
xor UO_78 (O_78,N_4912,N_4991);
or UO_79 (O_79,N_4934,N_4974);
nand UO_80 (O_80,N_4989,N_4994);
nand UO_81 (O_81,N_4946,N_4981);
xor UO_82 (O_82,N_4978,N_4958);
and UO_83 (O_83,N_4945,N_4949);
xor UO_84 (O_84,N_4915,N_4982);
or UO_85 (O_85,N_4916,N_4979);
and UO_86 (O_86,N_4995,N_4949);
and UO_87 (O_87,N_4931,N_4988);
and UO_88 (O_88,N_4958,N_4935);
nand UO_89 (O_89,N_4998,N_4935);
nand UO_90 (O_90,N_4978,N_4921);
or UO_91 (O_91,N_4981,N_4951);
nand UO_92 (O_92,N_4955,N_4902);
or UO_93 (O_93,N_4989,N_4986);
nand UO_94 (O_94,N_4927,N_4964);
xnor UO_95 (O_95,N_4989,N_4966);
nand UO_96 (O_96,N_4911,N_4999);
xor UO_97 (O_97,N_4958,N_4999);
nor UO_98 (O_98,N_4995,N_4978);
nor UO_99 (O_99,N_4988,N_4951);
nand UO_100 (O_100,N_4921,N_4924);
and UO_101 (O_101,N_4932,N_4978);
or UO_102 (O_102,N_4987,N_4926);
nand UO_103 (O_103,N_4974,N_4989);
or UO_104 (O_104,N_4945,N_4942);
or UO_105 (O_105,N_4948,N_4962);
xor UO_106 (O_106,N_4968,N_4985);
nor UO_107 (O_107,N_4937,N_4982);
nand UO_108 (O_108,N_4981,N_4977);
and UO_109 (O_109,N_4932,N_4902);
xor UO_110 (O_110,N_4916,N_4963);
or UO_111 (O_111,N_4965,N_4910);
nor UO_112 (O_112,N_4903,N_4949);
and UO_113 (O_113,N_4939,N_4966);
nand UO_114 (O_114,N_4977,N_4944);
nor UO_115 (O_115,N_4939,N_4920);
and UO_116 (O_116,N_4936,N_4932);
or UO_117 (O_117,N_4999,N_4905);
nand UO_118 (O_118,N_4932,N_4907);
or UO_119 (O_119,N_4992,N_4955);
or UO_120 (O_120,N_4982,N_4906);
nor UO_121 (O_121,N_4907,N_4908);
or UO_122 (O_122,N_4970,N_4907);
and UO_123 (O_123,N_4994,N_4905);
and UO_124 (O_124,N_4903,N_4930);
and UO_125 (O_125,N_4930,N_4957);
or UO_126 (O_126,N_4917,N_4976);
and UO_127 (O_127,N_4913,N_4957);
and UO_128 (O_128,N_4902,N_4907);
or UO_129 (O_129,N_4902,N_4979);
nand UO_130 (O_130,N_4973,N_4946);
or UO_131 (O_131,N_4987,N_4937);
or UO_132 (O_132,N_4920,N_4934);
nor UO_133 (O_133,N_4967,N_4924);
nand UO_134 (O_134,N_4910,N_4980);
nand UO_135 (O_135,N_4938,N_4965);
xnor UO_136 (O_136,N_4930,N_4929);
and UO_137 (O_137,N_4905,N_4961);
xnor UO_138 (O_138,N_4917,N_4978);
xnor UO_139 (O_139,N_4940,N_4911);
nand UO_140 (O_140,N_4932,N_4985);
nor UO_141 (O_141,N_4952,N_4974);
and UO_142 (O_142,N_4918,N_4999);
and UO_143 (O_143,N_4981,N_4901);
and UO_144 (O_144,N_4920,N_4987);
nand UO_145 (O_145,N_4924,N_4952);
and UO_146 (O_146,N_4946,N_4971);
nand UO_147 (O_147,N_4952,N_4910);
xnor UO_148 (O_148,N_4990,N_4989);
nand UO_149 (O_149,N_4950,N_4926);
and UO_150 (O_150,N_4928,N_4971);
nor UO_151 (O_151,N_4920,N_4990);
nor UO_152 (O_152,N_4940,N_4965);
or UO_153 (O_153,N_4968,N_4952);
or UO_154 (O_154,N_4945,N_4999);
nor UO_155 (O_155,N_4965,N_4987);
xnor UO_156 (O_156,N_4937,N_4936);
and UO_157 (O_157,N_4958,N_4970);
xnor UO_158 (O_158,N_4978,N_4940);
or UO_159 (O_159,N_4980,N_4977);
xnor UO_160 (O_160,N_4947,N_4911);
nand UO_161 (O_161,N_4966,N_4964);
or UO_162 (O_162,N_4920,N_4926);
or UO_163 (O_163,N_4994,N_4933);
nand UO_164 (O_164,N_4982,N_4920);
and UO_165 (O_165,N_4936,N_4988);
nand UO_166 (O_166,N_4958,N_4952);
nor UO_167 (O_167,N_4908,N_4934);
nand UO_168 (O_168,N_4909,N_4946);
nor UO_169 (O_169,N_4936,N_4974);
and UO_170 (O_170,N_4902,N_4903);
and UO_171 (O_171,N_4947,N_4909);
or UO_172 (O_172,N_4990,N_4996);
nor UO_173 (O_173,N_4933,N_4904);
or UO_174 (O_174,N_4986,N_4902);
xor UO_175 (O_175,N_4926,N_4948);
nor UO_176 (O_176,N_4936,N_4957);
or UO_177 (O_177,N_4975,N_4944);
nor UO_178 (O_178,N_4903,N_4978);
nor UO_179 (O_179,N_4960,N_4986);
or UO_180 (O_180,N_4917,N_4995);
xor UO_181 (O_181,N_4918,N_4972);
or UO_182 (O_182,N_4969,N_4995);
and UO_183 (O_183,N_4963,N_4966);
nand UO_184 (O_184,N_4957,N_4993);
nand UO_185 (O_185,N_4944,N_4990);
and UO_186 (O_186,N_4907,N_4929);
nand UO_187 (O_187,N_4992,N_4982);
and UO_188 (O_188,N_4951,N_4964);
nor UO_189 (O_189,N_4943,N_4981);
nor UO_190 (O_190,N_4995,N_4954);
and UO_191 (O_191,N_4950,N_4921);
nor UO_192 (O_192,N_4978,N_4992);
nor UO_193 (O_193,N_4953,N_4962);
nand UO_194 (O_194,N_4932,N_4905);
and UO_195 (O_195,N_4945,N_4975);
xnor UO_196 (O_196,N_4955,N_4944);
and UO_197 (O_197,N_4921,N_4934);
nand UO_198 (O_198,N_4989,N_4991);
and UO_199 (O_199,N_4900,N_4948);
nand UO_200 (O_200,N_4938,N_4919);
and UO_201 (O_201,N_4960,N_4952);
and UO_202 (O_202,N_4907,N_4977);
or UO_203 (O_203,N_4997,N_4965);
and UO_204 (O_204,N_4954,N_4975);
nand UO_205 (O_205,N_4921,N_4969);
and UO_206 (O_206,N_4991,N_4909);
and UO_207 (O_207,N_4943,N_4951);
nor UO_208 (O_208,N_4917,N_4932);
or UO_209 (O_209,N_4991,N_4930);
xor UO_210 (O_210,N_4991,N_4920);
and UO_211 (O_211,N_4970,N_4998);
and UO_212 (O_212,N_4965,N_4998);
nor UO_213 (O_213,N_4956,N_4986);
and UO_214 (O_214,N_4932,N_4956);
nand UO_215 (O_215,N_4944,N_4925);
nor UO_216 (O_216,N_4939,N_4914);
or UO_217 (O_217,N_4997,N_4991);
xnor UO_218 (O_218,N_4901,N_4991);
nor UO_219 (O_219,N_4910,N_4973);
nand UO_220 (O_220,N_4969,N_4973);
and UO_221 (O_221,N_4900,N_4923);
nand UO_222 (O_222,N_4941,N_4909);
nor UO_223 (O_223,N_4904,N_4929);
or UO_224 (O_224,N_4958,N_4949);
and UO_225 (O_225,N_4914,N_4983);
nand UO_226 (O_226,N_4966,N_4957);
and UO_227 (O_227,N_4998,N_4911);
or UO_228 (O_228,N_4924,N_4908);
xnor UO_229 (O_229,N_4931,N_4990);
and UO_230 (O_230,N_4970,N_4964);
nor UO_231 (O_231,N_4967,N_4921);
nor UO_232 (O_232,N_4971,N_4951);
nand UO_233 (O_233,N_4991,N_4980);
nand UO_234 (O_234,N_4913,N_4974);
or UO_235 (O_235,N_4987,N_4912);
or UO_236 (O_236,N_4904,N_4922);
nand UO_237 (O_237,N_4926,N_4994);
and UO_238 (O_238,N_4977,N_4900);
and UO_239 (O_239,N_4921,N_4960);
nand UO_240 (O_240,N_4978,N_4913);
nor UO_241 (O_241,N_4931,N_4918);
and UO_242 (O_242,N_4910,N_4964);
nand UO_243 (O_243,N_4939,N_4988);
xor UO_244 (O_244,N_4902,N_4981);
or UO_245 (O_245,N_4912,N_4928);
nand UO_246 (O_246,N_4959,N_4991);
or UO_247 (O_247,N_4952,N_4932);
or UO_248 (O_248,N_4960,N_4932);
and UO_249 (O_249,N_4916,N_4947);
nand UO_250 (O_250,N_4944,N_4991);
nand UO_251 (O_251,N_4959,N_4982);
nand UO_252 (O_252,N_4954,N_4985);
xor UO_253 (O_253,N_4903,N_4974);
and UO_254 (O_254,N_4988,N_4949);
nand UO_255 (O_255,N_4908,N_4987);
nand UO_256 (O_256,N_4986,N_4971);
nand UO_257 (O_257,N_4969,N_4908);
nand UO_258 (O_258,N_4938,N_4909);
or UO_259 (O_259,N_4902,N_4952);
nand UO_260 (O_260,N_4940,N_4903);
or UO_261 (O_261,N_4967,N_4977);
nor UO_262 (O_262,N_4954,N_4983);
nor UO_263 (O_263,N_4913,N_4967);
nand UO_264 (O_264,N_4994,N_4906);
or UO_265 (O_265,N_4965,N_4966);
and UO_266 (O_266,N_4932,N_4951);
nand UO_267 (O_267,N_4967,N_4966);
or UO_268 (O_268,N_4925,N_4927);
and UO_269 (O_269,N_4990,N_4987);
nor UO_270 (O_270,N_4930,N_4946);
and UO_271 (O_271,N_4906,N_4970);
xor UO_272 (O_272,N_4971,N_4907);
and UO_273 (O_273,N_4953,N_4911);
nand UO_274 (O_274,N_4983,N_4950);
nor UO_275 (O_275,N_4927,N_4907);
nand UO_276 (O_276,N_4914,N_4945);
nor UO_277 (O_277,N_4956,N_4928);
nand UO_278 (O_278,N_4971,N_4993);
or UO_279 (O_279,N_4915,N_4959);
or UO_280 (O_280,N_4951,N_4998);
nor UO_281 (O_281,N_4922,N_4930);
and UO_282 (O_282,N_4977,N_4973);
or UO_283 (O_283,N_4930,N_4976);
or UO_284 (O_284,N_4914,N_4994);
or UO_285 (O_285,N_4978,N_4996);
nand UO_286 (O_286,N_4991,N_4975);
or UO_287 (O_287,N_4991,N_4999);
xor UO_288 (O_288,N_4944,N_4989);
xnor UO_289 (O_289,N_4997,N_4982);
xnor UO_290 (O_290,N_4979,N_4994);
nor UO_291 (O_291,N_4986,N_4945);
nand UO_292 (O_292,N_4928,N_4968);
or UO_293 (O_293,N_4968,N_4974);
xnor UO_294 (O_294,N_4913,N_4901);
nor UO_295 (O_295,N_4936,N_4907);
or UO_296 (O_296,N_4986,N_4933);
nor UO_297 (O_297,N_4905,N_4960);
xor UO_298 (O_298,N_4906,N_4953);
xnor UO_299 (O_299,N_4997,N_4948);
or UO_300 (O_300,N_4960,N_4964);
nor UO_301 (O_301,N_4917,N_4962);
or UO_302 (O_302,N_4954,N_4994);
or UO_303 (O_303,N_4925,N_4957);
nand UO_304 (O_304,N_4966,N_4914);
or UO_305 (O_305,N_4950,N_4914);
and UO_306 (O_306,N_4954,N_4936);
nand UO_307 (O_307,N_4921,N_4997);
nand UO_308 (O_308,N_4983,N_4924);
nand UO_309 (O_309,N_4990,N_4921);
and UO_310 (O_310,N_4956,N_4983);
nor UO_311 (O_311,N_4901,N_4920);
and UO_312 (O_312,N_4995,N_4901);
or UO_313 (O_313,N_4915,N_4952);
nand UO_314 (O_314,N_4956,N_4997);
and UO_315 (O_315,N_4973,N_4989);
or UO_316 (O_316,N_4979,N_4993);
and UO_317 (O_317,N_4940,N_4922);
nor UO_318 (O_318,N_4941,N_4925);
nor UO_319 (O_319,N_4976,N_4963);
and UO_320 (O_320,N_4922,N_4915);
and UO_321 (O_321,N_4967,N_4952);
or UO_322 (O_322,N_4970,N_4928);
nor UO_323 (O_323,N_4956,N_4954);
and UO_324 (O_324,N_4958,N_4957);
or UO_325 (O_325,N_4937,N_4991);
or UO_326 (O_326,N_4961,N_4958);
and UO_327 (O_327,N_4906,N_4940);
or UO_328 (O_328,N_4977,N_4984);
nand UO_329 (O_329,N_4915,N_4984);
and UO_330 (O_330,N_4985,N_4940);
nand UO_331 (O_331,N_4949,N_4904);
nand UO_332 (O_332,N_4999,N_4929);
and UO_333 (O_333,N_4970,N_4995);
nor UO_334 (O_334,N_4934,N_4942);
and UO_335 (O_335,N_4970,N_4901);
or UO_336 (O_336,N_4910,N_4909);
and UO_337 (O_337,N_4982,N_4964);
and UO_338 (O_338,N_4994,N_4998);
nor UO_339 (O_339,N_4975,N_4965);
nor UO_340 (O_340,N_4938,N_4990);
and UO_341 (O_341,N_4923,N_4974);
or UO_342 (O_342,N_4908,N_4973);
or UO_343 (O_343,N_4987,N_4911);
nand UO_344 (O_344,N_4955,N_4915);
nand UO_345 (O_345,N_4905,N_4900);
nand UO_346 (O_346,N_4954,N_4969);
nor UO_347 (O_347,N_4917,N_4970);
nand UO_348 (O_348,N_4920,N_4993);
nand UO_349 (O_349,N_4914,N_4927);
xnor UO_350 (O_350,N_4931,N_4933);
nand UO_351 (O_351,N_4988,N_4905);
and UO_352 (O_352,N_4929,N_4962);
nand UO_353 (O_353,N_4919,N_4924);
and UO_354 (O_354,N_4914,N_4985);
and UO_355 (O_355,N_4974,N_4977);
nand UO_356 (O_356,N_4950,N_4978);
xor UO_357 (O_357,N_4984,N_4992);
or UO_358 (O_358,N_4979,N_4907);
or UO_359 (O_359,N_4918,N_4988);
and UO_360 (O_360,N_4941,N_4979);
nand UO_361 (O_361,N_4952,N_4981);
or UO_362 (O_362,N_4938,N_4951);
or UO_363 (O_363,N_4972,N_4905);
or UO_364 (O_364,N_4959,N_4951);
nor UO_365 (O_365,N_4957,N_4998);
nor UO_366 (O_366,N_4909,N_4982);
or UO_367 (O_367,N_4982,N_4948);
nand UO_368 (O_368,N_4941,N_4973);
and UO_369 (O_369,N_4947,N_4932);
nand UO_370 (O_370,N_4976,N_4919);
or UO_371 (O_371,N_4916,N_4921);
nand UO_372 (O_372,N_4988,N_4975);
nor UO_373 (O_373,N_4925,N_4918);
and UO_374 (O_374,N_4987,N_4962);
and UO_375 (O_375,N_4935,N_4991);
nand UO_376 (O_376,N_4988,N_4979);
or UO_377 (O_377,N_4936,N_4903);
xor UO_378 (O_378,N_4904,N_4966);
nor UO_379 (O_379,N_4982,N_4967);
and UO_380 (O_380,N_4974,N_4910);
nor UO_381 (O_381,N_4923,N_4962);
nor UO_382 (O_382,N_4949,N_4913);
nand UO_383 (O_383,N_4924,N_4904);
nand UO_384 (O_384,N_4984,N_4912);
and UO_385 (O_385,N_4972,N_4927);
and UO_386 (O_386,N_4967,N_4915);
nor UO_387 (O_387,N_4957,N_4978);
or UO_388 (O_388,N_4921,N_4957);
nand UO_389 (O_389,N_4993,N_4978);
nand UO_390 (O_390,N_4960,N_4997);
xor UO_391 (O_391,N_4902,N_4954);
and UO_392 (O_392,N_4986,N_4953);
nor UO_393 (O_393,N_4948,N_4999);
or UO_394 (O_394,N_4914,N_4921);
and UO_395 (O_395,N_4994,N_4907);
nand UO_396 (O_396,N_4915,N_4934);
and UO_397 (O_397,N_4980,N_4967);
or UO_398 (O_398,N_4901,N_4974);
and UO_399 (O_399,N_4999,N_4931);
and UO_400 (O_400,N_4910,N_4900);
nand UO_401 (O_401,N_4986,N_4972);
xor UO_402 (O_402,N_4999,N_4967);
nand UO_403 (O_403,N_4924,N_4953);
nand UO_404 (O_404,N_4981,N_4989);
or UO_405 (O_405,N_4902,N_4926);
nand UO_406 (O_406,N_4961,N_4988);
and UO_407 (O_407,N_4972,N_4964);
and UO_408 (O_408,N_4967,N_4974);
nor UO_409 (O_409,N_4979,N_4923);
nand UO_410 (O_410,N_4933,N_4992);
nor UO_411 (O_411,N_4912,N_4926);
and UO_412 (O_412,N_4940,N_4983);
and UO_413 (O_413,N_4987,N_4963);
nand UO_414 (O_414,N_4906,N_4938);
nand UO_415 (O_415,N_4997,N_4971);
or UO_416 (O_416,N_4993,N_4940);
and UO_417 (O_417,N_4917,N_4942);
or UO_418 (O_418,N_4905,N_4987);
and UO_419 (O_419,N_4979,N_4915);
nand UO_420 (O_420,N_4937,N_4961);
or UO_421 (O_421,N_4904,N_4956);
or UO_422 (O_422,N_4956,N_4990);
or UO_423 (O_423,N_4975,N_4959);
or UO_424 (O_424,N_4986,N_4961);
nand UO_425 (O_425,N_4977,N_4958);
or UO_426 (O_426,N_4953,N_4978);
or UO_427 (O_427,N_4914,N_4984);
nand UO_428 (O_428,N_4943,N_4950);
nor UO_429 (O_429,N_4997,N_4917);
nand UO_430 (O_430,N_4904,N_4911);
or UO_431 (O_431,N_4985,N_4943);
or UO_432 (O_432,N_4973,N_4988);
nand UO_433 (O_433,N_4934,N_4929);
or UO_434 (O_434,N_4909,N_4970);
nor UO_435 (O_435,N_4922,N_4972);
or UO_436 (O_436,N_4949,N_4973);
nand UO_437 (O_437,N_4972,N_4957);
and UO_438 (O_438,N_4998,N_4968);
and UO_439 (O_439,N_4936,N_4951);
nor UO_440 (O_440,N_4915,N_4932);
or UO_441 (O_441,N_4969,N_4906);
nor UO_442 (O_442,N_4961,N_4998);
or UO_443 (O_443,N_4920,N_4974);
and UO_444 (O_444,N_4954,N_4931);
nor UO_445 (O_445,N_4992,N_4939);
and UO_446 (O_446,N_4989,N_4977);
and UO_447 (O_447,N_4924,N_4925);
nand UO_448 (O_448,N_4926,N_4976);
nor UO_449 (O_449,N_4929,N_4991);
or UO_450 (O_450,N_4972,N_4989);
and UO_451 (O_451,N_4940,N_4989);
and UO_452 (O_452,N_4961,N_4973);
nand UO_453 (O_453,N_4991,N_4953);
nor UO_454 (O_454,N_4914,N_4962);
and UO_455 (O_455,N_4985,N_4952);
or UO_456 (O_456,N_4936,N_4983);
nor UO_457 (O_457,N_4922,N_4931);
nor UO_458 (O_458,N_4999,N_4976);
or UO_459 (O_459,N_4954,N_4908);
and UO_460 (O_460,N_4961,N_4914);
or UO_461 (O_461,N_4967,N_4995);
and UO_462 (O_462,N_4925,N_4935);
or UO_463 (O_463,N_4976,N_4940);
or UO_464 (O_464,N_4953,N_4976);
nor UO_465 (O_465,N_4961,N_4936);
and UO_466 (O_466,N_4963,N_4955);
and UO_467 (O_467,N_4927,N_4908);
xor UO_468 (O_468,N_4952,N_4918);
nand UO_469 (O_469,N_4965,N_4918);
nand UO_470 (O_470,N_4957,N_4953);
or UO_471 (O_471,N_4959,N_4981);
nand UO_472 (O_472,N_4908,N_4965);
nor UO_473 (O_473,N_4982,N_4979);
and UO_474 (O_474,N_4939,N_4905);
or UO_475 (O_475,N_4977,N_4912);
nor UO_476 (O_476,N_4986,N_4913);
xor UO_477 (O_477,N_4942,N_4991);
nand UO_478 (O_478,N_4987,N_4931);
and UO_479 (O_479,N_4973,N_4975);
nand UO_480 (O_480,N_4940,N_4918);
and UO_481 (O_481,N_4924,N_4911);
and UO_482 (O_482,N_4985,N_4996);
and UO_483 (O_483,N_4975,N_4998);
and UO_484 (O_484,N_4956,N_4940);
nor UO_485 (O_485,N_4940,N_4904);
and UO_486 (O_486,N_4962,N_4978);
nand UO_487 (O_487,N_4994,N_4921);
and UO_488 (O_488,N_4973,N_4954);
and UO_489 (O_489,N_4996,N_4992);
and UO_490 (O_490,N_4900,N_4930);
or UO_491 (O_491,N_4946,N_4964);
or UO_492 (O_492,N_4983,N_4959);
and UO_493 (O_493,N_4942,N_4973);
xor UO_494 (O_494,N_4907,N_4974);
or UO_495 (O_495,N_4986,N_4959);
or UO_496 (O_496,N_4902,N_4939);
nand UO_497 (O_497,N_4902,N_4941);
and UO_498 (O_498,N_4965,N_4957);
or UO_499 (O_499,N_4946,N_4966);
or UO_500 (O_500,N_4909,N_4927);
nand UO_501 (O_501,N_4953,N_4983);
nand UO_502 (O_502,N_4921,N_4920);
nor UO_503 (O_503,N_4983,N_4969);
nor UO_504 (O_504,N_4916,N_4996);
xor UO_505 (O_505,N_4906,N_4936);
and UO_506 (O_506,N_4915,N_4937);
and UO_507 (O_507,N_4914,N_4919);
nand UO_508 (O_508,N_4951,N_4975);
nor UO_509 (O_509,N_4990,N_4952);
xor UO_510 (O_510,N_4923,N_4995);
nor UO_511 (O_511,N_4947,N_4997);
and UO_512 (O_512,N_4918,N_4979);
and UO_513 (O_513,N_4928,N_4931);
or UO_514 (O_514,N_4933,N_4948);
and UO_515 (O_515,N_4969,N_4997);
and UO_516 (O_516,N_4963,N_4901);
nand UO_517 (O_517,N_4968,N_4900);
nor UO_518 (O_518,N_4928,N_4906);
and UO_519 (O_519,N_4923,N_4935);
nor UO_520 (O_520,N_4949,N_4908);
nand UO_521 (O_521,N_4929,N_4968);
nor UO_522 (O_522,N_4924,N_4990);
and UO_523 (O_523,N_4959,N_4968);
nand UO_524 (O_524,N_4947,N_4936);
xor UO_525 (O_525,N_4958,N_4912);
nor UO_526 (O_526,N_4925,N_4949);
nor UO_527 (O_527,N_4952,N_4959);
and UO_528 (O_528,N_4901,N_4928);
xnor UO_529 (O_529,N_4937,N_4902);
or UO_530 (O_530,N_4924,N_4970);
xor UO_531 (O_531,N_4925,N_4904);
xor UO_532 (O_532,N_4956,N_4900);
nor UO_533 (O_533,N_4989,N_4992);
or UO_534 (O_534,N_4949,N_4922);
and UO_535 (O_535,N_4979,N_4909);
nand UO_536 (O_536,N_4919,N_4920);
and UO_537 (O_537,N_4925,N_4929);
nand UO_538 (O_538,N_4968,N_4934);
nand UO_539 (O_539,N_4964,N_4930);
nand UO_540 (O_540,N_4988,N_4953);
and UO_541 (O_541,N_4998,N_4962);
nor UO_542 (O_542,N_4971,N_4961);
nor UO_543 (O_543,N_4908,N_4967);
xor UO_544 (O_544,N_4939,N_4911);
nand UO_545 (O_545,N_4910,N_4985);
or UO_546 (O_546,N_4947,N_4901);
or UO_547 (O_547,N_4933,N_4921);
xor UO_548 (O_548,N_4976,N_4929);
or UO_549 (O_549,N_4909,N_4996);
xnor UO_550 (O_550,N_4983,N_4937);
nand UO_551 (O_551,N_4967,N_4996);
or UO_552 (O_552,N_4917,N_4969);
and UO_553 (O_553,N_4996,N_4936);
and UO_554 (O_554,N_4930,N_4960);
nand UO_555 (O_555,N_4993,N_4958);
or UO_556 (O_556,N_4934,N_4949);
nand UO_557 (O_557,N_4998,N_4902);
and UO_558 (O_558,N_4922,N_4943);
and UO_559 (O_559,N_4953,N_4920);
and UO_560 (O_560,N_4998,N_4926);
and UO_561 (O_561,N_4988,N_4921);
nor UO_562 (O_562,N_4938,N_4950);
or UO_563 (O_563,N_4957,N_4970);
xnor UO_564 (O_564,N_4963,N_4946);
nor UO_565 (O_565,N_4902,N_4904);
nand UO_566 (O_566,N_4913,N_4982);
or UO_567 (O_567,N_4980,N_4966);
or UO_568 (O_568,N_4946,N_4931);
nor UO_569 (O_569,N_4988,N_4944);
or UO_570 (O_570,N_4983,N_4938);
and UO_571 (O_571,N_4988,N_4903);
or UO_572 (O_572,N_4970,N_4905);
and UO_573 (O_573,N_4978,N_4966);
and UO_574 (O_574,N_4969,N_4904);
and UO_575 (O_575,N_4924,N_4955);
nor UO_576 (O_576,N_4915,N_4910);
or UO_577 (O_577,N_4934,N_4905);
nand UO_578 (O_578,N_4941,N_4953);
and UO_579 (O_579,N_4944,N_4924);
nand UO_580 (O_580,N_4968,N_4924);
nand UO_581 (O_581,N_4974,N_4998);
nand UO_582 (O_582,N_4964,N_4948);
nor UO_583 (O_583,N_4929,N_4900);
xnor UO_584 (O_584,N_4994,N_4910);
or UO_585 (O_585,N_4996,N_4922);
or UO_586 (O_586,N_4912,N_4998);
xnor UO_587 (O_587,N_4928,N_4967);
nand UO_588 (O_588,N_4983,N_4962);
or UO_589 (O_589,N_4987,N_4993);
xor UO_590 (O_590,N_4928,N_4926);
or UO_591 (O_591,N_4994,N_4993);
and UO_592 (O_592,N_4977,N_4965);
xor UO_593 (O_593,N_4964,N_4978);
nand UO_594 (O_594,N_4962,N_4974);
or UO_595 (O_595,N_4932,N_4971);
or UO_596 (O_596,N_4910,N_4954);
nor UO_597 (O_597,N_4932,N_4940);
nor UO_598 (O_598,N_4950,N_4927);
and UO_599 (O_599,N_4981,N_4975);
xnor UO_600 (O_600,N_4937,N_4957);
nor UO_601 (O_601,N_4952,N_4939);
nor UO_602 (O_602,N_4919,N_4971);
or UO_603 (O_603,N_4936,N_4943);
and UO_604 (O_604,N_4976,N_4913);
and UO_605 (O_605,N_4962,N_4922);
nor UO_606 (O_606,N_4970,N_4942);
and UO_607 (O_607,N_4999,N_4951);
xnor UO_608 (O_608,N_4959,N_4988);
or UO_609 (O_609,N_4993,N_4966);
and UO_610 (O_610,N_4926,N_4967);
nand UO_611 (O_611,N_4996,N_4938);
nor UO_612 (O_612,N_4958,N_4910);
xor UO_613 (O_613,N_4964,N_4900);
and UO_614 (O_614,N_4913,N_4919);
xnor UO_615 (O_615,N_4997,N_4909);
and UO_616 (O_616,N_4934,N_4927);
xor UO_617 (O_617,N_4994,N_4968);
nand UO_618 (O_618,N_4982,N_4923);
or UO_619 (O_619,N_4953,N_4948);
nand UO_620 (O_620,N_4922,N_4906);
or UO_621 (O_621,N_4930,N_4970);
and UO_622 (O_622,N_4959,N_4908);
xor UO_623 (O_623,N_4945,N_4912);
nand UO_624 (O_624,N_4994,N_4986);
or UO_625 (O_625,N_4941,N_4927);
nand UO_626 (O_626,N_4999,N_4944);
nor UO_627 (O_627,N_4909,N_4928);
nand UO_628 (O_628,N_4959,N_4974);
nand UO_629 (O_629,N_4903,N_4914);
and UO_630 (O_630,N_4960,N_4935);
or UO_631 (O_631,N_4917,N_4959);
nor UO_632 (O_632,N_4910,N_4922);
nand UO_633 (O_633,N_4960,N_4991);
nor UO_634 (O_634,N_4990,N_4979);
nand UO_635 (O_635,N_4922,N_4947);
or UO_636 (O_636,N_4937,N_4913);
nor UO_637 (O_637,N_4994,N_4960);
and UO_638 (O_638,N_4976,N_4949);
or UO_639 (O_639,N_4920,N_4922);
nor UO_640 (O_640,N_4986,N_4985);
nand UO_641 (O_641,N_4929,N_4903);
or UO_642 (O_642,N_4912,N_4917);
and UO_643 (O_643,N_4971,N_4914);
or UO_644 (O_644,N_4917,N_4982);
xnor UO_645 (O_645,N_4962,N_4944);
nand UO_646 (O_646,N_4987,N_4955);
or UO_647 (O_647,N_4947,N_4923);
and UO_648 (O_648,N_4973,N_4900);
nand UO_649 (O_649,N_4936,N_4976);
nand UO_650 (O_650,N_4947,N_4946);
or UO_651 (O_651,N_4985,N_4911);
and UO_652 (O_652,N_4929,N_4983);
and UO_653 (O_653,N_4938,N_4947);
or UO_654 (O_654,N_4932,N_4974);
nor UO_655 (O_655,N_4972,N_4909);
nand UO_656 (O_656,N_4915,N_4935);
and UO_657 (O_657,N_4961,N_4942);
nor UO_658 (O_658,N_4972,N_4952);
and UO_659 (O_659,N_4905,N_4912);
nor UO_660 (O_660,N_4983,N_4976);
nor UO_661 (O_661,N_4973,N_4980);
or UO_662 (O_662,N_4920,N_4924);
nor UO_663 (O_663,N_4982,N_4965);
and UO_664 (O_664,N_4901,N_4943);
or UO_665 (O_665,N_4975,N_4994);
and UO_666 (O_666,N_4943,N_4973);
nand UO_667 (O_667,N_4917,N_4949);
or UO_668 (O_668,N_4964,N_4954);
or UO_669 (O_669,N_4973,N_4922);
and UO_670 (O_670,N_4962,N_4908);
xnor UO_671 (O_671,N_4928,N_4939);
nand UO_672 (O_672,N_4906,N_4911);
nor UO_673 (O_673,N_4960,N_4965);
or UO_674 (O_674,N_4958,N_4941);
or UO_675 (O_675,N_4978,N_4918);
nand UO_676 (O_676,N_4998,N_4922);
nand UO_677 (O_677,N_4917,N_4923);
nand UO_678 (O_678,N_4976,N_4906);
nor UO_679 (O_679,N_4966,N_4941);
xor UO_680 (O_680,N_4989,N_4980);
nor UO_681 (O_681,N_4938,N_4911);
or UO_682 (O_682,N_4986,N_4903);
and UO_683 (O_683,N_4925,N_4923);
nand UO_684 (O_684,N_4939,N_4916);
or UO_685 (O_685,N_4905,N_4949);
and UO_686 (O_686,N_4947,N_4955);
and UO_687 (O_687,N_4952,N_4971);
or UO_688 (O_688,N_4972,N_4931);
nand UO_689 (O_689,N_4999,N_4927);
nor UO_690 (O_690,N_4989,N_4933);
or UO_691 (O_691,N_4942,N_4943);
xnor UO_692 (O_692,N_4912,N_4981);
and UO_693 (O_693,N_4995,N_4994);
and UO_694 (O_694,N_4976,N_4959);
and UO_695 (O_695,N_4980,N_4927);
nand UO_696 (O_696,N_4965,N_4962);
nand UO_697 (O_697,N_4995,N_4900);
or UO_698 (O_698,N_4904,N_4978);
nand UO_699 (O_699,N_4985,N_4964);
nand UO_700 (O_700,N_4931,N_4989);
nor UO_701 (O_701,N_4985,N_4944);
nand UO_702 (O_702,N_4997,N_4979);
or UO_703 (O_703,N_4960,N_4920);
or UO_704 (O_704,N_4918,N_4976);
and UO_705 (O_705,N_4934,N_4999);
nor UO_706 (O_706,N_4966,N_4955);
nand UO_707 (O_707,N_4919,N_4961);
and UO_708 (O_708,N_4928,N_4951);
or UO_709 (O_709,N_4924,N_4909);
and UO_710 (O_710,N_4929,N_4961);
or UO_711 (O_711,N_4948,N_4994);
and UO_712 (O_712,N_4974,N_4975);
or UO_713 (O_713,N_4936,N_4952);
or UO_714 (O_714,N_4929,N_4994);
nand UO_715 (O_715,N_4968,N_4920);
nor UO_716 (O_716,N_4915,N_4993);
or UO_717 (O_717,N_4963,N_4981);
and UO_718 (O_718,N_4941,N_4906);
and UO_719 (O_719,N_4970,N_4967);
or UO_720 (O_720,N_4904,N_4916);
xor UO_721 (O_721,N_4933,N_4916);
or UO_722 (O_722,N_4989,N_4939);
nand UO_723 (O_723,N_4998,N_4979);
and UO_724 (O_724,N_4910,N_4942);
and UO_725 (O_725,N_4949,N_4932);
and UO_726 (O_726,N_4944,N_4958);
nand UO_727 (O_727,N_4937,N_4920);
and UO_728 (O_728,N_4952,N_4906);
nor UO_729 (O_729,N_4904,N_4991);
and UO_730 (O_730,N_4915,N_4942);
or UO_731 (O_731,N_4969,N_4914);
nand UO_732 (O_732,N_4929,N_4974);
nor UO_733 (O_733,N_4954,N_4945);
or UO_734 (O_734,N_4956,N_4957);
and UO_735 (O_735,N_4963,N_4998);
nor UO_736 (O_736,N_4968,N_4913);
and UO_737 (O_737,N_4943,N_4910);
or UO_738 (O_738,N_4956,N_4915);
nand UO_739 (O_739,N_4989,N_4952);
nor UO_740 (O_740,N_4949,N_4980);
xnor UO_741 (O_741,N_4921,N_4925);
nor UO_742 (O_742,N_4917,N_4964);
or UO_743 (O_743,N_4943,N_4982);
nor UO_744 (O_744,N_4977,N_4988);
nand UO_745 (O_745,N_4962,N_4976);
nand UO_746 (O_746,N_4985,N_4905);
and UO_747 (O_747,N_4904,N_4909);
or UO_748 (O_748,N_4976,N_4984);
nand UO_749 (O_749,N_4908,N_4942);
or UO_750 (O_750,N_4953,N_4918);
nand UO_751 (O_751,N_4915,N_4906);
or UO_752 (O_752,N_4930,N_4972);
nor UO_753 (O_753,N_4933,N_4957);
or UO_754 (O_754,N_4900,N_4921);
nand UO_755 (O_755,N_4945,N_4900);
or UO_756 (O_756,N_4950,N_4917);
xnor UO_757 (O_757,N_4926,N_4952);
nor UO_758 (O_758,N_4988,N_4964);
and UO_759 (O_759,N_4940,N_4949);
nand UO_760 (O_760,N_4991,N_4927);
and UO_761 (O_761,N_4946,N_4967);
nand UO_762 (O_762,N_4941,N_4931);
nand UO_763 (O_763,N_4990,N_4962);
nand UO_764 (O_764,N_4952,N_4982);
and UO_765 (O_765,N_4991,N_4957);
or UO_766 (O_766,N_4939,N_4938);
nor UO_767 (O_767,N_4990,N_4988);
nor UO_768 (O_768,N_4977,N_4978);
and UO_769 (O_769,N_4923,N_4944);
nor UO_770 (O_770,N_4991,N_4985);
nand UO_771 (O_771,N_4974,N_4995);
nand UO_772 (O_772,N_4905,N_4935);
or UO_773 (O_773,N_4989,N_4903);
nand UO_774 (O_774,N_4906,N_4920);
nor UO_775 (O_775,N_4963,N_4900);
or UO_776 (O_776,N_4976,N_4946);
or UO_777 (O_777,N_4956,N_4943);
or UO_778 (O_778,N_4972,N_4904);
and UO_779 (O_779,N_4980,N_4921);
nor UO_780 (O_780,N_4932,N_4967);
nor UO_781 (O_781,N_4949,N_4972);
and UO_782 (O_782,N_4973,N_4986);
xor UO_783 (O_783,N_4931,N_4934);
nand UO_784 (O_784,N_4970,N_4913);
and UO_785 (O_785,N_4945,N_4997);
and UO_786 (O_786,N_4994,N_4917);
nand UO_787 (O_787,N_4951,N_4907);
and UO_788 (O_788,N_4937,N_4934);
and UO_789 (O_789,N_4953,N_4997);
or UO_790 (O_790,N_4984,N_4988);
xnor UO_791 (O_791,N_4996,N_4955);
nor UO_792 (O_792,N_4941,N_4968);
nand UO_793 (O_793,N_4922,N_4911);
and UO_794 (O_794,N_4968,N_4981);
nor UO_795 (O_795,N_4915,N_4951);
nand UO_796 (O_796,N_4976,N_4993);
nand UO_797 (O_797,N_4933,N_4969);
nor UO_798 (O_798,N_4966,N_4968);
xor UO_799 (O_799,N_4984,N_4920);
nor UO_800 (O_800,N_4948,N_4949);
or UO_801 (O_801,N_4977,N_4990);
nand UO_802 (O_802,N_4907,N_4941);
xor UO_803 (O_803,N_4930,N_4973);
xor UO_804 (O_804,N_4901,N_4993);
nand UO_805 (O_805,N_4951,N_4955);
and UO_806 (O_806,N_4946,N_4999);
nand UO_807 (O_807,N_4906,N_4932);
nor UO_808 (O_808,N_4902,N_4957);
and UO_809 (O_809,N_4964,N_4903);
nor UO_810 (O_810,N_4961,N_4939);
nand UO_811 (O_811,N_4901,N_4992);
nor UO_812 (O_812,N_4909,N_4921);
nand UO_813 (O_813,N_4941,N_4939);
or UO_814 (O_814,N_4998,N_4959);
and UO_815 (O_815,N_4907,N_4904);
or UO_816 (O_816,N_4946,N_4984);
or UO_817 (O_817,N_4941,N_4912);
xor UO_818 (O_818,N_4961,N_4901);
nand UO_819 (O_819,N_4905,N_4942);
and UO_820 (O_820,N_4999,N_4916);
nand UO_821 (O_821,N_4951,N_4993);
and UO_822 (O_822,N_4918,N_4904);
and UO_823 (O_823,N_4980,N_4957);
xor UO_824 (O_824,N_4911,N_4959);
nor UO_825 (O_825,N_4935,N_4949);
or UO_826 (O_826,N_4967,N_4909);
xor UO_827 (O_827,N_4978,N_4948);
nor UO_828 (O_828,N_4903,N_4957);
or UO_829 (O_829,N_4906,N_4903);
or UO_830 (O_830,N_4935,N_4912);
nor UO_831 (O_831,N_4986,N_4954);
nand UO_832 (O_832,N_4966,N_4909);
and UO_833 (O_833,N_4925,N_4945);
nand UO_834 (O_834,N_4906,N_4967);
or UO_835 (O_835,N_4962,N_4999);
and UO_836 (O_836,N_4993,N_4923);
nand UO_837 (O_837,N_4972,N_4924);
nand UO_838 (O_838,N_4944,N_4942);
nand UO_839 (O_839,N_4927,N_4979);
and UO_840 (O_840,N_4987,N_4971);
and UO_841 (O_841,N_4937,N_4900);
nand UO_842 (O_842,N_4928,N_4986);
nand UO_843 (O_843,N_4932,N_4998);
and UO_844 (O_844,N_4912,N_4908);
or UO_845 (O_845,N_4986,N_4908);
and UO_846 (O_846,N_4981,N_4933);
xnor UO_847 (O_847,N_4925,N_4986);
nand UO_848 (O_848,N_4922,N_4991);
nor UO_849 (O_849,N_4941,N_4997);
and UO_850 (O_850,N_4911,N_4932);
and UO_851 (O_851,N_4901,N_4953);
xor UO_852 (O_852,N_4909,N_4914);
and UO_853 (O_853,N_4955,N_4986);
and UO_854 (O_854,N_4995,N_4935);
and UO_855 (O_855,N_4951,N_4925);
or UO_856 (O_856,N_4942,N_4903);
nand UO_857 (O_857,N_4958,N_4992);
and UO_858 (O_858,N_4931,N_4948);
nand UO_859 (O_859,N_4973,N_4936);
or UO_860 (O_860,N_4984,N_4967);
nand UO_861 (O_861,N_4942,N_4921);
and UO_862 (O_862,N_4961,N_4954);
and UO_863 (O_863,N_4950,N_4992);
xor UO_864 (O_864,N_4996,N_4966);
nand UO_865 (O_865,N_4931,N_4902);
and UO_866 (O_866,N_4923,N_4988);
nor UO_867 (O_867,N_4911,N_4930);
xor UO_868 (O_868,N_4995,N_4933);
and UO_869 (O_869,N_4928,N_4954);
and UO_870 (O_870,N_4901,N_4916);
and UO_871 (O_871,N_4922,N_4908);
nand UO_872 (O_872,N_4993,N_4944);
or UO_873 (O_873,N_4959,N_4961);
nor UO_874 (O_874,N_4928,N_4933);
or UO_875 (O_875,N_4943,N_4932);
nand UO_876 (O_876,N_4932,N_4919);
nor UO_877 (O_877,N_4941,N_4965);
and UO_878 (O_878,N_4950,N_4900);
nand UO_879 (O_879,N_4951,N_4935);
and UO_880 (O_880,N_4961,N_4968);
or UO_881 (O_881,N_4940,N_4959);
or UO_882 (O_882,N_4990,N_4994);
nand UO_883 (O_883,N_4965,N_4942);
and UO_884 (O_884,N_4987,N_4901);
nand UO_885 (O_885,N_4983,N_4900);
and UO_886 (O_886,N_4959,N_4928);
nor UO_887 (O_887,N_4918,N_4946);
nor UO_888 (O_888,N_4966,N_4901);
or UO_889 (O_889,N_4909,N_4923);
nand UO_890 (O_890,N_4915,N_4970);
and UO_891 (O_891,N_4903,N_4951);
or UO_892 (O_892,N_4946,N_4956);
xor UO_893 (O_893,N_4960,N_4988);
xnor UO_894 (O_894,N_4957,N_4969);
nor UO_895 (O_895,N_4934,N_4983);
or UO_896 (O_896,N_4971,N_4983);
and UO_897 (O_897,N_4993,N_4986);
or UO_898 (O_898,N_4966,N_4984);
or UO_899 (O_899,N_4973,N_4950);
xor UO_900 (O_900,N_4931,N_4957);
nor UO_901 (O_901,N_4938,N_4994);
or UO_902 (O_902,N_4941,N_4917);
or UO_903 (O_903,N_4973,N_4904);
and UO_904 (O_904,N_4905,N_4904);
nand UO_905 (O_905,N_4948,N_4984);
and UO_906 (O_906,N_4907,N_4983);
nor UO_907 (O_907,N_4970,N_4952);
nor UO_908 (O_908,N_4975,N_4985);
or UO_909 (O_909,N_4948,N_4971);
or UO_910 (O_910,N_4932,N_4904);
nand UO_911 (O_911,N_4949,N_4989);
nand UO_912 (O_912,N_4931,N_4993);
and UO_913 (O_913,N_4917,N_4925);
nor UO_914 (O_914,N_4925,N_4926);
or UO_915 (O_915,N_4944,N_4976);
or UO_916 (O_916,N_4950,N_4966);
and UO_917 (O_917,N_4922,N_4999);
and UO_918 (O_918,N_4989,N_4976);
or UO_919 (O_919,N_4995,N_4941);
xnor UO_920 (O_920,N_4905,N_4954);
and UO_921 (O_921,N_4927,N_4946);
nor UO_922 (O_922,N_4913,N_4931);
or UO_923 (O_923,N_4914,N_4913);
and UO_924 (O_924,N_4972,N_4968);
xor UO_925 (O_925,N_4928,N_4932);
and UO_926 (O_926,N_4995,N_4937);
xor UO_927 (O_927,N_4946,N_4912);
and UO_928 (O_928,N_4928,N_4980);
nor UO_929 (O_929,N_4996,N_4913);
or UO_930 (O_930,N_4912,N_4925);
nand UO_931 (O_931,N_4969,N_4931);
nor UO_932 (O_932,N_4982,N_4941);
nor UO_933 (O_933,N_4924,N_4962);
or UO_934 (O_934,N_4989,N_4921);
and UO_935 (O_935,N_4930,N_4974);
nor UO_936 (O_936,N_4976,N_4998);
or UO_937 (O_937,N_4973,N_4994);
nor UO_938 (O_938,N_4977,N_4911);
nand UO_939 (O_939,N_4990,N_4964);
nand UO_940 (O_940,N_4984,N_4937);
and UO_941 (O_941,N_4949,N_4953);
nor UO_942 (O_942,N_4951,N_4976);
nor UO_943 (O_943,N_4983,N_4915);
or UO_944 (O_944,N_4921,N_4927);
xnor UO_945 (O_945,N_4993,N_4912);
nand UO_946 (O_946,N_4914,N_4982);
nand UO_947 (O_947,N_4964,N_4933);
and UO_948 (O_948,N_4958,N_4969);
nand UO_949 (O_949,N_4919,N_4952);
and UO_950 (O_950,N_4973,N_4976);
or UO_951 (O_951,N_4961,N_4962);
xnor UO_952 (O_952,N_4985,N_4918);
nand UO_953 (O_953,N_4900,N_4984);
or UO_954 (O_954,N_4910,N_4923);
nand UO_955 (O_955,N_4904,N_4957);
and UO_956 (O_956,N_4980,N_4963);
or UO_957 (O_957,N_4949,N_4924);
nor UO_958 (O_958,N_4917,N_4924);
and UO_959 (O_959,N_4932,N_4962);
and UO_960 (O_960,N_4950,N_4972);
nor UO_961 (O_961,N_4995,N_4922);
or UO_962 (O_962,N_4902,N_4976);
xnor UO_963 (O_963,N_4991,N_4905);
or UO_964 (O_964,N_4932,N_4983);
nor UO_965 (O_965,N_4987,N_4978);
or UO_966 (O_966,N_4906,N_4907);
nor UO_967 (O_967,N_4928,N_4977);
nor UO_968 (O_968,N_4962,N_4920);
nand UO_969 (O_969,N_4943,N_4948);
nor UO_970 (O_970,N_4979,N_4919);
nor UO_971 (O_971,N_4992,N_4934);
and UO_972 (O_972,N_4976,N_4903);
nor UO_973 (O_973,N_4938,N_4912);
and UO_974 (O_974,N_4952,N_4944);
or UO_975 (O_975,N_4913,N_4934);
and UO_976 (O_976,N_4983,N_4941);
and UO_977 (O_977,N_4936,N_4995);
xor UO_978 (O_978,N_4996,N_4993);
or UO_979 (O_979,N_4904,N_4964);
nand UO_980 (O_980,N_4930,N_4917);
and UO_981 (O_981,N_4995,N_4996);
or UO_982 (O_982,N_4959,N_4999);
or UO_983 (O_983,N_4990,N_4913);
and UO_984 (O_984,N_4955,N_4905);
xor UO_985 (O_985,N_4945,N_4935);
nor UO_986 (O_986,N_4983,N_4960);
xnor UO_987 (O_987,N_4981,N_4937);
nand UO_988 (O_988,N_4907,N_4944);
nand UO_989 (O_989,N_4985,N_4938);
nand UO_990 (O_990,N_4928,N_4921);
nor UO_991 (O_991,N_4992,N_4965);
nand UO_992 (O_992,N_4985,N_4917);
xnor UO_993 (O_993,N_4906,N_4924);
or UO_994 (O_994,N_4913,N_4964);
nor UO_995 (O_995,N_4913,N_4925);
nand UO_996 (O_996,N_4911,N_4976);
nor UO_997 (O_997,N_4997,N_4919);
and UO_998 (O_998,N_4948,N_4925);
xor UO_999 (O_999,N_4991,N_4981);
endmodule