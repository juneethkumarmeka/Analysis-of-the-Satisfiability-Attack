module basic_2500_25000_3000_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_278,In_371);
xor U1 (N_1,In_1457,In_1213);
and U2 (N_2,In_925,In_585);
xor U3 (N_3,In_1350,In_1897);
nor U4 (N_4,In_52,In_1300);
xor U5 (N_5,In_1811,In_1332);
xnor U6 (N_6,In_2367,In_1173);
and U7 (N_7,In_2412,In_13);
or U8 (N_8,In_1931,In_2229);
and U9 (N_9,In_2038,In_402);
xor U10 (N_10,In_2334,In_632);
and U11 (N_11,In_1680,In_1490);
nor U12 (N_12,In_1356,In_2043);
and U13 (N_13,In_1721,In_2170);
xnor U14 (N_14,In_1299,In_591);
nor U15 (N_15,In_1198,In_645);
nand U16 (N_16,In_336,In_1708);
xnor U17 (N_17,In_1822,In_1914);
nor U18 (N_18,In_1540,In_698);
nand U19 (N_19,In_1499,In_1288);
nor U20 (N_20,In_2460,In_1113);
or U21 (N_21,In_350,In_597);
xor U22 (N_22,In_2318,In_2143);
nor U23 (N_23,In_851,In_1701);
nor U24 (N_24,In_1364,In_1690);
or U25 (N_25,In_123,In_1329);
xnor U26 (N_26,In_1804,In_1163);
and U27 (N_27,In_2049,In_1625);
nor U28 (N_28,In_1517,In_1202);
or U29 (N_29,In_427,In_1063);
nand U30 (N_30,In_1469,In_385);
or U31 (N_31,In_2354,In_477);
and U32 (N_32,In_167,In_2188);
and U33 (N_33,In_193,In_855);
xnor U34 (N_34,In_599,In_2177);
or U35 (N_35,In_265,In_163);
xnor U36 (N_36,In_2374,In_2103);
and U37 (N_37,In_1197,In_2014);
or U38 (N_38,In_2108,In_2063);
and U39 (N_39,In_759,In_458);
or U40 (N_40,In_2,In_2194);
and U41 (N_41,In_2041,In_1659);
or U42 (N_42,In_1018,In_655);
xor U43 (N_43,In_2276,In_257);
or U44 (N_44,In_1311,In_2448);
and U45 (N_45,In_2060,In_1881);
nand U46 (N_46,In_1672,In_924);
nand U47 (N_47,In_229,In_786);
xor U48 (N_48,In_2204,In_974);
xnor U49 (N_49,In_1029,In_1973);
nor U50 (N_50,In_2489,In_830);
nand U51 (N_51,In_139,In_1575);
and U52 (N_52,In_369,In_45);
xor U53 (N_53,In_2456,In_2148);
nor U54 (N_54,In_1910,In_2392);
nor U55 (N_55,In_318,In_1);
xor U56 (N_56,In_611,In_1468);
nor U57 (N_57,In_1654,In_737);
nand U58 (N_58,In_684,In_1152);
or U59 (N_59,In_399,In_2347);
and U60 (N_60,In_135,In_991);
nor U61 (N_61,In_1111,In_908);
and U62 (N_62,In_362,In_69);
nand U63 (N_63,In_798,In_1144);
xor U64 (N_64,In_1840,In_1145);
nand U65 (N_65,In_279,In_256);
or U66 (N_66,In_1806,In_1940);
and U67 (N_67,In_212,In_2158);
nand U68 (N_68,In_2244,In_457);
or U69 (N_69,In_2307,In_242);
nand U70 (N_70,In_299,In_1962);
nand U71 (N_71,In_1926,In_1449);
nand U72 (N_72,In_253,In_1417);
xor U73 (N_73,In_848,In_2436);
nand U74 (N_74,In_865,In_1409);
nand U75 (N_75,In_1651,In_62);
and U76 (N_76,In_1408,In_2110);
or U77 (N_77,In_2168,In_281);
or U78 (N_78,In_1005,In_1866);
or U79 (N_79,In_1969,In_348);
nor U80 (N_80,In_587,In_2338);
and U81 (N_81,In_156,In_209);
nand U82 (N_82,In_1780,In_125);
or U83 (N_83,In_1883,In_692);
and U84 (N_84,In_63,In_2457);
nor U85 (N_85,In_1707,In_95);
nand U86 (N_86,In_1878,In_975);
nand U87 (N_87,In_1611,In_2268);
xor U88 (N_88,In_1838,In_659);
xor U89 (N_89,In_1121,In_1714);
nor U90 (N_90,In_165,In_1676);
or U91 (N_91,In_2074,In_1218);
nand U92 (N_92,In_1475,In_1412);
nand U93 (N_93,In_2284,In_779);
or U94 (N_94,In_1293,In_817);
nand U95 (N_95,In_1512,In_929);
and U96 (N_96,In_651,In_1204);
nand U97 (N_97,In_29,In_1856);
xor U98 (N_98,In_1428,In_2261);
nand U99 (N_99,In_1407,In_543);
and U100 (N_100,In_1894,In_1712);
or U101 (N_101,In_460,In_1433);
xnor U102 (N_102,In_2393,In_164);
nor U103 (N_103,In_1867,In_787);
xor U104 (N_104,In_839,In_1777);
nor U105 (N_105,In_596,In_1139);
nor U106 (N_106,In_482,In_792);
xnor U107 (N_107,In_1219,In_861);
or U108 (N_108,In_81,In_346);
xnor U109 (N_109,In_0,In_1232);
or U110 (N_110,In_1536,In_2100);
nand U111 (N_111,In_2112,In_967);
or U112 (N_112,In_1136,In_1283);
and U113 (N_113,In_1315,In_1990);
nand U114 (N_114,In_1285,In_2228);
nand U115 (N_115,In_1869,In_1538);
and U116 (N_116,In_2432,In_963);
nand U117 (N_117,In_1051,In_1934);
or U118 (N_118,In_858,In_405);
xor U119 (N_119,In_2441,In_1747);
or U120 (N_120,In_884,In_1996);
xnor U121 (N_121,In_283,In_1434);
or U122 (N_122,In_2211,In_237);
and U123 (N_123,In_1864,In_488);
xnor U124 (N_124,In_854,In_1321);
and U125 (N_125,In_834,In_1030);
nor U126 (N_126,In_1470,In_794);
nor U127 (N_127,In_829,In_1482);
xnor U128 (N_128,In_2493,In_1599);
nor U129 (N_129,In_1862,In_1770);
nor U130 (N_130,In_629,In_961);
nand U131 (N_131,In_774,In_329);
and U132 (N_132,In_1743,In_696);
and U133 (N_133,In_2189,In_1571);
nand U134 (N_134,In_697,In_753);
nand U135 (N_135,In_1622,In_2180);
xnor U136 (N_136,In_2282,In_274);
xnor U137 (N_137,In_2409,In_1704);
xnor U138 (N_138,In_1831,In_2256);
or U139 (N_139,In_2013,In_833);
xnor U140 (N_140,In_681,In_897);
or U141 (N_141,In_894,In_625);
or U142 (N_142,In_1636,In_1270);
xor U143 (N_143,In_749,In_2327);
nand U144 (N_144,In_2251,In_714);
or U145 (N_145,In_2126,In_2184);
nor U146 (N_146,In_1724,In_2086);
nor U147 (N_147,In_1410,In_1312);
xor U148 (N_148,In_1362,In_1090);
xnor U149 (N_149,In_1049,In_1422);
xor U150 (N_150,In_2023,In_2019);
nor U151 (N_151,In_97,In_1013);
xnor U152 (N_152,In_518,In_1391);
or U153 (N_153,In_2147,In_1923);
and U154 (N_154,In_472,In_1650);
and U155 (N_155,In_1871,In_745);
and U156 (N_156,In_91,In_316);
nor U157 (N_157,In_2285,In_1220);
nand U158 (N_158,In_2012,In_937);
xnor U159 (N_159,In_1754,In_1264);
xor U160 (N_160,In_354,In_1861);
or U161 (N_161,In_2141,In_1104);
or U162 (N_162,In_464,In_33);
nor U163 (N_163,In_2315,In_2447);
and U164 (N_164,In_159,In_1166);
nor U165 (N_165,In_2042,In_1079);
nor U166 (N_166,In_2187,In_491);
nor U167 (N_167,In_1038,In_570);
nor U168 (N_168,In_1206,In_1280);
or U169 (N_169,In_280,In_2222);
nand U170 (N_170,In_111,In_1933);
xor U171 (N_171,In_1752,In_1157);
nand U172 (N_172,In_1799,In_153);
or U173 (N_173,In_2004,In_1101);
and U174 (N_174,In_537,In_351);
xnor U175 (N_175,In_2465,In_309);
xor U176 (N_176,In_539,In_1546);
xor U177 (N_177,In_1455,In_1130);
xor U178 (N_178,In_2006,In_1401);
xnor U179 (N_179,In_307,In_1769);
xor U180 (N_180,In_1942,In_1813);
nand U181 (N_181,In_2478,In_738);
xor U182 (N_182,In_536,In_1214);
xnor U183 (N_183,In_2319,In_1994);
nor U184 (N_184,In_1430,In_1068);
xnor U185 (N_185,In_227,In_945);
xor U186 (N_186,In_529,In_412);
nor U187 (N_187,In_2291,In_2459);
xnor U188 (N_188,In_1638,In_1353);
xor U189 (N_189,In_1429,In_1039);
and U190 (N_190,In_810,In_1758);
and U191 (N_191,In_2281,In_1110);
nor U192 (N_192,In_2482,In_1573);
nor U193 (N_193,In_1185,In_347);
and U194 (N_194,In_1569,In_2137);
and U195 (N_195,In_999,In_2263);
and U196 (N_196,In_1367,In_509);
nand U197 (N_197,In_284,In_795);
xor U198 (N_198,In_888,In_879);
nand U199 (N_199,In_1785,In_871);
or U200 (N_200,In_564,In_2320);
nand U201 (N_201,In_1556,In_1949);
nand U202 (N_202,In_1054,In_1282);
or U203 (N_203,In_1075,In_1972);
nand U204 (N_204,In_1067,In_1193);
nand U205 (N_205,In_382,In_923);
nor U206 (N_206,In_1252,In_2283);
or U207 (N_207,In_188,In_941);
or U208 (N_208,In_2259,In_2348);
xnor U209 (N_209,In_1235,In_653);
nor U210 (N_210,In_1249,In_634);
nor U211 (N_211,In_406,In_1447);
nand U212 (N_212,In_1802,In_1782);
nand U213 (N_213,In_550,In_705);
and U214 (N_214,In_483,In_2429);
xor U215 (N_215,In_1195,In_828);
or U216 (N_216,In_2312,In_652);
nand U217 (N_217,In_1877,In_1760);
nand U218 (N_218,In_720,In_589);
and U219 (N_219,In_2255,In_946);
or U220 (N_220,In_985,In_2215);
and U221 (N_221,In_124,In_1384);
and U222 (N_222,In_1805,In_87);
nand U223 (N_223,In_2310,In_2323);
or U224 (N_224,In_1757,In_475);
xor U225 (N_225,In_1924,In_664);
or U226 (N_226,In_685,In_57);
xor U227 (N_227,In_1526,In_2084);
nand U228 (N_228,In_1539,In_2379);
xor U229 (N_229,In_627,In_1627);
xor U230 (N_230,In_1435,In_1903);
xor U231 (N_231,In_313,In_1810);
nor U232 (N_232,In_2349,In_765);
nand U233 (N_233,In_287,In_262);
nand U234 (N_234,In_986,In_300);
or U235 (N_235,In_145,In_2124);
xor U236 (N_236,In_1096,In_1022);
or U237 (N_237,In_895,In_270);
nand U238 (N_238,In_1858,In_980);
nand U239 (N_239,In_147,In_919);
xor U240 (N_240,In_34,In_1199);
nor U241 (N_241,In_2212,In_459);
or U242 (N_242,In_1008,In_1480);
or U243 (N_243,In_217,In_508);
nand U244 (N_244,In_1365,In_1247);
nand U245 (N_245,In_400,In_1445);
or U246 (N_246,In_751,In_977);
xnor U247 (N_247,In_1907,In_2249);
xor U248 (N_248,In_1558,In_531);
nor U249 (N_249,In_1471,In_1191);
nor U250 (N_250,In_1549,In_2088);
nand U251 (N_251,In_8,In_1233);
or U252 (N_252,In_1242,In_1523);
nor U253 (N_253,In_1901,In_1789);
xor U254 (N_254,In_1863,In_1560);
and U255 (N_255,In_1003,In_484);
or U256 (N_256,In_2499,In_733);
nor U257 (N_257,In_2160,In_1203);
and U258 (N_258,In_1084,In_2171);
or U259 (N_259,In_492,In_397);
xnor U260 (N_260,In_1043,In_1014);
xnor U261 (N_261,In_1713,In_958);
and U262 (N_262,In_1501,In_517);
and U263 (N_263,In_2302,In_1669);
or U264 (N_264,In_1089,In_847);
nor U265 (N_265,In_2361,In_1513);
or U266 (N_266,In_886,In_534);
or U267 (N_267,In_1146,In_2186);
nand U268 (N_268,In_31,In_2484);
nor U269 (N_269,In_1272,In_100);
and U270 (N_270,In_2237,In_1153);
and U271 (N_271,In_2421,In_388);
nor U272 (N_272,In_1454,In_70);
or U273 (N_273,In_2142,In_1221);
xnor U274 (N_274,In_1631,In_1685);
nand U275 (N_275,In_86,In_2450);
nand U276 (N_276,In_1462,In_2300);
or U277 (N_277,In_2010,In_1527);
or U278 (N_278,In_979,In_690);
or U279 (N_279,In_2156,In_2411);
nor U280 (N_280,In_2238,In_1617);
nand U281 (N_281,In_1621,In_776);
and U282 (N_282,In_114,In_2073);
nor U283 (N_283,In_1016,In_248);
or U284 (N_284,In_1913,In_746);
xor U285 (N_285,In_1053,In_1699);
xor U286 (N_286,In_571,In_1390);
or U287 (N_287,In_682,In_345);
nand U288 (N_288,In_729,In_2169);
xor U289 (N_289,In_505,In_558);
or U290 (N_290,In_821,In_1208);
or U291 (N_291,In_2383,In_359);
xor U292 (N_292,In_90,In_1269);
and U293 (N_293,In_301,In_218);
nor U294 (N_294,In_415,In_356);
or U295 (N_295,In_1187,In_88);
nor U296 (N_296,In_1587,In_18);
or U297 (N_297,In_2225,In_1892);
xnor U298 (N_298,In_85,In_292);
nand U299 (N_299,In_1301,In_141);
or U300 (N_300,In_2136,In_1413);
xor U301 (N_301,In_998,In_805);
and U302 (N_302,In_1953,In_1920);
nand U303 (N_303,In_376,In_936);
xnor U304 (N_304,In_50,In_1594);
and U305 (N_305,In_1223,In_379);
nor U306 (N_306,In_1492,In_321);
xnor U307 (N_307,In_1226,In_1879);
xor U308 (N_308,In_1547,In_1670);
nor U309 (N_309,In_1976,In_452);
and U310 (N_310,In_1960,In_541);
or U311 (N_311,In_14,In_981);
xor U312 (N_312,In_2192,In_918);
nand U313 (N_313,In_2306,In_2353);
or U314 (N_314,In_661,In_71);
or U315 (N_315,In_557,In_691);
or U316 (N_316,In_559,In_1023);
and U317 (N_317,In_2253,In_1438);
and U318 (N_318,In_339,In_902);
nor U319 (N_319,In_468,In_323);
nor U320 (N_320,In_1419,In_906);
xnor U321 (N_321,In_1331,In_2352);
xor U322 (N_322,In_832,In_2395);
xnor U323 (N_323,In_2332,In_732);
xnor U324 (N_324,In_1395,In_2471);
nand U325 (N_325,In_480,In_222);
xnor U326 (N_326,In_1290,In_1541);
nor U327 (N_327,In_731,In_1974);
and U328 (N_328,In_1776,In_1403);
and U329 (N_329,In_2005,In_1865);
nand U330 (N_330,In_173,In_984);
nor U331 (N_331,In_2366,In_556);
or U332 (N_332,In_411,In_1201);
xor U333 (N_333,In_435,In_577);
nor U334 (N_334,In_1653,In_1125);
nand U335 (N_335,In_1108,In_780);
nand U336 (N_336,In_1641,In_2166);
nor U337 (N_337,In_1306,In_380);
or U338 (N_338,In_221,In_1278);
or U339 (N_339,In_899,In_620);
or U340 (N_340,In_1619,In_211);
or U341 (N_341,In_1647,In_1916);
nand U342 (N_342,In_2199,In_2105);
and U343 (N_343,In_2350,In_580);
or U344 (N_344,In_2378,In_410);
and U345 (N_345,In_758,In_2297);
nor U346 (N_346,In_2000,In_2260);
nor U347 (N_347,In_2406,In_421);
and U348 (N_348,In_357,In_2339);
and U349 (N_349,In_743,In_643);
nor U350 (N_350,In_210,In_1963);
nor U351 (N_351,In_2464,In_319);
and U352 (N_352,In_2410,In_291);
and U353 (N_353,In_275,In_213);
xnor U354 (N_354,In_2027,In_2183);
or U355 (N_355,In_1815,In_880);
xnor U356 (N_356,In_1807,In_909);
nand U357 (N_357,In_453,In_1689);
or U358 (N_358,In_662,In_2321);
and U359 (N_359,In_1124,In_2033);
or U360 (N_360,In_1932,In_1336);
nor U361 (N_361,In_286,In_2317);
nand U362 (N_362,In_2446,In_2364);
xor U363 (N_363,In_717,In_660);
xnor U364 (N_364,In_710,In_2236);
nand U365 (N_365,In_568,In_1261);
and U366 (N_366,In_108,In_1886);
xor U367 (N_367,In_656,In_1086);
xnor U368 (N_368,In_101,In_1880);
nor U369 (N_369,In_1281,In_782);
nand U370 (N_370,In_2007,In_48);
or U371 (N_371,In_510,In_2162);
or U372 (N_372,In_1277,In_1786);
xor U373 (N_373,In_2051,In_1506);
or U374 (N_374,In_1602,In_1081);
and U375 (N_375,In_1465,In_1060);
nand U376 (N_376,In_1964,In_375);
nor U377 (N_377,In_1779,In_674);
xor U378 (N_378,In_1225,In_2381);
or U379 (N_379,In_812,In_1262);
or U380 (N_380,In_1093,In_1010);
xor U381 (N_381,In_1762,In_616);
or U382 (N_382,In_2483,In_387);
nand U383 (N_383,In_1504,In_424);
nand U384 (N_384,In_2359,In_395);
xnor U385 (N_385,In_1240,In_1098);
or U386 (N_386,In_404,In_1255);
xor U387 (N_387,In_2331,In_361);
and U388 (N_388,In_1692,In_451);
or U389 (N_389,In_1411,In_609);
nor U390 (N_390,In_874,In_791);
and U391 (N_391,In_131,In_1369);
xor U392 (N_392,In_1818,In_32);
xor U393 (N_393,In_302,In_26);
nand U394 (N_394,In_1943,In_1832);
xor U395 (N_395,In_140,In_1735);
nand U396 (N_396,In_2152,In_1525);
or U397 (N_397,In_1948,In_996);
xor U398 (N_398,In_2330,In_2239);
xor U399 (N_399,In_566,In_703);
nor U400 (N_400,In_2468,In_930);
nand U401 (N_401,In_1006,In_2064);
and U402 (N_402,In_1474,In_1154);
nand U403 (N_403,In_1908,In_586);
nand U404 (N_404,In_752,In_335);
or U405 (N_405,In_1129,In_1229);
nand U406 (N_406,In_2087,In_1600);
nor U407 (N_407,In_2071,In_1359);
xnor U408 (N_408,In_850,In_1246);
and U409 (N_409,In_1801,In_1115);
or U410 (N_410,In_504,In_143);
and U411 (N_411,In_1833,In_1478);
nand U412 (N_412,In_181,In_770);
xor U413 (N_413,In_706,In_957);
nand U414 (N_414,In_2208,In_119);
xnor U415 (N_415,In_2373,In_1341);
nand U416 (N_416,In_2178,In_1792);
nand U417 (N_417,In_133,In_27);
or U418 (N_418,In_254,In_1088);
nand U419 (N_419,In_920,In_1491);
and U420 (N_420,In_1716,In_1849);
and U421 (N_421,In_2149,In_2342);
nand U422 (N_422,In_636,In_2495);
nor U423 (N_423,In_324,In_1027);
and U424 (N_424,In_2217,In_264);
xor U425 (N_425,In_1693,In_2485);
or U426 (N_426,In_224,In_523);
xnor U427 (N_427,In_2104,In_463);
and U428 (N_428,In_2397,In_1303);
and U429 (N_429,In_1773,In_5);
nor U430 (N_430,In_964,In_2009);
nand U431 (N_431,In_1889,In_498);
or U432 (N_432,In_514,In_1566);
and U433 (N_433,In_311,In_538);
and U434 (N_434,In_337,In_2055);
nor U435 (N_435,In_2335,In_522);
and U436 (N_436,In_962,In_740);
nand U437 (N_437,In_940,In_2139);
nor U438 (N_438,In_19,In_988);
nand U439 (N_439,In_973,In_1464);
xor U440 (N_440,In_1925,In_947);
nor U441 (N_441,In_1772,In_1420);
nor U442 (N_442,In_870,In_613);
nand U443 (N_443,In_1230,In_485);
nand U444 (N_444,In_840,In_1893);
nor U445 (N_445,In_1114,In_983);
xnor U446 (N_446,In_1905,In_2479);
or U447 (N_447,In_1993,In_420);
nor U448 (N_448,In_116,In_1576);
xnor U449 (N_449,In_1510,In_1586);
xnor U450 (N_450,In_355,In_1660);
nor U451 (N_451,In_863,In_1755);
nand U452 (N_452,In_1657,In_2434);
xor U453 (N_453,In_814,In_654);
xor U454 (N_454,In_2266,In_1040);
nand U455 (N_455,In_519,In_1138);
xnor U456 (N_456,In_1565,In_515);
nor U457 (N_457,In_305,In_55);
nand U458 (N_458,In_1405,In_1705);
xor U459 (N_459,In_592,In_490);
nand U460 (N_460,In_1548,In_1292);
xnor U461 (N_461,In_1266,In_1256);
nand U462 (N_462,In_2277,In_1000);
and U463 (N_463,In_608,In_1644);
nand U464 (N_464,In_251,In_1936);
nor U465 (N_465,In_1372,In_588);
and U466 (N_466,In_842,In_852);
nor U467 (N_467,In_1921,In_2018);
or U468 (N_468,In_470,In_1874);
xnor U469 (N_469,In_174,In_252);
xnor U470 (N_470,In_285,In_1335);
xor U471 (N_471,In_234,In_158);
xnor U472 (N_472,In_1550,In_1992);
or U473 (N_473,In_1190,In_1851);
nand U474 (N_474,In_1959,In_968);
or U475 (N_475,In_1396,In_1048);
or U476 (N_476,In_1170,In_185);
xor U477 (N_477,In_1887,In_2206);
and U478 (N_478,In_2114,In_2032);
and U479 (N_479,In_2340,In_2427);
nor U480 (N_480,In_1590,In_1258);
and U481 (N_481,In_1212,In_1155);
and U482 (N_482,In_149,In_2414);
or U483 (N_483,In_409,In_73);
xor U484 (N_484,In_712,In_1828);
nand U485 (N_485,In_2449,In_450);
or U486 (N_486,In_293,In_511);
xnor U487 (N_487,In_203,In_670);
nand U488 (N_488,In_462,In_809);
nor U489 (N_489,In_2190,In_1977);
and U490 (N_490,In_836,In_1065);
nand U491 (N_491,In_2377,In_2454);
nand U492 (N_492,In_1906,In_1847);
or U493 (N_493,In_177,In_943);
nor U494 (N_494,In_934,In_1626);
xor U495 (N_495,In_1694,In_532);
xor U496 (N_496,In_1911,In_1749);
nand U497 (N_497,In_1683,In_1265);
xnor U498 (N_498,In_171,In_2119);
nor U499 (N_499,In_2274,In_2415);
xnor U500 (N_500,In_1995,In_443);
nor U501 (N_501,In_892,In_1450);
nor U502 (N_502,In_1437,In_1181);
nor U503 (N_503,In_1764,In_2247);
or U504 (N_504,In_1425,In_1273);
and U505 (N_505,In_39,In_763);
xor U506 (N_506,In_1530,In_1629);
nor U507 (N_507,In_30,In_2035);
nor U508 (N_508,In_1015,In_521);
or U509 (N_509,In_2314,In_2252);
xor U510 (N_510,In_1824,In_1071);
nor U511 (N_511,In_1354,In_1333);
xnor U512 (N_512,In_1623,In_994);
or U513 (N_513,In_1058,In_1616);
nand U514 (N_514,In_314,In_1318);
and U515 (N_515,In_772,In_2078);
xor U516 (N_516,In_2057,In_449);
or U517 (N_517,In_864,In_907);
nor U518 (N_518,In_2294,In_428);
or U519 (N_519,In_2404,In_819);
nand U520 (N_520,In_701,In_2492);
nor U521 (N_521,In_465,In_2355);
nor U522 (N_522,In_1718,In_1338);
and U523 (N_523,In_2469,In_912);
nor U524 (N_524,In_2102,In_294);
or U525 (N_525,In_1207,In_196);
and U526 (N_526,In_1736,In_425);
or U527 (N_527,In_150,In_1358);
or U528 (N_528,In_2047,In_1684);
xor U529 (N_529,In_1326,In_2385);
nand U530 (N_530,In_1046,In_1555);
xor U531 (N_531,In_496,In_1509);
nand U532 (N_532,In_2232,In_2090);
or U533 (N_533,In_647,In_1946);
or U534 (N_534,In_827,In_408);
nand U535 (N_535,In_360,In_144);
nand U536 (N_536,In_77,In_807);
or U537 (N_537,In_2230,In_1386);
nand U538 (N_538,In_1452,In_250);
or U539 (N_539,In_1885,In_1250);
xnor U540 (N_540,In_1286,In_1244);
or U541 (N_541,In_2157,In_1514);
and U542 (N_542,In_1648,In_2210);
xnor U543 (N_543,In_1105,In_1604);
xnor U544 (N_544,In_1162,In_1231);
xor U545 (N_545,In_1444,In_756);
xnor U546 (N_546,In_1106,In_2301);
nand U547 (N_547,In_1605,In_2197);
nand U548 (N_548,In_191,In_1937);
xnor U549 (N_549,In_2134,In_494);
nand U550 (N_550,In_1852,In_1825);
and U551 (N_551,In_604,In_2205);
or U552 (N_552,In_2396,In_1983);
or U553 (N_553,In_904,In_1361);
nand U554 (N_554,In_2207,In_2029);
or U555 (N_555,In_860,In_939);
nor U556 (N_556,In_328,In_1902);
nor U557 (N_557,In_1939,In_1888);
nand U558 (N_558,In_1222,In_2030);
xnor U559 (N_559,In_137,In_679);
nor U560 (N_560,In_1642,In_2054);
or U561 (N_561,In_1767,In_2262);
and U562 (N_562,In_2203,In_1733);
and U563 (N_563,In_2356,In_398);
xnor U564 (N_564,In_942,In_180);
or U565 (N_565,In_1328,In_1026);
nand U566 (N_566,In_680,In_40);
nand U567 (N_567,In_1418,In_1746);
nand U568 (N_568,In_2098,In_353);
and U569 (N_569,In_330,In_37);
xnor U570 (N_570,In_750,In_436);
or U571 (N_571,In_1095,In_99);
nand U572 (N_572,In_268,In_623);
and U573 (N_573,In_700,In_1578);
nand U574 (N_574,In_1238,In_128);
and U575 (N_575,In_553,In_104);
xnor U576 (N_576,In_1097,In_479);
nand U577 (N_577,In_3,In_2272);
nor U578 (N_578,In_1323,In_1044);
nand U579 (N_579,In_1728,In_663);
nor U580 (N_580,In_1663,In_430);
or U581 (N_581,In_927,In_438);
xnor U582 (N_582,In_2120,In_184);
and U583 (N_583,In_2431,In_2181);
and U584 (N_584,In_243,In_2453);
nor U585 (N_585,In_2389,In_755);
nand U586 (N_586,In_862,In_1563);
nor U587 (N_587,In_802,In_1756);
nand U588 (N_588,In_1451,In_562);
xor U589 (N_589,In_215,In_1087);
nor U590 (N_590,In_1662,In_1004);
or U591 (N_591,In_1632,In_1304);
and U592 (N_592,In_1287,In_2219);
nand U593 (N_593,In_734,In_722);
nand U594 (N_594,In_1343,In_1415);
xor U595 (N_595,In_1966,In_65);
xnor U596 (N_596,In_598,In_2059);
and U597 (N_597,In_2117,In_676);
nor U598 (N_598,In_1345,In_1533);
nor U599 (N_599,In_1703,In_2015);
or U600 (N_600,In_1399,In_1700);
or U601 (N_601,In_1846,In_971);
nand U602 (N_602,In_2036,In_7);
and U603 (N_603,In_2144,In_1416);
nor U604 (N_604,In_2002,In_2494);
nand U605 (N_605,In_1373,In_78);
xnor U606 (N_606,In_1376,In_2417);
xnor U607 (N_607,In_122,In_735);
xnor U608 (N_608,In_273,In_1289);
nor U609 (N_609,In_1614,In_688);
or U610 (N_610,In_1370,In_36);
nor U611 (N_611,In_2423,In_889);
nand U612 (N_612,In_1149,In_2167);
nand U613 (N_613,In_667,In_2050);
or U614 (N_614,In_481,In_417);
and U615 (N_615,In_615,In_1975);
nor U616 (N_616,In_573,In_1062);
and U617 (N_617,In_736,In_2405);
nand U618 (N_618,In_2094,In_1494);
nor U619 (N_619,In_320,In_695);
nor U620 (N_620,In_1073,In_1085);
nand U621 (N_621,In_1589,In_1519);
or U622 (N_622,In_1050,In_2221);
and U623 (N_623,In_474,In_2265);
nand U624 (N_624,In_2498,In_1164);
xor U625 (N_625,In_993,In_600);
nor U626 (N_626,In_2351,In_1673);
or U627 (N_627,In_2390,In_310);
nand U628 (N_628,In_1956,In_151);
nor U629 (N_629,In_1618,In_1309);
and U630 (N_630,In_2091,In_1980);
nand U631 (N_631,In_2269,In_2164);
and U632 (N_632,In_2303,In_240);
xnor U633 (N_633,In_1172,In_2155);
nor U634 (N_634,In_2153,In_584);
nor U635 (N_635,In_1045,In_102);
nand U636 (N_636,In_1796,In_675);
and U637 (N_637,In_1486,In_1774);
or U638 (N_638,In_1687,In_1398);
and U639 (N_639,In_447,In_1377);
and U640 (N_640,In_711,In_1317);
or U641 (N_641,In_1112,In_1823);
xor U642 (N_642,In_109,In_1165);
or U643 (N_643,In_1037,In_308);
nor U644 (N_644,In_1371,In_426);
nand U645 (N_645,In_2026,In_1957);
nand U646 (N_646,In_1140,In_2267);
nor U647 (N_647,In_1845,In_844);
nand U648 (N_648,In_1483,In_1378);
xor U649 (N_649,In_1986,In_1927);
nor U650 (N_650,In_1606,In_219);
and U651 (N_651,In_1055,In_2235);
nor U652 (N_652,In_2174,In_1790);
nor U653 (N_653,In_1123,In_2243);
nor U654 (N_654,In_707,In_1634);
nor U655 (N_655,In_2257,In_921);
or U656 (N_656,In_2288,In_1147);
nand U657 (N_657,In_2401,In_466);
nor U658 (N_658,In_2008,In_1128);
xnor U659 (N_659,In_1951,In_1518);
nor U660 (N_660,In_325,In_2173);
nand U661 (N_661,In_393,In_641);
or U662 (N_662,In_183,In_825);
nor U663 (N_663,In_192,In_2313);
nand U664 (N_664,In_642,In_2324);
or U665 (N_665,In_2433,In_1981);
xor U666 (N_666,In_2357,In_2343);
and U667 (N_667,In_2270,In_1691);
xnor U668 (N_668,In_226,In_785);
or U669 (N_669,In_823,In_2278);
or U670 (N_670,In_49,In_1327);
and U671 (N_671,In_804,In_1339);
or U672 (N_672,In_2254,In_1209);
and U673 (N_673,In_198,In_694);
nand U674 (N_674,In_877,In_1876);
nor U675 (N_675,In_2426,In_434);
or U676 (N_676,In_1307,In_607);
nand U677 (N_677,In_1553,In_1929);
nand U678 (N_678,In_959,In_194);
xnor U679 (N_679,In_105,In_1295);
and U680 (N_680,In_561,In_2079);
or U681 (N_681,In_2034,In_1064);
nand U682 (N_682,In_866,In_1019);
nand U683 (N_683,In_258,In_503);
and U684 (N_684,In_901,In_127);
xor U685 (N_685,In_1917,In_796);
or U686 (N_686,In_2227,In_1070);
xor U687 (N_687,In_803,In_1667);
xnor U688 (N_688,In_1583,In_1440);
xnor U689 (N_689,In_1349,In_113);
xnor U690 (N_690,In_1665,In_1524);
xor U691 (N_691,In_622,In_186);
or U692 (N_692,In_726,In_11);
nand U693 (N_693,In_952,In_1991);
xnor U694 (N_694,In_22,In_2496);
nor U695 (N_695,In_1696,In_835);
or U696 (N_696,In_2360,In_1947);
nor U697 (N_697,In_1271,In_1135);
and U698 (N_698,In_1508,In_2070);
xnor U699 (N_699,In_1854,In_1814);
and U700 (N_700,In_1351,In_693);
or U701 (N_701,In_686,In_190);
or U702 (N_702,In_2001,In_1406);
or U703 (N_703,In_363,In_1711);
nand U704 (N_704,In_172,In_2293);
and U705 (N_705,In_232,In_1859);
and U706 (N_706,In_915,In_1784);
xor U707 (N_707,In_1507,In_1117);
xnor U708 (N_708,In_715,In_2066);
and U709 (N_709,In_204,In_2109);
nor U710 (N_710,In_2376,In_1296);
and U711 (N_711,In_2371,In_1744);
and U712 (N_712,In_2214,In_121);
xor U713 (N_713,In_1729,In_1585);
nor U714 (N_714,In_1568,In_2438);
or U715 (N_715,In_2151,In_487);
nand U716 (N_716,In_633,In_2422);
nand U717 (N_717,In_1839,In_1502);
nand U718 (N_718,In_1387,In_2248);
or U719 (N_719,In_1593,In_130);
nand U720 (N_720,In_1768,In_157);
xor U721 (N_721,In_79,In_666);
xor U722 (N_722,In_1817,In_51);
and U723 (N_723,In_1723,In_2394);
nand U724 (N_724,In_1720,In_1997);
or U725 (N_725,In_1968,In_969);
nor U726 (N_726,In_2344,In_2474);
nand U727 (N_727,In_1809,In_2309);
nand U728 (N_728,In_724,In_867);
or U729 (N_729,In_1355,In_1922);
nand U730 (N_730,In_2154,In_1150);
or U731 (N_731,In_118,In_1347);
xor U732 (N_732,In_28,In_1884);
nand U733 (N_733,In_432,In_1596);
and U734 (N_734,In_1950,In_1674);
nor U735 (N_735,In_2486,In_134);
and U736 (N_736,In_1970,In_1584);
nor U737 (N_737,In_2345,In_1340);
and U738 (N_738,In_1383,In_554);
xnor U739 (N_739,In_671,In_235);
or U740 (N_740,In_1603,In_2216);
nand U741 (N_741,In_205,In_1572);
nand U742 (N_742,In_2362,In_2299);
or U743 (N_743,In_1196,In_2304);
nand U744 (N_744,In_2082,In_1002);
nand U745 (N_745,In_326,In_42);
xnor U746 (N_746,In_507,In_418);
and U747 (N_747,In_669,In_1380);
or U748 (N_748,In_1263,In_1564);
xor U749 (N_749,In_1609,In_885);
and U750 (N_750,In_2264,In_502);
or U751 (N_751,In_1116,In_2455);
or U752 (N_752,In_495,In_197);
and U753 (N_753,In_1741,In_64);
and U754 (N_754,In_767,In_60);
and U755 (N_755,In_757,In_766);
or U756 (N_756,In_520,In_811);
xor U757 (N_757,In_1612,In_1652);
nor U758 (N_758,In_304,In_1057);
and U759 (N_759,In_548,In_2037);
nor U760 (N_760,In_1254,In_1260);
xor U761 (N_761,In_1788,In_138);
nor U762 (N_762,In_881,In_2475);
nor U763 (N_763,In_657,In_298);
or U764 (N_764,In_718,In_2308);
xor U765 (N_765,In_989,In_893);
xnor U766 (N_766,In_790,In_72);
xor U767 (N_767,In_315,In_506);
xnor U768 (N_768,In_16,In_1241);
nor U769 (N_769,In_574,In_444);
xnor U770 (N_770,In_38,In_80);
and U771 (N_771,In_1182,In_1320);
and U772 (N_772,In_231,In_446);
or U773 (N_773,In_241,In_949);
xnor U774 (N_774,In_1857,In_1158);
nand U775 (N_775,In_2083,In_84);
xor U776 (N_776,In_1224,In_658);
xor U777 (N_777,In_489,In_312);
xor U778 (N_778,In_1601,In_1276);
and U779 (N_779,In_1890,In_220);
nand U780 (N_780,In_35,In_2135);
nand U781 (N_781,In_1082,In_1597);
nor U782 (N_782,In_1217,In_461);
nand U783 (N_783,In_1717,In_1771);
and U784 (N_784,In_1928,In_2161);
nor U785 (N_785,In_728,In_891);
xnor U786 (N_786,In_1414,In_951);
nand U787 (N_787,In_1985,In_1176);
nand U788 (N_788,In_1787,In_2290);
or U789 (N_789,In_1479,In_813);
and U790 (N_790,In_2127,In_2425);
xnor U791 (N_791,In_581,In_2470);
nand U792 (N_792,In_2025,In_20);
xnor U793 (N_793,In_2444,In_162);
nand U794 (N_794,In_4,In_2065);
nor U795 (N_795,In_486,In_2458);
xnor U796 (N_796,In_1179,In_2077);
nand U797 (N_797,In_365,In_225);
xnor U798 (N_798,In_1174,In_2106);
nor U799 (N_799,In_2138,In_2295);
or U800 (N_800,In_638,In_1918);
and U801 (N_801,In_1374,In_849);
or U802 (N_802,In_890,In_2391);
nor U803 (N_803,In_1730,In_579);
nor U804 (N_804,In_605,In_2311);
and U805 (N_805,In_46,In_2461);
xor U806 (N_806,In_1275,In_1069);
and U807 (N_807,In_1812,In_606);
and U808 (N_808,In_1167,In_953);
and U809 (N_809,In_2476,In_2011);
xor U810 (N_810,In_1516,In_249);
nor U811 (N_811,In_1967,In_214);
xnor U812 (N_812,In_1133,In_1633);
xor U813 (N_813,In_2382,In_1661);
nor U814 (N_814,In_1800,In_266);
xor U815 (N_815,In_2046,In_2424);
nor U816 (N_816,In_1025,In_900);
xor U817 (N_817,In_155,In_910);
and U818 (N_818,In_1382,In_1868);
or U819 (N_819,In_775,In_2133);
xor U820 (N_820,In_2130,In_601);
and U821 (N_821,In_2022,In_563);
or U822 (N_822,In_2150,In_1551);
and U823 (N_823,In_1909,In_760);
nor U824 (N_824,In_469,In_2440);
nand U825 (N_825,In_2341,In_1793);
and U826 (N_826,In_640,In_1915);
or U827 (N_827,In_1834,In_549);
nor U828 (N_828,In_1803,In_2329);
nor U829 (N_829,In_1719,In_372);
xor U830 (N_830,In_1821,In_338);
nand U831 (N_831,In_1697,In_903);
nor U832 (N_832,In_2193,In_59);
and U833 (N_833,In_987,In_841);
nor U834 (N_834,In_259,In_1177);
xor U835 (N_835,In_2419,In_1076);
xnor U836 (N_836,In_1753,In_1314);
and U837 (N_837,In_1511,In_1615);
and U838 (N_838,In_2031,In_1268);
or U839 (N_839,In_76,In_2363);
and U840 (N_840,In_896,In_9);
or U841 (N_841,In_1795,In_1935);
nand U842 (N_842,In_1151,In_1477);
or U843 (N_843,In_132,In_53);
xnor U844 (N_844,In_617,In_1357);
or U845 (N_845,In_1109,In_303);
nor U846 (N_846,In_637,In_1557);
xnor U847 (N_847,In_972,In_970);
and U848 (N_848,In_754,In_578);
or U849 (N_849,In_1554,In_2132);
and U850 (N_850,In_1459,In_2368);
nor U851 (N_851,In_93,In_1368);
nand U852 (N_852,In_818,In_883);
nor U853 (N_853,In_290,In_2003);
and U854 (N_854,In_1965,In_1702);
xor U855 (N_855,In_110,In_2039);
or U856 (N_856,In_1047,In_112);
nor U857 (N_857,In_1102,In_1431);
xnor U858 (N_858,In_75,In_1302);
or U859 (N_859,In_820,In_1895);
nand U860 (N_860,In_1522,In_713);
or U861 (N_861,In_2116,In_1192);
or U862 (N_862,In_1945,In_2163);
or U863 (N_863,In_2028,In_476);
and U864 (N_864,In_875,In_1591);
and U865 (N_865,In_2202,In_1375);
xor U866 (N_866,In_741,In_646);
and U867 (N_867,In_407,In_730);
nor U868 (N_868,In_1559,In_2145);
nand U869 (N_869,In_445,In_2159);
nand U870 (N_870,In_546,In_1808);
nor U871 (N_871,In_17,In_978);
nor U872 (N_872,In_744,In_2435);
nand U873 (N_873,In_2080,In_801);
nor U874 (N_874,In_364,In_524);
or U875 (N_875,In_115,In_761);
nor U876 (N_876,In_800,In_1971);
nor U877 (N_877,In_24,In_107);
and U878 (N_878,In_1346,In_2305);
nor U879 (N_879,In_678,In_126);
nor U880 (N_880,In_1498,In_1322);
or U881 (N_881,In_160,In_1798);
nor U882 (N_882,In_628,In_1987);
nand U883 (N_883,In_1456,In_1899);
and U884 (N_884,In_2497,In_2146);
and U885 (N_885,In_1216,In_331);
xor U886 (N_886,In_1186,In_2287);
xnor U887 (N_887,In_1161,In_1007);
and U888 (N_888,In_1706,In_665);
xnor U889 (N_889,In_1325,In_2245);
xor U890 (N_890,In_1184,In_358);
nor U891 (N_891,In_2016,In_859);
and U892 (N_892,In_567,In_1397);
xor U893 (N_893,In_2081,In_1678);
or U894 (N_894,In_742,In_2467);
and U895 (N_895,In_208,In_1819);
and U896 (N_896,In_2275,In_1253);
nor U897 (N_897,In_1671,In_1009);
and U898 (N_898,In_928,In_2490);
nor U899 (N_899,In_1620,In_440);
nor U900 (N_900,In_853,In_2076);
or U901 (N_901,In_1582,In_2388);
nor U902 (N_902,In_2384,In_552);
xor U903 (N_903,In_2118,In_535);
nand U904 (N_904,In_932,In_228);
or U905 (N_905,In_2328,In_1842);
xor U906 (N_906,In_1580,In_551);
and U907 (N_907,In_2407,In_1898);
nand U908 (N_908,In_282,In_368);
or U909 (N_909,In_263,In_189);
nor U910 (N_910,In_2200,In_2398);
nor U911 (N_911,In_2175,In_1820);
nand U912 (N_912,In_1682,In_1954);
and U913 (N_913,In_89,In_783);
nor U914 (N_914,In_1656,In_1982);
nand U915 (N_915,In_423,In_2418);
xor U916 (N_916,In_1481,In_593);
nand U917 (N_917,In_374,In_1001);
nor U918 (N_918,In_575,In_1882);
and U919 (N_919,In_2185,In_1131);
and U920 (N_920,In_1503,In_1279);
and U921 (N_921,In_2387,In_322);
and U922 (N_922,In_808,In_2058);
and U923 (N_923,In_202,In_478);
nand U924 (N_924,In_1134,In_1194);
or U925 (N_925,In_1726,In_2258);
nor U926 (N_926,In_1020,In_2316);
xor U927 (N_927,In_624,In_1912);
or U928 (N_928,In_672,In_378);
xor U929 (N_929,In_1393,In_1872);
nand U930 (N_930,In_2129,In_289);
and U931 (N_931,In_1577,In_168);
and U932 (N_932,In_1120,In_2487);
xnor U933 (N_933,In_223,In_630);
nor U934 (N_934,In_148,In_1952);
nand U935 (N_935,In_96,In_1267);
nand U936 (N_936,In_442,In_1637);
nand U937 (N_937,In_1245,In_201);
xnor U938 (N_938,In_547,In_1423);
or U939 (N_939,In_2336,In_723);
and U940 (N_940,In_2224,In_2096);
nor U941 (N_941,In_1542,In_1781);
nor U942 (N_942,In_689,In_649);
or U943 (N_943,In_267,In_725);
nor U944 (N_944,In_23,In_471);
and U945 (N_945,In_784,In_704);
xnor U946 (N_946,In_621,In_1178);
and U947 (N_947,In_1156,In_542);
and U948 (N_948,In_1313,In_1737);
nor U949 (N_949,In_384,In_2128);
nand U950 (N_950,In_1775,In_1143);
or U951 (N_951,In_1032,In_439);
xor U952 (N_952,In_1826,In_1236);
and U953 (N_953,In_1738,In_612);
or U954 (N_954,In_92,In_1794);
nand U955 (N_955,In_1761,In_873);
xnor U956 (N_956,In_306,In_1337);
xor U957 (N_957,In_1052,In_857);
or U958 (N_958,In_152,In_822);
or U959 (N_959,In_831,In_1200);
and U960 (N_960,In_544,In_1243);
nand U961 (N_961,In_1686,In_525);
xnor U962 (N_962,In_1366,In_142);
nor U963 (N_963,In_277,In_419);
nor U964 (N_964,In_2322,In_1443);
or U965 (N_965,In_1461,In_1466);
nand U966 (N_966,In_1463,In_2140);
xor U967 (N_967,In_244,In_2430);
nand U968 (N_968,In_297,In_2045);
xnor U969 (N_969,In_673,In_1783);
or U970 (N_970,In_1984,In_416);
nor U971 (N_971,In_1835,In_2400);
nand U972 (N_972,In_2380,In_255);
nand U973 (N_973,In_239,In_716);
or U974 (N_974,In_1552,In_938);
or U975 (N_975,In_2213,In_1715);
xnor U976 (N_976,In_422,In_799);
and U977 (N_977,In_1107,In_1042);
or U978 (N_978,In_403,In_83);
nand U979 (N_979,In_1436,In_352);
nor U980 (N_980,In_6,In_966);
and U981 (N_981,In_377,In_2220);
nand U982 (N_982,In_824,In_1215);
xor U983 (N_983,In_768,In_603);
xnor U984 (N_984,In_1142,In_2223);
nor U985 (N_985,In_762,In_1581);
or U986 (N_986,In_499,In_473);
or U987 (N_987,In_2271,In_1999);
and U988 (N_988,In_1251,In_1958);
xnor U989 (N_989,In_1141,In_1453);
nor U990 (N_990,In_2298,In_120);
or U991 (N_991,In_1126,In_1745);
or U992 (N_992,In_1751,In_1442);
and U993 (N_993,In_614,In_2131);
nand U994 (N_994,In_1298,In_1137);
nor U995 (N_995,In_1679,In_1677);
nand U996 (N_996,In_856,In_1850);
nand U997 (N_997,In_1989,In_1348);
and U998 (N_998,In_10,In_1392);
or U999 (N_999,In_576,In_230);
or U1000 (N_1000,In_1432,In_1658);
xnor U1001 (N_1001,In_1210,In_341);
xor U1002 (N_1002,In_2044,In_1860);
nand U1003 (N_1003,In_777,In_455);
or U1004 (N_1004,In_650,In_2452);
nand U1005 (N_1005,In_1344,In_1324);
nand U1006 (N_1006,In_207,In_342);
nand U1007 (N_1007,In_1535,In_1837);
nor U1008 (N_1008,In_2466,In_887);
and U1009 (N_1009,In_2481,In_1493);
nor U1010 (N_1010,In_1011,In_2241);
nor U1011 (N_1011,In_1031,In_2099);
nor U1012 (N_1012,In_788,In_233);
nand U1013 (N_1013,In_2093,In_1160);
xnor U1014 (N_1014,In_21,In_1476);
or U1015 (N_1015,In_2280,In_1520);
nand U1016 (N_1016,In_764,In_1148);
xor U1017 (N_1017,In_1078,In_1979);
and U1018 (N_1018,In_216,In_2372);
or U1019 (N_1019,In_1766,In_2346);
nor U1020 (N_1020,In_317,In_1649);
nor U1021 (N_1021,In_2068,In_454);
or U1022 (N_1022,In_401,In_739);
nor U1023 (N_1023,In_954,In_2123);
xor U1024 (N_1024,In_1424,In_527);
and U1025 (N_1025,In_648,In_2101);
xnor U1026 (N_1026,In_1330,In_129);
nand U1027 (N_1027,In_1579,In_456);
nor U1028 (N_1028,In_1896,In_433);
xor U1029 (N_1029,In_195,In_2020);
nor U1030 (N_1030,In_1829,In_497);
nor U1031 (N_1031,In_2402,In_2273);
nor U1032 (N_1032,In_1211,In_948);
and U1033 (N_1033,In_965,In_2333);
nand U1034 (N_1034,In_1574,In_1588);
nor U1035 (N_1035,In_771,In_1830);
nand U1036 (N_1036,In_1870,In_1844);
nor U1037 (N_1037,In_1472,In_1534);
nor U1038 (N_1038,In_1567,In_2231);
and U1039 (N_1039,In_1237,In_1610);
nor U1040 (N_1040,In_98,In_843);
nor U1041 (N_1041,In_187,In_1646);
or U1042 (N_1042,In_1035,In_1941);
and U1043 (N_1043,In_619,In_1797);
nor U1044 (N_1044,In_1645,In_635);
and U1045 (N_1045,In_2179,In_2292);
or U1046 (N_1046,In_396,In_1034);
or U1047 (N_1047,In_516,In_699);
or U1048 (N_1048,In_2358,In_1732);
or U1049 (N_1049,In_54,In_1316);
or U1050 (N_1050,In_1100,In_610);
xnor U1051 (N_1051,In_1608,In_56);
xnor U1052 (N_1052,In_702,In_2369);
nor U1053 (N_1053,In_815,In_1487);
nor U1054 (N_1054,In_1497,In_1695);
nor U1055 (N_1055,In_2234,In_781);
nand U1056 (N_1056,In_161,In_793);
nand U1057 (N_1057,In_1944,In_389);
nand U1058 (N_1058,In_1630,In_367);
xnor U1059 (N_1059,In_602,In_555);
nor U1060 (N_1060,In_1036,In_1904);
or U1061 (N_1061,In_1291,In_1092);
nand U1062 (N_1062,In_2111,In_719);
and U1063 (N_1063,In_2122,In_1763);
or U1064 (N_1064,In_1528,In_1094);
and U1065 (N_1065,In_1873,In_44);
nand U1066 (N_1066,In_618,In_1189);
and U1067 (N_1067,In_687,In_1938);
or U1068 (N_1068,In_381,In_1352);
nand U1069 (N_1069,In_1072,In_2052);
xor U1070 (N_1070,In_340,In_677);
xor U1071 (N_1071,In_2326,In_914);
xor U1072 (N_1072,In_1505,In_709);
nand U1073 (N_1073,In_837,In_1521);
nand U1074 (N_1074,In_2242,In_344);
nor U1075 (N_1075,In_2095,In_2442);
xor U1076 (N_1076,In_1544,In_2480);
xor U1077 (N_1077,In_2420,In_2472);
or U1078 (N_1078,In_876,In_1132);
and U1079 (N_1079,In_1739,In_1848);
xor U1080 (N_1080,In_1891,In_2191);
nor U1081 (N_1081,In_182,In_905);
and U1082 (N_1082,In_1021,In_260);
nand U1083 (N_1083,In_721,In_2196);
nor U1084 (N_1084,In_545,In_390);
or U1085 (N_1085,In_1778,In_1394);
or U1086 (N_1086,In_806,In_526);
or U1087 (N_1087,In_12,In_1841);
xnor U1088 (N_1088,In_74,In_2056);
xor U1089 (N_1089,In_2246,In_1675);
or U1090 (N_1090,In_992,In_1635);
xnor U1091 (N_1091,In_1426,In_1360);
nand U1092 (N_1092,In_995,In_1059);
nand U1093 (N_1093,In_1091,In_271);
nand U1094 (N_1094,In_917,In_1681);
or U1095 (N_1095,In_386,In_997);
nand U1096 (N_1096,In_1740,In_288);
xnor U1097 (N_1097,In_1484,In_2289);
or U1098 (N_1098,In_2365,In_1628);
nand U1099 (N_1099,In_2048,In_1122);
nor U1100 (N_1100,In_41,In_560);
nand U1101 (N_1101,In_246,In_1066);
nand U1102 (N_1102,In_2370,In_1731);
and U1103 (N_1103,In_2092,In_170);
nor U1104 (N_1104,In_1389,In_878);
nand U1105 (N_1105,In_845,In_2488);
nor U1106 (N_1106,In_2250,In_206);
nor U1107 (N_1107,In_528,In_1613);
nand U1108 (N_1108,In_590,In_935);
or U1109 (N_1109,In_1592,In_2125);
xor U1110 (N_1110,In_2085,In_1404);
nor U1111 (N_1111,In_708,In_373);
nand U1112 (N_1112,In_748,In_869);
xor U1113 (N_1113,In_1077,In_846);
and U1114 (N_1114,In_106,In_343);
or U1115 (N_1115,In_82,In_683);
and U1116 (N_1116,In_448,In_769);
or U1117 (N_1117,In_175,In_882);
xnor U1118 (N_1118,In_1308,In_1319);
and U1119 (N_1119,In_2437,In_1439);
nand U1120 (N_1120,In_146,In_1381);
nand U1121 (N_1121,In_2017,In_441);
xnor U1122 (N_1122,In_1228,In_2337);
or U1123 (N_1123,In_1448,In_1334);
and U1124 (N_1124,In_913,In_43);
and U1125 (N_1125,In_639,In_916);
nor U1126 (N_1126,In_2463,In_1169);
xor U1127 (N_1127,In_2445,In_245);
nor U1128 (N_1128,In_2062,In_366);
or U1129 (N_1129,In_594,In_1664);
and U1130 (N_1130,In_2172,In_1183);
and U1131 (N_1131,In_2040,In_1607);
nand U1132 (N_1132,In_1041,In_1961);
nor U1133 (N_1133,In_1836,In_25);
nor U1134 (N_1134,In_595,In_1561);
and U1135 (N_1135,In_1400,In_1257);
nand U1136 (N_1136,In_1033,In_2233);
nor U1137 (N_1137,In_1791,In_272);
nor U1138 (N_1138,In_2416,In_583);
xor U1139 (N_1139,In_2075,In_1188);
or U1140 (N_1140,In_1099,In_990);
nand U1141 (N_1141,In_1460,In_431);
nand U1142 (N_1142,In_1489,In_1500);
and U1143 (N_1143,In_778,In_1624);
and U1144 (N_1144,In_176,In_1446);
and U1145 (N_1145,In_2218,In_513);
nor U1146 (N_1146,In_1168,In_1725);
and U1147 (N_1147,In_826,In_68);
or U1148 (N_1148,In_1305,In_1855);
and U1149 (N_1149,In_2451,In_1543);
nor U1150 (N_1150,In_2107,In_1742);
and U1151 (N_1151,In_1061,In_199);
nand U1152 (N_1152,In_1496,In_2491);
nand U1153 (N_1153,In_1900,In_1488);
and U1154 (N_1154,In_933,In_1843);
nor U1155 (N_1155,In_1710,In_1080);
nor U1156 (N_1156,In_1363,In_2428);
nand U1157 (N_1157,In_1159,In_1274);
nand U1158 (N_1158,In_727,In_2209);
xor U1159 (N_1159,In_117,In_1570);
xor U1160 (N_1160,In_2176,In_166);
nand U1161 (N_1161,In_2386,In_236);
and U1162 (N_1162,In_1643,In_955);
nand U1163 (N_1163,In_922,In_1056);
and U1164 (N_1164,In_1537,In_2403);
nor U1165 (N_1165,In_2201,In_467);
xnor U1166 (N_1166,In_1284,In_1666);
nor U1167 (N_1167,In_394,In_1930);
and U1168 (N_1168,In_1227,In_2053);
nor U1169 (N_1169,In_1748,In_269);
nand U1170 (N_1170,In_2115,In_136);
xnor U1171 (N_1171,In_631,In_816);
nor U1172 (N_1172,In_103,In_1640);
nand U1173 (N_1173,In_200,In_429);
or U1174 (N_1174,In_66,In_2121);
nand U1175 (N_1175,In_644,In_1441);
nand U1176 (N_1176,In_1180,In_2240);
nand U1177 (N_1177,In_1118,In_1532);
nor U1178 (N_1178,In_1175,In_2413);
nor U1179 (N_1179,In_332,In_58);
nand U1180 (N_1180,In_926,In_333);
nand U1181 (N_1181,In_1668,In_261);
and U1182 (N_1182,In_1485,In_1103);
xor U1183 (N_1183,In_2067,In_797);
or U1184 (N_1184,In_1310,In_1827);
xor U1185 (N_1185,In_1562,In_540);
nand U1186 (N_1186,In_2198,In_1342);
nand U1187 (N_1187,In_533,In_1545);
xnor U1188 (N_1188,In_1639,In_626);
nand U1189 (N_1189,In_295,In_2443);
and U1190 (N_1190,In_1515,In_1998);
and U1191 (N_1191,In_1234,In_1759);
nand U1192 (N_1192,In_1259,In_2165);
nor U1193 (N_1193,In_931,In_1495);
and U1194 (N_1194,In_565,In_247);
and U1195 (N_1195,In_1119,In_1017);
nand U1196 (N_1196,In_414,In_1083);
or U1197 (N_1197,In_334,In_383);
or U1198 (N_1198,In_327,In_944);
xnor U1199 (N_1199,In_1875,In_773);
or U1200 (N_1200,In_47,In_1978);
xnor U1201 (N_1201,In_976,In_178);
xnor U1202 (N_1202,In_1427,In_296);
nor U1203 (N_1203,In_956,In_747);
or U1204 (N_1204,In_179,In_2325);
nand U1205 (N_1205,In_2279,In_1297);
or U1206 (N_1206,In_1816,In_2399);
and U1207 (N_1207,In_1598,In_370);
xnor U1208 (N_1208,In_2072,In_1688);
nor U1209 (N_1209,In_1722,In_2375);
nor U1210 (N_1210,In_169,In_1853);
nand U1211 (N_1211,In_2113,In_1529);
and U1212 (N_1212,In_1028,In_154);
and U1213 (N_1213,In_493,In_2408);
and U1214 (N_1214,In_500,In_2473);
nor U1215 (N_1215,In_276,In_911);
and U1216 (N_1216,In_950,In_2097);
xnor U1217 (N_1217,In_349,In_1127);
and U1218 (N_1218,In_2286,In_1750);
nor U1219 (N_1219,In_1379,In_1727);
or U1220 (N_1220,In_1248,In_2069);
or U1221 (N_1221,In_2439,In_982);
nand U1222 (N_1222,In_1473,In_413);
nor U1223 (N_1223,In_1709,In_1655);
or U1224 (N_1224,In_1171,In_2024);
nand U1225 (N_1225,In_2195,In_2021);
or U1226 (N_1226,In_2089,In_582);
nand U1227 (N_1227,In_2226,In_1955);
xor U1228 (N_1228,In_872,In_572);
or U1229 (N_1229,In_1294,In_1595);
xnor U1230 (N_1230,In_94,In_1205);
nand U1231 (N_1231,In_668,In_501);
nand U1232 (N_1232,In_1458,In_61);
and U1233 (N_1233,In_1467,In_2296);
xor U1234 (N_1234,In_1012,In_392);
nand U1235 (N_1235,In_238,In_1024);
or U1236 (N_1236,In_2182,In_15);
xnor U1237 (N_1237,In_898,In_1765);
xnor U1238 (N_1238,In_1698,In_512);
or U1239 (N_1239,In_1402,In_1919);
or U1240 (N_1240,In_569,In_789);
and U1241 (N_1241,In_530,In_960);
or U1242 (N_1242,In_2061,In_391);
xnor U1243 (N_1243,In_67,In_1388);
or U1244 (N_1244,In_2462,In_1385);
and U1245 (N_1245,In_437,In_868);
nand U1246 (N_1246,In_1734,In_1531);
xnor U1247 (N_1247,In_1074,In_1988);
nand U1248 (N_1248,In_1239,In_838);
xor U1249 (N_1249,In_2477,In_1421);
or U1250 (N_1250,In_89,In_1356);
and U1251 (N_1251,In_807,In_1650);
and U1252 (N_1252,In_1701,In_1623);
and U1253 (N_1253,In_147,In_2402);
nand U1254 (N_1254,In_1376,In_1127);
nor U1255 (N_1255,In_119,In_2179);
and U1256 (N_1256,In_1409,In_2227);
nand U1257 (N_1257,In_2265,In_1644);
and U1258 (N_1258,In_921,In_464);
nand U1259 (N_1259,In_1986,In_1246);
xnor U1260 (N_1260,In_147,In_1278);
or U1261 (N_1261,In_40,In_626);
nand U1262 (N_1262,In_313,In_2457);
nand U1263 (N_1263,In_1201,In_910);
nand U1264 (N_1264,In_1573,In_1535);
nor U1265 (N_1265,In_26,In_2103);
xor U1266 (N_1266,In_1685,In_643);
and U1267 (N_1267,In_436,In_2353);
or U1268 (N_1268,In_1819,In_2087);
nand U1269 (N_1269,In_1777,In_1780);
nor U1270 (N_1270,In_2042,In_285);
nand U1271 (N_1271,In_1887,In_228);
or U1272 (N_1272,In_2491,In_221);
and U1273 (N_1273,In_1639,In_58);
nand U1274 (N_1274,In_504,In_979);
and U1275 (N_1275,In_189,In_1925);
and U1276 (N_1276,In_1118,In_1336);
nor U1277 (N_1277,In_333,In_1980);
nand U1278 (N_1278,In_1369,In_1520);
or U1279 (N_1279,In_1305,In_2345);
nand U1280 (N_1280,In_1780,In_690);
nor U1281 (N_1281,In_632,In_745);
and U1282 (N_1282,In_402,In_233);
nor U1283 (N_1283,In_1768,In_1253);
nor U1284 (N_1284,In_975,In_1607);
nand U1285 (N_1285,In_1992,In_2361);
or U1286 (N_1286,In_1673,In_1493);
nor U1287 (N_1287,In_2247,In_2448);
xor U1288 (N_1288,In_1577,In_1938);
or U1289 (N_1289,In_2305,In_1222);
nor U1290 (N_1290,In_1741,In_1204);
nand U1291 (N_1291,In_9,In_2380);
xnor U1292 (N_1292,In_1614,In_1404);
xor U1293 (N_1293,In_281,In_1279);
and U1294 (N_1294,In_451,In_1228);
and U1295 (N_1295,In_1582,In_327);
nor U1296 (N_1296,In_1797,In_832);
nand U1297 (N_1297,In_1916,In_482);
or U1298 (N_1298,In_60,In_1869);
nand U1299 (N_1299,In_1388,In_982);
nand U1300 (N_1300,In_916,In_1691);
nor U1301 (N_1301,In_509,In_788);
nor U1302 (N_1302,In_1411,In_480);
and U1303 (N_1303,In_517,In_781);
nor U1304 (N_1304,In_135,In_453);
and U1305 (N_1305,In_1682,In_2297);
xor U1306 (N_1306,In_1207,In_2193);
and U1307 (N_1307,In_1484,In_1744);
nand U1308 (N_1308,In_1620,In_322);
and U1309 (N_1309,In_1232,In_1300);
xnor U1310 (N_1310,In_390,In_97);
xnor U1311 (N_1311,In_2042,In_1472);
or U1312 (N_1312,In_1178,In_1721);
nand U1313 (N_1313,In_1768,In_1649);
nor U1314 (N_1314,In_2499,In_1129);
nor U1315 (N_1315,In_1429,In_2298);
xnor U1316 (N_1316,In_1100,In_319);
nor U1317 (N_1317,In_1097,In_2013);
and U1318 (N_1318,In_1161,In_1998);
nor U1319 (N_1319,In_1311,In_1323);
nand U1320 (N_1320,In_856,In_456);
or U1321 (N_1321,In_55,In_728);
and U1322 (N_1322,In_1024,In_2142);
and U1323 (N_1323,In_647,In_1872);
or U1324 (N_1324,In_1541,In_923);
or U1325 (N_1325,In_734,In_1939);
xor U1326 (N_1326,In_339,In_2466);
xnor U1327 (N_1327,In_1050,In_564);
or U1328 (N_1328,In_39,In_681);
xor U1329 (N_1329,In_1953,In_1443);
nand U1330 (N_1330,In_557,In_1136);
nor U1331 (N_1331,In_879,In_1988);
nor U1332 (N_1332,In_1988,In_208);
and U1333 (N_1333,In_1402,In_1991);
nand U1334 (N_1334,In_1038,In_1606);
or U1335 (N_1335,In_172,In_122);
nand U1336 (N_1336,In_1004,In_1476);
nor U1337 (N_1337,In_46,In_2059);
nand U1338 (N_1338,In_1081,In_2316);
nor U1339 (N_1339,In_528,In_2410);
nand U1340 (N_1340,In_1197,In_937);
nand U1341 (N_1341,In_1817,In_375);
or U1342 (N_1342,In_572,In_496);
xnor U1343 (N_1343,In_2121,In_845);
or U1344 (N_1344,In_2119,In_922);
or U1345 (N_1345,In_806,In_1816);
nand U1346 (N_1346,In_1034,In_1064);
or U1347 (N_1347,In_1364,In_1844);
nor U1348 (N_1348,In_1690,In_1168);
nand U1349 (N_1349,In_1020,In_1956);
and U1350 (N_1350,In_922,In_558);
and U1351 (N_1351,In_583,In_49);
nand U1352 (N_1352,In_677,In_690);
nand U1353 (N_1353,In_2296,In_653);
xnor U1354 (N_1354,In_300,In_2248);
nand U1355 (N_1355,In_1068,In_1864);
nor U1356 (N_1356,In_2000,In_1622);
or U1357 (N_1357,In_361,In_2154);
or U1358 (N_1358,In_1784,In_1313);
xnor U1359 (N_1359,In_1775,In_307);
or U1360 (N_1360,In_1014,In_1202);
and U1361 (N_1361,In_1631,In_927);
xnor U1362 (N_1362,In_2433,In_1123);
nand U1363 (N_1363,In_2489,In_1758);
nand U1364 (N_1364,In_1859,In_87);
or U1365 (N_1365,In_1144,In_2383);
nand U1366 (N_1366,In_77,In_865);
xnor U1367 (N_1367,In_300,In_909);
or U1368 (N_1368,In_919,In_721);
nand U1369 (N_1369,In_1095,In_23);
and U1370 (N_1370,In_1381,In_1880);
nand U1371 (N_1371,In_625,In_2228);
nor U1372 (N_1372,In_899,In_2272);
or U1373 (N_1373,In_1934,In_683);
nor U1374 (N_1374,In_65,In_2448);
or U1375 (N_1375,In_22,In_326);
or U1376 (N_1376,In_1605,In_664);
and U1377 (N_1377,In_1020,In_1124);
or U1378 (N_1378,In_878,In_1134);
or U1379 (N_1379,In_1284,In_577);
nor U1380 (N_1380,In_233,In_2384);
xnor U1381 (N_1381,In_630,In_908);
xor U1382 (N_1382,In_914,In_860);
nand U1383 (N_1383,In_134,In_151);
xor U1384 (N_1384,In_691,In_2026);
xnor U1385 (N_1385,In_2134,In_949);
nand U1386 (N_1386,In_2367,In_2117);
nor U1387 (N_1387,In_1222,In_1810);
or U1388 (N_1388,In_2377,In_2084);
xor U1389 (N_1389,In_918,In_253);
xor U1390 (N_1390,In_690,In_2028);
or U1391 (N_1391,In_2009,In_1768);
xor U1392 (N_1392,In_2178,In_1919);
and U1393 (N_1393,In_1833,In_2286);
or U1394 (N_1394,In_1603,In_1388);
or U1395 (N_1395,In_1055,In_886);
or U1396 (N_1396,In_2239,In_328);
nand U1397 (N_1397,In_537,In_514);
nor U1398 (N_1398,In_44,In_1880);
and U1399 (N_1399,In_1835,In_1245);
and U1400 (N_1400,In_1234,In_2489);
nand U1401 (N_1401,In_1619,In_1472);
xnor U1402 (N_1402,In_964,In_1916);
xnor U1403 (N_1403,In_814,In_1206);
nand U1404 (N_1404,In_2472,In_1433);
nand U1405 (N_1405,In_1899,In_2269);
nor U1406 (N_1406,In_1676,In_555);
or U1407 (N_1407,In_2369,In_2139);
nor U1408 (N_1408,In_1745,In_2066);
nand U1409 (N_1409,In_1478,In_1509);
xor U1410 (N_1410,In_1185,In_1003);
and U1411 (N_1411,In_736,In_391);
or U1412 (N_1412,In_401,In_539);
xor U1413 (N_1413,In_942,In_1946);
nor U1414 (N_1414,In_2453,In_578);
and U1415 (N_1415,In_861,In_1869);
nand U1416 (N_1416,In_2166,In_1380);
or U1417 (N_1417,In_493,In_641);
or U1418 (N_1418,In_2001,In_1670);
nand U1419 (N_1419,In_1461,In_1404);
nand U1420 (N_1420,In_820,In_1447);
and U1421 (N_1421,In_377,In_1279);
nor U1422 (N_1422,In_1953,In_1284);
nor U1423 (N_1423,In_1557,In_1232);
nor U1424 (N_1424,In_472,In_562);
and U1425 (N_1425,In_2112,In_1778);
xor U1426 (N_1426,In_2465,In_1337);
nor U1427 (N_1427,In_133,In_1728);
nor U1428 (N_1428,In_2415,In_2148);
nand U1429 (N_1429,In_974,In_580);
and U1430 (N_1430,In_2426,In_1352);
or U1431 (N_1431,In_281,In_1179);
nand U1432 (N_1432,In_1978,In_2004);
and U1433 (N_1433,In_2484,In_100);
and U1434 (N_1434,In_1224,In_137);
or U1435 (N_1435,In_1850,In_551);
or U1436 (N_1436,In_1494,In_2179);
or U1437 (N_1437,In_944,In_2153);
or U1438 (N_1438,In_1365,In_1317);
and U1439 (N_1439,In_313,In_215);
and U1440 (N_1440,In_552,In_297);
xnor U1441 (N_1441,In_1013,In_1940);
or U1442 (N_1442,In_1932,In_1498);
nor U1443 (N_1443,In_767,In_1007);
xnor U1444 (N_1444,In_466,In_635);
and U1445 (N_1445,In_2496,In_397);
or U1446 (N_1446,In_1055,In_686);
nor U1447 (N_1447,In_1648,In_1160);
xnor U1448 (N_1448,In_407,In_2143);
nor U1449 (N_1449,In_1693,In_1058);
or U1450 (N_1450,In_2014,In_1980);
nand U1451 (N_1451,In_1730,In_609);
xnor U1452 (N_1452,In_370,In_1448);
xnor U1453 (N_1453,In_72,In_1484);
xor U1454 (N_1454,In_485,In_1696);
and U1455 (N_1455,In_2413,In_1593);
nand U1456 (N_1456,In_2458,In_279);
xor U1457 (N_1457,In_129,In_2409);
nand U1458 (N_1458,In_1812,In_1348);
or U1459 (N_1459,In_1318,In_1087);
xor U1460 (N_1460,In_79,In_2395);
nor U1461 (N_1461,In_11,In_1780);
nor U1462 (N_1462,In_2483,In_726);
xnor U1463 (N_1463,In_655,In_1911);
xnor U1464 (N_1464,In_165,In_658);
xnor U1465 (N_1465,In_443,In_1729);
nor U1466 (N_1466,In_1157,In_738);
and U1467 (N_1467,In_1009,In_1404);
nor U1468 (N_1468,In_1953,In_726);
xnor U1469 (N_1469,In_325,In_1620);
nor U1470 (N_1470,In_2277,In_500);
and U1471 (N_1471,In_217,In_1549);
nand U1472 (N_1472,In_2010,In_1585);
and U1473 (N_1473,In_1611,In_450);
xor U1474 (N_1474,In_572,In_1784);
or U1475 (N_1475,In_687,In_408);
xor U1476 (N_1476,In_2062,In_56);
and U1477 (N_1477,In_956,In_175);
or U1478 (N_1478,In_1895,In_900);
nor U1479 (N_1479,In_1589,In_1007);
xor U1480 (N_1480,In_845,In_1659);
or U1481 (N_1481,In_1835,In_2192);
nand U1482 (N_1482,In_798,In_1121);
and U1483 (N_1483,In_1350,In_158);
nand U1484 (N_1484,In_1859,In_2286);
and U1485 (N_1485,In_1126,In_1427);
or U1486 (N_1486,In_1378,In_2204);
nor U1487 (N_1487,In_1010,In_215);
nand U1488 (N_1488,In_1142,In_822);
xnor U1489 (N_1489,In_1406,In_1262);
nor U1490 (N_1490,In_1528,In_1355);
or U1491 (N_1491,In_2181,In_2146);
nor U1492 (N_1492,In_91,In_2328);
nor U1493 (N_1493,In_2197,In_1154);
or U1494 (N_1494,In_1533,In_850);
nand U1495 (N_1495,In_636,In_1929);
or U1496 (N_1496,In_1596,In_1009);
nor U1497 (N_1497,In_82,In_1633);
xnor U1498 (N_1498,In_1351,In_608);
nand U1499 (N_1499,In_1257,In_2206);
nor U1500 (N_1500,In_946,In_1979);
nor U1501 (N_1501,In_813,In_1277);
nor U1502 (N_1502,In_644,In_1600);
and U1503 (N_1503,In_1719,In_1305);
and U1504 (N_1504,In_34,In_1887);
nor U1505 (N_1505,In_2430,In_780);
and U1506 (N_1506,In_1995,In_191);
nand U1507 (N_1507,In_708,In_1755);
nand U1508 (N_1508,In_547,In_1398);
or U1509 (N_1509,In_2284,In_1026);
or U1510 (N_1510,In_1420,In_1864);
nor U1511 (N_1511,In_1975,In_775);
nor U1512 (N_1512,In_31,In_2265);
nor U1513 (N_1513,In_1988,In_2236);
and U1514 (N_1514,In_1397,In_238);
and U1515 (N_1515,In_2118,In_339);
nand U1516 (N_1516,In_1401,In_1095);
or U1517 (N_1517,In_946,In_1231);
nand U1518 (N_1518,In_361,In_310);
nor U1519 (N_1519,In_72,In_5);
nand U1520 (N_1520,In_162,In_48);
nand U1521 (N_1521,In_2156,In_1361);
and U1522 (N_1522,In_1865,In_2469);
xnor U1523 (N_1523,In_507,In_1488);
or U1524 (N_1524,In_1008,In_1899);
xor U1525 (N_1525,In_1527,In_632);
xnor U1526 (N_1526,In_1333,In_1853);
or U1527 (N_1527,In_2446,In_1942);
nor U1528 (N_1528,In_1189,In_1958);
nor U1529 (N_1529,In_937,In_1934);
xnor U1530 (N_1530,In_2435,In_2118);
nor U1531 (N_1531,In_1361,In_466);
xor U1532 (N_1532,In_316,In_574);
xor U1533 (N_1533,In_1459,In_2469);
xor U1534 (N_1534,In_953,In_614);
or U1535 (N_1535,In_2259,In_2);
xor U1536 (N_1536,In_85,In_2399);
nand U1537 (N_1537,In_2466,In_225);
nand U1538 (N_1538,In_2319,In_703);
and U1539 (N_1539,In_2427,In_1116);
nand U1540 (N_1540,In_516,In_68);
xnor U1541 (N_1541,In_1538,In_1295);
and U1542 (N_1542,In_1616,In_817);
and U1543 (N_1543,In_2036,In_1202);
xnor U1544 (N_1544,In_198,In_2273);
or U1545 (N_1545,In_2366,In_54);
nand U1546 (N_1546,In_984,In_291);
nor U1547 (N_1547,In_284,In_440);
nor U1548 (N_1548,In_1082,In_63);
nand U1549 (N_1549,In_114,In_660);
nor U1550 (N_1550,In_0,In_730);
or U1551 (N_1551,In_1676,In_2126);
xnor U1552 (N_1552,In_830,In_916);
nand U1553 (N_1553,In_1505,In_2002);
and U1554 (N_1554,In_573,In_1864);
nand U1555 (N_1555,In_1122,In_2047);
and U1556 (N_1556,In_976,In_67);
or U1557 (N_1557,In_1595,In_491);
or U1558 (N_1558,In_399,In_1576);
nand U1559 (N_1559,In_1222,In_2366);
xnor U1560 (N_1560,In_985,In_2397);
xor U1561 (N_1561,In_1881,In_794);
nor U1562 (N_1562,In_390,In_2177);
xnor U1563 (N_1563,In_1065,In_985);
nand U1564 (N_1564,In_1411,In_190);
nor U1565 (N_1565,In_411,In_1618);
xor U1566 (N_1566,In_48,In_335);
nand U1567 (N_1567,In_1889,In_349);
nand U1568 (N_1568,In_1552,In_2092);
and U1569 (N_1569,In_2412,In_1983);
nor U1570 (N_1570,In_1936,In_970);
and U1571 (N_1571,In_329,In_1159);
or U1572 (N_1572,In_407,In_1111);
and U1573 (N_1573,In_329,In_1670);
xor U1574 (N_1574,In_195,In_1322);
nor U1575 (N_1575,In_1765,In_2021);
and U1576 (N_1576,In_1892,In_1070);
and U1577 (N_1577,In_693,In_565);
and U1578 (N_1578,In_1887,In_2312);
nor U1579 (N_1579,In_545,In_1791);
and U1580 (N_1580,In_825,In_1124);
and U1581 (N_1581,In_728,In_1197);
and U1582 (N_1582,In_666,In_586);
xnor U1583 (N_1583,In_1101,In_1299);
or U1584 (N_1584,In_2118,In_520);
nand U1585 (N_1585,In_406,In_891);
or U1586 (N_1586,In_171,In_845);
xor U1587 (N_1587,In_2320,In_1995);
nor U1588 (N_1588,In_427,In_910);
and U1589 (N_1589,In_1884,In_2281);
and U1590 (N_1590,In_1589,In_1832);
xnor U1591 (N_1591,In_1236,In_298);
and U1592 (N_1592,In_197,In_1858);
nand U1593 (N_1593,In_120,In_322);
and U1594 (N_1594,In_2003,In_1487);
or U1595 (N_1595,In_2394,In_2406);
xnor U1596 (N_1596,In_224,In_976);
and U1597 (N_1597,In_1822,In_2307);
or U1598 (N_1598,In_1913,In_701);
nor U1599 (N_1599,In_1849,In_971);
and U1600 (N_1600,In_1359,In_1687);
or U1601 (N_1601,In_2022,In_488);
nor U1602 (N_1602,In_816,In_1281);
nor U1603 (N_1603,In_1813,In_257);
xor U1604 (N_1604,In_1337,In_2447);
or U1605 (N_1605,In_1298,In_2368);
or U1606 (N_1606,In_1016,In_906);
and U1607 (N_1607,In_362,In_569);
xnor U1608 (N_1608,In_1730,In_1903);
xor U1609 (N_1609,In_831,In_493);
xor U1610 (N_1610,In_2445,In_1739);
nor U1611 (N_1611,In_313,In_1107);
or U1612 (N_1612,In_1958,In_409);
xor U1613 (N_1613,In_1421,In_1767);
xnor U1614 (N_1614,In_2291,In_1712);
nor U1615 (N_1615,In_1780,In_2454);
xor U1616 (N_1616,In_417,In_1177);
xnor U1617 (N_1617,In_1021,In_1129);
or U1618 (N_1618,In_2455,In_877);
nand U1619 (N_1619,In_67,In_2032);
and U1620 (N_1620,In_1179,In_563);
xor U1621 (N_1621,In_705,In_2086);
xor U1622 (N_1622,In_1680,In_395);
and U1623 (N_1623,In_293,In_2356);
and U1624 (N_1624,In_2488,In_1406);
xor U1625 (N_1625,In_2159,In_1871);
xor U1626 (N_1626,In_1663,In_2274);
xnor U1627 (N_1627,In_2107,In_2001);
nor U1628 (N_1628,In_2053,In_583);
or U1629 (N_1629,In_1112,In_1298);
nor U1630 (N_1630,In_1786,In_1819);
and U1631 (N_1631,In_972,In_887);
xnor U1632 (N_1632,In_2255,In_1653);
and U1633 (N_1633,In_361,In_294);
xor U1634 (N_1634,In_655,In_2172);
nor U1635 (N_1635,In_216,In_1137);
nand U1636 (N_1636,In_2021,In_1725);
xor U1637 (N_1637,In_1164,In_1642);
xnor U1638 (N_1638,In_2296,In_2212);
or U1639 (N_1639,In_2241,In_647);
xor U1640 (N_1640,In_1367,In_848);
xnor U1641 (N_1641,In_82,In_2358);
and U1642 (N_1642,In_454,In_680);
nor U1643 (N_1643,In_1430,In_1252);
or U1644 (N_1644,In_2106,In_1826);
nand U1645 (N_1645,In_1092,In_430);
nand U1646 (N_1646,In_1056,In_2304);
and U1647 (N_1647,In_782,In_1988);
nand U1648 (N_1648,In_1260,In_495);
and U1649 (N_1649,In_2159,In_974);
nor U1650 (N_1650,In_2406,In_11);
or U1651 (N_1651,In_2450,In_1864);
and U1652 (N_1652,In_878,In_1522);
nand U1653 (N_1653,In_75,In_1487);
and U1654 (N_1654,In_1185,In_2057);
nand U1655 (N_1655,In_1382,In_335);
and U1656 (N_1656,In_1196,In_499);
xor U1657 (N_1657,In_816,In_670);
xnor U1658 (N_1658,In_805,In_334);
xnor U1659 (N_1659,In_611,In_561);
or U1660 (N_1660,In_1826,In_1532);
nor U1661 (N_1661,In_2475,In_1968);
or U1662 (N_1662,In_2451,In_1538);
or U1663 (N_1663,In_1704,In_119);
nand U1664 (N_1664,In_2201,In_90);
or U1665 (N_1665,In_198,In_868);
and U1666 (N_1666,In_34,In_113);
nor U1667 (N_1667,In_1025,In_2161);
xor U1668 (N_1668,In_2193,In_1579);
nor U1669 (N_1669,In_2248,In_446);
and U1670 (N_1670,In_1229,In_1475);
or U1671 (N_1671,In_1433,In_2357);
or U1672 (N_1672,In_2010,In_2483);
xor U1673 (N_1673,In_2486,In_159);
nor U1674 (N_1674,In_737,In_1943);
nor U1675 (N_1675,In_1667,In_689);
xor U1676 (N_1676,In_1330,In_887);
nand U1677 (N_1677,In_514,In_393);
and U1678 (N_1678,In_1710,In_749);
or U1679 (N_1679,In_917,In_45);
or U1680 (N_1680,In_871,In_1204);
and U1681 (N_1681,In_229,In_1075);
nor U1682 (N_1682,In_1532,In_506);
nand U1683 (N_1683,In_2025,In_1026);
nor U1684 (N_1684,In_205,In_793);
and U1685 (N_1685,In_247,In_609);
nor U1686 (N_1686,In_1483,In_2302);
xnor U1687 (N_1687,In_2081,In_338);
nor U1688 (N_1688,In_400,In_2482);
xor U1689 (N_1689,In_2210,In_1807);
nor U1690 (N_1690,In_1610,In_533);
and U1691 (N_1691,In_871,In_1140);
and U1692 (N_1692,In_2028,In_1801);
nor U1693 (N_1693,In_818,In_2298);
and U1694 (N_1694,In_1810,In_172);
and U1695 (N_1695,In_1089,In_1557);
nor U1696 (N_1696,In_2131,In_1309);
xnor U1697 (N_1697,In_2081,In_83);
nor U1698 (N_1698,In_16,In_465);
nor U1699 (N_1699,In_462,In_2222);
and U1700 (N_1700,In_2028,In_1138);
xnor U1701 (N_1701,In_909,In_1785);
xor U1702 (N_1702,In_1625,In_747);
and U1703 (N_1703,In_1677,In_401);
and U1704 (N_1704,In_1982,In_618);
nand U1705 (N_1705,In_1420,In_756);
nand U1706 (N_1706,In_1289,In_1123);
xnor U1707 (N_1707,In_981,In_2072);
and U1708 (N_1708,In_1451,In_2019);
and U1709 (N_1709,In_2037,In_1661);
and U1710 (N_1710,In_2202,In_179);
xor U1711 (N_1711,In_160,In_115);
or U1712 (N_1712,In_1828,In_2017);
xnor U1713 (N_1713,In_737,In_1346);
nor U1714 (N_1714,In_900,In_2149);
xnor U1715 (N_1715,In_558,In_2379);
and U1716 (N_1716,In_865,In_738);
or U1717 (N_1717,In_2172,In_548);
nor U1718 (N_1718,In_209,In_1470);
xor U1719 (N_1719,In_538,In_428);
or U1720 (N_1720,In_1358,In_1325);
and U1721 (N_1721,In_81,In_1034);
xor U1722 (N_1722,In_1598,In_2104);
and U1723 (N_1723,In_1035,In_296);
or U1724 (N_1724,In_1338,In_848);
or U1725 (N_1725,In_267,In_1811);
and U1726 (N_1726,In_118,In_751);
xor U1727 (N_1727,In_7,In_1830);
and U1728 (N_1728,In_1684,In_808);
xor U1729 (N_1729,In_2392,In_1365);
and U1730 (N_1730,In_368,In_2047);
xnor U1731 (N_1731,In_1855,In_2256);
nor U1732 (N_1732,In_505,In_1512);
and U1733 (N_1733,In_2427,In_1220);
and U1734 (N_1734,In_687,In_1948);
or U1735 (N_1735,In_903,In_2004);
or U1736 (N_1736,In_2126,In_2122);
nor U1737 (N_1737,In_863,In_2024);
xor U1738 (N_1738,In_1403,In_1195);
nor U1739 (N_1739,In_851,In_219);
or U1740 (N_1740,In_708,In_135);
and U1741 (N_1741,In_679,In_1930);
and U1742 (N_1742,In_359,In_1318);
nor U1743 (N_1743,In_1625,In_49);
xnor U1744 (N_1744,In_1375,In_239);
nand U1745 (N_1745,In_1052,In_2401);
xor U1746 (N_1746,In_2324,In_2007);
nand U1747 (N_1747,In_1882,In_2061);
and U1748 (N_1748,In_276,In_1313);
and U1749 (N_1749,In_284,In_2461);
nor U1750 (N_1750,In_399,In_842);
xor U1751 (N_1751,In_2317,In_1739);
and U1752 (N_1752,In_2065,In_938);
or U1753 (N_1753,In_2448,In_1527);
and U1754 (N_1754,In_1187,In_1041);
nand U1755 (N_1755,In_1743,In_895);
nand U1756 (N_1756,In_728,In_1830);
nor U1757 (N_1757,In_956,In_2217);
or U1758 (N_1758,In_228,In_2380);
or U1759 (N_1759,In_288,In_33);
and U1760 (N_1760,In_2103,In_1108);
nand U1761 (N_1761,In_1134,In_2272);
nor U1762 (N_1762,In_1904,In_2101);
nand U1763 (N_1763,In_1357,In_852);
or U1764 (N_1764,In_2254,In_70);
and U1765 (N_1765,In_813,In_1937);
xor U1766 (N_1766,In_936,In_401);
xnor U1767 (N_1767,In_448,In_133);
and U1768 (N_1768,In_1919,In_245);
xor U1769 (N_1769,In_2464,In_720);
nor U1770 (N_1770,In_770,In_1675);
nor U1771 (N_1771,In_2062,In_1245);
and U1772 (N_1772,In_2422,In_10);
or U1773 (N_1773,In_1040,In_261);
and U1774 (N_1774,In_2472,In_14);
xnor U1775 (N_1775,In_2004,In_296);
xor U1776 (N_1776,In_1238,In_1409);
nor U1777 (N_1777,In_702,In_731);
nor U1778 (N_1778,In_2343,In_243);
nand U1779 (N_1779,In_475,In_2412);
xnor U1780 (N_1780,In_2226,In_497);
nor U1781 (N_1781,In_936,In_2082);
xnor U1782 (N_1782,In_362,In_1532);
or U1783 (N_1783,In_2117,In_104);
and U1784 (N_1784,In_690,In_1331);
and U1785 (N_1785,In_2332,In_534);
xor U1786 (N_1786,In_738,In_2268);
xnor U1787 (N_1787,In_1899,In_1350);
and U1788 (N_1788,In_1299,In_334);
nand U1789 (N_1789,In_1296,In_47);
xor U1790 (N_1790,In_1383,In_320);
or U1791 (N_1791,In_350,In_2367);
and U1792 (N_1792,In_1533,In_1540);
and U1793 (N_1793,In_152,In_2163);
nand U1794 (N_1794,In_124,In_672);
nand U1795 (N_1795,In_920,In_2389);
xor U1796 (N_1796,In_295,In_973);
or U1797 (N_1797,In_1688,In_1744);
or U1798 (N_1798,In_1661,In_212);
xor U1799 (N_1799,In_656,In_260);
and U1800 (N_1800,In_997,In_1942);
and U1801 (N_1801,In_265,In_1556);
or U1802 (N_1802,In_672,In_1917);
or U1803 (N_1803,In_2228,In_1463);
and U1804 (N_1804,In_887,In_168);
xnor U1805 (N_1805,In_1715,In_668);
xor U1806 (N_1806,In_1901,In_1107);
and U1807 (N_1807,In_1854,In_1004);
and U1808 (N_1808,In_2324,In_1027);
nand U1809 (N_1809,In_962,In_2243);
xor U1810 (N_1810,In_729,In_95);
nor U1811 (N_1811,In_2151,In_1339);
xor U1812 (N_1812,In_16,In_1698);
nand U1813 (N_1813,In_724,In_549);
and U1814 (N_1814,In_3,In_1615);
or U1815 (N_1815,In_888,In_269);
nor U1816 (N_1816,In_2452,In_2467);
nand U1817 (N_1817,In_1167,In_759);
or U1818 (N_1818,In_1076,In_2116);
and U1819 (N_1819,In_1405,In_235);
or U1820 (N_1820,In_1875,In_2476);
nand U1821 (N_1821,In_1236,In_215);
xor U1822 (N_1822,In_867,In_808);
xor U1823 (N_1823,In_2191,In_757);
nor U1824 (N_1824,In_590,In_1470);
nand U1825 (N_1825,In_1999,In_171);
nand U1826 (N_1826,In_1226,In_2179);
nand U1827 (N_1827,In_2132,In_1510);
or U1828 (N_1828,In_339,In_2277);
nor U1829 (N_1829,In_1546,In_2088);
and U1830 (N_1830,In_518,In_2305);
nor U1831 (N_1831,In_270,In_590);
or U1832 (N_1832,In_239,In_16);
and U1833 (N_1833,In_1919,In_2008);
nor U1834 (N_1834,In_1666,In_1590);
nand U1835 (N_1835,In_191,In_1615);
or U1836 (N_1836,In_1847,In_2161);
xor U1837 (N_1837,In_1111,In_721);
or U1838 (N_1838,In_2387,In_26);
and U1839 (N_1839,In_1028,In_1693);
and U1840 (N_1840,In_627,In_2406);
and U1841 (N_1841,In_1701,In_591);
nand U1842 (N_1842,In_1886,In_1892);
xor U1843 (N_1843,In_1553,In_282);
and U1844 (N_1844,In_2046,In_1652);
and U1845 (N_1845,In_1691,In_1165);
xnor U1846 (N_1846,In_809,In_1291);
or U1847 (N_1847,In_2310,In_274);
nor U1848 (N_1848,In_1313,In_1442);
nor U1849 (N_1849,In_147,In_906);
or U1850 (N_1850,In_174,In_547);
xnor U1851 (N_1851,In_1104,In_165);
nor U1852 (N_1852,In_1375,In_1268);
nor U1853 (N_1853,In_226,In_2434);
or U1854 (N_1854,In_2204,In_1789);
xnor U1855 (N_1855,In_1105,In_2035);
xor U1856 (N_1856,In_1834,In_1138);
nand U1857 (N_1857,In_747,In_1080);
nand U1858 (N_1858,In_1558,In_2072);
nand U1859 (N_1859,In_163,In_2019);
nand U1860 (N_1860,In_1290,In_1030);
and U1861 (N_1861,In_1946,In_1693);
and U1862 (N_1862,In_1196,In_17);
xor U1863 (N_1863,In_594,In_1002);
nand U1864 (N_1864,In_2428,In_2440);
nand U1865 (N_1865,In_1681,In_1785);
nor U1866 (N_1866,In_1098,In_1138);
nor U1867 (N_1867,In_618,In_1759);
and U1868 (N_1868,In_1134,In_868);
nand U1869 (N_1869,In_1174,In_2109);
xnor U1870 (N_1870,In_2089,In_1014);
nor U1871 (N_1871,In_1504,In_919);
nand U1872 (N_1872,In_2157,In_416);
nand U1873 (N_1873,In_1299,In_2253);
nand U1874 (N_1874,In_2135,In_1397);
and U1875 (N_1875,In_228,In_2181);
and U1876 (N_1876,In_13,In_2447);
nor U1877 (N_1877,In_387,In_784);
and U1878 (N_1878,In_2434,In_642);
nor U1879 (N_1879,In_1444,In_78);
and U1880 (N_1880,In_1436,In_1108);
nor U1881 (N_1881,In_1102,In_1560);
and U1882 (N_1882,In_412,In_62);
nand U1883 (N_1883,In_744,In_1208);
and U1884 (N_1884,In_2493,In_1301);
xor U1885 (N_1885,In_2489,In_2322);
nand U1886 (N_1886,In_658,In_166);
nand U1887 (N_1887,In_2061,In_1509);
and U1888 (N_1888,In_474,In_1184);
and U1889 (N_1889,In_210,In_1053);
nand U1890 (N_1890,In_911,In_2244);
xor U1891 (N_1891,In_2472,In_179);
nor U1892 (N_1892,In_933,In_1156);
nand U1893 (N_1893,In_575,In_1412);
nor U1894 (N_1894,In_258,In_889);
xnor U1895 (N_1895,In_881,In_175);
nand U1896 (N_1896,In_478,In_2109);
and U1897 (N_1897,In_1155,In_63);
and U1898 (N_1898,In_1194,In_674);
and U1899 (N_1899,In_676,In_1639);
nor U1900 (N_1900,In_1576,In_1172);
xor U1901 (N_1901,In_1134,In_501);
or U1902 (N_1902,In_610,In_2139);
nor U1903 (N_1903,In_813,In_1669);
and U1904 (N_1904,In_424,In_1733);
or U1905 (N_1905,In_1065,In_583);
and U1906 (N_1906,In_1807,In_1068);
nor U1907 (N_1907,In_1944,In_1587);
or U1908 (N_1908,In_1232,In_1977);
or U1909 (N_1909,In_1290,In_2202);
and U1910 (N_1910,In_310,In_1011);
nor U1911 (N_1911,In_69,In_2229);
nor U1912 (N_1912,In_208,In_511);
and U1913 (N_1913,In_2388,In_915);
xnor U1914 (N_1914,In_514,In_109);
or U1915 (N_1915,In_2124,In_2363);
and U1916 (N_1916,In_385,In_1639);
xor U1917 (N_1917,In_582,In_1746);
xnor U1918 (N_1918,In_2195,In_434);
xnor U1919 (N_1919,In_2139,In_2141);
nor U1920 (N_1920,In_1605,In_2184);
nand U1921 (N_1921,In_1667,In_1415);
xnor U1922 (N_1922,In_2358,In_1916);
xnor U1923 (N_1923,In_1833,In_1851);
nor U1924 (N_1924,In_1657,In_1676);
xnor U1925 (N_1925,In_479,In_1975);
and U1926 (N_1926,In_2231,In_2187);
and U1927 (N_1927,In_540,In_1624);
or U1928 (N_1928,In_1204,In_2462);
nand U1929 (N_1929,In_901,In_2128);
or U1930 (N_1930,In_2447,In_862);
nor U1931 (N_1931,In_1492,In_1651);
nand U1932 (N_1932,In_1432,In_2251);
or U1933 (N_1933,In_2187,In_2225);
xnor U1934 (N_1934,In_778,In_941);
or U1935 (N_1935,In_129,In_1697);
or U1936 (N_1936,In_348,In_119);
and U1937 (N_1937,In_538,In_2222);
and U1938 (N_1938,In_574,In_162);
or U1939 (N_1939,In_1543,In_1912);
xor U1940 (N_1940,In_844,In_167);
and U1941 (N_1941,In_1183,In_1469);
and U1942 (N_1942,In_1488,In_1043);
and U1943 (N_1943,In_365,In_980);
nand U1944 (N_1944,In_38,In_1236);
and U1945 (N_1945,In_1453,In_2332);
nand U1946 (N_1946,In_2265,In_1421);
nand U1947 (N_1947,In_1453,In_2043);
nor U1948 (N_1948,In_1127,In_1950);
nand U1949 (N_1949,In_1042,In_1708);
nand U1950 (N_1950,In_1859,In_1415);
or U1951 (N_1951,In_2351,In_839);
nor U1952 (N_1952,In_2365,In_1224);
nor U1953 (N_1953,In_2142,In_203);
nand U1954 (N_1954,In_325,In_6);
and U1955 (N_1955,In_2400,In_1390);
nor U1956 (N_1956,In_1775,In_2255);
nor U1957 (N_1957,In_1366,In_848);
and U1958 (N_1958,In_1449,In_2042);
xor U1959 (N_1959,In_1557,In_1903);
or U1960 (N_1960,In_533,In_219);
nor U1961 (N_1961,In_968,In_218);
or U1962 (N_1962,In_2136,In_22);
nor U1963 (N_1963,In_1823,In_86);
xor U1964 (N_1964,In_2400,In_48);
nor U1965 (N_1965,In_1716,In_1582);
and U1966 (N_1966,In_2373,In_257);
nand U1967 (N_1967,In_462,In_1924);
xor U1968 (N_1968,In_1530,In_272);
nand U1969 (N_1969,In_1828,In_920);
xnor U1970 (N_1970,In_169,In_1706);
nor U1971 (N_1971,In_1751,In_2443);
or U1972 (N_1972,In_1026,In_2400);
xor U1973 (N_1973,In_113,In_2478);
nor U1974 (N_1974,In_1697,In_2294);
nor U1975 (N_1975,In_1156,In_1568);
nand U1976 (N_1976,In_2295,In_141);
nor U1977 (N_1977,In_482,In_1359);
and U1978 (N_1978,In_1237,In_1149);
nand U1979 (N_1979,In_1181,In_1571);
nand U1980 (N_1980,In_2268,In_1074);
nand U1981 (N_1981,In_279,In_609);
nand U1982 (N_1982,In_1264,In_195);
and U1983 (N_1983,In_671,In_1242);
nand U1984 (N_1984,In_1491,In_1086);
nand U1985 (N_1985,In_276,In_2381);
nand U1986 (N_1986,In_874,In_469);
or U1987 (N_1987,In_788,In_1790);
nor U1988 (N_1988,In_1305,In_629);
or U1989 (N_1989,In_270,In_1296);
xor U1990 (N_1990,In_180,In_1657);
nand U1991 (N_1991,In_1805,In_428);
nand U1992 (N_1992,In_336,In_107);
nand U1993 (N_1993,In_1704,In_1529);
and U1994 (N_1994,In_810,In_2015);
and U1995 (N_1995,In_1493,In_1250);
nor U1996 (N_1996,In_1889,In_27);
and U1997 (N_1997,In_2056,In_1738);
nor U1998 (N_1998,In_1941,In_1563);
nand U1999 (N_1999,In_2472,In_762);
and U2000 (N_2000,In_1571,In_1693);
nor U2001 (N_2001,In_937,In_2389);
nor U2002 (N_2002,In_2184,In_1551);
nor U2003 (N_2003,In_114,In_1894);
nor U2004 (N_2004,In_1799,In_2311);
nand U2005 (N_2005,In_406,In_741);
and U2006 (N_2006,In_177,In_1345);
or U2007 (N_2007,In_798,In_751);
nor U2008 (N_2008,In_768,In_747);
xor U2009 (N_2009,In_1424,In_1509);
xor U2010 (N_2010,In_1214,In_1537);
and U2011 (N_2011,In_439,In_933);
xnor U2012 (N_2012,In_2070,In_2090);
or U2013 (N_2013,In_608,In_1523);
and U2014 (N_2014,In_2017,In_582);
nand U2015 (N_2015,In_193,In_1448);
and U2016 (N_2016,In_1738,In_112);
or U2017 (N_2017,In_2003,In_1931);
xor U2018 (N_2018,In_2400,In_2132);
and U2019 (N_2019,In_123,In_1860);
or U2020 (N_2020,In_1472,In_1304);
and U2021 (N_2021,In_1,In_327);
nand U2022 (N_2022,In_908,In_1222);
nor U2023 (N_2023,In_2147,In_898);
xnor U2024 (N_2024,In_799,In_2198);
xor U2025 (N_2025,In_65,In_1674);
or U2026 (N_2026,In_2250,In_2189);
xnor U2027 (N_2027,In_1791,In_2056);
xor U2028 (N_2028,In_1341,In_2440);
nor U2029 (N_2029,In_859,In_234);
or U2030 (N_2030,In_1901,In_2273);
xnor U2031 (N_2031,In_838,In_474);
nand U2032 (N_2032,In_2153,In_2081);
nor U2033 (N_2033,In_472,In_485);
xnor U2034 (N_2034,In_1930,In_2281);
nor U2035 (N_2035,In_1072,In_1314);
and U2036 (N_2036,In_2190,In_1709);
nor U2037 (N_2037,In_1106,In_1758);
or U2038 (N_2038,In_1422,In_1989);
nand U2039 (N_2039,In_270,In_1772);
or U2040 (N_2040,In_1264,In_1402);
nor U2041 (N_2041,In_1741,In_1631);
xnor U2042 (N_2042,In_2315,In_2132);
nor U2043 (N_2043,In_1777,In_190);
xor U2044 (N_2044,In_1585,In_738);
and U2045 (N_2045,In_2368,In_1304);
nand U2046 (N_2046,In_2251,In_2464);
nor U2047 (N_2047,In_408,In_1195);
or U2048 (N_2048,In_1582,In_1462);
nand U2049 (N_2049,In_177,In_2384);
xnor U2050 (N_2050,In_1016,In_761);
and U2051 (N_2051,In_147,In_793);
or U2052 (N_2052,In_1496,In_1969);
xnor U2053 (N_2053,In_1489,In_1934);
nor U2054 (N_2054,In_473,In_2246);
nor U2055 (N_2055,In_361,In_761);
and U2056 (N_2056,In_2183,In_1564);
or U2057 (N_2057,In_612,In_982);
nor U2058 (N_2058,In_1230,In_1279);
xor U2059 (N_2059,In_1129,In_1165);
and U2060 (N_2060,In_2466,In_600);
xnor U2061 (N_2061,In_2456,In_990);
or U2062 (N_2062,In_170,In_865);
nor U2063 (N_2063,In_116,In_997);
and U2064 (N_2064,In_238,In_1921);
xnor U2065 (N_2065,In_1920,In_1151);
nand U2066 (N_2066,In_517,In_1277);
xor U2067 (N_2067,In_828,In_82);
nand U2068 (N_2068,In_272,In_1225);
nand U2069 (N_2069,In_2107,In_1373);
nand U2070 (N_2070,In_2365,In_535);
nand U2071 (N_2071,In_905,In_2064);
nor U2072 (N_2072,In_2351,In_1348);
or U2073 (N_2073,In_659,In_406);
xor U2074 (N_2074,In_2009,In_756);
or U2075 (N_2075,In_2127,In_1765);
nand U2076 (N_2076,In_1899,In_1058);
or U2077 (N_2077,In_2070,In_1060);
and U2078 (N_2078,In_1433,In_406);
xnor U2079 (N_2079,In_1057,In_2489);
nor U2080 (N_2080,In_465,In_1798);
or U2081 (N_2081,In_584,In_167);
or U2082 (N_2082,In_1517,In_1594);
nand U2083 (N_2083,In_455,In_2008);
nor U2084 (N_2084,In_540,In_1441);
nor U2085 (N_2085,In_583,In_773);
nor U2086 (N_2086,In_1670,In_1482);
and U2087 (N_2087,In_202,In_591);
nand U2088 (N_2088,In_1252,In_2435);
xor U2089 (N_2089,In_1964,In_386);
and U2090 (N_2090,In_1471,In_2252);
or U2091 (N_2091,In_1530,In_1599);
nor U2092 (N_2092,In_769,In_642);
and U2093 (N_2093,In_1889,In_329);
xnor U2094 (N_2094,In_404,In_1843);
nand U2095 (N_2095,In_2424,In_1580);
or U2096 (N_2096,In_2007,In_1417);
nor U2097 (N_2097,In_1732,In_894);
nor U2098 (N_2098,In_754,In_1811);
or U2099 (N_2099,In_98,In_1895);
nand U2100 (N_2100,In_1787,In_1469);
nand U2101 (N_2101,In_1973,In_837);
xnor U2102 (N_2102,In_1027,In_5);
and U2103 (N_2103,In_840,In_1376);
xnor U2104 (N_2104,In_1731,In_356);
or U2105 (N_2105,In_1506,In_158);
nor U2106 (N_2106,In_925,In_247);
and U2107 (N_2107,In_2260,In_764);
or U2108 (N_2108,In_2073,In_226);
nor U2109 (N_2109,In_427,In_739);
nor U2110 (N_2110,In_1328,In_563);
nor U2111 (N_2111,In_1094,In_379);
nand U2112 (N_2112,In_523,In_728);
xnor U2113 (N_2113,In_1892,In_1944);
nor U2114 (N_2114,In_274,In_503);
and U2115 (N_2115,In_326,In_277);
xor U2116 (N_2116,In_87,In_86);
xor U2117 (N_2117,In_1357,In_589);
xor U2118 (N_2118,In_239,In_1436);
xnor U2119 (N_2119,In_962,In_876);
nor U2120 (N_2120,In_1184,In_1943);
and U2121 (N_2121,In_703,In_1075);
xor U2122 (N_2122,In_308,In_958);
or U2123 (N_2123,In_296,In_2152);
nand U2124 (N_2124,In_1223,In_377);
nand U2125 (N_2125,In_1905,In_2022);
and U2126 (N_2126,In_885,In_1715);
nor U2127 (N_2127,In_2291,In_1327);
and U2128 (N_2128,In_272,In_1007);
and U2129 (N_2129,In_431,In_768);
nor U2130 (N_2130,In_786,In_86);
and U2131 (N_2131,In_1628,In_1994);
xnor U2132 (N_2132,In_1076,In_1654);
xor U2133 (N_2133,In_65,In_2480);
or U2134 (N_2134,In_1544,In_1475);
xnor U2135 (N_2135,In_1897,In_1467);
and U2136 (N_2136,In_2127,In_809);
or U2137 (N_2137,In_2156,In_1208);
and U2138 (N_2138,In_1893,In_1177);
nand U2139 (N_2139,In_1969,In_1619);
or U2140 (N_2140,In_1083,In_1248);
or U2141 (N_2141,In_1385,In_1083);
or U2142 (N_2142,In_1268,In_1798);
and U2143 (N_2143,In_1951,In_1213);
nand U2144 (N_2144,In_1223,In_1007);
xnor U2145 (N_2145,In_1252,In_1422);
or U2146 (N_2146,In_630,In_1501);
or U2147 (N_2147,In_2264,In_1428);
nor U2148 (N_2148,In_2110,In_1550);
or U2149 (N_2149,In_878,In_2021);
xnor U2150 (N_2150,In_1822,In_606);
or U2151 (N_2151,In_2308,In_1682);
and U2152 (N_2152,In_1261,In_1187);
or U2153 (N_2153,In_1943,In_1680);
nor U2154 (N_2154,In_1870,In_2402);
xor U2155 (N_2155,In_1848,In_1332);
nand U2156 (N_2156,In_616,In_2213);
nand U2157 (N_2157,In_22,In_1597);
xor U2158 (N_2158,In_746,In_1555);
xnor U2159 (N_2159,In_2111,In_673);
nor U2160 (N_2160,In_1750,In_2052);
xnor U2161 (N_2161,In_1119,In_695);
nand U2162 (N_2162,In_1831,In_473);
and U2163 (N_2163,In_20,In_1874);
or U2164 (N_2164,In_2001,In_657);
xor U2165 (N_2165,In_728,In_2191);
nand U2166 (N_2166,In_333,In_1697);
nor U2167 (N_2167,In_909,In_1695);
nand U2168 (N_2168,In_1035,In_1650);
nand U2169 (N_2169,In_1325,In_10);
xor U2170 (N_2170,In_2483,In_1244);
nor U2171 (N_2171,In_1699,In_343);
or U2172 (N_2172,In_1090,In_1389);
nor U2173 (N_2173,In_2140,In_181);
nor U2174 (N_2174,In_978,In_2335);
xor U2175 (N_2175,In_2426,In_2023);
and U2176 (N_2176,In_789,In_2172);
xor U2177 (N_2177,In_1304,In_945);
nor U2178 (N_2178,In_488,In_998);
nand U2179 (N_2179,In_859,In_1382);
xnor U2180 (N_2180,In_783,In_1820);
and U2181 (N_2181,In_892,In_2362);
nor U2182 (N_2182,In_1623,In_2099);
nor U2183 (N_2183,In_61,In_922);
xor U2184 (N_2184,In_377,In_2013);
xor U2185 (N_2185,In_1698,In_1758);
nand U2186 (N_2186,In_1720,In_2488);
nand U2187 (N_2187,In_1384,In_1132);
nand U2188 (N_2188,In_519,In_1745);
nor U2189 (N_2189,In_789,In_2128);
and U2190 (N_2190,In_1385,In_892);
and U2191 (N_2191,In_2340,In_150);
xor U2192 (N_2192,In_1266,In_1822);
nand U2193 (N_2193,In_1691,In_531);
or U2194 (N_2194,In_1159,In_1425);
or U2195 (N_2195,In_1042,In_482);
and U2196 (N_2196,In_1682,In_1505);
and U2197 (N_2197,In_260,In_2240);
and U2198 (N_2198,In_739,In_443);
xor U2199 (N_2199,In_841,In_2277);
or U2200 (N_2200,In_1071,In_2038);
nand U2201 (N_2201,In_1804,In_29);
or U2202 (N_2202,In_1507,In_2457);
xnor U2203 (N_2203,In_1152,In_1279);
and U2204 (N_2204,In_58,In_2241);
nor U2205 (N_2205,In_1179,In_690);
nand U2206 (N_2206,In_372,In_313);
or U2207 (N_2207,In_1757,In_1066);
and U2208 (N_2208,In_1215,In_399);
or U2209 (N_2209,In_590,In_2433);
xnor U2210 (N_2210,In_2021,In_2429);
xnor U2211 (N_2211,In_1540,In_199);
or U2212 (N_2212,In_564,In_1357);
nor U2213 (N_2213,In_768,In_1320);
or U2214 (N_2214,In_2128,In_504);
and U2215 (N_2215,In_1763,In_1760);
nand U2216 (N_2216,In_673,In_2297);
nor U2217 (N_2217,In_2489,In_2052);
nand U2218 (N_2218,In_1178,In_212);
nand U2219 (N_2219,In_812,In_1354);
or U2220 (N_2220,In_647,In_1527);
and U2221 (N_2221,In_832,In_1941);
nor U2222 (N_2222,In_2248,In_2377);
xor U2223 (N_2223,In_2017,In_450);
nor U2224 (N_2224,In_481,In_188);
nand U2225 (N_2225,In_2472,In_1628);
and U2226 (N_2226,In_487,In_2364);
nor U2227 (N_2227,In_663,In_1199);
and U2228 (N_2228,In_1533,In_694);
xnor U2229 (N_2229,In_2007,In_908);
and U2230 (N_2230,In_215,In_1438);
nand U2231 (N_2231,In_526,In_1251);
nand U2232 (N_2232,In_919,In_1535);
nand U2233 (N_2233,In_927,In_81);
nor U2234 (N_2234,In_978,In_1931);
or U2235 (N_2235,In_2248,In_1687);
nand U2236 (N_2236,In_759,In_818);
nor U2237 (N_2237,In_195,In_2361);
and U2238 (N_2238,In_1421,In_1115);
or U2239 (N_2239,In_1591,In_407);
nor U2240 (N_2240,In_724,In_905);
or U2241 (N_2241,In_2346,In_717);
nand U2242 (N_2242,In_511,In_2089);
nor U2243 (N_2243,In_1820,In_901);
nor U2244 (N_2244,In_694,In_236);
nand U2245 (N_2245,In_1633,In_2036);
nand U2246 (N_2246,In_1263,In_1512);
and U2247 (N_2247,In_1465,In_665);
nor U2248 (N_2248,In_2102,In_2371);
nor U2249 (N_2249,In_1415,In_1558);
and U2250 (N_2250,In_1981,In_2381);
nand U2251 (N_2251,In_1827,In_1863);
or U2252 (N_2252,In_2377,In_1188);
or U2253 (N_2253,In_1766,In_593);
nor U2254 (N_2254,In_122,In_1036);
nor U2255 (N_2255,In_714,In_2177);
xor U2256 (N_2256,In_51,In_2239);
nor U2257 (N_2257,In_63,In_516);
or U2258 (N_2258,In_321,In_850);
xor U2259 (N_2259,In_2027,In_216);
xnor U2260 (N_2260,In_482,In_848);
nor U2261 (N_2261,In_1806,In_1301);
or U2262 (N_2262,In_1122,In_289);
xor U2263 (N_2263,In_1435,In_67);
or U2264 (N_2264,In_1526,In_1812);
and U2265 (N_2265,In_2408,In_871);
or U2266 (N_2266,In_1339,In_1692);
or U2267 (N_2267,In_1830,In_1339);
and U2268 (N_2268,In_859,In_2000);
nor U2269 (N_2269,In_786,In_583);
xor U2270 (N_2270,In_1272,In_1757);
nand U2271 (N_2271,In_821,In_737);
nor U2272 (N_2272,In_1816,In_2408);
or U2273 (N_2273,In_1731,In_777);
nor U2274 (N_2274,In_648,In_2088);
or U2275 (N_2275,In_1032,In_1197);
nor U2276 (N_2276,In_1358,In_1471);
nand U2277 (N_2277,In_2006,In_1138);
and U2278 (N_2278,In_1113,In_1628);
xor U2279 (N_2279,In_627,In_1466);
and U2280 (N_2280,In_1927,In_643);
and U2281 (N_2281,In_1406,In_2128);
or U2282 (N_2282,In_421,In_1588);
and U2283 (N_2283,In_2121,In_2153);
xor U2284 (N_2284,In_888,In_404);
or U2285 (N_2285,In_1707,In_2154);
nor U2286 (N_2286,In_563,In_1033);
nor U2287 (N_2287,In_2449,In_808);
and U2288 (N_2288,In_1184,In_1076);
nor U2289 (N_2289,In_940,In_1456);
or U2290 (N_2290,In_1811,In_1885);
nand U2291 (N_2291,In_1900,In_880);
and U2292 (N_2292,In_692,In_2256);
and U2293 (N_2293,In_416,In_1292);
nand U2294 (N_2294,In_1526,In_2127);
or U2295 (N_2295,In_2424,In_1938);
or U2296 (N_2296,In_1793,In_1979);
or U2297 (N_2297,In_2042,In_1337);
or U2298 (N_2298,In_331,In_673);
and U2299 (N_2299,In_280,In_1302);
and U2300 (N_2300,In_1120,In_1626);
xnor U2301 (N_2301,In_1514,In_334);
nand U2302 (N_2302,In_1575,In_699);
nor U2303 (N_2303,In_349,In_359);
nor U2304 (N_2304,In_592,In_2085);
and U2305 (N_2305,In_1572,In_923);
nand U2306 (N_2306,In_677,In_1555);
nor U2307 (N_2307,In_1709,In_2091);
and U2308 (N_2308,In_259,In_977);
nand U2309 (N_2309,In_2243,In_878);
and U2310 (N_2310,In_2129,In_515);
nor U2311 (N_2311,In_2382,In_1655);
nor U2312 (N_2312,In_1517,In_1861);
and U2313 (N_2313,In_2257,In_763);
or U2314 (N_2314,In_955,In_1638);
or U2315 (N_2315,In_2107,In_966);
nor U2316 (N_2316,In_958,In_1297);
xnor U2317 (N_2317,In_1612,In_463);
xor U2318 (N_2318,In_1030,In_1962);
and U2319 (N_2319,In_1576,In_211);
nand U2320 (N_2320,In_918,In_1196);
or U2321 (N_2321,In_79,In_1992);
xor U2322 (N_2322,In_1653,In_2300);
nand U2323 (N_2323,In_1071,In_808);
nand U2324 (N_2324,In_2155,In_863);
nor U2325 (N_2325,In_331,In_942);
and U2326 (N_2326,In_2230,In_1007);
nor U2327 (N_2327,In_1416,In_1410);
nand U2328 (N_2328,In_356,In_2402);
and U2329 (N_2329,In_222,In_1176);
or U2330 (N_2330,In_1015,In_764);
and U2331 (N_2331,In_2468,In_1321);
and U2332 (N_2332,In_1684,In_1919);
xor U2333 (N_2333,In_1892,In_1437);
nand U2334 (N_2334,In_1690,In_2474);
and U2335 (N_2335,In_588,In_2494);
and U2336 (N_2336,In_2109,In_1061);
nand U2337 (N_2337,In_347,In_1342);
nand U2338 (N_2338,In_1518,In_2091);
xnor U2339 (N_2339,In_638,In_880);
xnor U2340 (N_2340,In_1006,In_1761);
nand U2341 (N_2341,In_1394,In_2366);
xor U2342 (N_2342,In_179,In_1401);
nor U2343 (N_2343,In_1372,In_479);
nor U2344 (N_2344,In_1098,In_1541);
nand U2345 (N_2345,In_2462,In_1582);
nor U2346 (N_2346,In_976,In_2050);
nand U2347 (N_2347,In_2046,In_124);
xor U2348 (N_2348,In_299,In_1694);
and U2349 (N_2349,In_926,In_1925);
xnor U2350 (N_2350,In_2464,In_836);
xnor U2351 (N_2351,In_1829,In_122);
or U2352 (N_2352,In_1281,In_1870);
and U2353 (N_2353,In_783,In_1867);
or U2354 (N_2354,In_1720,In_1291);
or U2355 (N_2355,In_356,In_2087);
and U2356 (N_2356,In_368,In_1178);
and U2357 (N_2357,In_468,In_1191);
nand U2358 (N_2358,In_1486,In_344);
xnor U2359 (N_2359,In_1024,In_593);
nor U2360 (N_2360,In_1202,In_1993);
nor U2361 (N_2361,In_641,In_1699);
nand U2362 (N_2362,In_21,In_138);
and U2363 (N_2363,In_78,In_668);
xnor U2364 (N_2364,In_2061,In_58);
and U2365 (N_2365,In_1103,In_308);
nor U2366 (N_2366,In_1799,In_199);
and U2367 (N_2367,In_1109,In_2430);
nand U2368 (N_2368,In_884,In_730);
nor U2369 (N_2369,In_148,In_2419);
nand U2370 (N_2370,In_758,In_501);
or U2371 (N_2371,In_1662,In_404);
or U2372 (N_2372,In_793,In_966);
nand U2373 (N_2373,In_1011,In_1651);
nor U2374 (N_2374,In_745,In_327);
nor U2375 (N_2375,In_434,In_477);
and U2376 (N_2376,In_1918,In_1530);
nor U2377 (N_2377,In_228,In_914);
nand U2378 (N_2378,In_1222,In_1789);
nor U2379 (N_2379,In_445,In_1867);
nor U2380 (N_2380,In_1947,In_1166);
or U2381 (N_2381,In_1405,In_1583);
nor U2382 (N_2382,In_1698,In_204);
nor U2383 (N_2383,In_1659,In_1115);
or U2384 (N_2384,In_247,In_966);
nand U2385 (N_2385,In_253,In_1586);
xnor U2386 (N_2386,In_2218,In_1873);
nand U2387 (N_2387,In_2461,In_1202);
nor U2388 (N_2388,In_899,In_804);
nand U2389 (N_2389,In_390,In_1408);
nor U2390 (N_2390,In_1223,In_493);
and U2391 (N_2391,In_466,In_2430);
nor U2392 (N_2392,In_1320,In_1840);
nand U2393 (N_2393,In_1000,In_497);
and U2394 (N_2394,In_48,In_2014);
xor U2395 (N_2395,In_1466,In_1854);
nor U2396 (N_2396,In_685,In_2093);
and U2397 (N_2397,In_2242,In_1677);
nand U2398 (N_2398,In_468,In_1689);
xor U2399 (N_2399,In_561,In_713);
xor U2400 (N_2400,In_2406,In_2071);
xor U2401 (N_2401,In_604,In_2495);
nor U2402 (N_2402,In_704,In_318);
or U2403 (N_2403,In_2201,In_1884);
xnor U2404 (N_2404,In_1055,In_1913);
xnor U2405 (N_2405,In_2271,In_2330);
xnor U2406 (N_2406,In_1088,In_1154);
xnor U2407 (N_2407,In_952,In_1266);
nand U2408 (N_2408,In_1874,In_82);
xor U2409 (N_2409,In_261,In_920);
xor U2410 (N_2410,In_109,In_2467);
and U2411 (N_2411,In_1828,In_1193);
xor U2412 (N_2412,In_39,In_417);
nor U2413 (N_2413,In_1337,In_2310);
xor U2414 (N_2414,In_1505,In_670);
or U2415 (N_2415,In_886,In_2394);
and U2416 (N_2416,In_1614,In_734);
nand U2417 (N_2417,In_182,In_575);
nand U2418 (N_2418,In_185,In_2062);
and U2419 (N_2419,In_1704,In_2126);
or U2420 (N_2420,In_1669,In_409);
and U2421 (N_2421,In_626,In_285);
or U2422 (N_2422,In_2339,In_1569);
or U2423 (N_2423,In_1008,In_534);
nor U2424 (N_2424,In_383,In_2215);
and U2425 (N_2425,In_475,In_61);
and U2426 (N_2426,In_913,In_1246);
nand U2427 (N_2427,In_1770,In_2077);
nand U2428 (N_2428,In_1247,In_400);
xnor U2429 (N_2429,In_98,In_1809);
xnor U2430 (N_2430,In_1823,In_1619);
and U2431 (N_2431,In_2183,In_136);
nand U2432 (N_2432,In_1145,In_572);
xor U2433 (N_2433,In_1588,In_1940);
nor U2434 (N_2434,In_777,In_2024);
or U2435 (N_2435,In_134,In_542);
or U2436 (N_2436,In_153,In_2308);
xor U2437 (N_2437,In_1752,In_2406);
xor U2438 (N_2438,In_2385,In_1472);
nand U2439 (N_2439,In_192,In_1420);
xnor U2440 (N_2440,In_51,In_331);
nor U2441 (N_2441,In_1709,In_2357);
nor U2442 (N_2442,In_944,In_926);
and U2443 (N_2443,In_1858,In_115);
and U2444 (N_2444,In_101,In_1890);
nor U2445 (N_2445,In_1535,In_1830);
xor U2446 (N_2446,In_2448,In_674);
or U2447 (N_2447,In_2155,In_2336);
or U2448 (N_2448,In_2238,In_1864);
and U2449 (N_2449,In_29,In_298);
nand U2450 (N_2450,In_1379,In_1034);
nand U2451 (N_2451,In_1830,In_1815);
or U2452 (N_2452,In_2399,In_1291);
xor U2453 (N_2453,In_2104,In_1823);
and U2454 (N_2454,In_2396,In_1924);
or U2455 (N_2455,In_911,In_672);
and U2456 (N_2456,In_516,In_2108);
and U2457 (N_2457,In_1786,In_584);
xor U2458 (N_2458,In_1414,In_1469);
and U2459 (N_2459,In_157,In_2356);
nor U2460 (N_2460,In_16,In_1112);
xnor U2461 (N_2461,In_1138,In_1559);
or U2462 (N_2462,In_1522,In_452);
and U2463 (N_2463,In_561,In_1149);
nand U2464 (N_2464,In_1415,In_1073);
or U2465 (N_2465,In_2276,In_2484);
and U2466 (N_2466,In_1247,In_612);
nor U2467 (N_2467,In_1891,In_615);
nand U2468 (N_2468,In_544,In_137);
or U2469 (N_2469,In_1398,In_2041);
and U2470 (N_2470,In_1139,In_1956);
or U2471 (N_2471,In_1091,In_391);
nand U2472 (N_2472,In_1601,In_1920);
and U2473 (N_2473,In_2201,In_41);
and U2474 (N_2474,In_1874,In_2305);
and U2475 (N_2475,In_1572,In_802);
or U2476 (N_2476,In_2057,In_949);
and U2477 (N_2477,In_201,In_1405);
nor U2478 (N_2478,In_392,In_1446);
and U2479 (N_2479,In_2042,In_850);
nand U2480 (N_2480,In_637,In_327);
nor U2481 (N_2481,In_1927,In_498);
xnor U2482 (N_2482,In_820,In_818);
and U2483 (N_2483,In_1386,In_1053);
nand U2484 (N_2484,In_1163,In_1558);
and U2485 (N_2485,In_1891,In_1418);
xor U2486 (N_2486,In_2204,In_1299);
xor U2487 (N_2487,In_2144,In_125);
xnor U2488 (N_2488,In_1877,In_1239);
or U2489 (N_2489,In_822,In_2383);
or U2490 (N_2490,In_1388,In_2041);
or U2491 (N_2491,In_2044,In_2354);
or U2492 (N_2492,In_916,In_140);
nand U2493 (N_2493,In_1467,In_1772);
nand U2494 (N_2494,In_2042,In_988);
nor U2495 (N_2495,In_931,In_296);
or U2496 (N_2496,In_2124,In_2054);
xnor U2497 (N_2497,In_962,In_889);
or U2498 (N_2498,In_977,In_2437);
and U2499 (N_2499,In_1350,In_2249);
or U2500 (N_2500,N_861,N_132);
nand U2501 (N_2501,N_1262,N_131);
nor U2502 (N_2502,N_659,N_1221);
xor U2503 (N_2503,N_2000,N_612);
nand U2504 (N_2504,N_1548,N_190);
nand U2505 (N_2505,N_1187,N_1703);
nand U2506 (N_2506,N_1294,N_462);
and U2507 (N_2507,N_2181,N_472);
or U2508 (N_2508,N_370,N_1957);
nand U2509 (N_2509,N_2058,N_389);
nand U2510 (N_2510,N_553,N_1227);
and U2511 (N_2511,N_1580,N_14);
nand U2512 (N_2512,N_195,N_308);
or U2513 (N_2513,N_499,N_1357);
or U2514 (N_2514,N_873,N_558);
nor U2515 (N_2515,N_885,N_2005);
nand U2516 (N_2516,N_2300,N_739);
xor U2517 (N_2517,N_1329,N_2362);
xor U2518 (N_2518,N_1612,N_2432);
xor U2519 (N_2519,N_1488,N_2187);
and U2520 (N_2520,N_563,N_1610);
or U2521 (N_2521,N_853,N_97);
nand U2522 (N_2522,N_762,N_653);
nor U2523 (N_2523,N_2,N_2280);
xnor U2524 (N_2524,N_1983,N_851);
or U2525 (N_2525,N_1729,N_2207);
xnor U2526 (N_2526,N_706,N_1731);
xnor U2527 (N_2527,N_1020,N_2335);
or U2528 (N_2528,N_1785,N_1219);
or U2529 (N_2529,N_2373,N_1486);
and U2530 (N_2530,N_928,N_1318);
nand U2531 (N_2531,N_1069,N_1196);
nand U2532 (N_2532,N_2338,N_382);
nor U2533 (N_2533,N_2385,N_1477);
and U2534 (N_2534,N_1896,N_108);
xnor U2535 (N_2535,N_1209,N_1953);
nor U2536 (N_2536,N_650,N_1251);
nand U2537 (N_2537,N_1324,N_1579);
and U2538 (N_2538,N_1934,N_2471);
or U2539 (N_2539,N_833,N_2415);
and U2540 (N_2540,N_465,N_2081);
or U2541 (N_2541,N_2480,N_198);
and U2542 (N_2542,N_1977,N_2115);
xor U2543 (N_2543,N_275,N_2424);
or U2544 (N_2544,N_1623,N_779);
nor U2545 (N_2545,N_997,N_1675);
and U2546 (N_2546,N_719,N_1239);
xnor U2547 (N_2547,N_60,N_1875);
xor U2548 (N_2548,N_317,N_1427);
or U2549 (N_2549,N_19,N_576);
and U2550 (N_2550,N_2410,N_1720);
xor U2551 (N_2551,N_404,N_2124);
nand U2552 (N_2552,N_2093,N_333);
nor U2553 (N_2553,N_749,N_575);
and U2554 (N_2554,N_2487,N_1863);
nand U2555 (N_2555,N_1442,N_1797);
and U2556 (N_2556,N_1871,N_2407);
nor U2557 (N_2557,N_1041,N_307);
nor U2558 (N_2558,N_713,N_2278);
or U2559 (N_2559,N_2245,N_524);
nor U2560 (N_2560,N_1824,N_1345);
nand U2561 (N_2561,N_1267,N_162);
nor U2562 (N_2562,N_792,N_663);
nand U2563 (N_2563,N_120,N_693);
or U2564 (N_2564,N_2165,N_1835);
xnor U2565 (N_2565,N_468,N_420);
or U2566 (N_2566,N_416,N_691);
nor U2567 (N_2567,N_1128,N_2073);
xor U2568 (N_2568,N_2046,N_822);
nor U2569 (N_2569,N_2074,N_2337);
xor U2570 (N_2570,N_996,N_1599);
nor U2571 (N_2571,N_2412,N_654);
nor U2572 (N_2572,N_365,N_2399);
nor U2573 (N_2573,N_805,N_116);
xor U2574 (N_2574,N_1667,N_388);
or U2575 (N_2575,N_1012,N_585);
nor U2576 (N_2576,N_734,N_1154);
xor U2577 (N_2577,N_874,N_572);
xnor U2578 (N_2578,N_1420,N_1100);
and U2579 (N_2579,N_1887,N_2052);
or U2580 (N_2580,N_2273,N_1003);
and U2581 (N_2581,N_989,N_1894);
and U2582 (N_2582,N_634,N_2376);
xnor U2583 (N_2583,N_2473,N_1690);
nor U2584 (N_2584,N_1560,N_0);
nand U2585 (N_2585,N_1382,N_1350);
or U2586 (N_2586,N_737,N_90);
nor U2587 (N_2587,N_398,N_770);
and U2588 (N_2588,N_1657,N_1862);
nand U2589 (N_2589,N_1163,N_574);
or U2590 (N_2590,N_1431,N_2174);
xor U2591 (N_2591,N_1426,N_126);
nand U2592 (N_2592,N_1047,N_1143);
and U2593 (N_2593,N_754,N_1320);
nand U2594 (N_2594,N_1620,N_2164);
nor U2595 (N_2595,N_1445,N_973);
and U2596 (N_2596,N_661,N_1592);
nand U2597 (N_2597,N_64,N_1521);
xor U2598 (N_2598,N_2214,N_1578);
nand U2599 (N_2599,N_1259,N_2226);
or U2600 (N_2600,N_474,N_497);
xor U2601 (N_2601,N_795,N_252);
nand U2602 (N_2602,N_1884,N_871);
nor U2603 (N_2603,N_1590,N_1528);
and U2604 (N_2604,N_1997,N_633);
and U2605 (N_2605,N_1039,N_1421);
nand U2606 (N_2606,N_2258,N_456);
nor U2607 (N_2607,N_1473,N_1091);
nor U2608 (N_2608,N_20,N_1790);
xor U2609 (N_2609,N_61,N_1561);
nand U2610 (N_2610,N_1933,N_1389);
and U2611 (N_2611,N_1193,N_1409);
and U2612 (N_2612,N_199,N_2326);
xor U2613 (N_2613,N_1479,N_1302);
nor U2614 (N_2614,N_1805,N_1954);
nor U2615 (N_2615,N_865,N_1391);
nor U2616 (N_2616,N_110,N_710);
or U2617 (N_2617,N_1168,N_2215);
nand U2618 (N_2618,N_1857,N_729);
and U2619 (N_2619,N_1822,N_1809);
and U2620 (N_2620,N_1016,N_2088);
and U2621 (N_2621,N_1996,N_2201);
nor U2622 (N_2622,N_615,N_945);
or U2623 (N_2623,N_2106,N_1352);
and U2624 (N_2624,N_148,N_1723);
or U2625 (N_2625,N_2315,N_1757);
nand U2626 (N_2626,N_2481,N_2395);
xnor U2627 (N_2627,N_1874,N_902);
or U2628 (N_2628,N_230,N_67);
or U2629 (N_2629,N_1543,N_915);
nor U2630 (N_2630,N_2220,N_2314);
nor U2631 (N_2631,N_2168,N_2047);
nand U2632 (N_2632,N_900,N_522);
xor U2633 (N_2633,N_1107,N_1779);
nand U2634 (N_2634,N_2072,N_239);
and U2635 (N_2635,N_1721,N_1718);
or U2636 (N_2636,N_1717,N_1183);
nand U2637 (N_2637,N_2411,N_590);
or U2638 (N_2638,N_30,N_500);
nor U2639 (N_2639,N_1529,N_123);
and U2640 (N_2640,N_243,N_2234);
xor U2641 (N_2641,N_545,N_2430);
and U2642 (N_2642,N_769,N_1913);
or U2643 (N_2643,N_1413,N_431);
and U2644 (N_2644,N_2116,N_1719);
nor U2645 (N_2645,N_2425,N_2062);
and U2646 (N_2646,N_1945,N_430);
or U2647 (N_2647,N_1429,N_104);
and U2648 (N_2648,N_2382,N_886);
nand U2649 (N_2649,N_877,N_670);
nand U2650 (N_2650,N_1565,N_1402);
and U2651 (N_2651,N_514,N_507);
nor U2652 (N_2652,N_2217,N_1990);
nand U2653 (N_2653,N_1353,N_668);
and U2654 (N_2654,N_56,N_2331);
or U2655 (N_2655,N_2169,N_820);
and U2656 (N_2656,N_10,N_1748);
or U2657 (N_2657,N_422,N_2344);
xnor U2658 (N_2658,N_1906,N_2449);
xnor U2659 (N_2659,N_2292,N_1938);
and U2660 (N_2660,N_2244,N_1483);
and U2661 (N_2661,N_28,N_1085);
or U2662 (N_2662,N_1129,N_1813);
or U2663 (N_2663,N_893,N_2434);
nand U2664 (N_2664,N_251,N_1727);
nand U2665 (N_2665,N_2299,N_1393);
nand U2666 (N_2666,N_2405,N_147);
xnor U2667 (N_2667,N_1075,N_931);
nand U2668 (N_2668,N_2421,N_606);
and U2669 (N_2669,N_2444,N_1747);
nand U2670 (N_2670,N_1484,N_669);
nor U2671 (N_2671,N_712,N_926);
and U2672 (N_2672,N_1551,N_964);
and U2673 (N_2673,N_717,N_335);
nand U2674 (N_2674,N_642,N_635);
and U2675 (N_2675,N_1546,N_478);
xnor U2676 (N_2676,N_178,N_1585);
or U2677 (N_2677,N_351,N_340);
and U2678 (N_2678,N_1304,N_761);
xor U2679 (N_2679,N_2262,N_2077);
or U2680 (N_2680,N_1760,N_2135);
nand U2681 (N_2681,N_735,N_2184);
and U2682 (N_2682,N_1705,N_2084);
or U2683 (N_2683,N_1013,N_2064);
or U2684 (N_2684,N_1433,N_2166);
or U2685 (N_2685,N_1698,N_2018);
nor U2686 (N_2686,N_616,N_1365);
nand U2687 (N_2687,N_1078,N_1342);
nor U2688 (N_2688,N_1347,N_971);
and U2689 (N_2689,N_350,N_1908);
or U2690 (N_2690,N_912,N_1632);
and U2691 (N_2691,N_2040,N_1313);
and U2692 (N_2692,N_714,N_825);
nand U2693 (N_2693,N_878,N_1914);
nand U2694 (N_2694,N_2371,N_1234);
and U2695 (N_2695,N_904,N_818);
nand U2696 (N_2696,N_667,N_589);
and U2697 (N_2697,N_1388,N_1334);
nor U2698 (N_2698,N_358,N_1138);
xor U2699 (N_2699,N_791,N_968);
nor U2700 (N_2700,N_1146,N_867);
nand U2701 (N_2701,N_1197,N_262);
nor U2702 (N_2702,N_1192,N_184);
and U2703 (N_2703,N_1072,N_1279);
nand U2704 (N_2704,N_1820,N_1216);
nor U2705 (N_2705,N_1394,N_2205);
or U2706 (N_2706,N_1186,N_1097);
xor U2707 (N_2707,N_341,N_677);
or U2708 (N_2708,N_1586,N_1935);
and U2709 (N_2709,N_1542,N_329);
nor U2710 (N_2710,N_1090,N_803);
xor U2711 (N_2711,N_1976,N_344);
and U2712 (N_2712,N_773,N_1205);
nand U2713 (N_2713,N_1482,N_2178);
and U2714 (N_2714,N_146,N_2329);
xnor U2715 (N_2715,N_119,N_527);
nor U2716 (N_2716,N_1450,N_1001);
xor U2717 (N_2717,N_751,N_1384);
and U2718 (N_2718,N_196,N_1801);
xnor U2719 (N_2719,N_1988,N_399);
and U2720 (N_2720,N_785,N_2409);
nor U2721 (N_2721,N_1792,N_994);
and U2722 (N_2722,N_1504,N_1510);
and U2723 (N_2723,N_2218,N_582);
nor U2724 (N_2724,N_2422,N_2130);
nand U2725 (N_2725,N_1301,N_555);
nor U2726 (N_2726,N_1787,N_2119);
nand U2727 (N_2727,N_356,N_854);
xor U2728 (N_2728,N_1812,N_46);
nand U2729 (N_2729,N_1856,N_1463);
nand U2730 (N_2730,N_1086,N_2283);
nor U2731 (N_2731,N_2206,N_657);
or U2732 (N_2732,N_709,N_1271);
nor U2733 (N_2733,N_1866,N_213);
and U2734 (N_2734,N_2039,N_766);
or U2735 (N_2735,N_927,N_629);
xor U2736 (N_2736,N_1541,N_2398);
nand U2737 (N_2737,N_730,N_1826);
or U2738 (N_2738,N_1722,N_2388);
and U2739 (N_2739,N_1103,N_2241);
or U2740 (N_2740,N_1702,N_45);
and U2741 (N_2741,N_2157,N_2374);
and U2742 (N_2742,N_1277,N_982);
or U2743 (N_2743,N_1597,N_2347);
or U2744 (N_2744,N_911,N_1923);
or U2745 (N_2745,N_917,N_2360);
or U2746 (N_2746,N_174,N_492);
or U2747 (N_2747,N_2033,N_1540);
and U2748 (N_2748,N_139,N_1607);
and U2749 (N_2749,N_1700,N_393);
or U2750 (N_2750,N_2054,N_1199);
nor U2751 (N_2751,N_491,N_66);
or U2752 (N_2752,N_1877,N_725);
or U2753 (N_2753,N_2287,N_71);
and U2754 (N_2754,N_1535,N_494);
nor U2755 (N_2755,N_2276,N_530);
nand U2756 (N_2756,N_1371,N_1293);
and U2757 (N_2757,N_2308,N_96);
and U2758 (N_2758,N_658,N_421);
xor U2759 (N_2759,N_620,N_306);
and U2760 (N_2760,N_81,N_1872);
or U2761 (N_2761,N_1788,N_441);
nand U2762 (N_2762,N_1740,N_540);
nor U2763 (N_2763,N_2336,N_2332);
and U2764 (N_2764,N_1596,N_2488);
nand U2765 (N_2765,N_2389,N_2490);
nor U2766 (N_2766,N_1410,N_1485);
xnor U2767 (N_2767,N_2423,N_726);
nand U2768 (N_2768,N_415,N_951);
or U2769 (N_2769,N_345,N_488);
nand U2770 (N_2770,N_1766,N_36);
and U2771 (N_2771,N_1400,N_1613);
or U2772 (N_2772,N_1156,N_1270);
or U2773 (N_2773,N_2357,N_984);
or U2774 (N_2774,N_316,N_1245);
or U2775 (N_2775,N_619,N_380);
nor U2776 (N_2776,N_1967,N_1307);
and U2777 (N_2777,N_1306,N_1349);
xor U2778 (N_2778,N_1194,N_767);
nor U2779 (N_2779,N_2167,N_2153);
nand U2780 (N_2780,N_1272,N_798);
or U2781 (N_2781,N_817,N_1099);
or U2782 (N_2782,N_1182,N_1140);
and U2783 (N_2783,N_1108,N_286);
nand U2784 (N_2784,N_839,N_932);
xor U2785 (N_2785,N_609,N_1115);
and U2786 (N_2786,N_1157,N_1358);
or U2787 (N_2787,N_477,N_1452);
xor U2788 (N_2788,N_281,N_211);
and U2789 (N_2789,N_695,N_357);
nand U2790 (N_2790,N_2274,N_602);
or U2791 (N_2791,N_68,N_684);
and U2792 (N_2792,N_2459,N_1855);
and U2793 (N_2793,N_549,N_1033);
nor U2794 (N_2794,N_2464,N_2312);
nor U2795 (N_2795,N_1584,N_896);
nor U2796 (N_2796,N_1767,N_1195);
nand U2797 (N_2797,N_2354,N_674);
nor U2798 (N_2798,N_1474,N_276);
xor U2799 (N_2799,N_1074,N_1124);
nand U2800 (N_2800,N_2105,N_2003);
nor U2801 (N_2801,N_2392,N_976);
xnor U2802 (N_2802,N_637,N_2125);
or U2803 (N_2803,N_581,N_122);
or U2804 (N_2804,N_63,N_151);
nor U2805 (N_2805,N_1985,N_2061);
nor U2806 (N_2806,N_1122,N_269);
nand U2807 (N_2807,N_1654,N_274);
xor U2808 (N_2808,N_740,N_1455);
nand U2809 (N_2809,N_1806,N_2247);
and U2810 (N_2810,N_93,N_1849);
nor U2811 (N_2811,N_806,N_840);
and U2812 (N_2812,N_566,N_2393);
xor U2813 (N_2813,N_2253,N_191);
nand U2814 (N_2814,N_107,N_1517);
xnor U2815 (N_2815,N_1598,N_1110);
and U2816 (N_2816,N_1519,N_137);
and U2817 (N_2817,N_2295,N_2243);
and U2818 (N_2818,N_1763,N_2024);
xnor U2819 (N_2819,N_1786,N_387);
or U2820 (N_2820,N_1575,N_2212);
xor U2821 (N_2821,N_2366,N_1602);
nor U2822 (N_2822,N_1252,N_259);
or U2823 (N_2823,N_2067,N_2097);
or U2824 (N_2824,N_2351,N_12);
or U2825 (N_2825,N_2460,N_2390);
and U2826 (N_2826,N_1776,N_2325);
nand U2827 (N_2827,N_809,N_2078);
xnor U2828 (N_2828,N_1113,N_630);
nor U2829 (N_2829,N_470,N_149);
or U2830 (N_2830,N_167,N_424);
xor U2831 (N_2831,N_58,N_1066);
nand U2832 (N_2832,N_1040,N_1537);
nand U2833 (N_2833,N_44,N_1478);
xnor U2834 (N_2834,N_417,N_807);
xor U2835 (N_2835,N_517,N_177);
xnor U2836 (N_2836,N_2196,N_1764);
xnor U2837 (N_2837,N_1018,N_1716);
nand U2838 (N_2838,N_1774,N_999);
nand U2839 (N_2839,N_1472,N_843);
nand U2840 (N_2840,N_686,N_91);
and U2841 (N_2841,N_1782,N_1803);
or U2842 (N_2842,N_1002,N_2118);
nand U2843 (N_2843,N_310,N_2445);
nor U2844 (N_2844,N_445,N_1768);
nor U2845 (N_2845,N_1116,N_336);
nand U2846 (N_2846,N_662,N_1593);
nor U2847 (N_2847,N_2457,N_1924);
nor U2848 (N_2848,N_2177,N_949);
nor U2849 (N_2849,N_1512,N_1637);
or U2850 (N_2850,N_2059,N_1708);
nor U2851 (N_2851,N_1925,N_300);
nor U2852 (N_2852,N_1201,N_856);
xnor U2853 (N_2853,N_1907,N_881);
nand U2854 (N_2854,N_249,N_437);
xor U2855 (N_2855,N_1754,N_34);
nand U2856 (N_2856,N_1694,N_1443);
nor U2857 (N_2857,N_614,N_23);
xnor U2858 (N_2858,N_1978,N_220);
and U2859 (N_2859,N_1715,N_988);
nor U2860 (N_2860,N_763,N_1589);
or U2861 (N_2861,N_2497,N_1340);
and U2862 (N_2862,N_322,N_83);
and U2863 (N_2863,N_694,N_359);
nand U2864 (N_2864,N_1995,N_1266);
nor U2865 (N_2865,N_2305,N_1980);
nand U2866 (N_2866,N_2045,N_1462);
and U2867 (N_2867,N_2396,N_479);
xnor U2868 (N_2868,N_2296,N_485);
xor U2869 (N_2869,N_2453,N_2346);
and U2870 (N_2870,N_1035,N_1022);
nor U2871 (N_2871,N_202,N_930);
xnor U2872 (N_2872,N_1366,N_112);
or U2873 (N_2873,N_2259,N_2266);
or U2874 (N_2874,N_921,N_745);
xnor U2875 (N_2875,N_1556,N_774);
nor U2876 (N_2876,N_1775,N_1498);
nor U2877 (N_2877,N_432,N_849);
nand U2878 (N_2878,N_2397,N_1330);
and U2879 (N_2879,N_743,N_13);
or U2880 (N_2880,N_117,N_205);
xor U2881 (N_2881,N_2448,N_1397);
and U2882 (N_2882,N_1756,N_24);
or U2883 (N_2883,N_1361,N_2420);
or U2884 (N_2884,N_458,N_114);
nand U2885 (N_2885,N_888,N_223);
xor U2886 (N_2886,N_100,N_1215);
xnor U2887 (N_2887,N_1164,N_1525);
nand U2888 (N_2888,N_1026,N_780);
or U2889 (N_2889,N_969,N_2086);
xor U2890 (N_2890,N_511,N_229);
and U2891 (N_2891,N_1253,N_2092);
and U2892 (N_2892,N_521,N_2144);
and U2893 (N_2893,N_1360,N_1633);
nor U2894 (N_2894,N_154,N_2239);
or U2895 (N_2895,N_2009,N_295);
or U2896 (N_2896,N_1846,N_1112);
xor U2897 (N_2897,N_1550,N_1656);
or U2898 (N_2898,N_938,N_2185);
xnor U2899 (N_2899,N_510,N_1832);
nor U2900 (N_2900,N_1847,N_789);
or U2901 (N_2901,N_315,N_385);
and U2902 (N_2902,N_2051,N_1819);
nor U2903 (N_2903,N_652,N_238);
or U2904 (N_2904,N_675,N_161);
or U2905 (N_2905,N_876,N_1618);
or U2906 (N_2906,N_1506,N_179);
nor U2907 (N_2907,N_11,N_1710);
and U2908 (N_2908,N_1966,N_537);
or U2909 (N_2909,N_1870,N_1346);
nor U2910 (N_2910,N_292,N_1761);
and U2911 (N_2911,N_1594,N_369);
nor U2912 (N_2912,N_444,N_1791);
and U2913 (N_2913,N_554,N_1059);
xor U2914 (N_2914,N_2343,N_1333);
nand U2915 (N_2915,N_2137,N_594);
or U2916 (N_2916,N_665,N_2189);
and U2917 (N_2917,N_1858,N_1029);
xor U2918 (N_2918,N_1897,N_194);
nand U2919 (N_2919,N_918,N_80);
nor U2920 (N_2920,N_1929,N_435);
and U2921 (N_2921,N_42,N_2282);
nor U2922 (N_2922,N_425,N_810);
or U2923 (N_2923,N_811,N_486);
and U2924 (N_2924,N_1595,N_692);
xnor U2925 (N_2925,N_2200,N_2013);
nor U2926 (N_2926,N_1601,N_848);
or U2927 (N_2927,N_82,N_1886);
nand U2928 (N_2928,N_1885,N_349);
nand U2929 (N_2929,N_1379,N_1475);
nor U2930 (N_2930,N_883,N_859);
or U2931 (N_2931,N_2002,N_2489);
xor U2932 (N_2932,N_940,N_1403);
xor U2933 (N_2933,N_1689,N_852);
or U2934 (N_2934,N_623,N_1899);
and U2935 (N_2935,N_272,N_2483);
xnor U2936 (N_2936,N_101,N_1674);
and U2937 (N_2937,N_2136,N_1987);
nor U2938 (N_2938,N_1359,N_450);
nor U2939 (N_2939,N_189,N_2152);
and U2940 (N_2940,N_1777,N_962);
nor U2941 (N_2941,N_498,N_2203);
nor U2942 (N_2942,N_323,N_1328);
or U2943 (N_2943,N_879,N_1276);
nor U2944 (N_2944,N_2228,N_624);
or U2945 (N_2945,N_1701,N_1821);
and U2946 (N_2946,N_1123,N_1448);
and U2947 (N_2947,N_1404,N_704);
or U2948 (N_2948,N_2307,N_1971);
nor U2949 (N_2949,N_846,N_1299);
and U2950 (N_2950,N_218,N_1557);
nor U2951 (N_2951,N_1481,N_1514);
nand U2952 (N_2952,N_2080,N_588);
xor U2953 (N_2953,N_2378,N_1172);
and U2954 (N_2954,N_1332,N_1067);
nand U2955 (N_2955,N_533,N_1152);
xnor U2956 (N_2956,N_1362,N_406);
and U2957 (N_2957,N_504,N_482);
nand U2958 (N_2958,N_1982,N_1920);
xor U2959 (N_2959,N_52,N_7);
or U2960 (N_2960,N_2289,N_831);
or U2961 (N_2961,N_1335,N_2145);
xnor U2962 (N_2962,N_875,N_2345);
nor U2963 (N_2963,N_1453,N_1456);
or U2964 (N_2964,N_2069,N_2204);
xnor U2965 (N_2965,N_1214,N_1852);
and U2966 (N_2966,N_844,N_1770);
xor U2967 (N_2967,N_2339,N_2493);
and U2968 (N_2968,N_1738,N_1843);
nand U2969 (N_2969,N_453,N_1895);
xor U2970 (N_2970,N_1261,N_375);
xnor U2971 (N_2971,N_1068,N_919);
nor U2972 (N_2972,N_397,N_815);
nand U2973 (N_2973,N_643,N_983);
or U2974 (N_2974,N_1077,N_1696);
or U2975 (N_2975,N_707,N_72);
nand U2976 (N_2976,N_475,N_1850);
nor U2977 (N_2977,N_2414,N_682);
or U2978 (N_2978,N_1080,N_133);
nor U2979 (N_2979,N_1208,N_1600);
and U2980 (N_2980,N_1502,N_22);
and U2981 (N_2981,N_1203,N_860);
xor U2982 (N_2982,N_2242,N_2330);
xnor U2983 (N_2983,N_438,N_1531);
and U2984 (N_2984,N_2147,N_604);
xnor U2985 (N_2985,N_887,N_2049);
nand U2986 (N_2986,N_105,N_207);
nor U2987 (N_2987,N_1231,N_1118);
and U2988 (N_2988,N_2163,N_1869);
nor U2989 (N_2989,N_950,N_1395);
or U2990 (N_2990,N_1975,N_1052);
and U2991 (N_2991,N_1892,N_1962);
and U2992 (N_2992,N_1523,N_138);
or U2993 (N_2993,N_1109,N_366);
nor U2994 (N_2994,N_1750,N_666);
or U2995 (N_2995,N_1538,N_2462);
or U2996 (N_2996,N_1730,N_2149);
nor U2997 (N_2997,N_639,N_640);
and U2998 (N_2998,N_50,N_1651);
nor U2999 (N_2999,N_2446,N_1247);
xnor U3000 (N_3000,N_2031,N_715);
nor U3001 (N_3001,N_1338,N_1746);
nand U3002 (N_3002,N_760,N_1286);
xnor U3003 (N_3003,N_247,N_2450);
nor U3004 (N_3004,N_1693,N_1237);
nand U3005 (N_3005,N_413,N_625);
nor U3006 (N_3006,N_2456,N_1513);
nor U3007 (N_3007,N_234,N_257);
and U3008 (N_3008,N_142,N_449);
xor U3009 (N_3009,N_1739,N_1348);
xnor U3010 (N_3010,N_1867,N_1762);
or U3011 (N_3011,N_644,N_1631);
and U3012 (N_3012,N_1626,N_1105);
nor U3013 (N_3013,N_2479,N_121);
nor U3014 (N_3014,N_1881,N_2126);
xnor U3015 (N_3015,N_565,N_216);
nor U3016 (N_3016,N_1058,N_483);
xor U3017 (N_3017,N_987,N_1179);
nand U3018 (N_3018,N_232,N_2286);
and U3019 (N_3019,N_363,N_1981);
nor U3020 (N_3020,N_689,N_1202);
xor U3021 (N_3021,N_319,N_1210);
or U3022 (N_3022,N_1783,N_2035);
xor U3023 (N_3023,N_2478,N_250);
nand U3024 (N_3024,N_1414,N_1518);
and U3025 (N_3025,N_1860,N_1225);
nand U3026 (N_3026,N_2380,N_1622);
and U3027 (N_3027,N_2291,N_991);
xnor U3028 (N_3028,N_35,N_2317);
xnor U3029 (N_3029,N_1744,N_778);
nand U3030 (N_3030,N_1679,N_1131);
nand U3031 (N_3031,N_183,N_1060);
and U3032 (N_3032,N_1950,N_957);
or U3033 (N_3033,N_872,N_1430);
and U3034 (N_3034,N_25,N_484);
xor U3035 (N_3035,N_970,N_1355);
nand U3036 (N_3036,N_2028,N_1369);
and U3037 (N_3037,N_501,N_1628);
or U3038 (N_3038,N_1851,N_2154);
and U3039 (N_3039,N_1755,N_793);
and U3040 (N_3040,N_2436,N_2441);
or U3041 (N_3041,N_277,N_2491);
or U3042 (N_3042,N_1439,N_960);
nand U3043 (N_3043,N_802,N_1605);
nand U3044 (N_3044,N_1255,N_1217);
or U3045 (N_3045,N_797,N_318);
or U3046 (N_3046,N_587,N_2233);
nor U3047 (N_3047,N_583,N_1142);
nor U3048 (N_3048,N_747,N_1295);
or U3049 (N_3049,N_1804,N_1148);
and U3050 (N_3050,N_1284,N_512);
nand U3051 (N_3051,N_2094,N_312);
nand U3052 (N_3052,N_313,N_1532);
nand U3053 (N_3053,N_160,N_864);
nand U3054 (N_3054,N_1256,N_2375);
or U3055 (N_3055,N_1063,N_1969);
nor U3056 (N_3056,N_2285,N_870);
and U3057 (N_3057,N_1027,N_1555);
or U3058 (N_3058,N_1742,N_1998);
xnor U3059 (N_3059,N_1668,N_2363);
or U3060 (N_3060,N_1469,N_1932);
and U3061 (N_3061,N_943,N_242);
xnor U3062 (N_3062,N_722,N_157);
and U3063 (N_3063,N_1562,N_1511);
xor U3064 (N_3064,N_974,N_1931);
nor U3065 (N_3065,N_225,N_2120);
and U3066 (N_3066,N_1568,N_2038);
xnor U3067 (N_3067,N_2056,N_892);
or U3068 (N_3068,N_1454,N_2055);
or U3069 (N_3069,N_1042,N_520);
nand U3070 (N_3070,N_2469,N_244);
or U3071 (N_3071,N_434,N_2216);
nand U3072 (N_3072,N_2439,N_1683);
xnor U3073 (N_3073,N_1386,N_155);
and U3074 (N_3074,N_1960,N_235);
nor U3075 (N_3075,N_2350,N_571);
nor U3076 (N_3076,N_1970,N_1007);
nor U3077 (N_3077,N_279,N_776);
and U3078 (N_3078,N_1891,N_203);
nand U3079 (N_3079,N_2452,N_998);
nand U3080 (N_3080,N_342,N_828);
xnor U3081 (N_3081,N_2101,N_426);
nand U3082 (N_3082,N_2004,N_990);
and U3083 (N_3083,N_127,N_1515);
nor U3084 (N_3084,N_1554,N_1139);
nand U3085 (N_3085,N_925,N_143);
nand U3086 (N_3086,N_1162,N_2404);
xnor U3087 (N_3087,N_2316,N_518);
nand U3088 (N_3088,N_1930,N_2109);
nor U3089 (N_3089,N_1278,N_2255);
and U3090 (N_3090,N_1396,N_1212);
nor U3091 (N_3091,N_40,N_3);
or U3092 (N_3092,N_2176,N_1048);
nand U3093 (N_3093,N_1243,N_1501);
nand U3094 (N_3094,N_961,N_1282);
nand U3095 (N_3095,N_327,N_1645);
nor U3096 (N_3096,N_2387,N_2113);
xnor U3097 (N_3097,N_891,N_1178);
nor U3098 (N_3098,N_1520,N_2089);
nor U3099 (N_3099,N_86,N_2159);
or U3100 (N_3100,N_2034,N_1385);
nor U3101 (N_3101,N_941,N_1327);
nand U3102 (N_3102,N_361,N_608);
or U3103 (N_3103,N_1796,N_1544);
or U3104 (N_3104,N_43,N_1671);
nand U3105 (N_3105,N_2361,N_771);
or U3106 (N_3106,N_1435,N_1494);
or U3107 (N_3107,N_2463,N_1576);
or U3108 (N_3108,N_621,N_1949);
nand U3109 (N_3109,N_2194,N_1288);
nor U3110 (N_3110,N_1564,N_801);
or U3111 (N_3111,N_77,N_2408);
nor U3112 (N_3112,N_782,N_1161);
xnor U3113 (N_3113,N_1054,N_2377);
or U3114 (N_3114,N_1991,N_2138);
and U3115 (N_3115,N_1095,N_209);
xnor U3116 (N_3116,N_54,N_290);
nor U3117 (N_3117,N_464,N_718);
nand U3118 (N_3118,N_741,N_1180);
nand U3119 (N_3119,N_1526,N_738);
or U3120 (N_3120,N_897,N_1527);
or U3121 (N_3121,N_702,N_578);
nand U3122 (N_3122,N_1036,N_1876);
or U3123 (N_3123,N_386,N_145);
or U3124 (N_3124,N_1692,N_1370);
or U3125 (N_3125,N_955,N_993);
and U3126 (N_3126,N_282,N_1451);
xor U3127 (N_3127,N_436,N_1432);
xor U3128 (N_3128,N_680,N_1006);
nor U3129 (N_3129,N_2256,N_460);
and U3130 (N_3130,N_542,N_1190);
nand U3131 (N_3131,N_1171,N_226);
nor U3132 (N_3132,N_1354,N_302);
or U3133 (N_3133,N_2223,N_1132);
xor U3134 (N_3134,N_1670,N_463);
or U3135 (N_3135,N_1553,N_1942);
nand U3136 (N_3136,N_808,N_185);
and U3137 (N_3137,N_1664,N_200);
xor U3138 (N_3138,N_118,N_297);
and U3139 (N_3139,N_690,N_580);
nand U3140 (N_3140,N_1743,N_2341);
nand U3141 (N_3141,N_1629,N_2284);
nor U3142 (N_3142,N_2108,N_89);
nor U3143 (N_3143,N_2440,N_837);
xnor U3144 (N_3144,N_206,N_2248);
xor U3145 (N_3145,N_909,N_1558);
or U3146 (N_3146,N_69,N_1021);
and U3147 (N_3147,N_33,N_419);
nand U3148 (N_3148,N_2114,N_890);
xnor U3149 (N_3149,N_490,N_2006);
and U3150 (N_3150,N_134,N_1184);
nand U3151 (N_3151,N_2091,N_1476);
and U3152 (N_3152,N_503,N_2232);
xor U3153 (N_3153,N_1341,N_1699);
and U3154 (N_3154,N_409,N_1380);
and U3155 (N_3155,N_448,N_889);
nor U3156 (N_3156,N_2435,N_1024);
nor U3157 (N_3157,N_289,N_1713);
nor U3158 (N_3158,N_1311,N_1011);
and U3159 (N_3159,N_1901,N_836);
or U3160 (N_3160,N_172,N_32);
xnor U3161 (N_3161,N_688,N_2087);
nand U3162 (N_3162,N_480,N_2367);
and U3163 (N_3163,N_1459,N_1250);
or U3164 (N_3164,N_1968,N_2224);
or U3165 (N_3165,N_1559,N_1466);
nor U3166 (N_3166,N_459,N_1902);
and U3167 (N_3167,N_2447,N_2270);
nand U3168 (N_3168,N_2015,N_1649);
xnor U3169 (N_3169,N_433,N_2195);
or U3170 (N_3170,N_1010,N_561);
xor U3171 (N_3171,N_775,N_2027);
and U3172 (N_3172,N_1841,N_481);
nor U3173 (N_3173,N_2281,N_2155);
and U3174 (N_3174,N_1794,N_1368);
nor U3175 (N_3175,N_1467,N_1308);
and U3176 (N_3176,N_2349,N_1292);
nand U3177 (N_3177,N_595,N_2188);
and U3178 (N_3178,N_2269,N_320);
and U3179 (N_3179,N_2128,N_1312);
xnor U3180 (N_3180,N_539,N_1094);
nand U3181 (N_3181,N_2499,N_392);
xnor U3182 (N_3182,N_2288,N_1973);
nor U3183 (N_3183,N_2007,N_298);
or U3184 (N_3184,N_2182,N_1571);
nand U3185 (N_3185,N_212,N_402);
or U3186 (N_3186,N_827,N_2017);
or U3187 (N_3187,N_2229,N_2265);
nor U3188 (N_3188,N_379,N_2042);
or U3189 (N_3189,N_362,N_1229);
xor U3190 (N_3190,N_377,N_2193);
and U3191 (N_3191,N_1583,N_1223);
nand U3192 (N_3192,N_197,N_1480);
xor U3193 (N_3193,N_1780,N_1507);
and U3194 (N_3194,N_48,N_752);
nand U3195 (N_3195,N_1898,N_1226);
or U3196 (N_3196,N_696,N_2032);
nor U3197 (N_3197,N_2133,N_1);
or U3198 (N_3198,N_1888,N_6);
xor U3199 (N_3199,N_267,N_1336);
nor U3200 (N_3200,N_1569,N_1017);
xnor U3201 (N_3201,N_1155,N_2260);
nor U3202 (N_3202,N_1563,N_1056);
xor U3203 (N_3203,N_1465,N_1189);
nand U3204 (N_3204,N_2107,N_164);
or U3205 (N_3205,N_2222,N_176);
or U3206 (N_3206,N_603,N_1724);
xnor U3207 (N_3207,N_966,N_2383);
or U3208 (N_3208,N_219,N_2309);
or U3209 (N_3209,N_49,N_270);
or U3210 (N_3210,N_1034,N_2475);
nand U3211 (N_3211,N_1655,N_1257);
or U3212 (N_3212,N_2044,N_2298);
or U3213 (N_3213,N_1254,N_346);
or U3214 (N_3214,N_1999,N_560);
and U3215 (N_3215,N_1815,N_1249);
nor U3216 (N_3216,N_237,N_2340);
and U3217 (N_3217,N_2401,N_1447);
nor U3218 (N_3218,N_414,N_1915);
nand U3219 (N_3219,N_2010,N_922);
nor U3220 (N_3220,N_2012,N_1198);
nor U3221 (N_3221,N_271,N_1167);
xnor U3222 (N_3222,N_2183,N_1644);
nand U3223 (N_3223,N_1373,N_1873);
or U3224 (N_3224,N_1297,N_187);
nor U3225 (N_3225,N_2454,N_1912);
xor U3226 (N_3226,N_210,N_1552);
nand U3227 (N_3227,N_2348,N_1088);
nand U3228 (N_3228,N_2472,N_898);
xor U3229 (N_3229,N_264,N_1102);
xnor U3230 (N_3230,N_1677,N_593);
nor U3231 (N_3231,N_2438,N_98);
and U3232 (N_3232,N_2117,N_626);
xnor U3233 (N_3233,N_1125,N_866);
nor U3234 (N_3234,N_467,N_204);
and U3235 (N_3235,N_1828,N_1943);
nand U3236 (N_3236,N_65,N_227);
nor U3237 (N_3237,N_1709,N_1955);
and U3238 (N_3238,N_130,N_182);
xor U3239 (N_3239,N_1446,N_338);
and U3240 (N_3240,N_109,N_678);
and U3241 (N_3241,N_1081,N_215);
and U3242 (N_3242,N_628,N_1992);
and U3243 (N_3243,N_2098,N_1606);
xor U3244 (N_3244,N_95,N_1200);
nand U3245 (N_3245,N_347,N_2261);
and U3246 (N_3246,N_2172,N_1289);
xnor U3247 (N_3247,N_2429,N_376);
xnor U3248 (N_3248,N_1408,N_2198);
or U3249 (N_3249,N_1309,N_618);
nand U3250 (N_3250,N_764,N_1503);
nor U3251 (N_3251,N_1882,N_1070);
and U3252 (N_3252,N_31,N_600);
and U3253 (N_3253,N_1117,N_2057);
nand U3254 (N_3254,N_967,N_2486);
and U3255 (N_3255,N_2334,N_1825);
and U3256 (N_3256,N_1917,N_523);
nand U3257 (N_3257,N_508,N_381);
nor U3258 (N_3258,N_443,N_442);
xor U3259 (N_3259,N_772,N_584);
and U3260 (N_3260,N_1865,N_1057);
or U3261 (N_3261,N_1516,N_1436);
nand U3262 (N_3262,N_1572,N_2066);
and U3263 (N_3263,N_516,N_2427);
xnor U3264 (N_3264,N_1158,N_750);
nor U3265 (N_3265,N_610,N_1269);
or U3266 (N_3266,N_1922,N_1496);
xor U3267 (N_3267,N_222,N_1500);
and U3268 (N_3268,N_1356,N_1280);
nor U3269 (N_3269,N_371,N_1539);
and U3270 (N_3270,N_2219,N_1603);
nor U3271 (N_3271,N_135,N_1807);
xor U3272 (N_3272,N_596,N_2485);
nand U3273 (N_3273,N_1678,N_2364);
nor U3274 (N_3274,N_1323,N_1681);
or U3275 (N_3275,N_1524,N_1611);
nand U3276 (N_3276,N_995,N_418);
xor U3277 (N_3277,N_192,N_408);
xor U3278 (N_3278,N_2437,N_1460);
and U3279 (N_3279,N_975,N_78);
or U3280 (N_3280,N_1816,N_1758);
xnor U3281 (N_3281,N_1641,N_2065);
and U3282 (N_3282,N_1993,N_1691);
xor U3283 (N_3283,N_170,N_744);
and U3284 (N_3284,N_273,N_228);
and U3285 (N_3285,N_2433,N_2304);
or U3286 (N_3286,N_923,N_777);
nand U3287 (N_3287,N_664,N_1236);
xnor U3288 (N_3288,N_920,N_2369);
or U3289 (N_3289,N_701,N_2498);
or U3290 (N_3290,N_1079,N_934);
and U3291 (N_3291,N_1989,N_1624);
or U3292 (N_3292,N_2210,N_169);
xor U3293 (N_3293,N_1497,N_1646);
nand U3294 (N_3294,N_2468,N_2254);
xor U3295 (N_3295,N_1136,N_858);
and U3296 (N_3296,N_2426,N_1418);
and U3297 (N_3297,N_1159,N_1880);
xor U3298 (N_3298,N_241,N_74);
and U3299 (N_3299,N_1581,N_727);
xor U3300 (N_3300,N_2096,N_700);
nor U3301 (N_3301,N_954,N_1405);
or U3302 (N_3302,N_2100,N_1573);
nand U3303 (N_3303,N_1879,N_573);
or U3304 (N_3304,N_1848,N_2209);
xor U3305 (N_3305,N_2442,N_1303);
and U3306 (N_3306,N_759,N_248);
and U3307 (N_3307,N_1956,N_193);
or U3308 (N_3308,N_1643,N_1533);
nor U3309 (N_3309,N_1491,N_1240);
nand U3310 (N_3310,N_1188,N_1061);
or U3311 (N_3311,N_824,N_1043);
and U3312 (N_3312,N_2016,N_1166);
or U3313 (N_3313,N_163,N_2022);
and U3314 (N_3314,N_1044,N_708);
nor U3315 (N_3315,N_753,N_617);
or U3316 (N_3316,N_1728,N_1853);
nor U3317 (N_3317,N_538,N_1642);
xor U3318 (N_3318,N_673,N_1051);
xor U3319 (N_3319,N_1204,N_2246);
xor U3320 (N_3320,N_1919,N_1840);
or U3321 (N_3321,N_280,N_246);
or U3322 (N_3322,N_324,N_1224);
or U3323 (N_3323,N_1688,N_1233);
xnor U3324 (N_3324,N_1936,N_755);
nand U3325 (N_3325,N_559,N_944);
nor U3326 (N_3326,N_756,N_2443);
or U3327 (N_3327,N_321,N_1133);
or U3328 (N_3328,N_1367,N_977);
nor U3329 (N_3329,N_1045,N_2050);
nand U3330 (N_3330,N_2238,N_99);
and U3331 (N_3331,N_1351,N_1799);
nand U3332 (N_3332,N_838,N_2023);
xnor U3333 (N_3333,N_1574,N_1604);
and U3334 (N_3334,N_781,N_1549);
and U3335 (N_3335,N_396,N_1752);
xor U3336 (N_3336,N_383,N_452);
nor U3337 (N_3337,N_173,N_2263);
nor U3338 (N_3338,N_233,N_1046);
xnor U3339 (N_3339,N_2227,N_1175);
xnor U3340 (N_3340,N_981,N_284);
xor U3341 (N_3341,N_332,N_231);
or U3342 (N_3342,N_2192,N_2202);
xnor U3343 (N_3343,N_1711,N_2146);
nor U3344 (N_3344,N_660,N_1412);
xor U3345 (N_3345,N_2143,N_461);
and U3346 (N_3346,N_2484,N_103);
and U3347 (N_3347,N_1014,N_2112);
xor U3348 (N_3348,N_299,N_1686);
nor U3349 (N_3349,N_4,N_287);
nand U3350 (N_3350,N_1392,N_2230);
xnor U3351 (N_3351,N_794,N_2095);
or U3352 (N_3352,N_1838,N_1889);
nand U3353 (N_3353,N_1053,N_788);
or U3354 (N_3354,N_1398,N_513);
nand U3355 (N_3355,N_111,N_908);
nand U3356 (N_3356,N_2180,N_2001);
nor U3357 (N_3357,N_236,N_87);
xor U3358 (N_3358,N_2368,N_605);
nand U3359 (N_3359,N_1795,N_2495);
or U3360 (N_3360,N_2060,N_1169);
xor U3361 (N_3361,N_1023,N_1878);
nand U3362 (N_3362,N_1468,N_1470);
nor U3363 (N_3363,N_1609,N_929);
nand U3364 (N_3364,N_528,N_2466);
nand U3365 (N_3365,N_855,N_1844);
xnor U3366 (N_3366,N_599,N_1265);
nand U3367 (N_3367,N_2297,N_384);
xor U3368 (N_3368,N_395,N_903);
and U3369 (N_3369,N_765,N_790);
nand U3370 (N_3370,N_1343,N_2279);
or U3371 (N_3371,N_1300,N_1378);
or U3372 (N_3372,N_331,N_1640);
nand U3373 (N_3373,N_1191,N_1666);
nand U3374 (N_3374,N_469,N_550);
and U3375 (N_3375,N_1173,N_1050);
nand U3376 (N_3376,N_153,N_687);
nand U3377 (N_3377,N_75,N_699);
nor U3378 (N_3378,N_1089,N_597);
xor U3379 (N_3379,N_268,N_355);
nand U3380 (N_3380,N_1111,N_1964);
nand U3381 (N_3381,N_314,N_724);
nor U3382 (N_3382,N_1984,N_1213);
or U3383 (N_3383,N_2213,N_1273);
and U3384 (N_3384,N_2123,N_175);
and U3385 (N_3385,N_1638,N_2384);
nand U3386 (N_3386,N_1291,N_2372);
nand U3387 (N_3387,N_2151,N_168);
xor U3388 (N_3388,N_2121,N_1176);
or U3389 (N_3389,N_1326,N_894);
xor U3390 (N_3390,N_1248,N_2162);
xor U3391 (N_3391,N_2175,N_2063);
nor U3392 (N_3392,N_947,N_607);
xor U3393 (N_3393,N_2179,N_88);
and U3394 (N_3394,N_2008,N_2406);
xor U3395 (N_3395,N_1417,N_2467);
xor U3396 (N_3396,N_84,N_1946);
and U3397 (N_3397,N_489,N_2102);
or U3398 (N_3398,N_913,N_1144);
or U3399 (N_3399,N_2082,N_2496);
nor U3400 (N_3400,N_428,N_1383);
nor U3401 (N_3401,N_1522,N_1331);
nand U3402 (N_3402,N_255,N_15);
nand U3403 (N_3403,N_171,N_294);
and U3404 (N_3404,N_1911,N_152);
or U3405 (N_3405,N_2400,N_800);
xnor U3406 (N_3406,N_2140,N_115);
and U3407 (N_3407,N_1416,N_515);
and U3408 (N_3408,N_2170,N_1663);
or U3409 (N_3409,N_429,N_2267);
xor U3410 (N_3410,N_2235,N_2328);
nand U3411 (N_3411,N_2036,N_2324);
nand U3412 (N_3412,N_159,N_532);
xnor U3413 (N_3413,N_1283,N_1281);
nor U3414 (N_3414,N_655,N_1147);
nand U3415 (N_3415,N_819,N_2381);
xnor U3416 (N_3416,N_2342,N_1153);
and U3417 (N_3417,N_1665,N_2268);
or U3418 (N_3418,N_2026,N_736);
and U3419 (N_3419,N_2303,N_1287);
or U3420 (N_3420,N_2173,N_165);
or U3421 (N_3421,N_1096,N_1424);
nand U3422 (N_3422,N_758,N_1619);
and U3423 (N_3423,N_1264,N_1019);
xnor U3424 (N_3424,N_591,N_53);
or U3425 (N_3425,N_907,N_2358);
nor U3426 (N_3426,N_1098,N_1582);
or U3427 (N_3427,N_676,N_2053);
xnor U3428 (N_3428,N_933,N_884);
or U3429 (N_3429,N_980,N_622);
nor U3430 (N_3430,N_1071,N_144);
nand U3431 (N_3431,N_914,N_1495);
xnor U3432 (N_3432,N_2394,N_939);
nor U3433 (N_3433,N_1444,N_1684);
or U3434 (N_3434,N_2477,N_1464);
nor U3435 (N_3435,N_38,N_1789);
nand U3436 (N_3436,N_1298,N_845);
or U3437 (N_3437,N_47,N_1963);
nor U3438 (N_3438,N_1005,N_1141);
xor U3439 (N_3439,N_188,N_309);
nand U3440 (N_3440,N_562,N_1793);
or U3441 (N_3441,N_1769,N_641);
or U3442 (N_3442,N_862,N_1419);
xnor U3443 (N_3443,N_956,N_224);
and U3444 (N_3444,N_412,N_423);
nand U3445 (N_3445,N_5,N_1837);
xor U3446 (N_3446,N_937,N_535);
or U3447 (N_3447,N_731,N_1268);
nor U3448 (N_3448,N_156,N_8);
nor U3449 (N_3449,N_2311,N_2079);
nand U3450 (N_3450,N_1890,N_1926);
xor U3451 (N_3451,N_1818,N_1808);
xnor U3452 (N_3452,N_1928,N_2103);
xnor U3453 (N_3453,N_2275,N_454);
xnor U3454 (N_3454,N_372,N_2306);
or U3455 (N_3455,N_705,N_679);
nand U3456 (N_3456,N_57,N_1948);
and U3457 (N_3457,N_1230,N_129);
or U3458 (N_3458,N_2327,N_1508);
xor U3459 (N_3459,N_1119,N_2318);
and U3460 (N_3460,N_1712,N_568);
nand U3461 (N_3461,N_487,N_1242);
and U3462 (N_3462,N_1461,N_645);
xnor U3463 (N_3463,N_2048,N_1939);
nand U3464 (N_3464,N_2037,N_1120);
nor U3465 (N_3465,N_1084,N_965);
nand U3466 (N_3466,N_683,N_529);
or U3467 (N_3467,N_1648,N_2416);
xnor U3468 (N_3468,N_2041,N_1979);
or U3469 (N_3469,N_493,N_1662);
xnor U3470 (N_3470,N_721,N_2301);
nor U3471 (N_3471,N_869,N_405);
and U3472 (N_3472,N_1490,N_367);
nand U3473 (N_3473,N_62,N_716);
nor U3474 (N_3474,N_946,N_2293);
nand U3475 (N_3475,N_260,N_681);
nand U3476 (N_3476,N_1814,N_1831);
xor U3477 (N_3477,N_2199,N_1315);
nand U3478 (N_3478,N_1441,N_1101);
or U3479 (N_3479,N_2208,N_541);
xor U3480 (N_3480,N_166,N_2323);
nand U3481 (N_3481,N_1530,N_2129);
or U3482 (N_3482,N_158,N_1614);
xor U3483 (N_3483,N_1536,N_882);
nor U3484 (N_3484,N_2190,N_1854);
nand U3485 (N_3485,N_1062,N_2320);
xnor U3486 (N_3486,N_1407,N_2020);
nor U3487 (N_3487,N_546,N_720);
xor U3488 (N_3488,N_1726,N_337);
nor U3489 (N_3489,N_2122,N_1008);
nand U3490 (N_3490,N_2470,N_2197);
or U3491 (N_3491,N_278,N_1958);
nand U3492 (N_3492,N_857,N_1290);
nor U3493 (N_3493,N_1244,N_1937);
and U3494 (N_3494,N_59,N_1317);
or U3495 (N_3495,N_648,N_1647);
nand U3496 (N_3496,N_958,N_611);
or U3497 (N_3497,N_1737,N_2111);
nor U3498 (N_3498,N_296,N_1706);
nor U3499 (N_3499,N_2257,N_1587);
or U3500 (N_3500,N_505,N_1137);
xnor U3501 (N_3501,N_1073,N_1220);
or U3502 (N_3502,N_1947,N_579);
or U3503 (N_3503,N_905,N_1087);
or U3504 (N_3504,N_1687,N_2211);
nor U3505 (N_3505,N_796,N_2075);
nand U3506 (N_3506,N_258,N_1802);
and U3507 (N_3507,N_2355,N_2379);
and U3508 (N_3508,N_1625,N_1411);
or U3509 (N_3509,N_304,N_569);
nand U3510 (N_3510,N_953,N_1617);
nand U3511 (N_3511,N_829,N_1800);
nand U3512 (N_3512,N_2068,N_698);
nor U3513 (N_3513,N_55,N_1121);
xor U3514 (N_3514,N_1834,N_1235);
xnor U3515 (N_3515,N_2127,N_2085);
nand U3516 (N_3516,N_2014,N_102);
nand U3517 (N_3517,N_1771,N_1547);
nand U3518 (N_3518,N_1093,N_586);
or U3519 (N_3519,N_1959,N_2030);
nand U3520 (N_3520,N_245,N_2370);
and U3521 (N_3521,N_1305,N_1364);
xnor U3522 (N_3522,N_2142,N_1207);
or U3523 (N_3523,N_1082,N_1065);
nand U3524 (N_3524,N_1076,N_136);
and U3525 (N_3525,N_140,N_646);
nor U3526 (N_3526,N_1735,N_254);
and U3527 (N_3527,N_221,N_1381);
or U3528 (N_3528,N_1126,N_2156);
and U3529 (N_3529,N_1499,N_390);
nor U3530 (N_3530,N_400,N_1425);
and U3531 (N_3531,N_1049,N_1577);
nor U3532 (N_3532,N_1545,N_1160);
xor U3533 (N_3533,N_656,N_1733);
xnor U3534 (N_3534,N_1650,N_1784);
nand U3535 (N_3535,N_519,N_73);
or U3536 (N_3536,N_391,N_1092);
xor U3537 (N_3537,N_1170,N_51);
or U3538 (N_3538,N_2321,N_1325);
nand U3539 (N_3539,N_293,N_1864);
and U3540 (N_3540,N_1258,N_942);
or U3541 (N_3541,N_1493,N_1185);
nand U3542 (N_3542,N_263,N_1630);
nor U3543 (N_3543,N_959,N_266);
and U3544 (N_3544,N_29,N_1009);
xor U3545 (N_3545,N_1339,N_826);
nand U3546 (N_3546,N_2494,N_2310);
xnor U3547 (N_3547,N_821,N_2070);
xnor U3548 (N_3548,N_343,N_141);
or U3549 (N_3549,N_2272,N_1363);
xnor U3550 (N_3550,N_842,N_451);
xor U3551 (N_3551,N_1672,N_2191);
and U3552 (N_3552,N_1621,N_2161);
nor U3553 (N_3553,N_407,N_1434);
xnor U3554 (N_3554,N_1028,N_2029);
and U3555 (N_3555,N_16,N_979);
nor U3556 (N_3556,N_125,N_439);
and U3557 (N_3557,N_948,N_240);
nor U3558 (N_3558,N_816,N_1134);
and U3559 (N_3559,N_631,N_1177);
and U3560 (N_3560,N_536,N_2352);
or U3561 (N_3561,N_401,N_1836);
xor U3562 (N_3562,N_17,N_1829);
nor U3563 (N_3563,N_748,N_1135);
nor U3564 (N_3564,N_1827,N_374);
and U3565 (N_3565,N_1032,N_1145);
nand U3566 (N_3566,N_1401,N_1673);
and U3567 (N_3567,N_394,N_711);
or U3568 (N_3568,N_1732,N_2271);
and U3569 (N_3569,N_214,N_364);
xnor U3570 (N_3570,N_1905,N_638);
nor U3571 (N_3571,N_1636,N_784);
nor U3572 (N_3572,N_2322,N_1751);
and U3573 (N_3573,N_1639,N_2090);
or U3574 (N_3574,N_632,N_972);
xnor U3575 (N_3575,N_1150,N_1375);
and U3576 (N_3576,N_863,N_835);
xnor U3577 (N_3577,N_685,N_547);
nand U3578 (N_3578,N_1387,N_2025);
or U3579 (N_3579,N_901,N_757);
xnor U3580 (N_3580,N_814,N_1372);
nand U3581 (N_3581,N_1206,N_1591);
nand U3582 (N_3582,N_1658,N_2099);
nand U3583 (N_3583,N_697,N_1669);
xor U3584 (N_3584,N_466,N_1322);
xnor U3585 (N_3585,N_1151,N_2391);
nor U3586 (N_3586,N_2110,N_526);
or U3587 (N_3587,N_543,N_1704);
nor U3588 (N_3588,N_2333,N_2158);
nor U3589 (N_3589,N_2139,N_1974);
xnor U3590 (N_3590,N_330,N_1174);
xnor U3591 (N_3591,N_1232,N_1064);
nor U3592 (N_3592,N_1773,N_570);
xor U3593 (N_3593,N_41,N_334);
and U3594 (N_3594,N_812,N_1685);
nor U3595 (N_3595,N_567,N_180);
nand U3596 (N_3596,N_1274,N_1275);
xor U3597 (N_3597,N_1944,N_1437);
and U3598 (N_3598,N_1660,N_531);
and U3599 (N_3599,N_1680,N_2402);
nand U3600 (N_3600,N_1422,N_2231);
nand U3601 (N_3601,N_1859,N_895);
nor U3602 (N_3602,N_1961,N_368);
xnor U3603 (N_3603,N_1316,N_2250);
and U3604 (N_3604,N_847,N_21);
or U3605 (N_3605,N_1918,N_1921);
nand U3606 (N_3606,N_1149,N_799);
and U3607 (N_3607,N_2240,N_899);
and U3608 (N_3608,N_1566,N_427);
nand U3609 (N_3609,N_786,N_2451);
or U3610 (N_3610,N_1031,N_1845);
nand U3611 (N_3611,N_1951,N_301);
nor U3612 (N_3612,N_2492,N_1986);
or U3613 (N_3613,N_495,N_1238);
or U3614 (N_3614,N_1741,N_1534);
nor U3615 (N_3615,N_496,N_2083);
and U3616 (N_3616,N_1374,N_2482);
or U3617 (N_3617,N_1337,N_1015);
nor U3618 (N_3618,N_534,N_2249);
xnor U3619 (N_3619,N_1246,N_2419);
and U3620 (N_3620,N_2428,N_2236);
or U3621 (N_3621,N_1759,N_1904);
nand U3622 (N_3622,N_1682,N_2141);
nand U3623 (N_3623,N_2251,N_2319);
and U3624 (N_3624,N_1438,N_1910);
or U3625 (N_3625,N_1634,N_552);
nand U3626 (N_3626,N_1749,N_2294);
nand U3627 (N_3627,N_2431,N_94);
and U3628 (N_3628,N_1772,N_85);
nand U3629 (N_3629,N_1321,N_601);
nor U3630 (N_3630,N_1659,N_1319);
nand U3631 (N_3631,N_1130,N_2313);
nor U3632 (N_3632,N_1817,N_832);
nor U3633 (N_3633,N_150,N_2418);
nand U3634 (N_3634,N_2461,N_1055);
and U3635 (N_3635,N_353,N_1661);
xor U3636 (N_3636,N_1916,N_1753);
xnor U3637 (N_3637,N_1570,N_1457);
xor U3638 (N_3638,N_2264,N_1377);
or U3639 (N_3639,N_76,N_440);
or U3640 (N_3640,N_471,N_27);
or U3641 (N_3641,N_113,N_577);
and U3642 (N_3642,N_868,N_1471);
xor U3643 (N_3643,N_992,N_1025);
nand U3644 (N_3644,N_1627,N_703);
nor U3645 (N_3645,N_834,N_2465);
nor U3646 (N_3646,N_1228,N_447);
and U3647 (N_3647,N_910,N_2076);
nand U3648 (N_3648,N_476,N_1376);
and U3649 (N_3649,N_37,N_1104);
nor U3650 (N_3650,N_1165,N_339);
and U3651 (N_3651,N_551,N_2458);
and U3652 (N_3652,N_348,N_1778);
and U3653 (N_3653,N_1505,N_1830);
nand U3654 (N_3654,N_285,N_1509);
xor U3655 (N_3655,N_265,N_2186);
or U3656 (N_3656,N_1440,N_2365);
nand U3657 (N_3657,N_2019,N_783);
nor U3658 (N_3658,N_548,N_985);
xor U3659 (N_3659,N_1004,N_2150);
nor U3660 (N_3660,N_1714,N_906);
nor U3661 (N_3661,N_1823,N_564);
nand U3662 (N_3662,N_1487,N_986);
nor U3663 (N_3663,N_1588,N_2252);
nand U3664 (N_3664,N_1927,N_1798);
xor U3665 (N_3665,N_2277,N_1181);
nor U3666 (N_3666,N_723,N_2131);
nor U3667 (N_3667,N_768,N_1781);
nand U3668 (N_3668,N_328,N_1263);
nor U3669 (N_3669,N_1296,N_2476);
nand U3670 (N_3670,N_672,N_1725);
nand U3671 (N_3671,N_1736,N_1839);
or U3672 (N_3672,N_978,N_457);
and U3673 (N_3673,N_2132,N_649);
nor U3674 (N_3674,N_850,N_303);
nand U3675 (N_3675,N_2455,N_1449);
or U3676 (N_3676,N_2356,N_1909);
or U3677 (N_3677,N_92,N_1868);
xor U3678 (N_3678,N_1893,N_1941);
and U3679 (N_3679,N_2011,N_186);
and U3680 (N_3680,N_360,N_1695);
xor U3681 (N_3681,N_2403,N_1037);
nand U3682 (N_3682,N_1811,N_1810);
or U3683 (N_3683,N_1734,N_841);
or U3684 (N_3684,N_106,N_1000);
and U3685 (N_3685,N_1765,N_2302);
nor U3686 (N_3686,N_804,N_830);
or U3687 (N_3687,N_1127,N_373);
or U3688 (N_3688,N_1707,N_18);
xnor U3689 (N_3689,N_2290,N_473);
or U3690 (N_3690,N_1222,N_201);
or U3691 (N_3691,N_1428,N_556);
nand U3692 (N_3692,N_253,N_1697);
and U3693 (N_3693,N_936,N_1900);
nand U3694 (N_3694,N_256,N_288);
nand U3695 (N_3695,N_9,N_217);
nand U3696 (N_3696,N_2413,N_1458);
xor U3697 (N_3697,N_455,N_2134);
nor U3698 (N_3698,N_2359,N_1861);
nor U3699 (N_3699,N_2417,N_733);
or U3700 (N_3700,N_1390,N_613);
nand U3701 (N_3701,N_1492,N_1241);
nor U3702 (N_3702,N_2071,N_311);
or U3703 (N_3703,N_411,N_410);
and U3704 (N_3704,N_1285,N_1940);
nand U3705 (N_3705,N_354,N_598);
nor U3706 (N_3706,N_557,N_2221);
xor U3707 (N_3707,N_627,N_636);
xor U3708 (N_3708,N_647,N_1883);
and U3709 (N_3709,N_1310,N_2474);
xor U3710 (N_3710,N_2148,N_671);
nor U3711 (N_3711,N_506,N_1965);
and U3712 (N_3712,N_181,N_823);
nand U3713 (N_3713,N_1218,N_1489);
or U3714 (N_3714,N_1903,N_1344);
xor U3715 (N_3715,N_1399,N_502);
and U3716 (N_3716,N_787,N_1114);
nor U3717 (N_3717,N_1972,N_1106);
nor U3718 (N_3718,N_352,N_1676);
nor U3719 (N_3719,N_2043,N_1030);
and U3720 (N_3720,N_728,N_924);
and U3721 (N_3721,N_742,N_2104);
nor U3722 (N_3722,N_305,N_446);
nand U3723 (N_3723,N_1406,N_1653);
or U3724 (N_3724,N_544,N_79);
or U3725 (N_3725,N_1615,N_2021);
and U3726 (N_3726,N_128,N_2160);
nand U3727 (N_3727,N_963,N_1842);
nand U3728 (N_3728,N_916,N_39);
nand U3729 (N_3729,N_1994,N_1635);
nand U3730 (N_3730,N_26,N_1260);
nor U3731 (N_3731,N_208,N_1415);
xnor U3732 (N_3732,N_1038,N_1211);
and U3733 (N_3733,N_2237,N_1567);
nand U3734 (N_3734,N_325,N_1833);
nand U3735 (N_3735,N_326,N_1652);
or U3736 (N_3736,N_592,N_1314);
and U3737 (N_3737,N_1745,N_1952);
and U3738 (N_3738,N_261,N_2225);
nor U3739 (N_3739,N_1423,N_291);
xnor U3740 (N_3740,N_952,N_124);
nor U3741 (N_3741,N_935,N_2171);
nand U3742 (N_3742,N_509,N_813);
nand U3743 (N_3743,N_2386,N_1616);
nand U3744 (N_3744,N_746,N_2353);
nor U3745 (N_3745,N_651,N_732);
xor U3746 (N_3746,N_283,N_403);
nand U3747 (N_3747,N_880,N_525);
or U3748 (N_3748,N_378,N_1608);
and U3749 (N_3749,N_70,N_1083);
xnor U3750 (N_3750,N_776,N_728);
xnor U3751 (N_3751,N_1859,N_2362);
or U3752 (N_3752,N_20,N_2304);
xor U3753 (N_3753,N_561,N_168);
and U3754 (N_3754,N_693,N_1023);
nand U3755 (N_3755,N_622,N_1912);
nand U3756 (N_3756,N_1084,N_942);
nand U3757 (N_3757,N_782,N_2175);
nor U3758 (N_3758,N_1398,N_1170);
nand U3759 (N_3759,N_2314,N_1315);
or U3760 (N_3760,N_17,N_190);
and U3761 (N_3761,N_1882,N_677);
nor U3762 (N_3762,N_714,N_683);
nor U3763 (N_3763,N_1454,N_1609);
or U3764 (N_3764,N_1243,N_1558);
nor U3765 (N_3765,N_940,N_1678);
xnor U3766 (N_3766,N_2352,N_472);
xor U3767 (N_3767,N_1383,N_2225);
or U3768 (N_3768,N_1174,N_1719);
and U3769 (N_3769,N_2103,N_842);
xnor U3770 (N_3770,N_1661,N_19);
and U3771 (N_3771,N_5,N_1703);
nand U3772 (N_3772,N_1668,N_70);
xor U3773 (N_3773,N_1363,N_1193);
and U3774 (N_3774,N_216,N_1182);
xnor U3775 (N_3775,N_352,N_2450);
and U3776 (N_3776,N_1469,N_1473);
nand U3777 (N_3777,N_1292,N_1739);
nor U3778 (N_3778,N_1167,N_960);
or U3779 (N_3779,N_481,N_73);
nor U3780 (N_3780,N_1851,N_666);
nand U3781 (N_3781,N_1530,N_44);
nand U3782 (N_3782,N_2334,N_2127);
nand U3783 (N_3783,N_141,N_445);
and U3784 (N_3784,N_604,N_2266);
nor U3785 (N_3785,N_944,N_840);
or U3786 (N_3786,N_1517,N_1799);
or U3787 (N_3787,N_2103,N_2267);
nor U3788 (N_3788,N_1184,N_1845);
or U3789 (N_3789,N_2303,N_640);
or U3790 (N_3790,N_1069,N_1002);
xor U3791 (N_3791,N_2393,N_2202);
nand U3792 (N_3792,N_49,N_1612);
or U3793 (N_3793,N_546,N_2419);
nor U3794 (N_3794,N_1449,N_2074);
xor U3795 (N_3795,N_75,N_2374);
or U3796 (N_3796,N_1542,N_815);
xor U3797 (N_3797,N_1945,N_330);
and U3798 (N_3798,N_989,N_1909);
and U3799 (N_3799,N_353,N_905);
and U3800 (N_3800,N_1899,N_167);
nor U3801 (N_3801,N_2028,N_697);
xnor U3802 (N_3802,N_184,N_1055);
xnor U3803 (N_3803,N_726,N_643);
and U3804 (N_3804,N_2012,N_1057);
or U3805 (N_3805,N_1011,N_27);
and U3806 (N_3806,N_461,N_1502);
nor U3807 (N_3807,N_234,N_1787);
nand U3808 (N_3808,N_1701,N_55);
nor U3809 (N_3809,N_1818,N_848);
and U3810 (N_3810,N_485,N_2012);
and U3811 (N_3811,N_67,N_2331);
and U3812 (N_3812,N_294,N_692);
xnor U3813 (N_3813,N_1818,N_1663);
nor U3814 (N_3814,N_870,N_150);
xor U3815 (N_3815,N_1544,N_191);
nand U3816 (N_3816,N_1447,N_831);
or U3817 (N_3817,N_1996,N_1864);
or U3818 (N_3818,N_2335,N_467);
nand U3819 (N_3819,N_711,N_438);
nand U3820 (N_3820,N_219,N_1316);
nand U3821 (N_3821,N_2300,N_2366);
nor U3822 (N_3822,N_1118,N_686);
nor U3823 (N_3823,N_2147,N_122);
nand U3824 (N_3824,N_1439,N_299);
or U3825 (N_3825,N_1289,N_1501);
and U3826 (N_3826,N_1749,N_2354);
or U3827 (N_3827,N_61,N_2011);
or U3828 (N_3828,N_743,N_214);
nor U3829 (N_3829,N_2094,N_1026);
nand U3830 (N_3830,N_1,N_909);
and U3831 (N_3831,N_830,N_1937);
xnor U3832 (N_3832,N_1132,N_2357);
or U3833 (N_3833,N_691,N_759);
or U3834 (N_3834,N_416,N_1803);
nor U3835 (N_3835,N_2179,N_486);
nor U3836 (N_3836,N_1866,N_479);
nand U3837 (N_3837,N_2164,N_1804);
nor U3838 (N_3838,N_1473,N_2477);
nor U3839 (N_3839,N_685,N_1172);
or U3840 (N_3840,N_2084,N_1983);
and U3841 (N_3841,N_1399,N_2428);
and U3842 (N_3842,N_636,N_582);
nand U3843 (N_3843,N_827,N_2498);
nor U3844 (N_3844,N_1856,N_1096);
or U3845 (N_3845,N_1498,N_2188);
and U3846 (N_3846,N_2253,N_460);
or U3847 (N_3847,N_1543,N_2271);
nor U3848 (N_3848,N_1717,N_2257);
and U3849 (N_3849,N_434,N_1057);
nor U3850 (N_3850,N_1393,N_1543);
nor U3851 (N_3851,N_2471,N_562);
or U3852 (N_3852,N_1696,N_824);
nor U3853 (N_3853,N_872,N_254);
and U3854 (N_3854,N_2289,N_2477);
and U3855 (N_3855,N_516,N_2477);
xnor U3856 (N_3856,N_1188,N_1755);
nor U3857 (N_3857,N_1198,N_113);
xor U3858 (N_3858,N_2415,N_212);
nor U3859 (N_3859,N_1715,N_314);
and U3860 (N_3860,N_1814,N_1156);
nand U3861 (N_3861,N_1049,N_420);
nor U3862 (N_3862,N_1784,N_2497);
or U3863 (N_3863,N_532,N_2437);
and U3864 (N_3864,N_2212,N_2);
and U3865 (N_3865,N_2385,N_1519);
or U3866 (N_3866,N_318,N_1398);
xor U3867 (N_3867,N_2452,N_2022);
or U3868 (N_3868,N_1578,N_42);
nor U3869 (N_3869,N_410,N_1846);
nand U3870 (N_3870,N_902,N_955);
nand U3871 (N_3871,N_822,N_998);
nand U3872 (N_3872,N_1024,N_899);
xor U3873 (N_3873,N_228,N_1885);
or U3874 (N_3874,N_1781,N_1262);
or U3875 (N_3875,N_401,N_283);
nor U3876 (N_3876,N_1173,N_1813);
xnor U3877 (N_3877,N_1913,N_587);
xor U3878 (N_3878,N_1893,N_1982);
and U3879 (N_3879,N_705,N_1714);
xor U3880 (N_3880,N_2089,N_1225);
nor U3881 (N_3881,N_1556,N_831);
or U3882 (N_3882,N_2149,N_2421);
or U3883 (N_3883,N_2065,N_1917);
nor U3884 (N_3884,N_756,N_1988);
or U3885 (N_3885,N_1116,N_2248);
xor U3886 (N_3886,N_2277,N_113);
nor U3887 (N_3887,N_741,N_2312);
or U3888 (N_3888,N_1082,N_895);
nor U3889 (N_3889,N_1481,N_722);
nor U3890 (N_3890,N_630,N_1296);
and U3891 (N_3891,N_1123,N_1565);
nand U3892 (N_3892,N_2309,N_2327);
xor U3893 (N_3893,N_1799,N_423);
nand U3894 (N_3894,N_188,N_1448);
xnor U3895 (N_3895,N_2301,N_1389);
and U3896 (N_3896,N_741,N_1160);
xnor U3897 (N_3897,N_1614,N_229);
nor U3898 (N_3898,N_2212,N_256);
or U3899 (N_3899,N_1567,N_869);
xor U3900 (N_3900,N_308,N_1635);
nor U3901 (N_3901,N_1975,N_1352);
or U3902 (N_3902,N_344,N_2413);
nand U3903 (N_3903,N_2184,N_288);
and U3904 (N_3904,N_728,N_678);
nor U3905 (N_3905,N_1548,N_248);
nor U3906 (N_3906,N_958,N_2490);
or U3907 (N_3907,N_1645,N_1661);
xnor U3908 (N_3908,N_1801,N_1787);
or U3909 (N_3909,N_558,N_2286);
and U3910 (N_3910,N_1597,N_1244);
nor U3911 (N_3911,N_136,N_1297);
and U3912 (N_3912,N_1685,N_546);
xor U3913 (N_3913,N_823,N_2324);
nor U3914 (N_3914,N_1770,N_308);
or U3915 (N_3915,N_1903,N_1831);
or U3916 (N_3916,N_1138,N_981);
nor U3917 (N_3917,N_2138,N_667);
xor U3918 (N_3918,N_11,N_1734);
xnor U3919 (N_3919,N_1931,N_442);
or U3920 (N_3920,N_2183,N_1943);
nand U3921 (N_3921,N_540,N_1383);
xor U3922 (N_3922,N_1128,N_1735);
or U3923 (N_3923,N_1073,N_137);
nor U3924 (N_3924,N_1033,N_228);
or U3925 (N_3925,N_955,N_1543);
or U3926 (N_3926,N_2087,N_1818);
nand U3927 (N_3927,N_899,N_790);
xnor U3928 (N_3928,N_789,N_1404);
or U3929 (N_3929,N_342,N_481);
or U3930 (N_3930,N_1872,N_2476);
nor U3931 (N_3931,N_2450,N_143);
or U3932 (N_3932,N_1715,N_176);
nor U3933 (N_3933,N_2143,N_1527);
and U3934 (N_3934,N_2082,N_247);
nand U3935 (N_3935,N_2039,N_2130);
nor U3936 (N_3936,N_1601,N_1805);
and U3937 (N_3937,N_1513,N_2055);
and U3938 (N_3938,N_142,N_1733);
nor U3939 (N_3939,N_1956,N_1700);
or U3940 (N_3940,N_63,N_1936);
xnor U3941 (N_3941,N_541,N_1685);
xor U3942 (N_3942,N_2178,N_480);
nor U3943 (N_3943,N_1481,N_696);
and U3944 (N_3944,N_2139,N_2236);
and U3945 (N_3945,N_513,N_92);
or U3946 (N_3946,N_1521,N_2087);
and U3947 (N_3947,N_2100,N_393);
xnor U3948 (N_3948,N_1100,N_832);
and U3949 (N_3949,N_1166,N_2330);
nor U3950 (N_3950,N_1505,N_1109);
nor U3951 (N_3951,N_732,N_2416);
nand U3952 (N_3952,N_1544,N_1481);
nand U3953 (N_3953,N_1175,N_2100);
nor U3954 (N_3954,N_1115,N_980);
nor U3955 (N_3955,N_1617,N_2489);
nand U3956 (N_3956,N_1217,N_768);
or U3957 (N_3957,N_284,N_526);
xnor U3958 (N_3958,N_2231,N_1623);
nand U3959 (N_3959,N_162,N_1614);
nor U3960 (N_3960,N_1604,N_1008);
nand U3961 (N_3961,N_1476,N_673);
nor U3962 (N_3962,N_183,N_1076);
nor U3963 (N_3963,N_1716,N_2202);
nor U3964 (N_3964,N_1808,N_347);
nand U3965 (N_3965,N_1047,N_2187);
nor U3966 (N_3966,N_1947,N_910);
or U3967 (N_3967,N_1315,N_1551);
xor U3968 (N_3968,N_1331,N_1304);
or U3969 (N_3969,N_581,N_1963);
or U3970 (N_3970,N_1319,N_2214);
nand U3971 (N_3971,N_501,N_1985);
and U3972 (N_3972,N_1830,N_1869);
and U3973 (N_3973,N_1668,N_977);
xor U3974 (N_3974,N_1304,N_36);
nand U3975 (N_3975,N_2156,N_2279);
xnor U3976 (N_3976,N_2493,N_1103);
or U3977 (N_3977,N_1025,N_126);
and U3978 (N_3978,N_2459,N_1934);
nor U3979 (N_3979,N_437,N_1185);
nor U3980 (N_3980,N_441,N_159);
nor U3981 (N_3981,N_961,N_1925);
and U3982 (N_3982,N_1587,N_923);
xor U3983 (N_3983,N_1674,N_414);
nor U3984 (N_3984,N_1589,N_1113);
or U3985 (N_3985,N_825,N_432);
nor U3986 (N_3986,N_1276,N_784);
or U3987 (N_3987,N_1523,N_2298);
xnor U3988 (N_3988,N_863,N_1316);
or U3989 (N_3989,N_2050,N_1506);
nor U3990 (N_3990,N_1674,N_2239);
or U3991 (N_3991,N_287,N_2371);
or U3992 (N_3992,N_2335,N_954);
xor U3993 (N_3993,N_2139,N_2028);
or U3994 (N_3994,N_13,N_1888);
nor U3995 (N_3995,N_1792,N_2004);
xnor U3996 (N_3996,N_2331,N_1960);
or U3997 (N_3997,N_1977,N_465);
or U3998 (N_3998,N_189,N_1787);
and U3999 (N_3999,N_63,N_154);
xnor U4000 (N_4000,N_1651,N_1418);
and U4001 (N_4001,N_71,N_1047);
nor U4002 (N_4002,N_493,N_757);
xor U4003 (N_4003,N_611,N_1246);
nor U4004 (N_4004,N_1867,N_384);
nand U4005 (N_4005,N_1848,N_2032);
and U4006 (N_4006,N_1337,N_1356);
nor U4007 (N_4007,N_2400,N_392);
or U4008 (N_4008,N_1578,N_643);
and U4009 (N_4009,N_281,N_1872);
and U4010 (N_4010,N_2496,N_1479);
or U4011 (N_4011,N_2076,N_860);
xor U4012 (N_4012,N_397,N_1930);
and U4013 (N_4013,N_1664,N_795);
nor U4014 (N_4014,N_1890,N_1325);
xor U4015 (N_4015,N_1018,N_195);
xor U4016 (N_4016,N_482,N_1723);
nor U4017 (N_4017,N_874,N_1939);
and U4018 (N_4018,N_548,N_2063);
xor U4019 (N_4019,N_2085,N_1605);
nand U4020 (N_4020,N_1397,N_2117);
nor U4021 (N_4021,N_1819,N_2308);
xnor U4022 (N_4022,N_474,N_2406);
nor U4023 (N_4023,N_1254,N_1124);
or U4024 (N_4024,N_901,N_1602);
nor U4025 (N_4025,N_1557,N_1793);
nand U4026 (N_4026,N_473,N_1648);
xor U4027 (N_4027,N_1705,N_2417);
and U4028 (N_4028,N_1811,N_1280);
or U4029 (N_4029,N_1027,N_1642);
and U4030 (N_4030,N_1758,N_1509);
nor U4031 (N_4031,N_2396,N_2395);
or U4032 (N_4032,N_2152,N_1802);
nor U4033 (N_4033,N_233,N_963);
xor U4034 (N_4034,N_1336,N_240);
nand U4035 (N_4035,N_1412,N_2048);
and U4036 (N_4036,N_187,N_1703);
and U4037 (N_4037,N_1685,N_456);
nand U4038 (N_4038,N_773,N_1979);
nor U4039 (N_4039,N_2306,N_776);
xor U4040 (N_4040,N_292,N_1368);
nor U4041 (N_4041,N_1497,N_1262);
nand U4042 (N_4042,N_1068,N_1318);
and U4043 (N_4043,N_2140,N_1363);
and U4044 (N_4044,N_917,N_2010);
or U4045 (N_4045,N_684,N_80);
or U4046 (N_4046,N_399,N_2464);
nor U4047 (N_4047,N_2125,N_880);
xor U4048 (N_4048,N_1234,N_2087);
xnor U4049 (N_4049,N_2331,N_415);
xor U4050 (N_4050,N_1770,N_188);
nand U4051 (N_4051,N_2437,N_875);
nor U4052 (N_4052,N_982,N_1583);
or U4053 (N_4053,N_2028,N_2278);
nand U4054 (N_4054,N_2448,N_517);
and U4055 (N_4055,N_547,N_174);
xor U4056 (N_4056,N_1424,N_1266);
nor U4057 (N_4057,N_1033,N_368);
xnor U4058 (N_4058,N_2160,N_2174);
and U4059 (N_4059,N_309,N_1557);
nand U4060 (N_4060,N_617,N_1281);
xnor U4061 (N_4061,N_1141,N_635);
nor U4062 (N_4062,N_2385,N_984);
and U4063 (N_4063,N_163,N_2332);
nand U4064 (N_4064,N_1159,N_2439);
nand U4065 (N_4065,N_793,N_2083);
nand U4066 (N_4066,N_1454,N_1762);
xnor U4067 (N_4067,N_1364,N_519);
nor U4068 (N_4068,N_1689,N_406);
or U4069 (N_4069,N_1303,N_576);
and U4070 (N_4070,N_1214,N_491);
or U4071 (N_4071,N_2191,N_1450);
and U4072 (N_4072,N_2290,N_374);
and U4073 (N_4073,N_1152,N_552);
xor U4074 (N_4074,N_2360,N_2064);
xnor U4075 (N_4075,N_1498,N_1834);
or U4076 (N_4076,N_2192,N_515);
or U4077 (N_4077,N_222,N_991);
nand U4078 (N_4078,N_1751,N_2073);
xnor U4079 (N_4079,N_1254,N_1506);
nand U4080 (N_4080,N_1400,N_855);
or U4081 (N_4081,N_2142,N_1664);
xnor U4082 (N_4082,N_1614,N_1073);
nor U4083 (N_4083,N_215,N_2473);
and U4084 (N_4084,N_1360,N_564);
nand U4085 (N_4085,N_120,N_1169);
nand U4086 (N_4086,N_62,N_1549);
nor U4087 (N_4087,N_552,N_973);
or U4088 (N_4088,N_311,N_2014);
nor U4089 (N_4089,N_2036,N_2469);
nor U4090 (N_4090,N_950,N_1347);
xnor U4091 (N_4091,N_25,N_606);
or U4092 (N_4092,N_1617,N_2250);
or U4093 (N_4093,N_2319,N_445);
nand U4094 (N_4094,N_1310,N_1753);
xnor U4095 (N_4095,N_645,N_1388);
nor U4096 (N_4096,N_1190,N_2234);
xor U4097 (N_4097,N_55,N_809);
nand U4098 (N_4098,N_1762,N_2204);
or U4099 (N_4099,N_1016,N_912);
and U4100 (N_4100,N_2412,N_1658);
xor U4101 (N_4101,N_73,N_924);
and U4102 (N_4102,N_1757,N_1726);
and U4103 (N_4103,N_699,N_1801);
xnor U4104 (N_4104,N_770,N_612);
nor U4105 (N_4105,N_1875,N_1652);
or U4106 (N_4106,N_327,N_1612);
nor U4107 (N_4107,N_1991,N_281);
nor U4108 (N_4108,N_43,N_1240);
nor U4109 (N_4109,N_2463,N_1822);
and U4110 (N_4110,N_2109,N_1006);
xor U4111 (N_4111,N_2023,N_1910);
and U4112 (N_4112,N_1082,N_21);
xor U4113 (N_4113,N_587,N_1905);
nand U4114 (N_4114,N_1841,N_2433);
nand U4115 (N_4115,N_164,N_1516);
or U4116 (N_4116,N_1813,N_1433);
or U4117 (N_4117,N_555,N_1268);
xnor U4118 (N_4118,N_1677,N_1208);
or U4119 (N_4119,N_450,N_2414);
and U4120 (N_4120,N_312,N_1258);
xnor U4121 (N_4121,N_1605,N_1782);
xor U4122 (N_4122,N_1811,N_298);
nor U4123 (N_4123,N_1406,N_654);
nand U4124 (N_4124,N_668,N_1567);
nor U4125 (N_4125,N_2146,N_978);
nand U4126 (N_4126,N_820,N_966);
and U4127 (N_4127,N_772,N_890);
and U4128 (N_4128,N_538,N_158);
and U4129 (N_4129,N_2126,N_2453);
nand U4130 (N_4130,N_1743,N_689);
nand U4131 (N_4131,N_226,N_358);
or U4132 (N_4132,N_767,N_740);
and U4133 (N_4133,N_3,N_2286);
xnor U4134 (N_4134,N_1083,N_1829);
and U4135 (N_4135,N_124,N_744);
and U4136 (N_4136,N_2159,N_449);
nor U4137 (N_4137,N_2067,N_1084);
nor U4138 (N_4138,N_2117,N_1587);
or U4139 (N_4139,N_1105,N_1540);
xnor U4140 (N_4140,N_309,N_1673);
nand U4141 (N_4141,N_674,N_1132);
and U4142 (N_4142,N_1929,N_2365);
or U4143 (N_4143,N_257,N_778);
xnor U4144 (N_4144,N_13,N_1117);
and U4145 (N_4145,N_1982,N_348);
xor U4146 (N_4146,N_941,N_1153);
nand U4147 (N_4147,N_1859,N_388);
nor U4148 (N_4148,N_359,N_228);
xnor U4149 (N_4149,N_793,N_2498);
or U4150 (N_4150,N_542,N_962);
xnor U4151 (N_4151,N_481,N_1147);
nor U4152 (N_4152,N_1364,N_594);
nand U4153 (N_4153,N_2481,N_514);
nor U4154 (N_4154,N_1785,N_2039);
nand U4155 (N_4155,N_865,N_360);
nor U4156 (N_4156,N_1547,N_2106);
nor U4157 (N_4157,N_2437,N_168);
xnor U4158 (N_4158,N_1282,N_1180);
nor U4159 (N_4159,N_1950,N_1436);
xnor U4160 (N_4160,N_2136,N_1665);
or U4161 (N_4161,N_10,N_2198);
or U4162 (N_4162,N_1548,N_1735);
nand U4163 (N_4163,N_1676,N_1534);
or U4164 (N_4164,N_509,N_1037);
xor U4165 (N_4165,N_609,N_1422);
nand U4166 (N_4166,N_1134,N_1264);
nor U4167 (N_4167,N_2328,N_1255);
xnor U4168 (N_4168,N_1378,N_968);
or U4169 (N_4169,N_2429,N_1559);
or U4170 (N_4170,N_514,N_488);
and U4171 (N_4171,N_535,N_12);
or U4172 (N_4172,N_2323,N_982);
xnor U4173 (N_4173,N_1973,N_814);
or U4174 (N_4174,N_2153,N_152);
nand U4175 (N_4175,N_1003,N_2290);
and U4176 (N_4176,N_1225,N_1226);
nand U4177 (N_4177,N_902,N_2396);
nor U4178 (N_4178,N_1268,N_584);
nor U4179 (N_4179,N_1148,N_1495);
nor U4180 (N_4180,N_1356,N_1830);
nor U4181 (N_4181,N_936,N_2157);
nor U4182 (N_4182,N_374,N_372);
or U4183 (N_4183,N_1846,N_2101);
and U4184 (N_4184,N_1529,N_1755);
nand U4185 (N_4185,N_27,N_81);
or U4186 (N_4186,N_920,N_1767);
xor U4187 (N_4187,N_2374,N_1654);
and U4188 (N_4188,N_1122,N_920);
and U4189 (N_4189,N_2000,N_1473);
or U4190 (N_4190,N_79,N_701);
nor U4191 (N_4191,N_2306,N_622);
xnor U4192 (N_4192,N_1377,N_2066);
xor U4193 (N_4193,N_279,N_1891);
or U4194 (N_4194,N_1076,N_1900);
or U4195 (N_4195,N_991,N_961);
or U4196 (N_4196,N_1202,N_758);
and U4197 (N_4197,N_544,N_818);
xnor U4198 (N_4198,N_1049,N_715);
and U4199 (N_4199,N_2210,N_1220);
xor U4200 (N_4200,N_1363,N_651);
nand U4201 (N_4201,N_595,N_1336);
xor U4202 (N_4202,N_1191,N_1709);
and U4203 (N_4203,N_398,N_258);
nor U4204 (N_4204,N_953,N_1753);
nor U4205 (N_4205,N_2165,N_2369);
xor U4206 (N_4206,N_323,N_2043);
xor U4207 (N_4207,N_1338,N_1346);
xor U4208 (N_4208,N_874,N_295);
xor U4209 (N_4209,N_1411,N_1498);
or U4210 (N_4210,N_1910,N_1755);
and U4211 (N_4211,N_354,N_385);
nor U4212 (N_4212,N_137,N_319);
nand U4213 (N_4213,N_883,N_1236);
or U4214 (N_4214,N_1279,N_450);
or U4215 (N_4215,N_209,N_1852);
nor U4216 (N_4216,N_465,N_617);
or U4217 (N_4217,N_1058,N_321);
and U4218 (N_4218,N_1831,N_2102);
or U4219 (N_4219,N_1163,N_1777);
nand U4220 (N_4220,N_2384,N_179);
nand U4221 (N_4221,N_410,N_1216);
nor U4222 (N_4222,N_805,N_1598);
or U4223 (N_4223,N_297,N_866);
xor U4224 (N_4224,N_1059,N_1864);
and U4225 (N_4225,N_228,N_2291);
xnor U4226 (N_4226,N_160,N_2166);
or U4227 (N_4227,N_931,N_1571);
xnor U4228 (N_4228,N_400,N_237);
xnor U4229 (N_4229,N_913,N_1492);
nand U4230 (N_4230,N_2279,N_2443);
nand U4231 (N_4231,N_982,N_41);
nand U4232 (N_4232,N_2087,N_1431);
xor U4233 (N_4233,N_819,N_1286);
nor U4234 (N_4234,N_271,N_1765);
and U4235 (N_4235,N_1405,N_3);
nand U4236 (N_4236,N_1944,N_1326);
nor U4237 (N_4237,N_1123,N_2413);
nand U4238 (N_4238,N_2432,N_1863);
and U4239 (N_4239,N_1784,N_1325);
or U4240 (N_4240,N_1842,N_499);
nor U4241 (N_4241,N_2071,N_1683);
or U4242 (N_4242,N_251,N_2470);
nor U4243 (N_4243,N_1622,N_180);
nor U4244 (N_4244,N_339,N_692);
xnor U4245 (N_4245,N_1514,N_2324);
nand U4246 (N_4246,N_2052,N_349);
or U4247 (N_4247,N_722,N_1819);
nand U4248 (N_4248,N_491,N_410);
xnor U4249 (N_4249,N_2202,N_1008);
and U4250 (N_4250,N_291,N_957);
nand U4251 (N_4251,N_1407,N_2420);
nor U4252 (N_4252,N_1002,N_2106);
xor U4253 (N_4253,N_1265,N_2304);
or U4254 (N_4254,N_1747,N_1057);
and U4255 (N_4255,N_2273,N_172);
nand U4256 (N_4256,N_123,N_2300);
nor U4257 (N_4257,N_468,N_775);
nand U4258 (N_4258,N_24,N_744);
nand U4259 (N_4259,N_817,N_1207);
or U4260 (N_4260,N_2253,N_1765);
and U4261 (N_4261,N_211,N_2451);
nor U4262 (N_4262,N_1710,N_1688);
nand U4263 (N_4263,N_2023,N_246);
nor U4264 (N_4264,N_1029,N_2345);
or U4265 (N_4265,N_1217,N_703);
or U4266 (N_4266,N_1403,N_1960);
and U4267 (N_4267,N_2105,N_27);
nor U4268 (N_4268,N_800,N_1851);
and U4269 (N_4269,N_1834,N_942);
nor U4270 (N_4270,N_1280,N_2039);
nor U4271 (N_4271,N_2061,N_1803);
xnor U4272 (N_4272,N_2039,N_288);
xnor U4273 (N_4273,N_1363,N_1257);
nor U4274 (N_4274,N_1188,N_2499);
nor U4275 (N_4275,N_1139,N_2420);
or U4276 (N_4276,N_1044,N_1502);
nor U4277 (N_4277,N_1223,N_1317);
and U4278 (N_4278,N_236,N_1276);
xor U4279 (N_4279,N_2475,N_108);
or U4280 (N_4280,N_1285,N_2484);
nor U4281 (N_4281,N_5,N_1880);
nand U4282 (N_4282,N_1583,N_459);
nor U4283 (N_4283,N_293,N_3);
or U4284 (N_4284,N_559,N_1589);
xnor U4285 (N_4285,N_47,N_2436);
and U4286 (N_4286,N_907,N_1372);
xnor U4287 (N_4287,N_297,N_1380);
nand U4288 (N_4288,N_998,N_1897);
xor U4289 (N_4289,N_1825,N_727);
or U4290 (N_4290,N_1665,N_2014);
nor U4291 (N_4291,N_1322,N_620);
and U4292 (N_4292,N_1496,N_1197);
and U4293 (N_4293,N_705,N_1374);
and U4294 (N_4294,N_1282,N_628);
or U4295 (N_4295,N_215,N_981);
nor U4296 (N_4296,N_1516,N_426);
xor U4297 (N_4297,N_2164,N_2105);
or U4298 (N_4298,N_591,N_635);
nor U4299 (N_4299,N_638,N_790);
xor U4300 (N_4300,N_561,N_143);
nor U4301 (N_4301,N_2465,N_810);
xor U4302 (N_4302,N_2181,N_934);
or U4303 (N_4303,N_2288,N_1781);
or U4304 (N_4304,N_1221,N_856);
nor U4305 (N_4305,N_2327,N_1920);
nand U4306 (N_4306,N_512,N_1464);
nand U4307 (N_4307,N_603,N_1580);
xnor U4308 (N_4308,N_1969,N_2081);
or U4309 (N_4309,N_594,N_1145);
nand U4310 (N_4310,N_257,N_469);
nand U4311 (N_4311,N_2313,N_1437);
xnor U4312 (N_4312,N_1363,N_502);
xor U4313 (N_4313,N_342,N_340);
or U4314 (N_4314,N_13,N_1833);
xor U4315 (N_4315,N_2393,N_539);
xnor U4316 (N_4316,N_841,N_799);
or U4317 (N_4317,N_1374,N_1991);
and U4318 (N_4318,N_2081,N_2066);
xnor U4319 (N_4319,N_1837,N_1432);
or U4320 (N_4320,N_2183,N_2281);
nand U4321 (N_4321,N_1269,N_952);
nor U4322 (N_4322,N_1246,N_733);
or U4323 (N_4323,N_1464,N_210);
nor U4324 (N_4324,N_794,N_1308);
xnor U4325 (N_4325,N_762,N_1327);
or U4326 (N_4326,N_868,N_140);
nand U4327 (N_4327,N_400,N_1840);
nor U4328 (N_4328,N_1603,N_1978);
nand U4329 (N_4329,N_1049,N_2178);
and U4330 (N_4330,N_811,N_2155);
xnor U4331 (N_4331,N_1279,N_1542);
nand U4332 (N_4332,N_1615,N_744);
or U4333 (N_4333,N_1257,N_2319);
nor U4334 (N_4334,N_2065,N_702);
and U4335 (N_4335,N_2283,N_16);
and U4336 (N_4336,N_2431,N_1453);
nor U4337 (N_4337,N_1314,N_1956);
and U4338 (N_4338,N_262,N_1326);
nor U4339 (N_4339,N_2495,N_2356);
or U4340 (N_4340,N_2223,N_536);
nor U4341 (N_4341,N_218,N_1644);
nand U4342 (N_4342,N_1334,N_2391);
and U4343 (N_4343,N_847,N_832);
and U4344 (N_4344,N_880,N_2020);
nor U4345 (N_4345,N_246,N_1750);
and U4346 (N_4346,N_2415,N_1235);
xor U4347 (N_4347,N_591,N_339);
xnor U4348 (N_4348,N_956,N_2207);
nor U4349 (N_4349,N_536,N_176);
and U4350 (N_4350,N_2143,N_624);
xnor U4351 (N_4351,N_598,N_1054);
nor U4352 (N_4352,N_771,N_2322);
nand U4353 (N_4353,N_707,N_2012);
xor U4354 (N_4354,N_1643,N_299);
nand U4355 (N_4355,N_952,N_700);
and U4356 (N_4356,N_1559,N_801);
or U4357 (N_4357,N_109,N_2358);
nor U4358 (N_4358,N_1777,N_693);
and U4359 (N_4359,N_2337,N_1449);
or U4360 (N_4360,N_1920,N_1519);
and U4361 (N_4361,N_2319,N_1420);
xnor U4362 (N_4362,N_1033,N_2244);
nand U4363 (N_4363,N_1468,N_2084);
xor U4364 (N_4364,N_2172,N_237);
nand U4365 (N_4365,N_2386,N_1464);
xor U4366 (N_4366,N_1669,N_1735);
and U4367 (N_4367,N_1903,N_1273);
and U4368 (N_4368,N_1531,N_43);
nand U4369 (N_4369,N_1401,N_438);
xor U4370 (N_4370,N_559,N_2266);
nand U4371 (N_4371,N_1733,N_2136);
or U4372 (N_4372,N_940,N_362);
and U4373 (N_4373,N_90,N_1334);
nand U4374 (N_4374,N_1124,N_1335);
nand U4375 (N_4375,N_609,N_2477);
or U4376 (N_4376,N_1344,N_2409);
nor U4377 (N_4377,N_795,N_479);
or U4378 (N_4378,N_1632,N_2000);
nand U4379 (N_4379,N_727,N_2297);
nand U4380 (N_4380,N_40,N_988);
and U4381 (N_4381,N_93,N_235);
or U4382 (N_4382,N_1738,N_1108);
nand U4383 (N_4383,N_1707,N_1239);
and U4384 (N_4384,N_1792,N_775);
nor U4385 (N_4385,N_2262,N_1860);
xor U4386 (N_4386,N_1469,N_585);
xnor U4387 (N_4387,N_2409,N_1508);
nor U4388 (N_4388,N_1402,N_127);
nor U4389 (N_4389,N_2319,N_2060);
and U4390 (N_4390,N_86,N_179);
or U4391 (N_4391,N_608,N_217);
xor U4392 (N_4392,N_2043,N_1643);
nor U4393 (N_4393,N_1049,N_1938);
nand U4394 (N_4394,N_1057,N_735);
xor U4395 (N_4395,N_695,N_382);
xor U4396 (N_4396,N_1728,N_303);
nand U4397 (N_4397,N_1360,N_1919);
nand U4398 (N_4398,N_1521,N_1006);
nor U4399 (N_4399,N_1234,N_1984);
xnor U4400 (N_4400,N_535,N_2448);
xor U4401 (N_4401,N_827,N_1867);
nor U4402 (N_4402,N_2266,N_16);
and U4403 (N_4403,N_2032,N_1491);
and U4404 (N_4404,N_1225,N_1213);
nor U4405 (N_4405,N_2325,N_2271);
and U4406 (N_4406,N_2326,N_1463);
or U4407 (N_4407,N_2027,N_556);
xnor U4408 (N_4408,N_1627,N_414);
nor U4409 (N_4409,N_2395,N_1211);
or U4410 (N_4410,N_1520,N_1457);
nor U4411 (N_4411,N_1846,N_1976);
nor U4412 (N_4412,N_812,N_629);
xor U4413 (N_4413,N_1393,N_1890);
nor U4414 (N_4414,N_39,N_2152);
nor U4415 (N_4415,N_560,N_947);
xnor U4416 (N_4416,N_399,N_1088);
nand U4417 (N_4417,N_228,N_1718);
and U4418 (N_4418,N_2194,N_2157);
or U4419 (N_4419,N_2035,N_2445);
and U4420 (N_4420,N_971,N_1216);
nor U4421 (N_4421,N_2217,N_787);
xor U4422 (N_4422,N_1229,N_1803);
and U4423 (N_4423,N_1392,N_1973);
and U4424 (N_4424,N_1025,N_1524);
and U4425 (N_4425,N_2324,N_1648);
or U4426 (N_4426,N_1484,N_674);
or U4427 (N_4427,N_548,N_1811);
nor U4428 (N_4428,N_2076,N_713);
nand U4429 (N_4429,N_184,N_2160);
nor U4430 (N_4430,N_2357,N_1503);
xnor U4431 (N_4431,N_2103,N_1528);
nor U4432 (N_4432,N_2113,N_501);
nor U4433 (N_4433,N_1090,N_2065);
xnor U4434 (N_4434,N_561,N_2195);
and U4435 (N_4435,N_1454,N_964);
nor U4436 (N_4436,N_209,N_1680);
or U4437 (N_4437,N_940,N_2229);
xnor U4438 (N_4438,N_1374,N_1889);
or U4439 (N_4439,N_364,N_2246);
and U4440 (N_4440,N_2223,N_573);
xnor U4441 (N_4441,N_625,N_1317);
nand U4442 (N_4442,N_375,N_1526);
nand U4443 (N_4443,N_336,N_535);
and U4444 (N_4444,N_1125,N_747);
nor U4445 (N_4445,N_502,N_2405);
nand U4446 (N_4446,N_1442,N_603);
and U4447 (N_4447,N_1380,N_166);
nor U4448 (N_4448,N_1958,N_1247);
and U4449 (N_4449,N_1955,N_293);
and U4450 (N_4450,N_80,N_1020);
nand U4451 (N_4451,N_2491,N_1788);
and U4452 (N_4452,N_434,N_2462);
nand U4453 (N_4453,N_715,N_246);
or U4454 (N_4454,N_1556,N_1672);
and U4455 (N_4455,N_925,N_873);
nor U4456 (N_4456,N_2341,N_383);
and U4457 (N_4457,N_802,N_1314);
xnor U4458 (N_4458,N_1106,N_2022);
or U4459 (N_4459,N_1799,N_528);
xnor U4460 (N_4460,N_263,N_400);
and U4461 (N_4461,N_1667,N_262);
xnor U4462 (N_4462,N_1196,N_1832);
xor U4463 (N_4463,N_1630,N_337);
or U4464 (N_4464,N_2008,N_2287);
nor U4465 (N_4465,N_834,N_133);
nor U4466 (N_4466,N_2323,N_144);
nor U4467 (N_4467,N_1152,N_401);
or U4468 (N_4468,N_1754,N_436);
xnor U4469 (N_4469,N_114,N_875);
and U4470 (N_4470,N_1747,N_1571);
nand U4471 (N_4471,N_159,N_508);
nor U4472 (N_4472,N_327,N_63);
and U4473 (N_4473,N_1839,N_777);
xor U4474 (N_4474,N_1238,N_876);
nand U4475 (N_4475,N_490,N_2245);
and U4476 (N_4476,N_1244,N_921);
and U4477 (N_4477,N_1737,N_675);
xnor U4478 (N_4478,N_212,N_610);
nor U4479 (N_4479,N_870,N_2326);
xor U4480 (N_4480,N_2437,N_567);
nand U4481 (N_4481,N_854,N_1434);
and U4482 (N_4482,N_385,N_438);
xor U4483 (N_4483,N_1591,N_1730);
xnor U4484 (N_4484,N_333,N_399);
or U4485 (N_4485,N_1928,N_291);
nand U4486 (N_4486,N_1563,N_824);
nor U4487 (N_4487,N_1409,N_549);
xnor U4488 (N_4488,N_90,N_1412);
xor U4489 (N_4489,N_1324,N_2389);
and U4490 (N_4490,N_611,N_570);
and U4491 (N_4491,N_500,N_1262);
nor U4492 (N_4492,N_67,N_93);
nand U4493 (N_4493,N_1311,N_390);
nand U4494 (N_4494,N_1042,N_942);
xnor U4495 (N_4495,N_2216,N_2409);
nand U4496 (N_4496,N_199,N_574);
or U4497 (N_4497,N_149,N_2077);
and U4498 (N_4498,N_427,N_1009);
nand U4499 (N_4499,N_275,N_1002);
nor U4500 (N_4500,N_1127,N_801);
or U4501 (N_4501,N_690,N_2115);
nand U4502 (N_4502,N_277,N_1458);
or U4503 (N_4503,N_2488,N_2253);
and U4504 (N_4504,N_577,N_1499);
nand U4505 (N_4505,N_625,N_345);
xnor U4506 (N_4506,N_833,N_1743);
xor U4507 (N_4507,N_724,N_2109);
or U4508 (N_4508,N_2041,N_1565);
nand U4509 (N_4509,N_2145,N_160);
xor U4510 (N_4510,N_343,N_1201);
nor U4511 (N_4511,N_784,N_2426);
and U4512 (N_4512,N_212,N_172);
and U4513 (N_4513,N_2082,N_1241);
and U4514 (N_4514,N_2346,N_2242);
or U4515 (N_4515,N_1552,N_530);
and U4516 (N_4516,N_2176,N_387);
nand U4517 (N_4517,N_2345,N_1274);
nor U4518 (N_4518,N_265,N_1694);
or U4519 (N_4519,N_1532,N_1618);
and U4520 (N_4520,N_872,N_1565);
nand U4521 (N_4521,N_1787,N_2315);
and U4522 (N_4522,N_1944,N_2333);
and U4523 (N_4523,N_1347,N_1095);
nand U4524 (N_4524,N_2321,N_1899);
nand U4525 (N_4525,N_614,N_1102);
xor U4526 (N_4526,N_273,N_2163);
xnor U4527 (N_4527,N_1782,N_618);
xor U4528 (N_4528,N_693,N_1690);
or U4529 (N_4529,N_1942,N_587);
nand U4530 (N_4530,N_1718,N_475);
nand U4531 (N_4531,N_2030,N_622);
and U4532 (N_4532,N_1786,N_1800);
xnor U4533 (N_4533,N_1535,N_52);
nand U4534 (N_4534,N_1537,N_70);
xor U4535 (N_4535,N_1256,N_1808);
and U4536 (N_4536,N_1523,N_1860);
nor U4537 (N_4537,N_317,N_1936);
nand U4538 (N_4538,N_2414,N_900);
or U4539 (N_4539,N_289,N_1373);
nor U4540 (N_4540,N_101,N_357);
nor U4541 (N_4541,N_651,N_1338);
xor U4542 (N_4542,N_2330,N_1509);
nand U4543 (N_4543,N_2035,N_2194);
xnor U4544 (N_4544,N_2317,N_1421);
and U4545 (N_4545,N_881,N_1374);
nor U4546 (N_4546,N_1325,N_2417);
nand U4547 (N_4547,N_1146,N_2031);
or U4548 (N_4548,N_1702,N_1438);
nor U4549 (N_4549,N_2117,N_494);
nand U4550 (N_4550,N_2254,N_1523);
or U4551 (N_4551,N_1698,N_234);
xnor U4552 (N_4552,N_1490,N_1173);
nor U4553 (N_4553,N_2374,N_2464);
nand U4554 (N_4554,N_195,N_1642);
and U4555 (N_4555,N_377,N_1360);
nor U4556 (N_4556,N_666,N_786);
nor U4557 (N_4557,N_107,N_1411);
nor U4558 (N_4558,N_511,N_1570);
or U4559 (N_4559,N_2370,N_1977);
nor U4560 (N_4560,N_2245,N_2468);
xor U4561 (N_4561,N_1867,N_819);
nor U4562 (N_4562,N_267,N_1502);
or U4563 (N_4563,N_2306,N_807);
nand U4564 (N_4564,N_1532,N_1788);
xnor U4565 (N_4565,N_765,N_1580);
or U4566 (N_4566,N_293,N_562);
nand U4567 (N_4567,N_861,N_1167);
xnor U4568 (N_4568,N_1459,N_772);
nand U4569 (N_4569,N_1543,N_2069);
or U4570 (N_4570,N_21,N_2418);
nand U4571 (N_4571,N_1642,N_80);
or U4572 (N_4572,N_1672,N_1759);
nand U4573 (N_4573,N_901,N_2363);
xor U4574 (N_4574,N_1280,N_457);
nand U4575 (N_4575,N_298,N_2183);
xnor U4576 (N_4576,N_379,N_2290);
xnor U4577 (N_4577,N_394,N_251);
or U4578 (N_4578,N_270,N_2115);
nand U4579 (N_4579,N_1275,N_1409);
nor U4580 (N_4580,N_308,N_759);
xnor U4581 (N_4581,N_1704,N_2217);
and U4582 (N_4582,N_1201,N_848);
xor U4583 (N_4583,N_487,N_770);
nand U4584 (N_4584,N_1440,N_1064);
nand U4585 (N_4585,N_2030,N_982);
nand U4586 (N_4586,N_576,N_943);
or U4587 (N_4587,N_1739,N_217);
or U4588 (N_4588,N_8,N_2323);
or U4589 (N_4589,N_1667,N_1924);
nor U4590 (N_4590,N_1253,N_1484);
and U4591 (N_4591,N_1829,N_1673);
xnor U4592 (N_4592,N_177,N_2165);
nor U4593 (N_4593,N_1059,N_150);
or U4594 (N_4594,N_1963,N_2266);
and U4595 (N_4595,N_181,N_2020);
or U4596 (N_4596,N_1187,N_1759);
and U4597 (N_4597,N_1212,N_2263);
or U4598 (N_4598,N_495,N_2363);
and U4599 (N_4599,N_2200,N_1312);
xor U4600 (N_4600,N_242,N_496);
nand U4601 (N_4601,N_2348,N_366);
nor U4602 (N_4602,N_1799,N_1997);
xor U4603 (N_4603,N_93,N_1069);
xor U4604 (N_4604,N_864,N_1290);
and U4605 (N_4605,N_1479,N_1334);
nor U4606 (N_4606,N_1054,N_1683);
nand U4607 (N_4607,N_215,N_325);
xnor U4608 (N_4608,N_1776,N_158);
nand U4609 (N_4609,N_1366,N_903);
xor U4610 (N_4610,N_173,N_675);
or U4611 (N_4611,N_1612,N_1364);
and U4612 (N_4612,N_1818,N_1609);
nor U4613 (N_4613,N_2154,N_879);
xnor U4614 (N_4614,N_1,N_416);
nand U4615 (N_4615,N_264,N_568);
nand U4616 (N_4616,N_1159,N_1986);
nor U4617 (N_4617,N_1168,N_1616);
and U4618 (N_4618,N_646,N_1396);
nand U4619 (N_4619,N_1146,N_1134);
and U4620 (N_4620,N_465,N_87);
nor U4621 (N_4621,N_781,N_1099);
or U4622 (N_4622,N_979,N_448);
nand U4623 (N_4623,N_1183,N_720);
nor U4624 (N_4624,N_1089,N_718);
or U4625 (N_4625,N_259,N_973);
and U4626 (N_4626,N_2021,N_562);
and U4627 (N_4627,N_2491,N_668);
and U4628 (N_4628,N_2132,N_138);
xor U4629 (N_4629,N_513,N_2410);
and U4630 (N_4630,N_1260,N_2176);
nand U4631 (N_4631,N_860,N_1677);
and U4632 (N_4632,N_1901,N_2034);
or U4633 (N_4633,N_2216,N_541);
nand U4634 (N_4634,N_1055,N_2478);
and U4635 (N_4635,N_577,N_1441);
nor U4636 (N_4636,N_1685,N_662);
nand U4637 (N_4637,N_1910,N_828);
and U4638 (N_4638,N_1604,N_1917);
and U4639 (N_4639,N_2380,N_2072);
nor U4640 (N_4640,N_1404,N_914);
nand U4641 (N_4641,N_1325,N_758);
nor U4642 (N_4642,N_2315,N_675);
nand U4643 (N_4643,N_2419,N_981);
and U4644 (N_4644,N_1597,N_223);
nand U4645 (N_4645,N_1987,N_1303);
nor U4646 (N_4646,N_745,N_979);
xor U4647 (N_4647,N_2037,N_1666);
or U4648 (N_4648,N_1902,N_442);
or U4649 (N_4649,N_487,N_846);
nand U4650 (N_4650,N_742,N_613);
nand U4651 (N_4651,N_1961,N_997);
nand U4652 (N_4652,N_1433,N_354);
or U4653 (N_4653,N_2001,N_1841);
or U4654 (N_4654,N_636,N_1545);
nand U4655 (N_4655,N_1113,N_214);
and U4656 (N_4656,N_944,N_83);
and U4657 (N_4657,N_690,N_2093);
nor U4658 (N_4658,N_1195,N_1528);
or U4659 (N_4659,N_1156,N_1996);
nand U4660 (N_4660,N_120,N_72);
or U4661 (N_4661,N_822,N_607);
nor U4662 (N_4662,N_1587,N_1397);
nand U4663 (N_4663,N_2450,N_520);
and U4664 (N_4664,N_1647,N_166);
nand U4665 (N_4665,N_1034,N_230);
nand U4666 (N_4666,N_349,N_466);
or U4667 (N_4667,N_2088,N_2275);
nor U4668 (N_4668,N_2075,N_1770);
nor U4669 (N_4669,N_1692,N_504);
nand U4670 (N_4670,N_2356,N_1274);
xor U4671 (N_4671,N_286,N_1100);
and U4672 (N_4672,N_1505,N_44);
xnor U4673 (N_4673,N_1382,N_1997);
or U4674 (N_4674,N_938,N_816);
nand U4675 (N_4675,N_140,N_1912);
or U4676 (N_4676,N_304,N_1258);
xnor U4677 (N_4677,N_2102,N_2319);
xnor U4678 (N_4678,N_2059,N_2377);
nor U4679 (N_4679,N_1711,N_162);
or U4680 (N_4680,N_331,N_543);
xnor U4681 (N_4681,N_742,N_2351);
xnor U4682 (N_4682,N_436,N_1326);
nand U4683 (N_4683,N_1448,N_2086);
xor U4684 (N_4684,N_1293,N_900);
xnor U4685 (N_4685,N_1946,N_459);
nor U4686 (N_4686,N_1480,N_1150);
xnor U4687 (N_4687,N_1444,N_2324);
and U4688 (N_4688,N_2094,N_2437);
xnor U4689 (N_4689,N_1976,N_1045);
xnor U4690 (N_4690,N_2099,N_1135);
nor U4691 (N_4691,N_1669,N_1539);
xor U4692 (N_4692,N_2324,N_616);
nand U4693 (N_4693,N_2276,N_809);
xnor U4694 (N_4694,N_1660,N_913);
nand U4695 (N_4695,N_566,N_1363);
nand U4696 (N_4696,N_1475,N_2204);
nor U4697 (N_4697,N_235,N_606);
and U4698 (N_4698,N_527,N_1827);
xnor U4699 (N_4699,N_10,N_1695);
nor U4700 (N_4700,N_906,N_2224);
nand U4701 (N_4701,N_760,N_2184);
nand U4702 (N_4702,N_2290,N_1260);
xor U4703 (N_4703,N_407,N_674);
nand U4704 (N_4704,N_2085,N_2310);
or U4705 (N_4705,N_877,N_1543);
nor U4706 (N_4706,N_410,N_1083);
nor U4707 (N_4707,N_552,N_472);
xor U4708 (N_4708,N_274,N_1596);
nand U4709 (N_4709,N_1733,N_2195);
xnor U4710 (N_4710,N_426,N_256);
nand U4711 (N_4711,N_876,N_2452);
nand U4712 (N_4712,N_1601,N_518);
nor U4713 (N_4713,N_1099,N_797);
or U4714 (N_4714,N_292,N_1282);
nor U4715 (N_4715,N_40,N_791);
or U4716 (N_4716,N_1372,N_170);
nor U4717 (N_4717,N_754,N_2189);
and U4718 (N_4718,N_371,N_2470);
or U4719 (N_4719,N_357,N_1800);
and U4720 (N_4720,N_1841,N_307);
nor U4721 (N_4721,N_1569,N_1982);
or U4722 (N_4722,N_1095,N_1444);
and U4723 (N_4723,N_451,N_889);
xor U4724 (N_4724,N_1218,N_1015);
nand U4725 (N_4725,N_1355,N_2428);
nand U4726 (N_4726,N_1590,N_1105);
and U4727 (N_4727,N_1047,N_1408);
nand U4728 (N_4728,N_1213,N_594);
nand U4729 (N_4729,N_2285,N_1504);
nor U4730 (N_4730,N_1022,N_2006);
nor U4731 (N_4731,N_630,N_664);
or U4732 (N_4732,N_417,N_1871);
xnor U4733 (N_4733,N_129,N_2007);
and U4734 (N_4734,N_1503,N_50);
and U4735 (N_4735,N_1904,N_1591);
nor U4736 (N_4736,N_1531,N_233);
or U4737 (N_4737,N_543,N_1697);
and U4738 (N_4738,N_2465,N_2274);
and U4739 (N_4739,N_905,N_1224);
nand U4740 (N_4740,N_2117,N_938);
nor U4741 (N_4741,N_358,N_825);
or U4742 (N_4742,N_263,N_1148);
and U4743 (N_4743,N_223,N_236);
xor U4744 (N_4744,N_188,N_504);
and U4745 (N_4745,N_2020,N_922);
or U4746 (N_4746,N_2221,N_2458);
or U4747 (N_4747,N_1117,N_2377);
or U4748 (N_4748,N_2488,N_546);
and U4749 (N_4749,N_2157,N_265);
and U4750 (N_4750,N_811,N_2473);
xnor U4751 (N_4751,N_552,N_2080);
nor U4752 (N_4752,N_2317,N_1925);
nor U4753 (N_4753,N_138,N_1311);
xnor U4754 (N_4754,N_2023,N_1314);
or U4755 (N_4755,N_576,N_2038);
and U4756 (N_4756,N_2332,N_1805);
nor U4757 (N_4757,N_1317,N_1950);
nor U4758 (N_4758,N_830,N_5);
nand U4759 (N_4759,N_2238,N_335);
or U4760 (N_4760,N_1469,N_982);
xor U4761 (N_4761,N_1876,N_1406);
or U4762 (N_4762,N_768,N_2280);
nand U4763 (N_4763,N_1868,N_1076);
or U4764 (N_4764,N_1327,N_2121);
nor U4765 (N_4765,N_1551,N_1072);
and U4766 (N_4766,N_1689,N_2044);
or U4767 (N_4767,N_1956,N_466);
or U4768 (N_4768,N_2044,N_130);
and U4769 (N_4769,N_1469,N_583);
and U4770 (N_4770,N_917,N_217);
and U4771 (N_4771,N_55,N_240);
nand U4772 (N_4772,N_1340,N_1053);
nor U4773 (N_4773,N_2247,N_1029);
or U4774 (N_4774,N_29,N_738);
nor U4775 (N_4775,N_1539,N_1445);
and U4776 (N_4776,N_1377,N_2092);
xor U4777 (N_4777,N_956,N_638);
or U4778 (N_4778,N_2123,N_1855);
xnor U4779 (N_4779,N_215,N_714);
and U4780 (N_4780,N_614,N_1428);
xor U4781 (N_4781,N_1393,N_1058);
or U4782 (N_4782,N_2230,N_1465);
or U4783 (N_4783,N_1504,N_49);
nor U4784 (N_4784,N_146,N_689);
or U4785 (N_4785,N_1216,N_1312);
and U4786 (N_4786,N_1674,N_2435);
xnor U4787 (N_4787,N_2010,N_377);
nor U4788 (N_4788,N_2274,N_1059);
xnor U4789 (N_4789,N_1458,N_1057);
and U4790 (N_4790,N_791,N_2054);
and U4791 (N_4791,N_774,N_1814);
and U4792 (N_4792,N_1549,N_1126);
and U4793 (N_4793,N_1407,N_1201);
xnor U4794 (N_4794,N_500,N_1219);
and U4795 (N_4795,N_1681,N_1932);
nand U4796 (N_4796,N_702,N_1571);
xnor U4797 (N_4797,N_2020,N_1222);
or U4798 (N_4798,N_1599,N_1946);
and U4799 (N_4799,N_527,N_2488);
nand U4800 (N_4800,N_732,N_908);
nor U4801 (N_4801,N_267,N_2155);
nor U4802 (N_4802,N_1528,N_1955);
xor U4803 (N_4803,N_302,N_996);
xnor U4804 (N_4804,N_702,N_1254);
xor U4805 (N_4805,N_250,N_1343);
nor U4806 (N_4806,N_794,N_929);
and U4807 (N_4807,N_46,N_1717);
or U4808 (N_4808,N_2303,N_1232);
nor U4809 (N_4809,N_900,N_1458);
nand U4810 (N_4810,N_2220,N_22);
nand U4811 (N_4811,N_1298,N_2001);
nand U4812 (N_4812,N_768,N_1752);
nor U4813 (N_4813,N_2348,N_353);
or U4814 (N_4814,N_1040,N_1833);
and U4815 (N_4815,N_543,N_2215);
or U4816 (N_4816,N_527,N_99);
and U4817 (N_4817,N_473,N_1965);
xnor U4818 (N_4818,N_425,N_621);
and U4819 (N_4819,N_2165,N_206);
or U4820 (N_4820,N_768,N_2416);
or U4821 (N_4821,N_2081,N_1632);
or U4822 (N_4822,N_2309,N_636);
or U4823 (N_4823,N_1411,N_355);
nor U4824 (N_4824,N_1663,N_2255);
nor U4825 (N_4825,N_589,N_2373);
and U4826 (N_4826,N_2188,N_1623);
nand U4827 (N_4827,N_729,N_734);
nor U4828 (N_4828,N_1003,N_323);
and U4829 (N_4829,N_1570,N_1812);
nand U4830 (N_4830,N_368,N_1376);
nor U4831 (N_4831,N_1336,N_1293);
nand U4832 (N_4832,N_722,N_505);
nand U4833 (N_4833,N_890,N_842);
or U4834 (N_4834,N_1552,N_2405);
nand U4835 (N_4835,N_1104,N_881);
nor U4836 (N_4836,N_2214,N_1102);
xor U4837 (N_4837,N_2117,N_1284);
and U4838 (N_4838,N_645,N_10);
or U4839 (N_4839,N_223,N_1260);
xor U4840 (N_4840,N_1259,N_828);
nor U4841 (N_4841,N_261,N_453);
and U4842 (N_4842,N_637,N_1497);
nand U4843 (N_4843,N_2317,N_981);
and U4844 (N_4844,N_52,N_907);
and U4845 (N_4845,N_16,N_771);
or U4846 (N_4846,N_147,N_1921);
nand U4847 (N_4847,N_2024,N_1209);
xor U4848 (N_4848,N_2428,N_1827);
xnor U4849 (N_4849,N_2464,N_752);
nor U4850 (N_4850,N_102,N_1672);
nand U4851 (N_4851,N_477,N_1861);
and U4852 (N_4852,N_627,N_1213);
nand U4853 (N_4853,N_2047,N_1939);
nor U4854 (N_4854,N_934,N_34);
nor U4855 (N_4855,N_230,N_20);
xnor U4856 (N_4856,N_483,N_1135);
nor U4857 (N_4857,N_713,N_199);
or U4858 (N_4858,N_1672,N_1677);
xor U4859 (N_4859,N_2127,N_1316);
and U4860 (N_4860,N_1774,N_843);
nand U4861 (N_4861,N_1442,N_945);
xor U4862 (N_4862,N_1401,N_2044);
or U4863 (N_4863,N_498,N_646);
nand U4864 (N_4864,N_1226,N_1305);
xnor U4865 (N_4865,N_1848,N_633);
and U4866 (N_4866,N_806,N_329);
nand U4867 (N_4867,N_583,N_847);
or U4868 (N_4868,N_986,N_481);
nor U4869 (N_4869,N_4,N_1437);
nand U4870 (N_4870,N_974,N_2286);
nand U4871 (N_4871,N_1817,N_464);
or U4872 (N_4872,N_1491,N_2262);
nor U4873 (N_4873,N_1259,N_1283);
or U4874 (N_4874,N_928,N_523);
nor U4875 (N_4875,N_2275,N_2305);
xor U4876 (N_4876,N_107,N_2498);
xnor U4877 (N_4877,N_2208,N_1707);
nand U4878 (N_4878,N_158,N_259);
or U4879 (N_4879,N_1528,N_2233);
and U4880 (N_4880,N_468,N_1154);
nand U4881 (N_4881,N_1365,N_1298);
nor U4882 (N_4882,N_2051,N_2050);
xnor U4883 (N_4883,N_2188,N_701);
or U4884 (N_4884,N_1644,N_2104);
or U4885 (N_4885,N_657,N_1278);
nand U4886 (N_4886,N_1888,N_93);
or U4887 (N_4887,N_1424,N_1418);
or U4888 (N_4888,N_130,N_2096);
nand U4889 (N_4889,N_841,N_1722);
and U4890 (N_4890,N_1372,N_423);
and U4891 (N_4891,N_40,N_832);
nor U4892 (N_4892,N_1169,N_635);
nand U4893 (N_4893,N_1783,N_2159);
nor U4894 (N_4894,N_658,N_992);
or U4895 (N_4895,N_1758,N_1622);
and U4896 (N_4896,N_1451,N_500);
nand U4897 (N_4897,N_296,N_1301);
or U4898 (N_4898,N_862,N_1296);
xor U4899 (N_4899,N_532,N_563);
and U4900 (N_4900,N_1889,N_193);
or U4901 (N_4901,N_1255,N_426);
or U4902 (N_4902,N_1913,N_1977);
or U4903 (N_4903,N_1662,N_1375);
or U4904 (N_4904,N_1593,N_2288);
and U4905 (N_4905,N_2111,N_1404);
nor U4906 (N_4906,N_554,N_411);
and U4907 (N_4907,N_1734,N_223);
or U4908 (N_4908,N_833,N_1260);
and U4909 (N_4909,N_1298,N_632);
nor U4910 (N_4910,N_417,N_801);
nor U4911 (N_4911,N_135,N_1546);
xnor U4912 (N_4912,N_407,N_103);
xor U4913 (N_4913,N_813,N_1687);
and U4914 (N_4914,N_1482,N_85);
nand U4915 (N_4915,N_161,N_1403);
xnor U4916 (N_4916,N_1442,N_1638);
or U4917 (N_4917,N_2251,N_2167);
nand U4918 (N_4918,N_1061,N_2485);
nand U4919 (N_4919,N_680,N_467);
and U4920 (N_4920,N_1872,N_1248);
nand U4921 (N_4921,N_2115,N_2377);
nor U4922 (N_4922,N_831,N_961);
nand U4923 (N_4923,N_1483,N_1499);
xnor U4924 (N_4924,N_1357,N_797);
nand U4925 (N_4925,N_660,N_2016);
and U4926 (N_4926,N_687,N_634);
nand U4927 (N_4927,N_612,N_1633);
nand U4928 (N_4928,N_332,N_29);
nor U4929 (N_4929,N_1262,N_1683);
nand U4930 (N_4930,N_727,N_512);
nand U4931 (N_4931,N_2011,N_1543);
nor U4932 (N_4932,N_1948,N_959);
nand U4933 (N_4933,N_22,N_1557);
and U4934 (N_4934,N_549,N_1742);
nor U4935 (N_4935,N_140,N_2422);
nand U4936 (N_4936,N_372,N_1987);
nor U4937 (N_4937,N_1744,N_2431);
nor U4938 (N_4938,N_2074,N_634);
and U4939 (N_4939,N_1044,N_429);
or U4940 (N_4940,N_350,N_363);
and U4941 (N_4941,N_959,N_2406);
xor U4942 (N_4942,N_2105,N_2298);
and U4943 (N_4943,N_396,N_603);
and U4944 (N_4944,N_2038,N_2311);
and U4945 (N_4945,N_1905,N_1000);
or U4946 (N_4946,N_1394,N_1164);
or U4947 (N_4947,N_708,N_1922);
xor U4948 (N_4948,N_2010,N_1013);
nor U4949 (N_4949,N_1125,N_849);
and U4950 (N_4950,N_1665,N_1507);
nand U4951 (N_4951,N_1178,N_712);
xnor U4952 (N_4952,N_314,N_1819);
xor U4953 (N_4953,N_2177,N_83);
or U4954 (N_4954,N_164,N_2317);
xnor U4955 (N_4955,N_1751,N_913);
and U4956 (N_4956,N_1778,N_1864);
nand U4957 (N_4957,N_166,N_2345);
nor U4958 (N_4958,N_905,N_941);
nor U4959 (N_4959,N_2251,N_1274);
or U4960 (N_4960,N_934,N_1861);
nor U4961 (N_4961,N_2224,N_581);
nand U4962 (N_4962,N_2202,N_37);
nor U4963 (N_4963,N_1692,N_432);
nor U4964 (N_4964,N_1650,N_2212);
nand U4965 (N_4965,N_1344,N_1880);
nand U4966 (N_4966,N_1339,N_443);
or U4967 (N_4967,N_60,N_1375);
or U4968 (N_4968,N_2393,N_192);
and U4969 (N_4969,N_2462,N_268);
and U4970 (N_4970,N_908,N_524);
and U4971 (N_4971,N_734,N_344);
nand U4972 (N_4972,N_1307,N_314);
xor U4973 (N_4973,N_992,N_1071);
xnor U4974 (N_4974,N_1427,N_1720);
nand U4975 (N_4975,N_1167,N_1630);
and U4976 (N_4976,N_2038,N_2134);
xnor U4977 (N_4977,N_2486,N_2154);
nor U4978 (N_4978,N_173,N_34);
or U4979 (N_4979,N_1648,N_1623);
and U4980 (N_4980,N_406,N_838);
nor U4981 (N_4981,N_1653,N_1297);
or U4982 (N_4982,N_1162,N_1674);
xor U4983 (N_4983,N_695,N_650);
and U4984 (N_4984,N_1149,N_1862);
and U4985 (N_4985,N_2336,N_2307);
or U4986 (N_4986,N_2289,N_853);
xor U4987 (N_4987,N_185,N_2100);
nor U4988 (N_4988,N_1844,N_213);
or U4989 (N_4989,N_2437,N_2351);
nor U4990 (N_4990,N_1694,N_25);
nand U4991 (N_4991,N_1069,N_503);
xor U4992 (N_4992,N_1084,N_325);
xor U4993 (N_4993,N_230,N_129);
xnor U4994 (N_4994,N_863,N_2169);
nand U4995 (N_4995,N_2047,N_598);
or U4996 (N_4996,N_496,N_55);
nor U4997 (N_4997,N_659,N_551);
xor U4998 (N_4998,N_1035,N_2362);
nor U4999 (N_4999,N_2264,N_808);
nand U5000 (N_5000,N_3998,N_3773);
xor U5001 (N_5001,N_3921,N_4434);
nand U5002 (N_5002,N_3538,N_4129);
nand U5003 (N_5003,N_2929,N_3276);
nand U5004 (N_5004,N_3487,N_4515);
and U5005 (N_5005,N_3503,N_3172);
nor U5006 (N_5006,N_3547,N_4939);
nand U5007 (N_5007,N_3979,N_4297);
and U5008 (N_5008,N_2744,N_4527);
or U5009 (N_5009,N_3382,N_2642);
nor U5010 (N_5010,N_3127,N_4153);
xor U5011 (N_5011,N_4985,N_4122);
nand U5012 (N_5012,N_2962,N_4531);
nor U5013 (N_5013,N_2707,N_4069);
xnor U5014 (N_5014,N_4646,N_2723);
nor U5015 (N_5015,N_4348,N_4758);
xnor U5016 (N_5016,N_4132,N_4102);
nand U5017 (N_5017,N_4441,N_4312);
or U5018 (N_5018,N_4231,N_4601);
and U5019 (N_5019,N_3575,N_3534);
xor U5020 (N_5020,N_3201,N_4130);
xnor U5021 (N_5021,N_2540,N_2607);
or U5022 (N_5022,N_2724,N_3595);
nor U5023 (N_5023,N_3543,N_3114);
nor U5024 (N_5024,N_4540,N_3782);
nand U5025 (N_5025,N_2823,N_3606);
or U5026 (N_5026,N_3411,N_4038);
xor U5027 (N_5027,N_4792,N_2660);
or U5028 (N_5028,N_4086,N_3392);
or U5029 (N_5029,N_3742,N_4697);
or U5030 (N_5030,N_3357,N_3031);
nand U5031 (N_5031,N_3147,N_3510);
or U5032 (N_5032,N_2507,N_2534);
and U5033 (N_5033,N_4876,N_3666);
and U5034 (N_5034,N_3884,N_4575);
and U5035 (N_5035,N_4980,N_4561);
and U5036 (N_5036,N_2947,N_3309);
xor U5037 (N_5037,N_4744,N_3369);
xor U5038 (N_5038,N_3540,N_4478);
and U5039 (N_5039,N_3067,N_3371);
nand U5040 (N_5040,N_4649,N_4904);
or U5041 (N_5041,N_3154,N_3511);
nor U5042 (N_5042,N_3610,N_3525);
nor U5043 (N_5043,N_4075,N_4556);
xor U5044 (N_5044,N_4570,N_3683);
and U5045 (N_5045,N_2579,N_4372);
nand U5046 (N_5046,N_4352,N_3562);
or U5047 (N_5047,N_3173,N_2572);
nor U5048 (N_5048,N_2968,N_2844);
xor U5049 (N_5049,N_4919,N_4710);
nor U5050 (N_5050,N_4375,N_2879);
xnor U5051 (N_5051,N_4334,N_3462);
or U5052 (N_5052,N_4296,N_4731);
or U5053 (N_5053,N_3139,N_3393);
xnor U5054 (N_5054,N_2632,N_3317);
and U5055 (N_5055,N_4573,N_3598);
xor U5056 (N_5056,N_4936,N_3810);
or U5057 (N_5057,N_4123,N_3966);
or U5058 (N_5058,N_4250,N_3638);
nand U5059 (N_5059,N_3484,N_2667);
nor U5060 (N_5060,N_4812,N_3596);
or U5061 (N_5061,N_3426,N_3640);
nand U5062 (N_5062,N_4030,N_4131);
or U5063 (N_5063,N_3539,N_2628);
and U5064 (N_5064,N_4551,N_4383);
nand U5065 (N_5065,N_3529,N_3809);
or U5066 (N_5066,N_3068,N_2917);
xor U5067 (N_5067,N_4977,N_4817);
nor U5068 (N_5068,N_2796,N_3004);
nand U5069 (N_5069,N_3675,N_4923);
xnor U5070 (N_5070,N_2626,N_4274);
and U5071 (N_5071,N_3234,N_4847);
nor U5072 (N_5072,N_4032,N_3479);
xnor U5073 (N_5073,N_4967,N_4167);
nand U5074 (N_5074,N_3604,N_3796);
nor U5075 (N_5075,N_2676,N_4475);
or U5076 (N_5076,N_4462,N_2689);
nor U5077 (N_5077,N_4143,N_4874);
or U5078 (N_5078,N_4180,N_3791);
or U5079 (N_5079,N_4740,N_3594);
nand U5080 (N_5080,N_2996,N_2564);
xor U5081 (N_5081,N_3224,N_2523);
and U5082 (N_5082,N_4076,N_3478);
xor U5083 (N_5083,N_3631,N_2892);
and U5084 (N_5084,N_4499,N_2623);
nand U5085 (N_5085,N_4861,N_4071);
and U5086 (N_5086,N_3340,N_3817);
nand U5087 (N_5087,N_2558,N_4880);
and U5088 (N_5088,N_4260,N_3203);
xor U5089 (N_5089,N_4047,N_3134);
xnor U5090 (N_5090,N_4060,N_3591);
xor U5091 (N_5091,N_2686,N_3522);
nand U5092 (N_5092,N_4626,N_3619);
nor U5093 (N_5093,N_4829,N_3308);
and U5094 (N_5094,N_3498,N_2903);
or U5095 (N_5095,N_4735,N_3280);
xor U5096 (N_5096,N_3560,N_3179);
or U5097 (N_5097,N_2663,N_3652);
nand U5098 (N_5098,N_4949,N_2598);
nand U5099 (N_5099,N_2687,N_3946);
and U5100 (N_5100,N_3999,N_2515);
and U5101 (N_5101,N_2593,N_3686);
or U5102 (N_5102,N_3326,N_2780);
xnor U5103 (N_5103,N_2567,N_2560);
xor U5104 (N_5104,N_3523,N_4893);
nand U5105 (N_5105,N_3010,N_4745);
nor U5106 (N_5106,N_3930,N_4189);
and U5107 (N_5107,N_4109,N_4748);
and U5108 (N_5108,N_3269,N_3559);
and U5109 (N_5109,N_2652,N_2910);
and U5110 (N_5110,N_3211,N_3096);
or U5111 (N_5111,N_4721,N_4222);
and U5112 (N_5112,N_4110,N_3303);
and U5113 (N_5113,N_2805,N_4770);
nor U5114 (N_5114,N_3243,N_4090);
and U5115 (N_5115,N_3993,N_4376);
and U5116 (N_5116,N_3585,N_4756);
nand U5117 (N_5117,N_4227,N_2922);
xor U5118 (N_5118,N_4835,N_3361);
and U5119 (N_5119,N_2822,N_4871);
nor U5120 (N_5120,N_3592,N_3120);
xor U5121 (N_5121,N_3703,N_3037);
or U5122 (N_5122,N_4628,N_3707);
xor U5123 (N_5123,N_3329,N_3839);
nand U5124 (N_5124,N_4544,N_3660);
and U5125 (N_5125,N_3048,N_4686);
and U5126 (N_5126,N_4908,N_4564);
xor U5127 (N_5127,N_2789,N_4722);
nand U5128 (N_5128,N_4488,N_3074);
and U5129 (N_5129,N_4332,N_4000);
and U5130 (N_5130,N_3316,N_3814);
or U5131 (N_5131,N_2672,N_3716);
or U5132 (N_5132,N_3777,N_4896);
xor U5133 (N_5133,N_4256,N_4002);
or U5134 (N_5134,N_3546,N_3358);
nand U5135 (N_5135,N_4245,N_4465);
and U5136 (N_5136,N_4738,N_3073);
xor U5137 (N_5137,N_3516,N_3651);
xor U5138 (N_5138,N_3249,N_3496);
xor U5139 (N_5139,N_4941,N_3226);
nor U5140 (N_5140,N_4307,N_4303);
and U5141 (N_5141,N_4025,N_4451);
and U5142 (N_5142,N_4327,N_4717);
or U5143 (N_5143,N_3415,N_3500);
and U5144 (N_5144,N_3821,N_4450);
nand U5145 (N_5145,N_2594,N_3138);
nand U5146 (N_5146,N_4088,N_3105);
xnor U5147 (N_5147,N_4202,N_3365);
and U5148 (N_5148,N_3701,N_3053);
or U5149 (N_5149,N_3548,N_3363);
nor U5150 (N_5150,N_4708,N_4553);
or U5151 (N_5151,N_4892,N_4435);
nand U5152 (N_5152,N_2666,N_4248);
nor U5153 (N_5153,N_3854,N_3488);
and U5154 (N_5154,N_3557,N_3163);
or U5155 (N_5155,N_4278,N_3518);
and U5156 (N_5156,N_4446,N_2920);
xor U5157 (N_5157,N_3285,N_3404);
nand U5158 (N_5158,N_2975,N_3607);
nor U5159 (N_5159,N_4747,N_2784);
xnor U5160 (N_5160,N_3008,N_3458);
xor U5161 (N_5161,N_4767,N_2927);
xor U5162 (N_5162,N_2983,N_3617);
xor U5163 (N_5163,N_4599,N_3236);
or U5164 (N_5164,N_2700,N_4331);
or U5165 (N_5165,N_4467,N_4403);
nor U5166 (N_5166,N_3279,N_4582);
or U5167 (N_5167,N_4347,N_4905);
and U5168 (N_5168,N_2706,N_4329);
xor U5169 (N_5169,N_4656,N_3865);
nor U5170 (N_5170,N_3117,N_3255);
xor U5171 (N_5171,N_3141,N_4356);
or U5172 (N_5172,N_4857,N_4511);
xnor U5173 (N_5173,N_3566,N_3264);
nand U5174 (N_5174,N_3792,N_3337);
nor U5175 (N_5175,N_3295,N_4999);
or U5176 (N_5176,N_4270,N_3808);
xnor U5177 (N_5177,N_4693,N_2646);
or U5178 (N_5178,N_4214,N_4267);
nand U5179 (N_5179,N_3251,N_4091);
or U5180 (N_5180,N_2788,N_2522);
nand U5181 (N_5181,N_4037,N_3018);
xor U5182 (N_5182,N_2682,N_4225);
nand U5183 (N_5183,N_2541,N_2504);
or U5184 (N_5184,N_2839,N_2810);
and U5185 (N_5185,N_4173,N_3876);
nor U5186 (N_5186,N_4391,N_4682);
xnor U5187 (N_5187,N_4098,N_4678);
or U5188 (N_5188,N_3978,N_4703);
nor U5189 (N_5189,N_3111,N_2872);
nand U5190 (N_5190,N_4918,N_2889);
nor U5191 (N_5191,N_2749,N_3844);
and U5192 (N_5192,N_2905,N_2665);
or U5193 (N_5193,N_4191,N_3795);
xor U5194 (N_5194,N_3681,N_4724);
nor U5195 (N_5195,N_3281,N_4164);
xnor U5196 (N_5196,N_3637,N_3881);
xor U5197 (N_5197,N_4469,N_4317);
xor U5198 (N_5198,N_4925,N_3212);
and U5199 (N_5199,N_2800,N_2685);
xnor U5200 (N_5200,N_4175,N_3204);
xnor U5201 (N_5201,N_2817,N_4978);
or U5202 (N_5202,N_2596,N_2502);
nand U5203 (N_5203,N_3167,N_3571);
xor U5204 (N_5204,N_4759,N_3233);
nor U5205 (N_5205,N_4765,N_4557);
nor U5206 (N_5206,N_3840,N_3324);
nor U5207 (N_5207,N_2690,N_4818);
xnor U5208 (N_5208,N_2843,N_4138);
or U5209 (N_5209,N_3313,N_3833);
nor U5210 (N_5210,N_3685,N_2783);
and U5211 (N_5211,N_2738,N_3104);
xnor U5212 (N_5212,N_4146,N_3422);
and U5213 (N_5213,N_3100,N_4583);
xnor U5214 (N_5214,N_3932,N_4423);
xnor U5215 (N_5215,N_4846,N_3784);
nand U5216 (N_5216,N_2831,N_4613);
or U5217 (N_5217,N_3649,N_4990);
xnor U5218 (N_5218,N_4491,N_3480);
nor U5219 (N_5219,N_3697,N_3629);
or U5220 (N_5220,N_3612,N_3661);
nand U5221 (N_5221,N_4359,N_3193);
and U5222 (N_5222,N_2734,N_4221);
nor U5223 (N_5223,N_3475,N_4052);
nand U5224 (N_5224,N_2737,N_4773);
nor U5225 (N_5225,N_4407,N_3659);
xnor U5226 (N_5226,N_2754,N_2832);
nand U5227 (N_5227,N_2520,N_3085);
nand U5228 (N_5228,N_4704,N_2824);
nor U5229 (N_5229,N_2945,N_4877);
nor U5230 (N_5230,N_2543,N_4714);
and U5231 (N_5231,N_4833,N_3799);
nand U5232 (N_5232,N_2926,N_4503);
xnor U5233 (N_5233,N_4785,N_4989);
nand U5234 (N_5234,N_4661,N_4257);
and U5235 (N_5235,N_2691,N_2739);
and U5236 (N_5236,N_3869,N_4156);
nor U5237 (N_5237,N_2852,N_2661);
and U5238 (N_5238,N_4080,N_4169);
or U5239 (N_5239,N_4067,N_4793);
or U5240 (N_5240,N_3396,N_4794);
xnor U5241 (N_5241,N_3941,N_3454);
and U5242 (N_5242,N_3191,N_2919);
xor U5243 (N_5243,N_4365,N_4866);
nor U5244 (N_5244,N_3901,N_3258);
nor U5245 (N_5245,N_4659,N_4059);
and U5246 (N_5246,N_4466,N_4652);
and U5247 (N_5247,N_3845,N_2787);
nand U5248 (N_5248,N_4565,N_4360);
and U5249 (N_5249,N_3835,N_3438);
and U5250 (N_5250,N_4720,N_3259);
nand U5251 (N_5251,N_4284,N_3348);
or U5252 (N_5252,N_3904,N_4955);
or U5253 (N_5253,N_3723,N_2894);
nor U5254 (N_5254,N_3726,N_2984);
or U5255 (N_5255,N_4473,N_4926);
and U5256 (N_5256,N_3145,N_4015);
or U5257 (N_5257,N_2518,N_4428);
and U5258 (N_5258,N_4120,N_4444);
xor U5259 (N_5259,N_3816,N_4909);
xnor U5260 (N_5260,N_3870,N_4276);
nand U5261 (N_5261,N_4101,N_3667);
nor U5262 (N_5262,N_2882,N_3239);
and U5263 (N_5263,N_4004,N_2753);
nand U5264 (N_5264,N_4723,N_3265);
nand U5265 (N_5265,N_3463,N_3729);
and U5266 (N_5266,N_3356,N_4886);
or U5267 (N_5267,N_4337,N_3984);
and U5268 (N_5268,N_4675,N_4070);
nor U5269 (N_5269,N_2538,N_3646);
or U5270 (N_5270,N_4290,N_4614);
xor U5271 (N_5271,N_4867,N_4524);
nor U5272 (N_5272,N_3272,N_3322);
nor U5273 (N_5273,N_4483,N_3058);
xor U5274 (N_5274,N_2509,N_4029);
nand U5275 (N_5275,N_4308,N_2804);
and U5276 (N_5276,N_3501,N_4558);
nor U5277 (N_5277,N_4392,N_4078);
nor U5278 (N_5278,N_2770,N_4568);
nand U5279 (N_5279,N_3602,N_4287);
and U5280 (N_5280,N_3070,N_4519);
xor U5281 (N_5281,N_2742,N_4298);
and U5282 (N_5282,N_2743,N_4803);
xnor U5283 (N_5283,N_3806,N_4969);
nor U5284 (N_5284,N_3207,N_4026);
or U5285 (N_5285,N_3938,N_3763);
xnor U5286 (N_5286,N_4258,N_2611);
or U5287 (N_5287,N_3164,N_4345);
or U5288 (N_5288,N_2684,N_4150);
or U5289 (N_5289,N_4041,N_3877);
xnor U5290 (N_5290,N_4823,N_3820);
xor U5291 (N_5291,N_4760,N_2512);
or U5292 (N_5292,N_4114,N_4368);
nand U5293 (N_5293,N_2828,N_4135);
nand U5294 (N_5294,N_4574,N_3132);
nand U5295 (N_5295,N_3097,N_4860);
and U5296 (N_5296,N_2932,N_3950);
nand U5297 (N_5297,N_3441,N_4916);
or U5298 (N_5298,N_3531,N_2972);
and U5299 (N_5299,N_4677,N_2500);
nor U5300 (N_5300,N_4636,N_3344);
nand U5301 (N_5301,N_4163,N_2931);
or U5302 (N_5302,N_4053,N_2536);
or U5303 (N_5303,N_2758,N_4580);
or U5304 (N_5304,N_3916,N_4242);
nand U5305 (N_5305,N_4160,N_3958);
xor U5306 (N_5306,N_4838,N_4797);
and U5307 (N_5307,N_2930,N_4801);
nand U5308 (N_5308,N_4679,N_3634);
or U5309 (N_5309,N_4313,N_2732);
nor U5310 (N_5310,N_4879,N_3020);
and U5311 (N_5311,N_4594,N_4251);
xor U5312 (N_5312,N_3116,N_3395);
and U5313 (N_5313,N_2835,N_4022);
nor U5314 (N_5314,N_3373,N_3533);
xnor U5315 (N_5315,N_4046,N_3714);
xnor U5316 (N_5316,N_3628,N_4044);
nor U5317 (N_5317,N_4578,N_2802);
xor U5318 (N_5318,N_4964,N_3811);
xor U5319 (N_5319,N_4863,N_3266);
xor U5320 (N_5320,N_3467,N_2547);
xnor U5321 (N_5321,N_3910,N_2963);
xor U5322 (N_5322,N_4903,N_2988);
and U5323 (N_5323,N_2830,N_2629);
xor U5324 (N_5324,N_2971,N_3323);
or U5325 (N_5325,N_3936,N_4219);
nand U5326 (N_5326,N_4431,N_3244);
and U5327 (N_5327,N_4255,N_4291);
nand U5328 (N_5328,N_3288,N_4726);
nor U5329 (N_5329,N_3033,N_3945);
xor U5330 (N_5330,N_4539,N_3248);
and U5331 (N_5331,N_2883,N_2748);
xnor U5332 (N_5332,N_4489,N_3692);
and U5333 (N_5333,N_3444,N_4453);
nor U5334 (N_5334,N_4836,N_4021);
and U5335 (N_5335,N_2938,N_3857);
or U5336 (N_5336,N_2631,N_2568);
or U5337 (N_5337,N_3690,N_4326);
nand U5338 (N_5338,N_2714,N_4933);
and U5339 (N_5339,N_3094,N_3178);
or U5340 (N_5340,N_2952,N_4358);
nand U5341 (N_5341,N_3732,N_3549);
xnor U5342 (N_5342,N_3042,N_4931);
xnor U5343 (N_5343,N_4597,N_3245);
and U5344 (N_5344,N_3554,N_3642);
nor U5345 (N_5345,N_4048,N_3747);
and U5346 (N_5346,N_4085,N_3694);
nor U5347 (N_5347,N_3590,N_3960);
nand U5348 (N_5348,N_2976,N_3355);
xor U5349 (N_5349,N_3861,N_3304);
and U5350 (N_5350,N_4424,N_2746);
and U5351 (N_5351,N_3988,N_3035);
xor U5352 (N_5352,N_3140,N_2811);
xnor U5353 (N_5353,N_2759,N_4800);
nand U5354 (N_5354,N_4897,N_2845);
nand U5355 (N_5355,N_2605,N_2985);
and U5356 (N_5356,N_4671,N_4822);
or U5357 (N_5357,N_3663,N_2969);
or U5358 (N_5358,N_3831,N_3536);
xnor U5359 (N_5359,N_4438,N_4429);
xor U5360 (N_5360,N_4657,N_4814);
nand U5361 (N_5361,N_4956,N_2840);
nor U5362 (N_5362,N_2636,N_3556);
and U5363 (N_5363,N_4463,N_2688);
and U5364 (N_5364,N_4777,N_4608);
and U5365 (N_5365,N_4912,N_3996);
or U5366 (N_5366,N_2978,N_3563);
nor U5367 (N_5367,N_4393,N_3748);
nand U5368 (N_5368,N_4602,N_3582);
or U5369 (N_5369,N_4330,N_2549);
and U5370 (N_5370,N_3768,N_3007);
nand U5371 (N_5371,N_4741,N_4304);
or U5372 (N_5372,N_3658,N_3704);
or U5373 (N_5373,N_2591,N_4145);
or U5374 (N_5374,N_4739,N_3750);
and U5375 (N_5375,N_4875,N_2981);
xnor U5376 (N_5376,N_3066,N_4286);
or U5377 (N_5377,N_3115,N_2939);
or U5378 (N_5378,N_3828,N_4713);
xnor U5379 (N_5379,N_3797,N_3353);
and U5380 (N_5380,N_3762,N_4302);
or U5381 (N_5381,N_3805,N_4269);
nor U5382 (N_5382,N_4209,N_3963);
xor U5383 (N_5383,N_4631,N_3247);
nor U5384 (N_5384,N_2608,N_3890);
xnor U5385 (N_5385,N_2681,N_4968);
xor U5386 (N_5386,N_4315,N_4552);
or U5387 (N_5387,N_2836,N_3013);
or U5388 (N_5388,N_3362,N_3072);
xor U5389 (N_5389,N_3133,N_2552);
or U5390 (N_5390,N_4292,N_4676);
nor U5391 (N_5391,N_4901,N_3453);
nor U5392 (N_5392,N_3435,N_3584);
nor U5393 (N_5393,N_2516,N_4344);
or U5394 (N_5394,N_4013,N_4295);
xnor U5395 (N_5395,N_2878,N_3919);
and U5396 (N_5396,N_2774,N_3880);
and U5397 (N_5397,N_3011,N_3914);
and U5398 (N_5398,N_3907,N_4154);
xor U5399 (N_5399,N_4957,N_3601);
nor U5400 (N_5400,N_4674,N_3195);
nor U5401 (N_5401,N_4077,N_4917);
and U5402 (N_5402,N_4839,N_4367);
nand U5403 (N_5403,N_3520,N_2812);
nor U5404 (N_5404,N_4415,N_3779);
nor U5405 (N_5405,N_3029,N_3951);
nor U5406 (N_5406,N_3026,N_3586);
and U5407 (N_5407,N_4653,N_4899);
nor U5408 (N_5408,N_3184,N_2888);
or U5409 (N_5409,N_3994,N_4484);
nor U5410 (N_5410,N_3627,N_4516);
nand U5411 (N_5411,N_2833,N_4318);
and U5412 (N_5412,N_2943,N_2948);
nor U5413 (N_5413,N_2992,N_4394);
nor U5414 (N_5414,N_3399,N_4010);
and U5415 (N_5415,N_4187,N_4033);
nor U5416 (N_5416,N_3928,N_4324);
nor U5417 (N_5417,N_4397,N_3232);
or U5418 (N_5418,N_3222,N_4878);
and U5419 (N_5419,N_4247,N_3664);
nor U5420 (N_5420,N_3108,N_4426);
or U5421 (N_5421,N_2586,N_2771);
nor U5422 (N_5422,N_4196,N_2600);
nand U5423 (N_5423,N_4548,N_3564);
xor U5424 (N_5424,N_3793,N_2864);
nor U5425 (N_5425,N_4910,N_2779);
and U5426 (N_5426,N_3380,N_4279);
xnor U5427 (N_5427,N_4709,N_4730);
nor U5428 (N_5428,N_4333,N_4854);
and U5429 (N_5429,N_2803,N_3170);
xor U5430 (N_5430,N_2793,N_3215);
or U5431 (N_5431,N_4981,N_2813);
nand U5432 (N_5432,N_3071,N_3824);
nor U5433 (N_5433,N_3146,N_3765);
and U5434 (N_5434,N_3188,N_3225);
nor U5435 (N_5435,N_3328,N_3902);
and U5436 (N_5436,N_4525,N_4668);
and U5437 (N_5437,N_3391,N_3746);
nand U5438 (N_5438,N_4537,N_3158);
xnor U5439 (N_5439,N_3064,N_4328);
nand U5440 (N_5440,N_3194,N_3032);
or U5441 (N_5441,N_4830,N_3565);
and U5442 (N_5442,N_2550,N_3431);
xnor U5443 (N_5443,N_3034,N_4152);
or U5444 (N_5444,N_3156,N_3267);
or U5445 (N_5445,N_4244,N_4927);
nand U5446 (N_5446,N_4864,N_3962);
and U5447 (N_5447,N_3384,N_3455);
or U5448 (N_5448,N_3069,N_3579);
xor U5449 (N_5449,N_3130,N_3812);
or U5450 (N_5450,N_4549,N_4210);
xor U5451 (N_5451,N_4600,N_4220);
nand U5452 (N_5452,N_3045,N_4335);
and U5453 (N_5453,N_3443,N_3088);
and U5454 (N_5454,N_3110,N_3491);
xnor U5455 (N_5455,N_4036,N_4182);
xor U5456 (N_5456,N_3470,N_2622);
and U5457 (N_5457,N_3524,N_2965);
and U5458 (N_5458,N_3494,N_3860);
and U5459 (N_5459,N_4121,N_4051);
nand U5460 (N_5460,N_3465,N_4294);
and U5461 (N_5461,N_2589,N_4508);
nor U5462 (N_5462,N_2821,N_3761);
nand U5463 (N_5463,N_2643,N_4213);
and U5464 (N_5464,N_4206,N_4766);
nor U5465 (N_5465,N_3587,N_3050);
xnor U5466 (N_5466,N_3753,N_3937);
and U5467 (N_5467,N_4610,N_2573);
and U5468 (N_5468,N_2933,N_2797);
and U5469 (N_5469,N_3403,N_2880);
nor U5470 (N_5470,N_3949,N_3414);
nor U5471 (N_5471,N_3157,N_3802);
nand U5472 (N_5472,N_3298,N_4732);
nor U5473 (N_5473,N_4859,N_4805);
nand U5474 (N_5474,N_2761,N_4117);
nor U5475 (N_5475,N_4468,N_3442);
or U5476 (N_5476,N_2935,N_4983);
xor U5477 (N_5477,N_3231,N_2993);
and U5478 (N_5478,N_4433,N_4405);
and U5479 (N_5479,N_4159,N_2987);
nor U5480 (N_5480,N_4984,N_4079);
or U5481 (N_5481,N_3553,N_4408);
and U5482 (N_5482,N_2826,N_4486);
nand U5483 (N_5483,N_4663,N_4828);
or U5484 (N_5484,N_3083,N_2525);
nor U5485 (N_5485,N_3933,N_2859);
xnor U5486 (N_5486,N_4590,N_3780);
and U5487 (N_5487,N_3128,N_3630);
nor U5488 (N_5488,N_2959,N_2548);
xor U5489 (N_5489,N_4856,N_3873);
or U5490 (N_5490,N_4973,N_4865);
nand U5491 (N_5491,N_4692,N_4343);
xor U5492 (N_5492,N_3213,N_4843);
xor U5493 (N_5493,N_3878,N_3062);
nand U5494 (N_5494,N_3052,N_4577);
or U5495 (N_5495,N_2944,N_4593);
and U5496 (N_5496,N_3800,N_3990);
or U5497 (N_5497,N_3647,N_3098);
nand U5498 (N_5498,N_2875,N_3474);
and U5499 (N_5499,N_4223,N_4736);
or U5500 (N_5500,N_3731,N_4056);
nor U5501 (N_5501,N_2953,N_4137);
nand U5502 (N_5502,N_3210,N_3137);
nor U5503 (N_5503,N_4382,N_2982);
nor U5504 (N_5504,N_3229,N_3160);
and U5505 (N_5505,N_3764,N_4226);
nor U5506 (N_5506,N_3774,N_4447);
xor U5507 (N_5507,N_3874,N_2955);
and U5508 (N_5508,N_3648,N_3014);
or U5509 (N_5509,N_4535,N_4831);
nand U5510 (N_5510,N_3489,N_4596);
nand U5511 (N_5511,N_4961,N_2635);
nand U5512 (N_5512,N_3620,N_2995);
nor U5513 (N_5513,N_4396,N_3228);
or U5514 (N_5514,N_3499,N_3680);
xnor U5515 (N_5515,N_2649,N_4824);
nand U5516 (N_5516,N_3719,N_4641);
and U5517 (N_5517,N_3103,N_3864);
or U5518 (N_5518,N_3819,N_4546);
and U5519 (N_5519,N_4340,N_2529);
nand U5520 (N_5520,N_4325,N_3333);
nor U5521 (N_5521,N_2751,N_4715);
nor U5522 (N_5522,N_4734,N_2713);
nor U5523 (N_5523,N_3532,N_2757);
xor U5524 (N_5524,N_2657,N_3693);
nor U5525 (N_5525,N_4197,N_4808);
or U5526 (N_5526,N_2966,N_2697);
xor U5527 (N_5527,N_4798,N_4211);
and U5528 (N_5528,N_2721,N_4390);
and U5529 (N_5529,N_4684,N_3788);
xor U5530 (N_5530,N_3855,N_3180);
or U5531 (N_5531,N_3485,N_4559);
nor U5532 (N_5532,N_4982,N_2901);
nor U5533 (N_5533,N_2679,N_3674);
and U5534 (N_5534,N_4476,N_3186);
nand U5535 (N_5535,N_3786,N_4224);
xnor U5536 (N_5536,N_4894,N_2818);
xor U5537 (N_5537,N_4644,N_4139);
and U5538 (N_5538,N_3364,N_3223);
and U5539 (N_5539,N_4254,N_4263);
nand U5540 (N_5540,N_3040,N_4351);
or U5541 (N_5541,N_2669,N_3397);
xor U5542 (N_5542,N_3335,N_3162);
xor U5543 (N_5543,N_4712,N_3198);
xor U5544 (N_5544,N_2532,N_2695);
nand U5545 (N_5545,N_2777,N_2842);
nand U5546 (N_5546,N_4401,N_3389);
or U5547 (N_5547,N_2767,N_4639);
nand U5548 (N_5548,N_3025,N_2856);
nor U5549 (N_5549,N_2610,N_4913);
nand U5550 (N_5550,N_4868,N_3360);
or U5551 (N_5551,N_2730,N_3508);
or U5552 (N_5552,N_4545,N_4458);
xnor U5553 (N_5553,N_3577,N_4752);
xor U5554 (N_5554,N_4914,N_3940);
xnor U5555 (N_5555,N_2881,N_2979);
nor U5556 (N_5556,N_4695,N_3541);
nand U5557 (N_5557,N_3394,N_2595);
xor U5558 (N_5558,N_3875,N_4786);
nand U5559 (N_5559,N_3668,N_4778);
xnor U5560 (N_5560,N_4618,N_3220);
nand U5561 (N_5561,N_2825,N_4772);
nor U5562 (N_5562,N_3418,N_3942);
or U5563 (N_5563,N_2637,N_3889);
nor U5564 (N_5564,N_3082,N_2768);
nand U5565 (N_5565,N_2627,N_3273);
or U5566 (N_5566,N_3580,N_4181);
nand U5567 (N_5567,N_2798,N_2571);
xor U5568 (N_5568,N_4411,N_4588);
nor U5569 (N_5569,N_3850,N_4374);
nand U5570 (N_5570,N_3754,N_3843);
nand U5571 (N_5571,N_3829,N_4144);
and U5572 (N_5572,N_2801,N_3118);
nor U5573 (N_5573,N_4494,N_2986);
xor U5574 (N_5574,N_3572,N_2924);
and U5575 (N_5575,N_4068,N_2913);
and U5576 (N_5576,N_4262,N_4366);
nor U5577 (N_5577,N_3987,N_2819);
or U5578 (N_5578,N_3155,N_4665);
nor U5579 (N_5579,N_4963,N_4825);
or U5580 (N_5580,N_3131,N_3165);
or U5581 (N_5581,N_2645,N_3803);
xor U5582 (N_5582,N_2705,N_4142);
nand U5583 (N_5583,N_2760,N_4355);
nor U5584 (N_5584,N_3903,N_3113);
xnor U5585 (N_5585,N_3406,N_4207);
nor U5586 (N_5586,N_2750,N_2702);
or U5587 (N_5587,N_2782,N_4997);
nand U5588 (N_5588,N_3240,N_3838);
or U5589 (N_5589,N_4095,N_4509);
and U5590 (N_5590,N_3515,N_4791);
or U5591 (N_5591,N_2861,N_3402);
nand U5592 (N_5592,N_3856,N_4994);
or U5593 (N_5593,N_3551,N_3567);
and U5594 (N_5594,N_2556,N_4788);
nor U5595 (N_5595,N_2765,N_3804);
xor U5596 (N_5596,N_4113,N_4520);
nor U5597 (N_5597,N_4115,N_3775);
nand U5598 (N_5598,N_3202,N_3284);
or U5599 (N_5599,N_3989,N_4502);
nor U5600 (N_5600,N_3078,N_4935);
and U5601 (N_5601,N_4073,N_4342);
and U5602 (N_5602,N_3770,N_3625);
and U5603 (N_5603,N_3268,N_2863);
nand U5604 (N_5604,N_4986,N_3918);
and U5605 (N_5605,N_2592,N_4495);
and U5606 (N_5606,N_4199,N_4413);
or U5607 (N_5607,N_3934,N_2816);
and U5608 (N_5608,N_3975,N_4259);
xnor U5609 (N_5609,N_3905,N_4065);
nor U5610 (N_5610,N_3262,N_4057);
and U5611 (N_5611,N_3433,N_3076);
and U5612 (N_5612,N_4461,N_4834);
nor U5613 (N_5613,N_4338,N_4100);
or U5614 (N_5614,N_3851,N_2735);
and U5615 (N_5615,N_3457,N_3908);
nand U5616 (N_5616,N_3182,N_4457);
nor U5617 (N_5617,N_3460,N_4399);
and U5618 (N_5618,N_3842,N_4119);
nand U5619 (N_5619,N_3818,N_3679);
or U5620 (N_5620,N_3336,N_3175);
nor U5621 (N_5621,N_4719,N_4034);
nand U5622 (N_5622,N_3558,N_3574);
xor U5623 (N_5623,N_4606,N_2918);
and U5624 (N_5624,N_4104,N_4603);
nor U5625 (N_5625,N_4445,N_2728);
nand U5626 (N_5626,N_2950,N_3325);
nor U5627 (N_5627,N_4176,N_4107);
or U5628 (N_5628,N_3787,N_3971);
nand U5629 (N_5629,N_3187,N_3722);
xnor U5630 (N_5630,N_3862,N_4815);
or U5631 (N_5631,N_4586,N_4707);
and U5632 (N_5632,N_3408,N_4971);
nand U5633 (N_5633,N_4112,N_2624);
nor U5634 (N_5634,N_3370,N_2555);
nand U5635 (N_5635,N_4097,N_4240);
nor U5636 (N_5636,N_2874,N_4289);
or U5637 (N_5637,N_3057,N_3238);
and U5638 (N_5638,N_3124,N_3471);
nor U5639 (N_5639,N_4323,N_4311);
nor U5640 (N_5640,N_3696,N_4930);
nor U5641 (N_5641,N_3603,N_4900);
xor U5642 (N_5642,N_2650,N_2890);
nand U5643 (N_5643,N_4230,N_3003);
and U5644 (N_5644,N_3935,N_3982);
xor U5645 (N_5645,N_3961,N_3717);
xor U5646 (N_5646,N_4430,N_2912);
and U5647 (N_5647,N_4094,N_4655);
nor U5648 (N_5648,N_4008,N_3036);
and U5649 (N_5649,N_3079,N_4960);
or U5650 (N_5650,N_4201,N_4650);
nor U5651 (N_5651,N_3206,N_3286);
nand U5652 (N_5652,N_2618,N_3509);
nor U5653 (N_5653,N_2887,N_2647);
and U5654 (N_5654,N_4007,N_3912);
nand U5655 (N_5655,N_4522,N_3388);
and U5656 (N_5656,N_3473,N_4689);
or U5657 (N_5657,N_4554,N_3429);
and U5658 (N_5658,N_4288,N_2958);
xnor U5659 (N_5659,N_3605,N_4911);
xor U5660 (N_5660,N_3655,N_4379);
nor U5661 (N_5661,N_2641,N_4996);
and U5662 (N_5662,N_2980,N_3450);
nand U5663 (N_5663,N_3006,N_2991);
and U5664 (N_5664,N_2906,N_3305);
xor U5665 (N_5665,N_3695,N_2673);
and U5666 (N_5666,N_3778,N_4093);
or U5667 (N_5667,N_4377,N_4809);
nor U5668 (N_5668,N_4023,N_4517);
and U5669 (N_5669,N_4412,N_4281);
nor U5670 (N_5670,N_3713,N_3507);
and U5671 (N_5671,N_3923,N_3636);
nand U5672 (N_5672,N_4099,N_4543);
or U5673 (N_5673,N_2583,N_3366);
nand U5674 (N_5674,N_3641,N_4774);
xnor U5675 (N_5675,N_3046,N_4363);
and U5676 (N_5676,N_4779,N_4638);
or U5677 (N_5677,N_3801,N_4195);
nand U5678 (N_5678,N_3001,N_2876);
nor U5679 (N_5679,N_4481,N_2514);
nor U5680 (N_5680,N_3283,N_4253);
xor U5681 (N_5681,N_2763,N_4124);
or U5682 (N_5682,N_3711,N_3315);
nor U5683 (N_5683,N_3621,N_4660);
xnor U5684 (N_5684,N_3836,N_4648);
and U5685 (N_5685,N_2625,N_3521);
nor U5686 (N_5686,N_4929,N_4306);
nand U5687 (N_5687,N_4208,N_4532);
nor U5688 (N_5688,N_4542,N_3623);
or U5689 (N_5689,N_4921,N_4706);
nand U5690 (N_5690,N_3997,N_4699);
and U5691 (N_5691,N_2701,N_4581);
xor U5692 (N_5692,N_4161,N_3611);
nor U5693 (N_5693,N_2527,N_3502);
xor U5694 (N_5694,N_3282,N_3688);
nand U5695 (N_5695,N_3759,N_3024);
nand U5696 (N_5696,N_3955,N_4538);
or U5697 (N_5697,N_4615,N_3409);
and U5698 (N_5698,N_2506,N_4193);
and U5699 (N_5699,N_4460,N_3334);
xor U5700 (N_5700,N_2606,N_4536);
nand U5701 (N_5701,N_4849,N_2900);
nor U5702 (N_5702,N_3926,N_3506);
and U5703 (N_5703,N_4157,N_3447);
nand U5704 (N_5704,N_4009,N_3419);
and U5705 (N_5705,N_3209,N_2778);
nor U5706 (N_5706,N_3871,N_2587);
xnor U5707 (N_5707,N_4621,N_3060);
or U5708 (N_5708,N_4204,N_2530);
or U5709 (N_5709,N_3720,N_4234);
xnor U5710 (N_5710,N_3956,N_4796);
and U5711 (N_5711,N_2849,N_3112);
xor U5712 (N_5712,N_2741,N_3527);
or U5713 (N_5713,N_4992,N_3600);
nand U5714 (N_5714,N_4512,N_3832);
nand U5715 (N_5715,N_3174,N_2615);
and U5716 (N_5716,N_3519,N_3084);
or U5717 (N_5717,N_3448,N_4906);
xnor U5718 (N_5718,N_2868,N_4178);
or U5719 (N_5719,N_3841,N_4518);
xnor U5720 (N_5720,N_2940,N_3376);
nor U5721 (N_5721,N_4229,N_4504);
xnor U5722 (N_5722,N_3689,N_2696);
and U5723 (N_5723,N_3665,N_3481);
nor U5724 (N_5724,N_4237,N_3639);
xor U5725 (N_5725,N_4485,N_2597);
xnor U5726 (N_5726,N_2851,N_3119);
xor U5727 (N_5727,N_4106,N_2756);
or U5728 (N_5728,N_3466,N_4687);
or U5729 (N_5729,N_3166,N_2510);
or U5730 (N_5730,N_3662,N_2535);
nand U5731 (N_5731,N_3030,N_3657);
or U5732 (N_5732,N_2582,N_4887);
nand U5733 (N_5733,N_3924,N_3049);
nand U5734 (N_5734,N_3387,N_4349);
and U5735 (N_5735,N_3256,N_3410);
or U5736 (N_5736,N_4369,N_2717);
nor U5737 (N_5737,N_3512,N_4922);
xnor U5738 (N_5738,N_3785,N_2620);
or U5739 (N_5739,N_4126,N_2893);
nand U5740 (N_5740,N_4371,N_3917);
xnor U5741 (N_5741,N_3743,N_4228);
or U5742 (N_5742,N_4948,N_4762);
xor U5743 (N_5743,N_2997,N_3294);
nand U5744 (N_5744,N_4243,N_3656);
or U5745 (N_5745,N_3277,N_4934);
or U5746 (N_5746,N_4872,N_4380);
or U5747 (N_5747,N_3367,N_3437);
nand U5748 (N_5748,N_2674,N_4958);
or U5749 (N_5749,N_4541,N_3985);
nand U5750 (N_5750,N_4386,N_4001);
nor U5751 (N_5751,N_4625,N_3321);
or U5752 (N_5752,N_4776,N_3517);
nand U5753 (N_5753,N_4319,N_2569);
nor U5754 (N_5754,N_4218,N_4148);
nand U5755 (N_5755,N_2921,N_3129);
and U5756 (N_5756,N_2640,N_4592);
nor U5757 (N_5757,N_2846,N_3297);
xor U5758 (N_5758,N_2873,N_2908);
or U5759 (N_5759,N_4136,N_4705);
and U5760 (N_5760,N_3090,N_3401);
xnor U5761 (N_5761,N_3483,N_2867);
or U5762 (N_5762,N_3745,N_3086);
and U5763 (N_5763,N_3087,N_4569);
xor U5764 (N_5764,N_4664,N_4804);
nand U5765 (N_5765,N_3350,N_2693);
nand U5766 (N_5766,N_2899,N_4216);
or U5767 (N_5767,N_2577,N_2588);
and U5768 (N_5768,N_3991,N_3897);
or U5769 (N_5769,N_4534,N_4995);
and U5770 (N_5770,N_3189,N_4236);
and U5771 (N_5771,N_4395,N_4604);
xnor U5772 (N_5772,N_3530,N_3739);
xor U5773 (N_5773,N_2616,N_3235);
nor U5774 (N_5774,N_4769,N_2941);
nand U5775 (N_5775,N_4127,N_3973);
nor U5776 (N_5776,N_3981,N_2662);
xnor U5777 (N_5777,N_2675,N_2961);
and U5778 (N_5778,N_4579,N_4198);
or U5779 (N_5779,N_2513,N_3253);
nand U5780 (N_5780,N_3849,N_3915);
and U5781 (N_5781,N_3177,N_2764);
nor U5782 (N_5782,N_3214,N_3834);
or U5783 (N_5783,N_4273,N_3459);
or U5784 (N_5784,N_4743,N_3301);
nand U5785 (N_5785,N_4174,N_4826);
or U5786 (N_5786,N_3737,N_4998);
xnor U5787 (N_5787,N_4378,N_2658);
nand U5788 (N_5788,N_3299,N_4232);
and U5789 (N_5789,N_3432,N_4662);
and U5790 (N_5790,N_2858,N_3866);
or U5791 (N_5791,N_4238,N_4976);
or U5792 (N_5792,N_3867,N_3767);
xnor U5793 (N_5793,N_2574,N_3221);
nor U5794 (N_5794,N_3171,N_2542);
xor U5795 (N_5795,N_2590,N_3772);
nor U5796 (N_5796,N_4975,N_2829);
and U5797 (N_5797,N_4533,N_3196);
and U5798 (N_5798,N_2973,N_3092);
nand U5799 (N_5799,N_4420,N_3751);
nor U5800 (N_5800,N_3733,N_3123);
xnor U5801 (N_5801,N_3526,N_2809);
nand U5802 (N_5802,N_2671,N_3913);
nand U5803 (N_5803,N_3813,N_2517);
and U5804 (N_5804,N_2736,N_3755);
xor U5805 (N_5805,N_3972,N_4584);
and U5806 (N_5806,N_4011,N_4885);
or U5807 (N_5807,N_3614,N_4888);
xor U5808 (N_5808,N_2578,N_4322);
nor U5809 (N_5809,N_2954,N_3227);
nand U5810 (N_5810,N_4750,N_3699);
nand U5811 (N_5811,N_3965,N_2837);
nor U5812 (N_5812,N_4116,N_4842);
xnor U5813 (N_5813,N_4920,N_4072);
nor U5814 (N_5814,N_4783,N_2698);
nor U5815 (N_5815,N_4272,N_2915);
or U5816 (N_5816,N_2806,N_4436);
nand U5817 (N_5817,N_4118,N_2928);
or U5818 (N_5818,N_4691,N_4035);
and U5819 (N_5819,N_4498,N_4373);
xnor U5820 (N_5820,N_3218,N_4249);
and U5821 (N_5821,N_2722,N_3216);
nand U5822 (N_5822,N_2923,N_3341);
xor U5823 (N_5823,N_4853,N_4179);
xnor U5824 (N_5824,N_4300,N_4045);
nor U5825 (N_5825,N_4275,N_4953);
nand U5826 (N_5826,N_3920,N_4084);
nand U5827 (N_5827,N_2820,N_2699);
xnor U5828 (N_5828,N_2790,N_2781);
or U5829 (N_5829,N_4852,N_4816);
xnor U5830 (N_5830,N_2847,N_4733);
or U5831 (N_5831,N_4789,N_4477);
xnor U5832 (N_5832,N_3671,N_4685);
or U5833 (N_5833,N_2848,N_4265);
xor U5834 (N_5834,N_4669,N_3368);
nand U5835 (N_5835,N_3017,N_2565);
nor U5836 (N_5836,N_2559,N_3756);
xor U5837 (N_5837,N_4321,N_3126);
nand U5838 (N_5838,N_4576,N_4282);
xor U5839 (N_5839,N_4806,N_4902);
nor U5840 (N_5840,N_2869,N_2519);
nor U5841 (N_5841,N_3807,N_4133);
or U5842 (N_5842,N_3537,N_4629);
or U5843 (N_5843,N_4299,N_2807);
nand U5844 (N_5844,N_3039,N_2727);
nand U5845 (N_5845,N_4521,N_4168);
nand U5846 (N_5846,N_4645,N_4683);
xnor U5847 (N_5847,N_2576,N_3900);
and U5848 (N_5848,N_3237,N_3390);
nor U5849 (N_5849,N_4974,N_3853);
xor U5850 (N_5850,N_3676,N_4346);
and U5851 (N_5851,N_2566,N_3896);
nor U5852 (N_5852,N_4844,N_3486);
nor U5853 (N_5853,N_3449,N_2841);
nor U5854 (N_5854,N_2659,N_3250);
nor U5855 (N_5855,N_3065,N_3677);
nand U5856 (N_5856,N_3497,N_3080);
nand U5857 (N_5857,N_4184,N_4514);
or U5858 (N_5858,N_3758,N_2602);
nor U5859 (N_5859,N_3514,N_3544);
nor U5860 (N_5860,N_4884,N_4666);
or U5861 (N_5861,N_4402,N_2785);
or U5862 (N_5862,N_3708,N_4510);
or U5863 (N_5863,N_4310,N_2865);
nand U5864 (N_5864,N_4718,N_2942);
nor U5865 (N_5865,N_4361,N_2654);
and U5866 (N_5866,N_3143,N_4018);
nor U5867 (N_5867,N_2731,N_3091);
xor U5868 (N_5868,N_3477,N_4314);
nor U5869 (N_5869,N_3135,N_4353);
xnor U5870 (N_5870,N_2773,N_4749);
or U5871 (N_5871,N_3476,N_2561);
nor U5872 (N_5872,N_3205,N_3597);
or U5873 (N_5873,N_3482,N_4480);
xnor U5874 (N_5874,N_3730,N_3106);
and U5875 (N_5875,N_3847,N_3290);
or U5876 (N_5876,N_4725,N_2655);
nand U5877 (N_5877,N_2668,N_2537);
nor U5878 (N_5878,N_4694,N_3495);
nor U5879 (N_5879,N_2692,N_3456);
nor U5880 (N_5880,N_4681,N_2814);
nor U5881 (N_5881,N_3102,N_4562);
nand U5882 (N_5882,N_3898,N_4419);
nor U5883 (N_5883,N_4063,N_4364);
nor U5884 (N_5884,N_2562,N_4239);
xnor U5885 (N_5885,N_3469,N_3593);
or U5886 (N_5886,N_3825,N_2795);
or U5887 (N_5887,N_3650,N_2563);
and U5888 (N_5888,N_3242,N_4493);
nor U5889 (N_5889,N_4140,N_4414);
xor U5890 (N_5890,N_3721,N_4607);
or U5891 (N_5891,N_4404,N_3948);
or U5892 (N_5892,N_4459,N_3109);
or U5893 (N_5893,N_2630,N_3047);
nor U5894 (N_5894,N_2521,N_4632);
and U5895 (N_5895,N_3528,N_2956);
nor U5896 (N_5896,N_4742,N_3306);
or U5897 (N_5897,N_3504,N_4452);
and U5898 (N_5898,N_4024,N_2554);
or U5899 (N_5899,N_3826,N_4066);
nand U5900 (N_5900,N_4889,N_3275);
and U5901 (N_5901,N_3152,N_4965);
nor U5902 (N_5902,N_3254,N_3678);
and U5903 (N_5903,N_3883,N_3330);
and U5904 (N_5904,N_3021,N_3561);
xnor U5905 (N_5905,N_3752,N_2853);
or U5906 (N_5906,N_4943,N_2854);
nand U5907 (N_5907,N_3425,N_3347);
nand U5908 (N_5908,N_3947,N_3569);
and U5909 (N_5909,N_2539,N_4673);
and U5910 (N_5910,N_2581,N_2639);
xor U5911 (N_5911,N_3252,N_4185);
or U5912 (N_5912,N_4507,N_4855);
nand U5913 (N_5913,N_2896,N_2904);
nand U5914 (N_5914,N_3944,N_3413);
nand U5915 (N_5915,N_2694,N_3859);
nor U5916 (N_5916,N_4690,N_3552);
nand U5917 (N_5917,N_3911,N_3706);
nand U5918 (N_5918,N_3827,N_4050);
nor U5919 (N_5919,N_3766,N_3142);
xnor U5920 (N_5920,N_3359,N_3957);
nor U5921 (N_5921,N_4932,N_2545);
or U5922 (N_5922,N_2998,N_3888);
nor U5923 (N_5923,N_4111,N_4764);
nor U5924 (N_5924,N_4790,N_3176);
and U5925 (N_5925,N_4039,N_3217);
xnor U5926 (N_5926,N_3776,N_3012);
or U5927 (N_5927,N_2677,N_4716);
xor U5928 (N_5928,N_4427,N_3343);
nand U5929 (N_5929,N_3246,N_4555);
nand U5930 (N_5930,N_4799,N_3434);
xor U5931 (N_5931,N_3009,N_4907);
and U5932 (N_5932,N_4437,N_4696);
or U5933 (N_5933,N_2551,N_3725);
or U5934 (N_5934,N_4566,N_3626);
or U5935 (N_5935,N_3670,N_4820);
nand U5936 (N_5936,N_3342,N_4040);
xnor U5937 (N_5937,N_3608,N_4819);
nor U5938 (N_5938,N_4370,N_3015);
xor U5939 (N_5939,N_4737,N_2791);
nor U5940 (N_5940,N_3943,N_4841);
xnor U5941 (N_5941,N_3099,N_3043);
or U5942 (N_5942,N_4280,N_4064);
nor U5943 (N_5943,N_4246,N_3063);
or U5944 (N_5944,N_4339,N_3439);
xnor U5945 (N_5945,N_2960,N_3891);
and U5946 (N_5946,N_3331,N_2974);
nor U5947 (N_5947,N_2916,N_3122);
nor U5948 (N_5948,N_4261,N_2557);
nand U5949 (N_5949,N_4354,N_2718);
xor U5950 (N_5950,N_4305,N_3107);
and U5951 (N_5951,N_2871,N_2508);
xor U5952 (N_5952,N_4456,N_2644);
xnor U5953 (N_5953,N_2570,N_4928);
and U5954 (N_5954,N_4028,N_3925);
or U5955 (N_5955,N_3101,N_3794);
nor U5956 (N_5956,N_4881,N_2855);
xnor U5957 (N_5957,N_3744,N_4108);
xor U5958 (N_5958,N_4617,N_3909);
or U5959 (N_5959,N_4784,N_3682);
xor U5960 (N_5960,N_2716,N_4620);
and U5961 (N_5961,N_2653,N_3954);
nand U5962 (N_5962,N_3150,N_4087);
and U5963 (N_5963,N_3492,N_2914);
nor U5964 (N_5964,N_3624,N_4585);
nor U5965 (N_5965,N_2712,N_3576);
or U5966 (N_5966,N_4285,N_3420);
or U5967 (N_5967,N_3310,N_3879);
xnor U5968 (N_5968,N_2633,N_2680);
nand U5969 (N_5969,N_4350,N_3339);
nor U5970 (N_5970,N_4074,N_4500);
nand U5971 (N_5971,N_2951,N_4547);
or U5972 (N_5972,N_3848,N_2524);
nor U5973 (N_5973,N_2747,N_4200);
xor U5974 (N_5974,N_4151,N_3241);
nor U5975 (N_5975,N_3798,N_2990);
or U5976 (N_5976,N_3199,N_4640);
and U5977 (N_5977,N_3445,N_3332);
and U5978 (N_5978,N_4268,N_4858);
and U5979 (N_5979,N_4627,N_4755);
xnor U5980 (N_5980,N_4751,N_4560);
xnor U5981 (N_5981,N_3669,N_2634);
nand U5982 (N_5982,N_3976,N_3822);
xnor U5983 (N_5983,N_3724,N_4727);
or U5984 (N_5984,N_2651,N_2533);
nor U5985 (N_5985,N_4821,N_4417);
nor U5986 (N_5986,N_4103,N_4398);
nand U5987 (N_5987,N_2884,N_4205);
or U5988 (N_5988,N_3159,N_3644);
or U5989 (N_5989,N_3314,N_3440);
and U5990 (N_5990,N_2862,N_3741);
nor U5991 (N_5991,N_3992,N_4496);
nand U5992 (N_5992,N_4012,N_4530);
and U5993 (N_5993,N_3581,N_4432);
or U5994 (N_5994,N_4166,N_4529);
xnor U5995 (N_5995,N_3589,N_2815);
xnor U5996 (N_5996,N_3421,N_2838);
xnor U5997 (N_5997,N_4634,N_3263);
xnor U5998 (N_5998,N_3261,N_4252);
and U5999 (N_5999,N_3852,N_4440);
nor U6000 (N_6000,N_4506,N_4016);
nor U6001 (N_6001,N_3041,N_4054);
nand U6002 (N_6002,N_3632,N_4439);
or U6003 (N_6003,N_2740,N_4563);
or U6004 (N_6004,N_3892,N_3830);
nor U6005 (N_6005,N_3749,N_2619);
or U6006 (N_6006,N_4271,N_4155);
and U6007 (N_6007,N_2584,N_3378);
and U6008 (N_6008,N_3002,N_3710);
or U6009 (N_6009,N_3728,N_2526);
nor U6010 (N_6010,N_3312,N_2531);
nor U6011 (N_6011,N_2720,N_4869);
nand U6012 (N_6012,N_3691,N_2601);
and U6013 (N_6013,N_3570,N_3757);
or U6014 (N_6014,N_2704,N_4388);
or U6015 (N_6015,N_3684,N_4528);
and U6016 (N_6016,N_2794,N_2575);
nor U6017 (N_6017,N_4092,N_2664);
nand U6018 (N_6018,N_3700,N_2870);
xor U6019 (N_6019,N_3882,N_2585);
xor U6020 (N_6020,N_2909,N_4763);
nor U6021 (N_6021,N_3318,N_3136);
nand U6022 (N_6022,N_3144,N_3653);
xor U6023 (N_6023,N_3023,N_3643);
nor U6024 (N_6024,N_2719,N_3846);
xor U6025 (N_6025,N_2776,N_2715);
nor U6026 (N_6026,N_2877,N_4017);
nand U6027 (N_6027,N_2612,N_4505);
xor U6028 (N_6028,N_4171,N_4389);
xnor U6029 (N_6029,N_4651,N_3377);
or U6030 (N_6030,N_3181,N_3687);
nor U6031 (N_6031,N_4970,N_3952);
nor U6032 (N_6032,N_2621,N_4771);
nor U6033 (N_6033,N_3974,N_3028);
nor U6034 (N_6034,N_4598,N_4497);
and U6035 (N_6035,N_2711,N_3760);
nand U6036 (N_6036,N_4192,N_4061);
nor U6037 (N_6037,N_3970,N_3735);
or U6038 (N_6038,N_3790,N_3185);
and U6039 (N_6039,N_3769,N_3000);
nor U6040 (N_6040,N_4523,N_2503);
or U6041 (N_6041,N_2772,N_3464);
nand U6042 (N_6042,N_3709,N_2580);
nor U6043 (N_6043,N_2957,N_3059);
and U6044 (N_6044,N_4979,N_4134);
or U6045 (N_6045,N_3296,N_3615);
or U6046 (N_6046,N_4938,N_4951);
xnor U6047 (N_6047,N_3823,N_3583);
nand U6048 (N_6048,N_2850,N_3931);
nand U6049 (N_6049,N_4950,N_3044);
and U6050 (N_6050,N_3715,N_3352);
xor U6051 (N_6051,N_3051,N_4915);
xnor U6052 (N_6052,N_4630,N_4357);
nand U6053 (N_6053,N_2911,N_2609);
or U6054 (N_6054,N_3789,N_3738);
nand U6055 (N_6055,N_3346,N_3461);
and U6056 (N_6056,N_4782,N_2544);
nor U6057 (N_6057,N_3868,N_4947);
nor U6058 (N_6058,N_3542,N_3505);
and U6059 (N_6059,N_3654,N_4616);
or U6060 (N_6060,N_2683,N_4058);
xnor U6061 (N_6061,N_3490,N_3599);
and U6062 (N_6062,N_4567,N_4049);
and U6063 (N_6063,N_3054,N_4487);
or U6064 (N_6064,N_4513,N_4027);
or U6065 (N_6065,N_4031,N_4611);
or U6066 (N_6066,N_3906,N_3190);
and U6067 (N_6067,N_4811,N_4442);
nand U6068 (N_6068,N_3320,N_2946);
or U6069 (N_6069,N_2902,N_4474);
and U6070 (N_6070,N_4924,N_4945);
and U6071 (N_6071,N_4991,N_3405);
nand U6072 (N_6072,N_3428,N_3969);
or U6073 (N_6073,N_4501,N_2599);
nor U6074 (N_6074,N_4754,N_3858);
xnor U6075 (N_6075,N_2886,N_3673);
xor U6076 (N_6076,N_4768,N_3125);
xor U6077 (N_6077,N_3345,N_4081);
xnor U6078 (N_6078,N_3300,N_4472);
nor U6079 (N_6079,N_3452,N_4571);
nor U6080 (N_6080,N_3588,N_4624);
nand U6081 (N_6081,N_3372,N_4410);
and U6082 (N_6082,N_4188,N_4055);
or U6083 (N_6083,N_2603,N_4384);
xnor U6084 (N_6084,N_3430,N_4105);
nor U6085 (N_6085,N_3886,N_2656);
nand U6086 (N_6086,N_4572,N_4320);
nand U6087 (N_6087,N_2511,N_4089);
or U6088 (N_6088,N_3121,N_4125);
nand U6089 (N_6089,N_3837,N_4381);
xnor U6090 (N_6090,N_3929,N_4890);
nor U6091 (N_6091,N_2866,N_4406);
nor U6092 (N_6092,N_2834,N_3168);
nand U6093 (N_6093,N_3383,N_3056);
and U6094 (N_6094,N_4019,N_3148);
nand U6095 (N_6095,N_4848,N_3734);
or U6096 (N_6096,N_4972,N_3278);
and U6097 (N_6097,N_3986,N_3922);
nand U6098 (N_6098,N_3635,N_2766);
and U6099 (N_6099,N_4622,N_2709);
and U6100 (N_6100,N_3271,N_3959);
nor U6101 (N_6101,N_3400,N_3354);
nor U6102 (N_6102,N_2885,N_4183);
or U6103 (N_6103,N_4891,N_2614);
xor U6104 (N_6104,N_4882,N_3885);
nor U6105 (N_6105,N_3712,N_4471);
xor U6106 (N_6106,N_4761,N_2808);
xnor U6107 (N_6107,N_4217,N_4635);
xnor U6108 (N_6108,N_2907,N_2501);
and U6109 (N_6109,N_4862,N_3019);
and U6110 (N_6110,N_2857,N_4233);
or U6111 (N_6111,N_4688,N_4595);
nand U6112 (N_6112,N_3983,N_3702);
or U6113 (N_6113,N_2769,N_4966);
and U6114 (N_6114,N_3287,N_3578);
and U6115 (N_6115,N_4895,N_3386);
and U6116 (N_6116,N_2895,N_2762);
nand U6117 (N_6117,N_3927,N_3740);
xor U6118 (N_6118,N_4654,N_4162);
or U6119 (N_6119,N_3894,N_3815);
and U6120 (N_6120,N_3980,N_4309);
nand U6121 (N_6121,N_2977,N_4873);
and U6122 (N_6122,N_4165,N_4845);
or U6123 (N_6123,N_3964,N_3291);
and U6124 (N_6124,N_4942,N_3727);
nand U6125 (N_6125,N_4042,N_4062);
nand U6126 (N_6126,N_4959,N_4526);
xnor U6127 (N_6127,N_3412,N_2546);
xor U6128 (N_6128,N_4944,N_2786);
and U6129 (N_6129,N_4416,N_3005);
or U6130 (N_6130,N_4946,N_4005);
and U6131 (N_6131,N_3618,N_4454);
xnor U6132 (N_6132,N_3061,N_3307);
and U6133 (N_6133,N_4840,N_3385);
nor U6134 (N_6134,N_3977,N_4186);
nor U6135 (N_6135,N_3545,N_4647);
xnor U6136 (N_6136,N_3872,N_3200);
nor U6137 (N_6137,N_3398,N_4470);
xnor U6138 (N_6138,N_4729,N_3260);
xor U6139 (N_6139,N_3416,N_4482);
xnor U6140 (N_6140,N_4807,N_4425);
or U6141 (N_6141,N_3718,N_3446);
nor U6142 (N_6142,N_4795,N_2994);
nor U6143 (N_6143,N_2745,N_4387);
or U6144 (N_6144,N_4455,N_2755);
nand U6145 (N_6145,N_4194,N_4810);
or U6146 (N_6146,N_4190,N_4448);
or U6147 (N_6147,N_2528,N_2648);
and U6148 (N_6148,N_2638,N_4658);
nor U6149 (N_6149,N_4746,N_3089);
and U6150 (N_6150,N_4385,N_4605);
xor U6151 (N_6151,N_3183,N_4832);
xnor U6152 (N_6152,N_4449,N_3609);
xor U6153 (N_6153,N_2725,N_4667);
and U6154 (N_6154,N_4293,N_3192);
and U6155 (N_6155,N_3161,N_4619);
nand U6156 (N_6156,N_2678,N_3077);
nand U6157 (N_6157,N_2970,N_4096);
or U6158 (N_6158,N_4014,N_4813);
or U6159 (N_6159,N_4802,N_4421);
xnor U6160 (N_6160,N_3899,N_4043);
and U6161 (N_6161,N_4728,N_3781);
nor U6162 (N_6162,N_4141,N_4336);
nand U6163 (N_6163,N_4409,N_4203);
and U6164 (N_6164,N_3095,N_2604);
xor U6165 (N_6165,N_4623,N_4643);
xnor U6166 (N_6166,N_3153,N_4479);
nand U6167 (N_6167,N_3895,N_4870);
nor U6168 (N_6168,N_3381,N_4837);
xnor U6169 (N_6169,N_4277,N_3887);
or U6170 (N_6170,N_3351,N_2752);
xor U6171 (N_6171,N_4591,N_3672);
nand U6172 (N_6172,N_3893,N_3257);
and U6173 (N_6173,N_4264,N_4128);
or U6174 (N_6174,N_2726,N_3622);
and U6175 (N_6175,N_2613,N_3513);
or U6176 (N_6176,N_4701,N_4177);
nand U6177 (N_6177,N_3550,N_2897);
nand U6178 (N_6178,N_3197,N_3995);
or U6179 (N_6179,N_3568,N_4787);
nand U6180 (N_6180,N_3783,N_3374);
xnor U6181 (N_6181,N_3292,N_3327);
or U6182 (N_6182,N_3417,N_3270);
nor U6183 (N_6183,N_4215,N_3451);
nor U6184 (N_6184,N_2505,N_3645);
xor U6185 (N_6185,N_4952,N_3472);
and U6186 (N_6186,N_4954,N_2670);
nand U6187 (N_6187,N_3468,N_4589);
nand U6188 (N_6188,N_4172,N_4464);
xnor U6189 (N_6189,N_3698,N_3705);
nand U6190 (N_6190,N_3407,N_2617);
or U6191 (N_6191,N_4083,N_4962);
xor U6192 (N_6192,N_4698,N_3151);
or U6193 (N_6193,N_4612,N_3075);
and U6194 (N_6194,N_3573,N_2775);
nor U6195 (N_6195,N_3424,N_3613);
xnor U6196 (N_6196,N_4609,N_3016);
xnor U6197 (N_6197,N_4587,N_4781);
and U6198 (N_6198,N_4212,N_2949);
or U6199 (N_6199,N_4341,N_4993);
and U6200 (N_6200,N_3208,N_4827);
or U6201 (N_6201,N_4637,N_3027);
nand U6202 (N_6202,N_4006,N_4757);
xnor U6203 (N_6203,N_3093,N_3968);
nor U6204 (N_6204,N_2860,N_3616);
nand U6205 (N_6205,N_3939,N_3555);
nor U6206 (N_6206,N_3771,N_3022);
or U6207 (N_6207,N_4850,N_2999);
nor U6208 (N_6208,N_2934,N_3633);
nor U6209 (N_6209,N_4700,N_3349);
or U6210 (N_6210,N_2792,N_3379);
xnor U6211 (N_6211,N_4780,N_3493);
xor U6212 (N_6212,N_4550,N_4158);
or U6213 (N_6213,N_3436,N_3423);
nor U6214 (N_6214,N_3736,N_4672);
and U6215 (N_6215,N_4940,N_2710);
or U6216 (N_6216,N_4147,N_4490);
or U6217 (N_6217,N_3427,N_3149);
nand U6218 (N_6218,N_4633,N_4988);
nand U6219 (N_6219,N_2891,N_2967);
xor U6220 (N_6220,N_2799,N_4283);
nand U6221 (N_6221,N_4170,N_4492);
nand U6222 (N_6222,N_4642,N_2553);
and U6223 (N_6223,N_4702,N_4149);
xor U6224 (N_6224,N_4898,N_2708);
nand U6225 (N_6225,N_3319,N_4418);
nand U6226 (N_6226,N_2729,N_4670);
or U6227 (N_6227,N_3169,N_3055);
or U6228 (N_6228,N_3219,N_2898);
nor U6229 (N_6229,N_4235,N_3289);
nand U6230 (N_6230,N_4422,N_4316);
nand U6231 (N_6231,N_3230,N_2989);
nor U6232 (N_6232,N_4400,N_3274);
nand U6233 (N_6233,N_2827,N_2936);
or U6234 (N_6234,N_4082,N_3535);
nor U6235 (N_6235,N_2964,N_2733);
or U6236 (N_6236,N_4266,N_4775);
nand U6237 (N_6237,N_3953,N_3038);
or U6238 (N_6238,N_4987,N_3967);
nand U6239 (N_6239,N_4003,N_3293);
and U6240 (N_6240,N_4362,N_2703);
or U6241 (N_6241,N_3311,N_4753);
nor U6242 (N_6242,N_3302,N_3081);
nor U6243 (N_6243,N_4937,N_3338);
xnor U6244 (N_6244,N_4301,N_3375);
nor U6245 (N_6245,N_4020,N_4851);
xnor U6246 (N_6246,N_4443,N_2925);
xnor U6247 (N_6247,N_4711,N_4680);
xnor U6248 (N_6248,N_4883,N_4241);
xor U6249 (N_6249,N_3863,N_2937);
nor U6250 (N_6250,N_4572,N_3937);
xor U6251 (N_6251,N_3377,N_4092);
nor U6252 (N_6252,N_3397,N_4358);
nand U6253 (N_6253,N_2506,N_4164);
xnor U6254 (N_6254,N_4005,N_3546);
nand U6255 (N_6255,N_2808,N_3171);
nand U6256 (N_6256,N_3258,N_4278);
nor U6257 (N_6257,N_2542,N_3270);
or U6258 (N_6258,N_4264,N_3744);
xor U6259 (N_6259,N_3133,N_3040);
or U6260 (N_6260,N_4458,N_3565);
xor U6261 (N_6261,N_3997,N_3446);
and U6262 (N_6262,N_2843,N_4989);
or U6263 (N_6263,N_4595,N_3821);
nand U6264 (N_6264,N_3624,N_4761);
nor U6265 (N_6265,N_4062,N_3655);
nand U6266 (N_6266,N_4172,N_2609);
nor U6267 (N_6267,N_2665,N_3750);
nor U6268 (N_6268,N_4738,N_2709);
and U6269 (N_6269,N_3365,N_3022);
xnor U6270 (N_6270,N_3628,N_4337);
xnor U6271 (N_6271,N_4281,N_4576);
xor U6272 (N_6272,N_2600,N_4336);
nor U6273 (N_6273,N_2871,N_3804);
nand U6274 (N_6274,N_4667,N_2711);
or U6275 (N_6275,N_4585,N_3878);
or U6276 (N_6276,N_4565,N_3801);
nand U6277 (N_6277,N_2720,N_3600);
nand U6278 (N_6278,N_3642,N_4939);
nand U6279 (N_6279,N_2890,N_4870);
nor U6280 (N_6280,N_4689,N_4649);
or U6281 (N_6281,N_4672,N_2873);
nor U6282 (N_6282,N_3389,N_3194);
nand U6283 (N_6283,N_3473,N_3202);
or U6284 (N_6284,N_2891,N_4331);
or U6285 (N_6285,N_3823,N_4325);
and U6286 (N_6286,N_4150,N_4175);
nand U6287 (N_6287,N_3725,N_2627);
nand U6288 (N_6288,N_4984,N_3316);
or U6289 (N_6289,N_3986,N_3705);
or U6290 (N_6290,N_4862,N_2811);
and U6291 (N_6291,N_4614,N_3303);
nor U6292 (N_6292,N_3288,N_4746);
or U6293 (N_6293,N_3488,N_4203);
xnor U6294 (N_6294,N_2696,N_3261);
xor U6295 (N_6295,N_4206,N_4495);
or U6296 (N_6296,N_4558,N_3498);
or U6297 (N_6297,N_3275,N_3990);
xor U6298 (N_6298,N_3541,N_2796);
nand U6299 (N_6299,N_2930,N_3583);
nand U6300 (N_6300,N_4863,N_3696);
nor U6301 (N_6301,N_3887,N_4261);
xnor U6302 (N_6302,N_3134,N_2906);
nand U6303 (N_6303,N_4453,N_4567);
nor U6304 (N_6304,N_3393,N_2582);
nand U6305 (N_6305,N_4065,N_4900);
or U6306 (N_6306,N_3488,N_4583);
or U6307 (N_6307,N_2920,N_3940);
and U6308 (N_6308,N_2704,N_3472);
and U6309 (N_6309,N_4229,N_4984);
nand U6310 (N_6310,N_2736,N_3094);
nor U6311 (N_6311,N_3260,N_3577);
and U6312 (N_6312,N_3171,N_4352);
or U6313 (N_6313,N_3983,N_4299);
and U6314 (N_6314,N_3979,N_3428);
nand U6315 (N_6315,N_3865,N_3408);
nand U6316 (N_6316,N_3630,N_4250);
and U6317 (N_6317,N_3148,N_3397);
nand U6318 (N_6318,N_3549,N_3401);
xor U6319 (N_6319,N_3373,N_3201);
nand U6320 (N_6320,N_4478,N_4854);
nand U6321 (N_6321,N_4868,N_3682);
nor U6322 (N_6322,N_4439,N_2916);
and U6323 (N_6323,N_3274,N_4238);
and U6324 (N_6324,N_4279,N_3595);
nand U6325 (N_6325,N_4215,N_2809);
or U6326 (N_6326,N_4042,N_3443);
xor U6327 (N_6327,N_2543,N_4965);
or U6328 (N_6328,N_3286,N_3773);
nand U6329 (N_6329,N_3319,N_3164);
xnor U6330 (N_6330,N_4346,N_3683);
and U6331 (N_6331,N_2991,N_3525);
xor U6332 (N_6332,N_4817,N_4516);
xor U6333 (N_6333,N_4381,N_3086);
xor U6334 (N_6334,N_2910,N_3032);
nor U6335 (N_6335,N_2697,N_3650);
and U6336 (N_6336,N_4417,N_2794);
nand U6337 (N_6337,N_3812,N_2501);
or U6338 (N_6338,N_2819,N_2512);
and U6339 (N_6339,N_3154,N_4442);
or U6340 (N_6340,N_4543,N_3881);
and U6341 (N_6341,N_4618,N_3624);
or U6342 (N_6342,N_2903,N_4200);
nand U6343 (N_6343,N_4199,N_4144);
nor U6344 (N_6344,N_4683,N_3965);
nand U6345 (N_6345,N_3613,N_4970);
and U6346 (N_6346,N_3320,N_3493);
nor U6347 (N_6347,N_3556,N_2558);
or U6348 (N_6348,N_3501,N_4809);
nor U6349 (N_6349,N_2543,N_4036);
xnor U6350 (N_6350,N_2952,N_4187);
xnor U6351 (N_6351,N_4572,N_4805);
nand U6352 (N_6352,N_2784,N_3361);
nand U6353 (N_6353,N_4710,N_4656);
and U6354 (N_6354,N_3643,N_4626);
xnor U6355 (N_6355,N_4774,N_4569);
nand U6356 (N_6356,N_3918,N_3683);
nor U6357 (N_6357,N_4485,N_3323);
nor U6358 (N_6358,N_4287,N_4203);
nor U6359 (N_6359,N_3592,N_2659);
nand U6360 (N_6360,N_3461,N_4907);
xnor U6361 (N_6361,N_4971,N_4722);
or U6362 (N_6362,N_3460,N_3057);
or U6363 (N_6363,N_4929,N_3110);
nor U6364 (N_6364,N_2638,N_4641);
or U6365 (N_6365,N_2597,N_3897);
or U6366 (N_6366,N_3483,N_4813);
and U6367 (N_6367,N_4435,N_4464);
or U6368 (N_6368,N_4109,N_3579);
and U6369 (N_6369,N_4796,N_3252);
and U6370 (N_6370,N_4158,N_3579);
nand U6371 (N_6371,N_4775,N_4174);
and U6372 (N_6372,N_3250,N_4687);
nor U6373 (N_6373,N_3537,N_3834);
nor U6374 (N_6374,N_2501,N_4567);
and U6375 (N_6375,N_3554,N_4432);
nor U6376 (N_6376,N_4086,N_3422);
nand U6377 (N_6377,N_2682,N_4613);
xnor U6378 (N_6378,N_4234,N_2723);
xnor U6379 (N_6379,N_3128,N_3311);
or U6380 (N_6380,N_3550,N_4285);
xnor U6381 (N_6381,N_3439,N_4649);
nand U6382 (N_6382,N_3736,N_3660);
and U6383 (N_6383,N_3643,N_3654);
xnor U6384 (N_6384,N_4046,N_4773);
nor U6385 (N_6385,N_3942,N_3094);
nand U6386 (N_6386,N_4421,N_3205);
or U6387 (N_6387,N_3873,N_3772);
or U6388 (N_6388,N_4112,N_3172);
and U6389 (N_6389,N_3473,N_2949);
xnor U6390 (N_6390,N_4981,N_4635);
nand U6391 (N_6391,N_4998,N_4971);
nor U6392 (N_6392,N_2976,N_4827);
nor U6393 (N_6393,N_3674,N_2930);
and U6394 (N_6394,N_3137,N_4650);
or U6395 (N_6395,N_4963,N_3967);
nand U6396 (N_6396,N_4837,N_2593);
xnor U6397 (N_6397,N_3298,N_3405);
xor U6398 (N_6398,N_3659,N_3892);
xnor U6399 (N_6399,N_3849,N_3709);
and U6400 (N_6400,N_3414,N_3230);
nand U6401 (N_6401,N_3618,N_3343);
nor U6402 (N_6402,N_4391,N_2950);
and U6403 (N_6403,N_3124,N_2735);
nor U6404 (N_6404,N_2547,N_3417);
nor U6405 (N_6405,N_2658,N_3821);
nor U6406 (N_6406,N_4965,N_3422);
nand U6407 (N_6407,N_3742,N_4119);
nand U6408 (N_6408,N_3647,N_3509);
xnor U6409 (N_6409,N_4357,N_3468);
nand U6410 (N_6410,N_3256,N_4789);
xnor U6411 (N_6411,N_4694,N_3332);
or U6412 (N_6412,N_3087,N_4283);
nand U6413 (N_6413,N_3918,N_4002);
and U6414 (N_6414,N_4374,N_3197);
xnor U6415 (N_6415,N_4405,N_3782);
xnor U6416 (N_6416,N_3144,N_2500);
nand U6417 (N_6417,N_3912,N_2585);
or U6418 (N_6418,N_2743,N_3249);
and U6419 (N_6419,N_4493,N_3922);
nand U6420 (N_6420,N_2531,N_2895);
xnor U6421 (N_6421,N_3112,N_3731);
nand U6422 (N_6422,N_4265,N_3815);
and U6423 (N_6423,N_2926,N_4242);
and U6424 (N_6424,N_3532,N_4026);
nand U6425 (N_6425,N_2679,N_4147);
or U6426 (N_6426,N_3568,N_3667);
nor U6427 (N_6427,N_4119,N_3264);
nor U6428 (N_6428,N_3424,N_4635);
xor U6429 (N_6429,N_3902,N_2963);
nor U6430 (N_6430,N_4098,N_2568);
and U6431 (N_6431,N_3439,N_4591);
nand U6432 (N_6432,N_4792,N_2712);
nand U6433 (N_6433,N_2671,N_4829);
nor U6434 (N_6434,N_3838,N_2896);
nor U6435 (N_6435,N_4464,N_2861);
xnor U6436 (N_6436,N_3500,N_4266);
or U6437 (N_6437,N_2950,N_2780);
nor U6438 (N_6438,N_4641,N_4056);
xor U6439 (N_6439,N_3205,N_3757);
xor U6440 (N_6440,N_4788,N_4257);
nand U6441 (N_6441,N_4342,N_4376);
or U6442 (N_6442,N_4291,N_3560);
nand U6443 (N_6443,N_2631,N_4357);
xnor U6444 (N_6444,N_4200,N_3951);
and U6445 (N_6445,N_3369,N_3425);
or U6446 (N_6446,N_3208,N_3817);
and U6447 (N_6447,N_4398,N_3777);
nand U6448 (N_6448,N_2685,N_4287);
or U6449 (N_6449,N_3945,N_3972);
nor U6450 (N_6450,N_4935,N_2768);
nand U6451 (N_6451,N_4358,N_3526);
or U6452 (N_6452,N_4115,N_3526);
and U6453 (N_6453,N_4989,N_2505);
and U6454 (N_6454,N_2528,N_4099);
or U6455 (N_6455,N_2905,N_4904);
nor U6456 (N_6456,N_3049,N_3421);
or U6457 (N_6457,N_4085,N_4961);
xor U6458 (N_6458,N_4005,N_2823);
nand U6459 (N_6459,N_4861,N_2787);
nand U6460 (N_6460,N_3203,N_3435);
nor U6461 (N_6461,N_3856,N_3980);
nand U6462 (N_6462,N_4055,N_4122);
nand U6463 (N_6463,N_3176,N_4820);
nand U6464 (N_6464,N_4824,N_3806);
xnor U6465 (N_6465,N_4162,N_4196);
nor U6466 (N_6466,N_4849,N_4495);
nor U6467 (N_6467,N_3569,N_2774);
xnor U6468 (N_6468,N_3900,N_3904);
nor U6469 (N_6469,N_4381,N_3016);
or U6470 (N_6470,N_2855,N_4761);
xor U6471 (N_6471,N_3459,N_3265);
nor U6472 (N_6472,N_4602,N_4085);
nand U6473 (N_6473,N_2547,N_3110);
nand U6474 (N_6474,N_4258,N_3935);
xnor U6475 (N_6475,N_3827,N_3820);
and U6476 (N_6476,N_4768,N_4257);
and U6477 (N_6477,N_4455,N_4380);
nand U6478 (N_6478,N_3302,N_4831);
nor U6479 (N_6479,N_4963,N_4806);
xor U6480 (N_6480,N_2917,N_4039);
or U6481 (N_6481,N_3952,N_2816);
nand U6482 (N_6482,N_4707,N_3596);
or U6483 (N_6483,N_4505,N_4175);
xnor U6484 (N_6484,N_2862,N_4011);
nand U6485 (N_6485,N_4832,N_2898);
or U6486 (N_6486,N_3393,N_4865);
nand U6487 (N_6487,N_3680,N_2930);
or U6488 (N_6488,N_4600,N_2901);
or U6489 (N_6489,N_3117,N_3993);
nand U6490 (N_6490,N_2947,N_3134);
or U6491 (N_6491,N_3187,N_3065);
nor U6492 (N_6492,N_4333,N_4477);
and U6493 (N_6493,N_4745,N_3222);
nand U6494 (N_6494,N_3217,N_3246);
xnor U6495 (N_6495,N_4966,N_4052);
nor U6496 (N_6496,N_4520,N_4009);
or U6497 (N_6497,N_3829,N_3023);
nand U6498 (N_6498,N_2978,N_3347);
nor U6499 (N_6499,N_2815,N_4185);
xor U6500 (N_6500,N_2883,N_4285);
nand U6501 (N_6501,N_3779,N_4802);
xnor U6502 (N_6502,N_4573,N_4672);
or U6503 (N_6503,N_2623,N_2677);
nor U6504 (N_6504,N_2634,N_3062);
or U6505 (N_6505,N_2964,N_4917);
nor U6506 (N_6506,N_3752,N_4034);
or U6507 (N_6507,N_3987,N_3894);
nand U6508 (N_6508,N_3721,N_3712);
nand U6509 (N_6509,N_4370,N_3818);
nand U6510 (N_6510,N_3724,N_3255);
or U6511 (N_6511,N_3084,N_3635);
nor U6512 (N_6512,N_4719,N_4309);
or U6513 (N_6513,N_3499,N_3453);
or U6514 (N_6514,N_4046,N_3740);
and U6515 (N_6515,N_3476,N_2782);
and U6516 (N_6516,N_2859,N_3540);
or U6517 (N_6517,N_4797,N_3228);
and U6518 (N_6518,N_3430,N_2816);
nor U6519 (N_6519,N_3411,N_2827);
nand U6520 (N_6520,N_4149,N_3790);
or U6521 (N_6521,N_3571,N_3454);
xnor U6522 (N_6522,N_2604,N_2669);
nor U6523 (N_6523,N_4839,N_3340);
and U6524 (N_6524,N_4690,N_2663);
nand U6525 (N_6525,N_4994,N_4979);
xor U6526 (N_6526,N_4491,N_3599);
or U6527 (N_6527,N_4288,N_3034);
xnor U6528 (N_6528,N_4326,N_3399);
and U6529 (N_6529,N_3042,N_3838);
and U6530 (N_6530,N_2509,N_2790);
nand U6531 (N_6531,N_2692,N_4888);
nor U6532 (N_6532,N_3281,N_4242);
nand U6533 (N_6533,N_4133,N_2762);
xor U6534 (N_6534,N_4869,N_4571);
nand U6535 (N_6535,N_4970,N_3854);
and U6536 (N_6536,N_3761,N_3224);
and U6537 (N_6537,N_3968,N_3747);
nand U6538 (N_6538,N_3257,N_3255);
or U6539 (N_6539,N_4781,N_3578);
xnor U6540 (N_6540,N_4004,N_4043);
or U6541 (N_6541,N_4189,N_4566);
nand U6542 (N_6542,N_3383,N_3596);
xor U6543 (N_6543,N_4363,N_4021);
xor U6544 (N_6544,N_4656,N_3574);
nand U6545 (N_6545,N_4509,N_4394);
and U6546 (N_6546,N_4067,N_4045);
xnor U6547 (N_6547,N_4757,N_3815);
nand U6548 (N_6548,N_4599,N_3373);
or U6549 (N_6549,N_4689,N_2772);
and U6550 (N_6550,N_4888,N_4842);
nor U6551 (N_6551,N_3994,N_2650);
nand U6552 (N_6552,N_4212,N_4796);
nor U6553 (N_6553,N_2623,N_2529);
nor U6554 (N_6554,N_2982,N_3793);
nor U6555 (N_6555,N_4849,N_3870);
and U6556 (N_6556,N_4130,N_3133);
or U6557 (N_6557,N_2651,N_4028);
nor U6558 (N_6558,N_2678,N_2590);
nand U6559 (N_6559,N_2651,N_3112);
or U6560 (N_6560,N_3902,N_3865);
xor U6561 (N_6561,N_4639,N_4996);
nor U6562 (N_6562,N_3063,N_3991);
nand U6563 (N_6563,N_4309,N_2768);
or U6564 (N_6564,N_4241,N_4596);
xnor U6565 (N_6565,N_2588,N_4312);
or U6566 (N_6566,N_3990,N_3856);
xor U6567 (N_6567,N_3976,N_3140);
and U6568 (N_6568,N_3082,N_2537);
and U6569 (N_6569,N_3588,N_3513);
and U6570 (N_6570,N_4690,N_4277);
and U6571 (N_6571,N_4644,N_4733);
nand U6572 (N_6572,N_2965,N_3243);
xnor U6573 (N_6573,N_2689,N_3290);
or U6574 (N_6574,N_4899,N_4321);
nor U6575 (N_6575,N_4147,N_4952);
and U6576 (N_6576,N_3883,N_2835);
nand U6577 (N_6577,N_4277,N_2692);
nand U6578 (N_6578,N_4484,N_3127);
xnor U6579 (N_6579,N_3400,N_3520);
and U6580 (N_6580,N_2947,N_2835);
xnor U6581 (N_6581,N_3775,N_4180);
or U6582 (N_6582,N_2687,N_4387);
nand U6583 (N_6583,N_4622,N_4292);
or U6584 (N_6584,N_4851,N_3557);
and U6585 (N_6585,N_3876,N_3379);
xnor U6586 (N_6586,N_4549,N_3792);
or U6587 (N_6587,N_4322,N_3404);
nand U6588 (N_6588,N_4200,N_2941);
nor U6589 (N_6589,N_2934,N_4861);
and U6590 (N_6590,N_2695,N_4504);
nand U6591 (N_6591,N_3957,N_3556);
xnor U6592 (N_6592,N_2512,N_4858);
and U6593 (N_6593,N_4378,N_2737);
and U6594 (N_6594,N_4275,N_4466);
and U6595 (N_6595,N_3628,N_2899);
nand U6596 (N_6596,N_4318,N_4918);
or U6597 (N_6597,N_4027,N_4201);
nor U6598 (N_6598,N_2888,N_3592);
xnor U6599 (N_6599,N_4928,N_4725);
and U6600 (N_6600,N_2908,N_3565);
nor U6601 (N_6601,N_4202,N_3581);
and U6602 (N_6602,N_4654,N_4261);
xor U6603 (N_6603,N_4258,N_2970);
and U6604 (N_6604,N_4942,N_3709);
xor U6605 (N_6605,N_2634,N_4109);
xnor U6606 (N_6606,N_3118,N_3067);
xor U6607 (N_6607,N_2622,N_3295);
nand U6608 (N_6608,N_2710,N_4910);
or U6609 (N_6609,N_3999,N_3524);
and U6610 (N_6610,N_2629,N_4554);
nor U6611 (N_6611,N_3087,N_3700);
and U6612 (N_6612,N_3551,N_4441);
and U6613 (N_6613,N_2706,N_4806);
nand U6614 (N_6614,N_4600,N_2592);
xnor U6615 (N_6615,N_4814,N_3068);
nor U6616 (N_6616,N_4912,N_3579);
or U6617 (N_6617,N_3862,N_3078);
xnor U6618 (N_6618,N_4117,N_2739);
and U6619 (N_6619,N_2694,N_3306);
and U6620 (N_6620,N_3661,N_3902);
nand U6621 (N_6621,N_4762,N_4139);
nor U6622 (N_6622,N_3288,N_2913);
and U6623 (N_6623,N_2717,N_4691);
or U6624 (N_6624,N_2934,N_3496);
or U6625 (N_6625,N_4513,N_3550);
and U6626 (N_6626,N_3719,N_3224);
and U6627 (N_6627,N_3434,N_2629);
nor U6628 (N_6628,N_4210,N_3966);
or U6629 (N_6629,N_2576,N_2708);
nor U6630 (N_6630,N_3829,N_2869);
xor U6631 (N_6631,N_3325,N_4297);
and U6632 (N_6632,N_4794,N_3345);
nand U6633 (N_6633,N_4419,N_4953);
or U6634 (N_6634,N_3355,N_3221);
and U6635 (N_6635,N_4826,N_3514);
or U6636 (N_6636,N_4782,N_4840);
nor U6637 (N_6637,N_3084,N_2567);
or U6638 (N_6638,N_2956,N_4759);
xnor U6639 (N_6639,N_3856,N_4083);
and U6640 (N_6640,N_4250,N_3885);
or U6641 (N_6641,N_2635,N_3156);
or U6642 (N_6642,N_4441,N_2938);
and U6643 (N_6643,N_4970,N_3713);
or U6644 (N_6644,N_4157,N_3908);
nor U6645 (N_6645,N_3687,N_2888);
nor U6646 (N_6646,N_4347,N_4435);
nor U6647 (N_6647,N_4228,N_3783);
and U6648 (N_6648,N_4344,N_4839);
or U6649 (N_6649,N_3718,N_4564);
nor U6650 (N_6650,N_3311,N_2768);
xor U6651 (N_6651,N_4844,N_4789);
or U6652 (N_6652,N_2522,N_3268);
and U6653 (N_6653,N_4034,N_3510);
or U6654 (N_6654,N_3058,N_3495);
nand U6655 (N_6655,N_4004,N_3191);
nor U6656 (N_6656,N_2991,N_4429);
xnor U6657 (N_6657,N_4096,N_2747);
nor U6658 (N_6658,N_2568,N_2936);
nor U6659 (N_6659,N_4312,N_3673);
nor U6660 (N_6660,N_2776,N_3877);
nand U6661 (N_6661,N_3126,N_4593);
xor U6662 (N_6662,N_3328,N_3961);
and U6663 (N_6663,N_3913,N_2515);
and U6664 (N_6664,N_2999,N_4279);
or U6665 (N_6665,N_4295,N_4346);
xnor U6666 (N_6666,N_4620,N_2507);
nand U6667 (N_6667,N_3008,N_3266);
xor U6668 (N_6668,N_2993,N_3536);
and U6669 (N_6669,N_2528,N_2962);
or U6670 (N_6670,N_3887,N_4259);
or U6671 (N_6671,N_4981,N_2929);
xor U6672 (N_6672,N_4523,N_3601);
and U6673 (N_6673,N_4677,N_4002);
and U6674 (N_6674,N_3650,N_3169);
and U6675 (N_6675,N_4912,N_3943);
or U6676 (N_6676,N_4606,N_4451);
nor U6677 (N_6677,N_4825,N_2740);
nor U6678 (N_6678,N_3513,N_2677);
or U6679 (N_6679,N_2989,N_4158);
xor U6680 (N_6680,N_3981,N_3307);
nor U6681 (N_6681,N_3101,N_3861);
xnor U6682 (N_6682,N_4207,N_3488);
nand U6683 (N_6683,N_3824,N_4897);
nor U6684 (N_6684,N_3276,N_3207);
and U6685 (N_6685,N_2632,N_3026);
nor U6686 (N_6686,N_4449,N_2686);
or U6687 (N_6687,N_3991,N_3109);
nand U6688 (N_6688,N_4452,N_2551);
and U6689 (N_6689,N_3666,N_4827);
xor U6690 (N_6690,N_3732,N_4248);
xnor U6691 (N_6691,N_3461,N_4660);
nand U6692 (N_6692,N_4422,N_4113);
xnor U6693 (N_6693,N_2656,N_4532);
or U6694 (N_6694,N_4319,N_4260);
xor U6695 (N_6695,N_2820,N_4413);
nand U6696 (N_6696,N_2600,N_4279);
nor U6697 (N_6697,N_4985,N_4071);
and U6698 (N_6698,N_4031,N_4348);
nand U6699 (N_6699,N_4259,N_4119);
nor U6700 (N_6700,N_3574,N_3896);
and U6701 (N_6701,N_2599,N_4886);
nor U6702 (N_6702,N_4139,N_3692);
and U6703 (N_6703,N_2787,N_3982);
nor U6704 (N_6704,N_4345,N_4507);
nor U6705 (N_6705,N_4456,N_3863);
and U6706 (N_6706,N_4293,N_4798);
and U6707 (N_6707,N_4225,N_4304);
xnor U6708 (N_6708,N_3051,N_3973);
or U6709 (N_6709,N_4020,N_4126);
and U6710 (N_6710,N_2954,N_4715);
nand U6711 (N_6711,N_4902,N_4515);
nor U6712 (N_6712,N_3875,N_3807);
or U6713 (N_6713,N_2712,N_4606);
xor U6714 (N_6714,N_4414,N_3420);
and U6715 (N_6715,N_2687,N_2649);
nor U6716 (N_6716,N_2680,N_3187);
xnor U6717 (N_6717,N_3658,N_2754);
nor U6718 (N_6718,N_4790,N_2998);
and U6719 (N_6719,N_3989,N_3644);
and U6720 (N_6720,N_3319,N_2907);
nand U6721 (N_6721,N_3511,N_4790);
xnor U6722 (N_6722,N_3259,N_3632);
or U6723 (N_6723,N_2927,N_3712);
nor U6724 (N_6724,N_3873,N_3263);
or U6725 (N_6725,N_4775,N_2942);
or U6726 (N_6726,N_2684,N_4610);
xor U6727 (N_6727,N_3126,N_3655);
nand U6728 (N_6728,N_3901,N_4386);
nand U6729 (N_6729,N_4226,N_3074);
or U6730 (N_6730,N_3414,N_4718);
nor U6731 (N_6731,N_3760,N_4589);
nor U6732 (N_6732,N_2649,N_4349);
xnor U6733 (N_6733,N_4668,N_2679);
or U6734 (N_6734,N_3130,N_3083);
xor U6735 (N_6735,N_4961,N_2975);
nor U6736 (N_6736,N_4993,N_4743);
nor U6737 (N_6737,N_3976,N_2626);
and U6738 (N_6738,N_4836,N_4667);
nand U6739 (N_6739,N_2699,N_3366);
nand U6740 (N_6740,N_3795,N_3046);
nor U6741 (N_6741,N_3461,N_4628);
nand U6742 (N_6742,N_3700,N_4836);
and U6743 (N_6743,N_3484,N_2653);
xnor U6744 (N_6744,N_4622,N_4984);
nor U6745 (N_6745,N_3186,N_3993);
nor U6746 (N_6746,N_4704,N_3677);
nand U6747 (N_6747,N_3560,N_2591);
nand U6748 (N_6748,N_3896,N_3287);
xor U6749 (N_6749,N_3105,N_4056);
or U6750 (N_6750,N_3780,N_3091);
nand U6751 (N_6751,N_3304,N_3799);
and U6752 (N_6752,N_2915,N_3960);
xnor U6753 (N_6753,N_2729,N_2508);
nand U6754 (N_6754,N_3107,N_3698);
xor U6755 (N_6755,N_3397,N_3428);
and U6756 (N_6756,N_3634,N_3409);
or U6757 (N_6757,N_2563,N_3924);
nand U6758 (N_6758,N_4136,N_3844);
xnor U6759 (N_6759,N_4994,N_3093);
or U6760 (N_6760,N_4518,N_2586);
nor U6761 (N_6761,N_3029,N_4813);
xor U6762 (N_6762,N_2807,N_3379);
nor U6763 (N_6763,N_3336,N_3573);
and U6764 (N_6764,N_2500,N_2650);
nor U6765 (N_6765,N_4284,N_3217);
xor U6766 (N_6766,N_4230,N_4540);
xnor U6767 (N_6767,N_4479,N_2989);
nor U6768 (N_6768,N_2932,N_3543);
nand U6769 (N_6769,N_4259,N_3839);
or U6770 (N_6770,N_4074,N_3988);
nor U6771 (N_6771,N_3269,N_4514);
xnor U6772 (N_6772,N_4293,N_4358);
xnor U6773 (N_6773,N_4296,N_3647);
nand U6774 (N_6774,N_3246,N_2601);
or U6775 (N_6775,N_3109,N_2797);
or U6776 (N_6776,N_3007,N_3783);
nor U6777 (N_6777,N_4945,N_4143);
nand U6778 (N_6778,N_4149,N_4599);
and U6779 (N_6779,N_3912,N_3451);
nand U6780 (N_6780,N_2719,N_3958);
and U6781 (N_6781,N_3811,N_4954);
nor U6782 (N_6782,N_4830,N_2877);
xnor U6783 (N_6783,N_4661,N_3096);
xnor U6784 (N_6784,N_3759,N_4121);
or U6785 (N_6785,N_3676,N_3908);
xor U6786 (N_6786,N_3138,N_4991);
or U6787 (N_6787,N_4266,N_3548);
xor U6788 (N_6788,N_3893,N_4740);
and U6789 (N_6789,N_3391,N_4084);
and U6790 (N_6790,N_3295,N_3585);
or U6791 (N_6791,N_4280,N_3330);
nor U6792 (N_6792,N_2961,N_3344);
and U6793 (N_6793,N_3901,N_3277);
or U6794 (N_6794,N_2629,N_4880);
xnor U6795 (N_6795,N_3251,N_4429);
nor U6796 (N_6796,N_2880,N_2911);
and U6797 (N_6797,N_3779,N_4461);
and U6798 (N_6798,N_4171,N_2929);
or U6799 (N_6799,N_4488,N_4826);
xor U6800 (N_6800,N_2812,N_4740);
nand U6801 (N_6801,N_4050,N_4171);
nand U6802 (N_6802,N_4194,N_4494);
or U6803 (N_6803,N_4356,N_3368);
nand U6804 (N_6804,N_3575,N_3731);
or U6805 (N_6805,N_2857,N_4230);
xor U6806 (N_6806,N_3926,N_2966);
xnor U6807 (N_6807,N_2935,N_3343);
nor U6808 (N_6808,N_2729,N_4099);
and U6809 (N_6809,N_4497,N_4946);
nand U6810 (N_6810,N_3064,N_2930);
nor U6811 (N_6811,N_4389,N_4532);
nor U6812 (N_6812,N_3287,N_4180);
nand U6813 (N_6813,N_4304,N_4955);
or U6814 (N_6814,N_3264,N_2566);
xor U6815 (N_6815,N_4238,N_2672);
xnor U6816 (N_6816,N_4714,N_3933);
nand U6817 (N_6817,N_3095,N_2856);
and U6818 (N_6818,N_2873,N_4980);
or U6819 (N_6819,N_3637,N_2532);
xor U6820 (N_6820,N_2811,N_3275);
nor U6821 (N_6821,N_4400,N_4435);
nor U6822 (N_6822,N_4511,N_3413);
nor U6823 (N_6823,N_3788,N_4054);
nor U6824 (N_6824,N_4206,N_3349);
nand U6825 (N_6825,N_4289,N_2652);
nor U6826 (N_6826,N_3004,N_2903);
and U6827 (N_6827,N_2811,N_4071);
xor U6828 (N_6828,N_3140,N_3657);
and U6829 (N_6829,N_3938,N_3862);
nand U6830 (N_6830,N_3477,N_2999);
and U6831 (N_6831,N_4547,N_4455);
nand U6832 (N_6832,N_3056,N_4947);
nor U6833 (N_6833,N_4744,N_4833);
nor U6834 (N_6834,N_2866,N_3681);
nor U6835 (N_6835,N_3419,N_3100);
xor U6836 (N_6836,N_4143,N_4015);
nand U6837 (N_6837,N_4655,N_2586);
nor U6838 (N_6838,N_3931,N_3293);
and U6839 (N_6839,N_4161,N_4122);
nand U6840 (N_6840,N_2764,N_4841);
nor U6841 (N_6841,N_3377,N_2864);
and U6842 (N_6842,N_3322,N_3306);
xnor U6843 (N_6843,N_3096,N_3466);
or U6844 (N_6844,N_2542,N_2769);
nor U6845 (N_6845,N_3003,N_3347);
and U6846 (N_6846,N_4644,N_3003);
and U6847 (N_6847,N_4629,N_4568);
nor U6848 (N_6848,N_3889,N_4887);
or U6849 (N_6849,N_4523,N_2715);
and U6850 (N_6850,N_4856,N_3457);
nor U6851 (N_6851,N_3429,N_4467);
or U6852 (N_6852,N_4108,N_4595);
and U6853 (N_6853,N_2837,N_4376);
nand U6854 (N_6854,N_3946,N_3442);
nor U6855 (N_6855,N_3560,N_3730);
or U6856 (N_6856,N_3932,N_4536);
and U6857 (N_6857,N_2984,N_4358);
or U6858 (N_6858,N_2902,N_3307);
xor U6859 (N_6859,N_2678,N_3488);
xnor U6860 (N_6860,N_4434,N_3193);
xor U6861 (N_6861,N_3020,N_4185);
or U6862 (N_6862,N_3003,N_3414);
nor U6863 (N_6863,N_4745,N_4259);
and U6864 (N_6864,N_3594,N_4782);
nand U6865 (N_6865,N_3708,N_4999);
or U6866 (N_6866,N_4774,N_2616);
and U6867 (N_6867,N_3926,N_4813);
nand U6868 (N_6868,N_4254,N_4173);
nand U6869 (N_6869,N_2653,N_4528);
xnor U6870 (N_6870,N_3042,N_4069);
and U6871 (N_6871,N_3301,N_3540);
and U6872 (N_6872,N_4848,N_3726);
and U6873 (N_6873,N_4857,N_3619);
or U6874 (N_6874,N_2573,N_2742);
or U6875 (N_6875,N_3853,N_3962);
xnor U6876 (N_6876,N_2991,N_4755);
nor U6877 (N_6877,N_3940,N_3359);
xor U6878 (N_6878,N_3511,N_2537);
xor U6879 (N_6879,N_4917,N_3492);
xnor U6880 (N_6880,N_3018,N_3200);
or U6881 (N_6881,N_2564,N_2794);
or U6882 (N_6882,N_4299,N_3404);
xor U6883 (N_6883,N_4309,N_3983);
nor U6884 (N_6884,N_4729,N_2935);
xor U6885 (N_6885,N_3876,N_3522);
xnor U6886 (N_6886,N_2881,N_2581);
or U6887 (N_6887,N_2961,N_4591);
or U6888 (N_6888,N_3261,N_2939);
nor U6889 (N_6889,N_3003,N_3819);
or U6890 (N_6890,N_3102,N_3211);
nor U6891 (N_6891,N_2671,N_3126);
or U6892 (N_6892,N_4054,N_4714);
and U6893 (N_6893,N_3762,N_3436);
nor U6894 (N_6894,N_3733,N_4499);
or U6895 (N_6895,N_4161,N_3030);
nor U6896 (N_6896,N_3660,N_2530);
or U6897 (N_6897,N_4949,N_3716);
or U6898 (N_6898,N_3361,N_3507);
or U6899 (N_6899,N_2873,N_2519);
nor U6900 (N_6900,N_4407,N_4258);
and U6901 (N_6901,N_3902,N_4512);
nand U6902 (N_6902,N_3862,N_3327);
nor U6903 (N_6903,N_3790,N_3053);
or U6904 (N_6904,N_4406,N_3863);
and U6905 (N_6905,N_3669,N_2630);
xnor U6906 (N_6906,N_4804,N_3716);
or U6907 (N_6907,N_2838,N_3413);
xnor U6908 (N_6908,N_2683,N_4545);
xnor U6909 (N_6909,N_4827,N_2557);
and U6910 (N_6910,N_2942,N_4470);
xnor U6911 (N_6911,N_4118,N_4406);
nor U6912 (N_6912,N_4536,N_3384);
and U6913 (N_6913,N_2876,N_4029);
or U6914 (N_6914,N_4756,N_2892);
xnor U6915 (N_6915,N_4253,N_3544);
nor U6916 (N_6916,N_3079,N_4696);
nor U6917 (N_6917,N_4810,N_2626);
nor U6918 (N_6918,N_3359,N_4237);
nand U6919 (N_6919,N_4716,N_2830);
or U6920 (N_6920,N_3745,N_2832);
or U6921 (N_6921,N_2774,N_4234);
and U6922 (N_6922,N_2837,N_2527);
nand U6923 (N_6923,N_4808,N_4635);
xnor U6924 (N_6924,N_4310,N_4710);
xor U6925 (N_6925,N_2621,N_3545);
nand U6926 (N_6926,N_3982,N_4071);
nand U6927 (N_6927,N_3876,N_3820);
nand U6928 (N_6928,N_4342,N_2995);
or U6929 (N_6929,N_4134,N_4823);
xor U6930 (N_6930,N_4413,N_3465);
or U6931 (N_6931,N_4439,N_2612);
and U6932 (N_6932,N_4083,N_3212);
or U6933 (N_6933,N_3051,N_3255);
xnor U6934 (N_6934,N_3919,N_2570);
and U6935 (N_6935,N_3800,N_2599);
and U6936 (N_6936,N_4225,N_3909);
or U6937 (N_6937,N_3079,N_3586);
nand U6938 (N_6938,N_3933,N_3399);
nand U6939 (N_6939,N_3274,N_3228);
and U6940 (N_6940,N_2699,N_3803);
xor U6941 (N_6941,N_4727,N_4703);
and U6942 (N_6942,N_3806,N_4902);
and U6943 (N_6943,N_3798,N_3059);
or U6944 (N_6944,N_4323,N_4858);
nand U6945 (N_6945,N_3582,N_4182);
and U6946 (N_6946,N_2863,N_3549);
or U6947 (N_6947,N_3455,N_2725);
xor U6948 (N_6948,N_3890,N_2720);
and U6949 (N_6949,N_3008,N_3271);
and U6950 (N_6950,N_4057,N_4300);
xnor U6951 (N_6951,N_4038,N_4098);
xnor U6952 (N_6952,N_4327,N_4829);
nand U6953 (N_6953,N_3820,N_4367);
xor U6954 (N_6954,N_4472,N_4597);
nand U6955 (N_6955,N_4480,N_3845);
nor U6956 (N_6956,N_3938,N_3625);
nor U6957 (N_6957,N_4249,N_4068);
xnor U6958 (N_6958,N_3219,N_4500);
xnor U6959 (N_6959,N_2507,N_4002);
or U6960 (N_6960,N_3391,N_4599);
nand U6961 (N_6961,N_4777,N_3661);
nor U6962 (N_6962,N_4714,N_4951);
nor U6963 (N_6963,N_4590,N_2787);
xor U6964 (N_6964,N_3473,N_4154);
nand U6965 (N_6965,N_4148,N_3312);
or U6966 (N_6966,N_3759,N_4047);
or U6967 (N_6967,N_2635,N_3510);
nor U6968 (N_6968,N_4917,N_3350);
or U6969 (N_6969,N_3927,N_4505);
or U6970 (N_6970,N_3792,N_2800);
and U6971 (N_6971,N_2608,N_2901);
nand U6972 (N_6972,N_3959,N_3557);
xor U6973 (N_6973,N_2940,N_4430);
and U6974 (N_6974,N_3178,N_2654);
nand U6975 (N_6975,N_4801,N_4401);
nand U6976 (N_6976,N_4418,N_4642);
nor U6977 (N_6977,N_4816,N_4480);
or U6978 (N_6978,N_2942,N_3448);
nand U6979 (N_6979,N_3909,N_2628);
xor U6980 (N_6980,N_3277,N_3587);
or U6981 (N_6981,N_3403,N_2574);
or U6982 (N_6982,N_4704,N_2699);
nor U6983 (N_6983,N_4363,N_2911);
or U6984 (N_6984,N_4296,N_4493);
nor U6985 (N_6985,N_4278,N_4187);
nor U6986 (N_6986,N_3355,N_3790);
and U6987 (N_6987,N_3994,N_3373);
nor U6988 (N_6988,N_4691,N_3133);
xnor U6989 (N_6989,N_4664,N_4260);
xor U6990 (N_6990,N_4575,N_4280);
xor U6991 (N_6991,N_3804,N_3246);
xor U6992 (N_6992,N_3750,N_4799);
nor U6993 (N_6993,N_3546,N_3009);
xor U6994 (N_6994,N_3527,N_4122);
and U6995 (N_6995,N_2577,N_3903);
xor U6996 (N_6996,N_4645,N_3348);
or U6997 (N_6997,N_3415,N_4315);
nand U6998 (N_6998,N_4846,N_4472);
or U6999 (N_6999,N_3769,N_3103);
nand U7000 (N_7000,N_3482,N_4537);
nand U7001 (N_7001,N_3254,N_4248);
and U7002 (N_7002,N_4045,N_3230);
xnor U7003 (N_7003,N_3773,N_3308);
nor U7004 (N_7004,N_3544,N_4554);
nand U7005 (N_7005,N_2646,N_4941);
nor U7006 (N_7006,N_4631,N_4543);
or U7007 (N_7007,N_4751,N_3741);
nand U7008 (N_7008,N_3474,N_4701);
xnor U7009 (N_7009,N_2985,N_4619);
nor U7010 (N_7010,N_4410,N_3259);
and U7011 (N_7011,N_3077,N_3002);
or U7012 (N_7012,N_3474,N_3649);
xor U7013 (N_7013,N_3817,N_4911);
and U7014 (N_7014,N_3335,N_4886);
nor U7015 (N_7015,N_3287,N_4259);
nand U7016 (N_7016,N_3824,N_4820);
nor U7017 (N_7017,N_4000,N_2729);
and U7018 (N_7018,N_4278,N_4527);
xnor U7019 (N_7019,N_3255,N_4026);
and U7020 (N_7020,N_3568,N_3032);
xor U7021 (N_7021,N_4524,N_3931);
nor U7022 (N_7022,N_2982,N_3596);
or U7023 (N_7023,N_2658,N_3148);
xnor U7024 (N_7024,N_3112,N_2755);
or U7025 (N_7025,N_4793,N_3355);
and U7026 (N_7026,N_4788,N_4787);
nor U7027 (N_7027,N_4612,N_4824);
or U7028 (N_7028,N_4676,N_4958);
and U7029 (N_7029,N_4037,N_4186);
xnor U7030 (N_7030,N_3949,N_4635);
and U7031 (N_7031,N_3525,N_3570);
nor U7032 (N_7032,N_2736,N_3791);
nand U7033 (N_7033,N_3513,N_3468);
xor U7034 (N_7034,N_4277,N_4312);
or U7035 (N_7035,N_4096,N_3362);
or U7036 (N_7036,N_4316,N_4785);
and U7037 (N_7037,N_3402,N_4324);
or U7038 (N_7038,N_2517,N_2594);
or U7039 (N_7039,N_4742,N_3780);
and U7040 (N_7040,N_3972,N_3301);
nor U7041 (N_7041,N_3198,N_2582);
nand U7042 (N_7042,N_4287,N_3921);
xor U7043 (N_7043,N_4487,N_2953);
xnor U7044 (N_7044,N_4462,N_3157);
nor U7045 (N_7045,N_4583,N_2602);
xor U7046 (N_7046,N_3314,N_3007);
and U7047 (N_7047,N_4539,N_4652);
xnor U7048 (N_7048,N_2779,N_3739);
or U7049 (N_7049,N_3496,N_2794);
nand U7050 (N_7050,N_4868,N_4335);
nor U7051 (N_7051,N_2598,N_3309);
and U7052 (N_7052,N_4505,N_2735);
nor U7053 (N_7053,N_3847,N_4688);
xor U7054 (N_7054,N_3524,N_4304);
and U7055 (N_7055,N_2988,N_3384);
nand U7056 (N_7056,N_2637,N_4922);
or U7057 (N_7057,N_4268,N_2772);
nor U7058 (N_7058,N_3449,N_2819);
and U7059 (N_7059,N_4296,N_3765);
or U7060 (N_7060,N_2550,N_3236);
nor U7061 (N_7061,N_4113,N_2750);
or U7062 (N_7062,N_4771,N_4408);
or U7063 (N_7063,N_2688,N_3282);
or U7064 (N_7064,N_3497,N_3368);
and U7065 (N_7065,N_4166,N_3032);
xnor U7066 (N_7066,N_2529,N_3991);
nor U7067 (N_7067,N_2883,N_2543);
and U7068 (N_7068,N_2936,N_2866);
or U7069 (N_7069,N_2710,N_3911);
nor U7070 (N_7070,N_4541,N_3040);
xnor U7071 (N_7071,N_4383,N_3811);
nor U7072 (N_7072,N_4526,N_4985);
xor U7073 (N_7073,N_3037,N_3048);
nor U7074 (N_7074,N_3496,N_2906);
or U7075 (N_7075,N_4917,N_3528);
xor U7076 (N_7076,N_4718,N_4828);
and U7077 (N_7077,N_3691,N_3659);
nor U7078 (N_7078,N_2924,N_3058);
and U7079 (N_7079,N_2972,N_3037);
and U7080 (N_7080,N_4035,N_3820);
and U7081 (N_7081,N_4604,N_3637);
or U7082 (N_7082,N_3777,N_4922);
nor U7083 (N_7083,N_2556,N_4070);
and U7084 (N_7084,N_2859,N_4647);
nor U7085 (N_7085,N_3516,N_3139);
nor U7086 (N_7086,N_2765,N_3171);
and U7087 (N_7087,N_4316,N_4623);
and U7088 (N_7088,N_3933,N_4527);
and U7089 (N_7089,N_4437,N_4038);
and U7090 (N_7090,N_3455,N_4702);
nor U7091 (N_7091,N_3829,N_4239);
xor U7092 (N_7092,N_3576,N_3967);
nand U7093 (N_7093,N_4655,N_3798);
xnor U7094 (N_7094,N_4084,N_4384);
nand U7095 (N_7095,N_3378,N_2624);
or U7096 (N_7096,N_3972,N_4614);
and U7097 (N_7097,N_2935,N_3625);
and U7098 (N_7098,N_3349,N_4391);
xnor U7099 (N_7099,N_3391,N_4988);
or U7100 (N_7100,N_4566,N_3975);
xnor U7101 (N_7101,N_4108,N_3820);
nor U7102 (N_7102,N_3309,N_3319);
nor U7103 (N_7103,N_2538,N_3685);
nor U7104 (N_7104,N_2807,N_4487);
xor U7105 (N_7105,N_4734,N_3778);
and U7106 (N_7106,N_2645,N_4154);
or U7107 (N_7107,N_3695,N_4946);
xnor U7108 (N_7108,N_3316,N_4915);
nor U7109 (N_7109,N_4835,N_3202);
and U7110 (N_7110,N_4354,N_2575);
xor U7111 (N_7111,N_4892,N_4794);
xnor U7112 (N_7112,N_4806,N_3664);
and U7113 (N_7113,N_2601,N_4991);
xor U7114 (N_7114,N_3451,N_3446);
nor U7115 (N_7115,N_2860,N_2732);
or U7116 (N_7116,N_3272,N_4432);
and U7117 (N_7117,N_3801,N_4927);
and U7118 (N_7118,N_3385,N_3740);
or U7119 (N_7119,N_4219,N_4554);
xor U7120 (N_7120,N_4616,N_4008);
and U7121 (N_7121,N_3417,N_3723);
nor U7122 (N_7122,N_2656,N_4681);
xnor U7123 (N_7123,N_3476,N_3604);
and U7124 (N_7124,N_2589,N_3968);
nand U7125 (N_7125,N_2662,N_4904);
nor U7126 (N_7126,N_2985,N_4516);
nand U7127 (N_7127,N_3371,N_2855);
xnor U7128 (N_7128,N_4612,N_4730);
nand U7129 (N_7129,N_2842,N_3530);
and U7130 (N_7130,N_4397,N_3544);
and U7131 (N_7131,N_4928,N_3280);
or U7132 (N_7132,N_2665,N_4085);
or U7133 (N_7133,N_3104,N_4313);
nor U7134 (N_7134,N_4317,N_4814);
nor U7135 (N_7135,N_2537,N_3844);
nand U7136 (N_7136,N_4462,N_2501);
or U7137 (N_7137,N_4306,N_2593);
and U7138 (N_7138,N_3523,N_4689);
or U7139 (N_7139,N_4006,N_4608);
and U7140 (N_7140,N_3230,N_4396);
and U7141 (N_7141,N_3077,N_4496);
and U7142 (N_7142,N_4666,N_3218);
nor U7143 (N_7143,N_2962,N_2937);
nand U7144 (N_7144,N_4630,N_3901);
or U7145 (N_7145,N_3398,N_4796);
or U7146 (N_7146,N_2687,N_4368);
or U7147 (N_7147,N_4884,N_3895);
xor U7148 (N_7148,N_4464,N_2652);
and U7149 (N_7149,N_2853,N_3297);
nor U7150 (N_7150,N_3093,N_4548);
nor U7151 (N_7151,N_3508,N_3110);
or U7152 (N_7152,N_4755,N_3860);
and U7153 (N_7153,N_3660,N_3841);
xor U7154 (N_7154,N_4960,N_3200);
nand U7155 (N_7155,N_4450,N_3221);
or U7156 (N_7156,N_3373,N_4611);
nand U7157 (N_7157,N_3834,N_3806);
and U7158 (N_7158,N_3444,N_3495);
or U7159 (N_7159,N_4095,N_3419);
or U7160 (N_7160,N_4007,N_2659);
xnor U7161 (N_7161,N_4161,N_2701);
xor U7162 (N_7162,N_2832,N_2527);
nand U7163 (N_7163,N_4781,N_3583);
nor U7164 (N_7164,N_3367,N_3450);
xnor U7165 (N_7165,N_4149,N_2982);
xnor U7166 (N_7166,N_4764,N_2702);
xnor U7167 (N_7167,N_3211,N_3996);
xor U7168 (N_7168,N_4800,N_2602);
nand U7169 (N_7169,N_4955,N_3493);
xnor U7170 (N_7170,N_2788,N_3545);
and U7171 (N_7171,N_3288,N_4799);
xor U7172 (N_7172,N_3517,N_2547);
or U7173 (N_7173,N_4174,N_3382);
or U7174 (N_7174,N_4204,N_4187);
and U7175 (N_7175,N_4307,N_4146);
nor U7176 (N_7176,N_4440,N_3270);
and U7177 (N_7177,N_2530,N_3264);
or U7178 (N_7178,N_4689,N_3547);
nand U7179 (N_7179,N_4177,N_3721);
xor U7180 (N_7180,N_3301,N_2775);
nor U7181 (N_7181,N_4206,N_2745);
nand U7182 (N_7182,N_2736,N_3552);
nand U7183 (N_7183,N_3783,N_3057);
nand U7184 (N_7184,N_3627,N_2697);
xnor U7185 (N_7185,N_3562,N_3216);
and U7186 (N_7186,N_4805,N_2854);
or U7187 (N_7187,N_4543,N_4758);
nand U7188 (N_7188,N_4032,N_3079);
xor U7189 (N_7189,N_3149,N_3931);
or U7190 (N_7190,N_2754,N_3238);
nand U7191 (N_7191,N_4643,N_2816);
and U7192 (N_7192,N_3481,N_4410);
nand U7193 (N_7193,N_4309,N_4161);
xor U7194 (N_7194,N_3067,N_3923);
and U7195 (N_7195,N_4739,N_3299);
and U7196 (N_7196,N_4844,N_4765);
xor U7197 (N_7197,N_4314,N_3777);
and U7198 (N_7198,N_2577,N_3160);
and U7199 (N_7199,N_4325,N_4474);
nand U7200 (N_7200,N_4643,N_3883);
xor U7201 (N_7201,N_3404,N_2859);
nand U7202 (N_7202,N_4520,N_4541);
or U7203 (N_7203,N_3126,N_3548);
and U7204 (N_7204,N_4736,N_3759);
xor U7205 (N_7205,N_4619,N_4603);
or U7206 (N_7206,N_4848,N_4618);
xor U7207 (N_7207,N_3004,N_3289);
xor U7208 (N_7208,N_4078,N_3659);
nand U7209 (N_7209,N_2933,N_3900);
xnor U7210 (N_7210,N_2606,N_3672);
or U7211 (N_7211,N_4069,N_4603);
xnor U7212 (N_7212,N_3137,N_4019);
and U7213 (N_7213,N_4028,N_4659);
nor U7214 (N_7214,N_2712,N_3636);
or U7215 (N_7215,N_3896,N_3991);
or U7216 (N_7216,N_4511,N_3113);
nand U7217 (N_7217,N_4964,N_4022);
nand U7218 (N_7218,N_2983,N_2784);
or U7219 (N_7219,N_4439,N_4619);
xor U7220 (N_7220,N_4935,N_3752);
nor U7221 (N_7221,N_4829,N_3132);
or U7222 (N_7222,N_3663,N_3955);
nand U7223 (N_7223,N_2583,N_4281);
nor U7224 (N_7224,N_4928,N_2989);
nand U7225 (N_7225,N_4786,N_3949);
nor U7226 (N_7226,N_3496,N_2992);
nand U7227 (N_7227,N_2819,N_3782);
and U7228 (N_7228,N_3131,N_4443);
and U7229 (N_7229,N_4903,N_3791);
nor U7230 (N_7230,N_3898,N_3785);
nand U7231 (N_7231,N_2536,N_3734);
xor U7232 (N_7232,N_4191,N_3349);
nand U7233 (N_7233,N_3800,N_3606);
nand U7234 (N_7234,N_2957,N_4701);
nand U7235 (N_7235,N_4337,N_4849);
nor U7236 (N_7236,N_4991,N_3731);
or U7237 (N_7237,N_3463,N_2914);
nor U7238 (N_7238,N_4033,N_3925);
xor U7239 (N_7239,N_3481,N_3941);
nor U7240 (N_7240,N_2741,N_3321);
nand U7241 (N_7241,N_2691,N_4275);
xor U7242 (N_7242,N_3199,N_4166);
xor U7243 (N_7243,N_2760,N_3500);
or U7244 (N_7244,N_4545,N_3504);
and U7245 (N_7245,N_4883,N_3825);
or U7246 (N_7246,N_3688,N_4021);
and U7247 (N_7247,N_3491,N_4607);
nand U7248 (N_7248,N_3166,N_4723);
or U7249 (N_7249,N_2766,N_2935);
xnor U7250 (N_7250,N_3853,N_2970);
nor U7251 (N_7251,N_4002,N_3465);
nand U7252 (N_7252,N_4476,N_4945);
nor U7253 (N_7253,N_2797,N_3229);
xor U7254 (N_7254,N_4072,N_4035);
nor U7255 (N_7255,N_4924,N_3800);
nand U7256 (N_7256,N_4253,N_4705);
nor U7257 (N_7257,N_3995,N_4750);
nand U7258 (N_7258,N_2702,N_3002);
xnor U7259 (N_7259,N_4892,N_2966);
xor U7260 (N_7260,N_2582,N_3354);
or U7261 (N_7261,N_3511,N_4909);
nand U7262 (N_7262,N_4981,N_4831);
nor U7263 (N_7263,N_4230,N_4262);
and U7264 (N_7264,N_4223,N_2587);
xor U7265 (N_7265,N_2937,N_3058);
or U7266 (N_7266,N_4846,N_2915);
or U7267 (N_7267,N_4758,N_2688);
and U7268 (N_7268,N_3046,N_3703);
or U7269 (N_7269,N_3332,N_4614);
and U7270 (N_7270,N_4275,N_3525);
nand U7271 (N_7271,N_3109,N_4138);
xnor U7272 (N_7272,N_2557,N_3491);
nor U7273 (N_7273,N_4973,N_4411);
xor U7274 (N_7274,N_4912,N_3042);
nor U7275 (N_7275,N_2884,N_2576);
nand U7276 (N_7276,N_4647,N_2845);
and U7277 (N_7277,N_3221,N_3057);
xnor U7278 (N_7278,N_4384,N_4398);
nand U7279 (N_7279,N_3778,N_3409);
and U7280 (N_7280,N_3097,N_3104);
or U7281 (N_7281,N_3873,N_3910);
or U7282 (N_7282,N_3636,N_3348);
and U7283 (N_7283,N_4521,N_4088);
nand U7284 (N_7284,N_3569,N_2799);
nand U7285 (N_7285,N_3840,N_3153);
nor U7286 (N_7286,N_4947,N_4389);
or U7287 (N_7287,N_3538,N_3824);
nand U7288 (N_7288,N_4734,N_2586);
or U7289 (N_7289,N_4506,N_3334);
and U7290 (N_7290,N_4797,N_4105);
nand U7291 (N_7291,N_3457,N_2732);
or U7292 (N_7292,N_2523,N_3263);
and U7293 (N_7293,N_2915,N_3528);
nand U7294 (N_7294,N_4376,N_3098);
nor U7295 (N_7295,N_4898,N_4374);
xor U7296 (N_7296,N_3385,N_3707);
nand U7297 (N_7297,N_3792,N_2768);
nor U7298 (N_7298,N_3795,N_2899);
and U7299 (N_7299,N_4413,N_3075);
or U7300 (N_7300,N_3481,N_2530);
nor U7301 (N_7301,N_2939,N_3998);
xnor U7302 (N_7302,N_4369,N_2995);
xor U7303 (N_7303,N_2699,N_4075);
xor U7304 (N_7304,N_3327,N_2825);
nor U7305 (N_7305,N_3789,N_2766);
and U7306 (N_7306,N_4107,N_2534);
nand U7307 (N_7307,N_2893,N_2936);
nor U7308 (N_7308,N_2554,N_2790);
xor U7309 (N_7309,N_3342,N_3226);
and U7310 (N_7310,N_3737,N_3933);
or U7311 (N_7311,N_4646,N_4700);
or U7312 (N_7312,N_4945,N_4898);
nor U7313 (N_7313,N_3823,N_3686);
xnor U7314 (N_7314,N_2585,N_4685);
nand U7315 (N_7315,N_4607,N_3334);
nor U7316 (N_7316,N_3141,N_3885);
nand U7317 (N_7317,N_4117,N_3906);
nor U7318 (N_7318,N_4790,N_3493);
and U7319 (N_7319,N_3343,N_3454);
or U7320 (N_7320,N_4201,N_2704);
and U7321 (N_7321,N_4081,N_4477);
and U7322 (N_7322,N_4197,N_4982);
xor U7323 (N_7323,N_2637,N_4414);
or U7324 (N_7324,N_4588,N_3127);
or U7325 (N_7325,N_3423,N_4733);
or U7326 (N_7326,N_4583,N_3631);
nand U7327 (N_7327,N_4816,N_3123);
and U7328 (N_7328,N_4443,N_4877);
xnor U7329 (N_7329,N_3162,N_4473);
and U7330 (N_7330,N_4558,N_3884);
nand U7331 (N_7331,N_2951,N_4450);
or U7332 (N_7332,N_3521,N_3415);
nand U7333 (N_7333,N_4169,N_4102);
and U7334 (N_7334,N_3949,N_4625);
nor U7335 (N_7335,N_4260,N_2793);
nand U7336 (N_7336,N_3397,N_3208);
nor U7337 (N_7337,N_4474,N_4341);
or U7338 (N_7338,N_4669,N_2688);
xor U7339 (N_7339,N_3627,N_2817);
and U7340 (N_7340,N_3378,N_3333);
nand U7341 (N_7341,N_4870,N_3726);
xnor U7342 (N_7342,N_4310,N_2781);
nor U7343 (N_7343,N_3774,N_3801);
nand U7344 (N_7344,N_4199,N_4167);
or U7345 (N_7345,N_4770,N_4478);
nand U7346 (N_7346,N_4407,N_4411);
xnor U7347 (N_7347,N_3238,N_3395);
and U7348 (N_7348,N_3536,N_3575);
xnor U7349 (N_7349,N_4002,N_4431);
nand U7350 (N_7350,N_2541,N_4330);
xnor U7351 (N_7351,N_4889,N_4347);
xor U7352 (N_7352,N_3496,N_3827);
nor U7353 (N_7353,N_4241,N_4864);
or U7354 (N_7354,N_3877,N_3302);
xnor U7355 (N_7355,N_4415,N_3829);
and U7356 (N_7356,N_4020,N_3055);
and U7357 (N_7357,N_4367,N_4476);
nor U7358 (N_7358,N_3851,N_3312);
xnor U7359 (N_7359,N_4206,N_2601);
and U7360 (N_7360,N_2961,N_4028);
or U7361 (N_7361,N_4690,N_3520);
or U7362 (N_7362,N_3531,N_4400);
nor U7363 (N_7363,N_4396,N_4005);
nor U7364 (N_7364,N_2722,N_3904);
and U7365 (N_7365,N_3645,N_3659);
or U7366 (N_7366,N_4778,N_2950);
nand U7367 (N_7367,N_2989,N_4023);
and U7368 (N_7368,N_4684,N_4727);
and U7369 (N_7369,N_3346,N_3600);
nor U7370 (N_7370,N_3721,N_2803);
nand U7371 (N_7371,N_4833,N_2658);
nor U7372 (N_7372,N_4620,N_2718);
nand U7373 (N_7373,N_3294,N_3005);
and U7374 (N_7374,N_3600,N_3512);
nor U7375 (N_7375,N_2581,N_4480);
nand U7376 (N_7376,N_2671,N_3680);
or U7377 (N_7377,N_2877,N_3696);
nor U7378 (N_7378,N_2513,N_4437);
and U7379 (N_7379,N_3671,N_4962);
nor U7380 (N_7380,N_3872,N_2815);
nand U7381 (N_7381,N_4903,N_3572);
or U7382 (N_7382,N_2765,N_4413);
or U7383 (N_7383,N_3283,N_4610);
nand U7384 (N_7384,N_4010,N_4632);
xor U7385 (N_7385,N_3949,N_3432);
or U7386 (N_7386,N_4881,N_3116);
xor U7387 (N_7387,N_3211,N_3399);
xnor U7388 (N_7388,N_4549,N_4177);
and U7389 (N_7389,N_4460,N_3590);
nand U7390 (N_7390,N_4624,N_4235);
and U7391 (N_7391,N_3358,N_3089);
or U7392 (N_7392,N_4716,N_3931);
or U7393 (N_7393,N_2856,N_3432);
nand U7394 (N_7394,N_2724,N_2949);
nand U7395 (N_7395,N_3273,N_2751);
and U7396 (N_7396,N_3181,N_4759);
and U7397 (N_7397,N_3204,N_4029);
nand U7398 (N_7398,N_4920,N_4702);
or U7399 (N_7399,N_4652,N_3251);
nor U7400 (N_7400,N_2660,N_4044);
xor U7401 (N_7401,N_3726,N_4203);
and U7402 (N_7402,N_3748,N_4892);
or U7403 (N_7403,N_3800,N_2806);
nand U7404 (N_7404,N_3604,N_4061);
xnor U7405 (N_7405,N_2877,N_3849);
nor U7406 (N_7406,N_3418,N_4890);
xor U7407 (N_7407,N_3767,N_3445);
nor U7408 (N_7408,N_2800,N_4972);
or U7409 (N_7409,N_3274,N_4661);
xnor U7410 (N_7410,N_3193,N_3366);
nand U7411 (N_7411,N_3123,N_3514);
nand U7412 (N_7412,N_3824,N_3714);
nor U7413 (N_7413,N_3799,N_3149);
xor U7414 (N_7414,N_2642,N_4269);
or U7415 (N_7415,N_3691,N_3376);
xnor U7416 (N_7416,N_2709,N_3234);
and U7417 (N_7417,N_4902,N_4853);
nor U7418 (N_7418,N_4525,N_3990);
xor U7419 (N_7419,N_3726,N_4668);
xnor U7420 (N_7420,N_4116,N_4854);
nor U7421 (N_7421,N_2837,N_4890);
nand U7422 (N_7422,N_2951,N_4344);
nor U7423 (N_7423,N_3508,N_3179);
xor U7424 (N_7424,N_2514,N_4108);
nor U7425 (N_7425,N_4606,N_4616);
and U7426 (N_7426,N_4368,N_2900);
nand U7427 (N_7427,N_3191,N_4833);
and U7428 (N_7428,N_4140,N_4179);
nor U7429 (N_7429,N_3871,N_3408);
xor U7430 (N_7430,N_2819,N_4435);
nor U7431 (N_7431,N_2869,N_4123);
nor U7432 (N_7432,N_3314,N_4874);
nor U7433 (N_7433,N_4047,N_4185);
and U7434 (N_7434,N_4226,N_4702);
nand U7435 (N_7435,N_4693,N_4359);
nor U7436 (N_7436,N_4850,N_3283);
or U7437 (N_7437,N_2833,N_3928);
xnor U7438 (N_7438,N_4316,N_4646);
or U7439 (N_7439,N_4787,N_3849);
xor U7440 (N_7440,N_4813,N_4215);
and U7441 (N_7441,N_4951,N_4087);
or U7442 (N_7442,N_2625,N_3082);
or U7443 (N_7443,N_3380,N_3695);
nand U7444 (N_7444,N_3536,N_3116);
or U7445 (N_7445,N_3535,N_2940);
xor U7446 (N_7446,N_4873,N_4542);
nor U7447 (N_7447,N_2851,N_3577);
nor U7448 (N_7448,N_2949,N_3519);
nand U7449 (N_7449,N_3696,N_4740);
and U7450 (N_7450,N_2766,N_2890);
or U7451 (N_7451,N_4004,N_3454);
xor U7452 (N_7452,N_4926,N_3236);
or U7453 (N_7453,N_4622,N_4845);
nand U7454 (N_7454,N_4601,N_3403);
or U7455 (N_7455,N_3949,N_4765);
or U7456 (N_7456,N_2984,N_4243);
nand U7457 (N_7457,N_4244,N_4727);
and U7458 (N_7458,N_3517,N_3914);
nor U7459 (N_7459,N_3531,N_4026);
and U7460 (N_7460,N_4149,N_3928);
nor U7461 (N_7461,N_3026,N_4248);
nor U7462 (N_7462,N_3797,N_3448);
nor U7463 (N_7463,N_3574,N_3788);
or U7464 (N_7464,N_3663,N_4344);
nand U7465 (N_7465,N_3317,N_3340);
nand U7466 (N_7466,N_2770,N_3309);
xor U7467 (N_7467,N_4806,N_4161);
or U7468 (N_7468,N_2701,N_2843);
xnor U7469 (N_7469,N_2993,N_3497);
and U7470 (N_7470,N_2723,N_2977);
xnor U7471 (N_7471,N_4898,N_2740);
or U7472 (N_7472,N_3013,N_3587);
or U7473 (N_7473,N_3540,N_4101);
or U7474 (N_7474,N_4116,N_2797);
nand U7475 (N_7475,N_4073,N_4797);
nand U7476 (N_7476,N_4822,N_3066);
or U7477 (N_7477,N_3653,N_4042);
xor U7478 (N_7478,N_3758,N_4665);
xor U7479 (N_7479,N_3822,N_2765);
nand U7480 (N_7480,N_2737,N_4420);
nand U7481 (N_7481,N_4067,N_4932);
and U7482 (N_7482,N_3213,N_2915);
and U7483 (N_7483,N_4140,N_2507);
nor U7484 (N_7484,N_4098,N_4977);
xnor U7485 (N_7485,N_3206,N_4860);
nor U7486 (N_7486,N_2884,N_2766);
or U7487 (N_7487,N_3748,N_3726);
and U7488 (N_7488,N_4084,N_4250);
xor U7489 (N_7489,N_4470,N_4210);
nor U7490 (N_7490,N_2946,N_3998);
and U7491 (N_7491,N_3519,N_3063);
nor U7492 (N_7492,N_4281,N_4481);
nor U7493 (N_7493,N_4048,N_4148);
or U7494 (N_7494,N_4211,N_3956);
xnor U7495 (N_7495,N_3877,N_3027);
or U7496 (N_7496,N_4249,N_2716);
or U7497 (N_7497,N_4107,N_3721);
and U7498 (N_7498,N_3517,N_2654);
nor U7499 (N_7499,N_4512,N_4326);
and U7500 (N_7500,N_5298,N_7307);
or U7501 (N_7501,N_7461,N_6365);
or U7502 (N_7502,N_6686,N_6375);
nor U7503 (N_7503,N_7399,N_6250);
and U7504 (N_7504,N_6011,N_5612);
nand U7505 (N_7505,N_6346,N_7357);
or U7506 (N_7506,N_5498,N_6502);
nand U7507 (N_7507,N_6040,N_5427);
nor U7508 (N_7508,N_7250,N_5341);
nor U7509 (N_7509,N_5509,N_7288);
and U7510 (N_7510,N_5724,N_6036);
or U7511 (N_7511,N_6195,N_5883);
or U7512 (N_7512,N_7369,N_5809);
or U7513 (N_7513,N_6157,N_5895);
and U7514 (N_7514,N_5260,N_5853);
and U7515 (N_7515,N_7085,N_6003);
nand U7516 (N_7516,N_7016,N_5748);
nor U7517 (N_7517,N_7295,N_6410);
xnor U7518 (N_7518,N_6903,N_5152);
or U7519 (N_7519,N_6837,N_5219);
and U7520 (N_7520,N_6715,N_5258);
nor U7521 (N_7521,N_6906,N_6597);
nand U7522 (N_7522,N_5868,N_5459);
nand U7523 (N_7523,N_6785,N_6997);
or U7524 (N_7524,N_7074,N_5441);
or U7525 (N_7525,N_5326,N_6475);
xnor U7526 (N_7526,N_5127,N_5848);
and U7527 (N_7527,N_5819,N_5079);
nor U7528 (N_7528,N_5769,N_6666);
nor U7529 (N_7529,N_5606,N_6849);
and U7530 (N_7530,N_6136,N_5083);
xor U7531 (N_7531,N_7107,N_5799);
and U7532 (N_7532,N_5491,N_7488);
nand U7533 (N_7533,N_6457,N_6590);
or U7534 (N_7534,N_6249,N_5806);
nand U7535 (N_7535,N_5948,N_5150);
xnor U7536 (N_7536,N_7019,N_5175);
xor U7537 (N_7537,N_6207,N_5858);
nand U7538 (N_7538,N_6438,N_6147);
or U7539 (N_7539,N_5942,N_6587);
nor U7540 (N_7540,N_6662,N_6319);
xnor U7541 (N_7541,N_5979,N_5771);
or U7542 (N_7542,N_5081,N_5843);
nor U7543 (N_7543,N_5148,N_7304);
xor U7544 (N_7544,N_5082,N_6265);
and U7545 (N_7545,N_5654,N_7396);
nand U7546 (N_7546,N_6167,N_7262);
and U7547 (N_7547,N_7240,N_6300);
nand U7548 (N_7548,N_5450,N_6835);
and U7549 (N_7549,N_6152,N_6066);
nand U7550 (N_7550,N_6325,N_7320);
and U7551 (N_7551,N_5707,N_5695);
nor U7552 (N_7552,N_6196,N_7064);
xor U7553 (N_7553,N_5741,N_5835);
and U7554 (N_7554,N_7395,N_5328);
nor U7555 (N_7555,N_5930,N_5734);
xor U7556 (N_7556,N_5121,N_5090);
nand U7557 (N_7557,N_6853,N_6809);
nor U7558 (N_7558,N_5627,N_5779);
and U7559 (N_7559,N_6830,N_6576);
or U7560 (N_7560,N_5305,N_6838);
xnor U7561 (N_7561,N_5009,N_7028);
xor U7562 (N_7562,N_7342,N_7470);
nand U7563 (N_7563,N_6071,N_6347);
xor U7564 (N_7564,N_7466,N_5413);
nor U7565 (N_7565,N_7386,N_5301);
nor U7566 (N_7566,N_6540,N_5006);
xnor U7567 (N_7567,N_5875,N_6428);
nor U7568 (N_7568,N_6851,N_6098);
or U7569 (N_7569,N_5193,N_6240);
or U7570 (N_7570,N_5797,N_6450);
or U7571 (N_7571,N_7242,N_6001);
or U7572 (N_7572,N_7473,N_7227);
or U7573 (N_7573,N_6269,N_5681);
and U7574 (N_7574,N_5173,N_5003);
xor U7575 (N_7575,N_5343,N_6092);
and U7576 (N_7576,N_6627,N_6018);
xnor U7577 (N_7577,N_6914,N_5332);
nor U7578 (N_7578,N_5200,N_6336);
or U7579 (N_7579,N_6205,N_5807);
and U7580 (N_7580,N_5689,N_5302);
nor U7581 (N_7581,N_6416,N_6584);
xnor U7582 (N_7582,N_6977,N_5666);
or U7583 (N_7583,N_6631,N_5608);
nor U7584 (N_7584,N_7257,N_5093);
and U7585 (N_7585,N_6174,N_5635);
nand U7586 (N_7586,N_5557,N_6959);
nor U7587 (N_7587,N_6206,N_5760);
nand U7588 (N_7588,N_6562,N_7026);
or U7589 (N_7589,N_6934,N_5803);
and U7590 (N_7590,N_6060,N_5692);
xor U7591 (N_7591,N_7283,N_6716);
or U7592 (N_7592,N_6923,N_5710);
nand U7593 (N_7593,N_5804,N_6727);
nand U7594 (N_7594,N_7467,N_5656);
or U7595 (N_7595,N_6312,N_6583);
xor U7596 (N_7596,N_7346,N_5435);
nand U7597 (N_7597,N_7476,N_5956);
nor U7598 (N_7598,N_7172,N_6955);
or U7599 (N_7599,N_5368,N_7049);
nor U7600 (N_7600,N_5639,N_6548);
or U7601 (N_7601,N_6537,N_5841);
nand U7602 (N_7602,N_6986,N_5316);
nand U7603 (N_7603,N_6689,N_5629);
and U7604 (N_7604,N_5688,N_6677);
and U7605 (N_7605,N_5837,N_7034);
nor U7606 (N_7606,N_6754,N_7429);
and U7607 (N_7607,N_6799,N_7426);
nand U7608 (N_7608,N_5617,N_5044);
or U7609 (N_7609,N_7224,N_6202);
and U7610 (N_7610,N_6455,N_6027);
nor U7611 (N_7611,N_5560,N_7344);
or U7612 (N_7612,N_6088,N_6432);
nand U7613 (N_7613,N_6637,N_7267);
xnor U7614 (N_7614,N_6035,N_6772);
nand U7615 (N_7615,N_5699,N_6225);
or U7616 (N_7616,N_5691,N_6840);
nor U7617 (N_7617,N_7382,N_5570);
xor U7618 (N_7618,N_7214,N_5318);
or U7619 (N_7619,N_7319,N_6616);
nor U7620 (N_7620,N_5628,N_5477);
nor U7621 (N_7621,N_6013,N_6067);
and U7622 (N_7622,N_6116,N_7389);
and U7623 (N_7623,N_6289,N_5236);
nor U7624 (N_7624,N_5567,N_6952);
xnor U7625 (N_7625,N_6429,N_6151);
xor U7626 (N_7626,N_7316,N_5242);
nand U7627 (N_7627,N_7206,N_6773);
or U7628 (N_7628,N_6413,N_7359);
or U7629 (N_7629,N_5231,N_5733);
nand U7630 (N_7630,N_5890,N_6973);
nand U7631 (N_7631,N_5180,N_6588);
or U7632 (N_7632,N_5167,N_7194);
xnor U7633 (N_7633,N_6976,N_6126);
nor U7634 (N_7634,N_5047,N_7237);
nand U7635 (N_7635,N_5631,N_5888);
and U7636 (N_7636,N_5506,N_5754);
xor U7637 (N_7637,N_5387,N_5214);
nand U7638 (N_7638,N_6551,N_6466);
nand U7639 (N_7639,N_6102,N_6443);
and U7640 (N_7640,N_7139,N_7037);
nand U7641 (N_7641,N_6259,N_5663);
nand U7642 (N_7642,N_6814,N_6002);
or U7643 (N_7643,N_5511,N_7373);
or U7644 (N_7644,N_5962,N_6639);
nand U7645 (N_7645,N_6882,N_5789);
and U7646 (N_7646,N_5985,N_6270);
or U7647 (N_7647,N_6056,N_5537);
xor U7648 (N_7648,N_6385,N_6142);
nor U7649 (N_7649,N_5008,N_6076);
and U7650 (N_7650,N_6471,N_6957);
nor U7651 (N_7651,N_6915,N_7286);
or U7652 (N_7652,N_5622,N_6982);
xor U7653 (N_7653,N_5582,N_5233);
nand U7654 (N_7654,N_6039,N_5542);
nand U7655 (N_7655,N_5857,N_6953);
nor U7656 (N_7656,N_5422,N_6185);
nor U7657 (N_7657,N_5181,N_5208);
or U7658 (N_7658,N_6841,N_6184);
nor U7659 (N_7659,N_7315,N_5292);
or U7660 (N_7660,N_7383,N_6761);
and U7661 (N_7661,N_6258,N_5348);
and U7662 (N_7662,N_5021,N_5675);
nor U7663 (N_7663,N_7090,N_6508);
nand U7664 (N_7664,N_5907,N_6006);
nor U7665 (N_7665,N_5275,N_7308);
and U7666 (N_7666,N_7495,N_5667);
nor U7667 (N_7667,N_5482,N_6424);
or U7668 (N_7668,N_7173,N_6296);
and U7669 (N_7669,N_5201,N_5244);
nor U7670 (N_7670,N_5241,N_7123);
and U7671 (N_7671,N_6379,N_6941);
and U7672 (N_7672,N_7013,N_6777);
nor U7673 (N_7673,N_7329,N_7324);
nand U7674 (N_7674,N_7217,N_6740);
nand U7675 (N_7675,N_5988,N_6722);
nand U7676 (N_7676,N_6218,N_6489);
or U7677 (N_7677,N_6030,N_6504);
nand U7678 (N_7678,N_7287,N_6893);
and U7679 (N_7679,N_6494,N_7441);
and U7680 (N_7680,N_6924,N_5794);
or U7681 (N_7681,N_7118,N_7143);
or U7682 (N_7682,N_6491,N_6931);
xor U7683 (N_7683,N_6978,N_7478);
nand U7684 (N_7684,N_6238,N_6546);
nand U7685 (N_7685,N_5598,N_6658);
xnor U7686 (N_7686,N_5320,N_6598);
or U7687 (N_7687,N_6956,N_5410);
xnor U7688 (N_7688,N_7141,N_5307);
nor U7689 (N_7689,N_7185,N_6527);
nand U7690 (N_7690,N_7100,N_5209);
and U7691 (N_7691,N_6589,N_7481);
nor U7692 (N_7692,N_7387,N_5863);
nand U7693 (N_7693,N_6900,N_5994);
nand U7694 (N_7694,N_5869,N_6372);
xor U7695 (N_7695,N_7174,N_5762);
or U7696 (N_7696,N_5404,N_6887);
xor U7697 (N_7697,N_5614,N_6493);
nor U7698 (N_7698,N_5932,N_5892);
and U7699 (N_7699,N_7246,N_6163);
nor U7700 (N_7700,N_5960,N_6612);
nor U7701 (N_7701,N_6282,N_6768);
and U7702 (N_7702,N_7079,N_5155);
and U7703 (N_7703,N_5945,N_7021);
nand U7704 (N_7704,N_5703,N_7380);
or U7705 (N_7705,N_6848,N_6257);
xnor U7706 (N_7706,N_7269,N_5507);
or U7707 (N_7707,N_6353,N_5362);
or U7708 (N_7708,N_6842,N_5553);
and U7709 (N_7709,N_6520,N_5177);
or U7710 (N_7710,N_7397,N_5522);
and U7711 (N_7711,N_6580,N_6525);
and U7712 (N_7712,N_6005,N_6125);
xnor U7713 (N_7713,N_6171,N_7419);
xor U7714 (N_7714,N_6180,N_6912);
xnor U7715 (N_7715,N_6884,N_6401);
nor U7716 (N_7716,N_6788,N_5329);
or U7717 (N_7717,N_7440,N_7213);
nor U7718 (N_7718,N_6779,N_5935);
and U7719 (N_7719,N_7136,N_7303);
nand U7720 (N_7720,N_5034,N_5494);
or U7721 (N_7721,N_5451,N_6097);
and U7722 (N_7722,N_6950,N_5564);
nand U7723 (N_7723,N_6419,N_7198);
nand U7724 (N_7724,N_7444,N_5687);
xor U7725 (N_7725,N_5538,N_6405);
nand U7726 (N_7726,N_5102,N_5030);
nand U7727 (N_7727,N_6750,N_6753);
or U7728 (N_7728,N_5073,N_5153);
xor U7729 (N_7729,N_6690,N_7219);
nand U7730 (N_7730,N_7105,N_7375);
nand U7731 (N_7731,N_5176,N_6642);
xor U7732 (N_7732,N_6684,N_5709);
xnor U7733 (N_7733,N_5203,N_5775);
and U7734 (N_7734,N_5097,N_5665);
or U7735 (N_7735,N_5826,N_7263);
nand U7736 (N_7736,N_6256,N_6996);
or U7737 (N_7737,N_7483,N_6963);
nor U7738 (N_7738,N_6267,N_7372);
nor U7739 (N_7739,N_5322,N_6513);
nor U7740 (N_7740,N_7042,N_6127);
nand U7741 (N_7741,N_6665,N_6942);
nor U7742 (N_7742,N_7111,N_6488);
nor U7743 (N_7743,N_6515,N_7443);
and U7744 (N_7744,N_5284,N_7068);
xor U7745 (N_7745,N_5955,N_6625);
nand U7746 (N_7746,N_5727,N_5984);
nand U7747 (N_7747,N_5142,N_5221);
or U7748 (N_7748,N_5766,N_5504);
and U7749 (N_7749,N_6691,N_5597);
nand U7750 (N_7750,N_5917,N_6767);
and U7751 (N_7751,N_5070,N_6749);
nand U7752 (N_7752,N_6200,N_7158);
and U7753 (N_7753,N_5376,N_5723);
xnor U7754 (N_7754,N_5212,N_5908);
xor U7755 (N_7755,N_6212,N_5356);
nand U7756 (N_7756,N_5293,N_5109);
nor U7757 (N_7757,N_6993,N_5901);
and U7758 (N_7758,N_7363,N_6723);
nor U7759 (N_7759,N_6254,N_5415);
nand U7760 (N_7760,N_5836,N_6641);
xor U7761 (N_7761,N_7184,N_5026);
and U7762 (N_7762,N_7255,N_5473);
and U7763 (N_7763,N_6468,N_6605);
and U7764 (N_7764,N_7349,N_5630);
xor U7765 (N_7765,N_6281,N_6521);
and U7766 (N_7766,N_5334,N_5669);
and U7767 (N_7767,N_5573,N_5434);
and U7768 (N_7768,N_5678,N_6861);
or U7769 (N_7769,N_6738,N_5920);
xnor U7770 (N_7770,N_7428,N_5999);
nor U7771 (N_7771,N_6949,N_7417);
nor U7772 (N_7772,N_6037,N_7088);
xor U7773 (N_7773,N_6038,N_6181);
nor U7774 (N_7774,N_6463,N_6057);
or U7775 (N_7775,N_7264,N_7345);
or U7776 (N_7776,N_5829,N_7390);
or U7777 (N_7777,N_5572,N_5157);
and U7778 (N_7778,N_6310,N_5753);
or U7779 (N_7779,N_7080,N_5261);
nand U7780 (N_7780,N_7017,N_5299);
nor U7781 (N_7781,N_6823,N_7254);
xnor U7782 (N_7782,N_5425,N_6918);
xnor U7783 (N_7783,N_5449,N_5374);
nor U7784 (N_7784,N_5549,N_7289);
xor U7785 (N_7785,N_6330,N_5736);
or U7786 (N_7786,N_6131,N_6119);
xnor U7787 (N_7787,N_6467,N_5717);
nor U7788 (N_7788,N_5478,N_5981);
and U7789 (N_7789,N_5772,N_7492);
xor U7790 (N_7790,N_7146,N_6436);
or U7791 (N_7791,N_6129,N_5162);
or U7792 (N_7792,N_5038,N_7196);
and U7793 (N_7793,N_7234,N_5353);
nand U7794 (N_7794,N_7048,N_6922);
nand U7795 (N_7795,N_6190,N_7140);
xnor U7796 (N_7796,N_6178,N_6549);
nand U7797 (N_7797,N_6247,N_5308);
nor U7798 (N_7798,N_7299,N_5787);
xor U7799 (N_7799,N_7258,N_7355);
or U7800 (N_7800,N_6813,N_5497);
nor U7801 (N_7801,N_6573,N_6411);
xor U7802 (N_7802,N_5202,N_5972);
or U7803 (N_7803,N_5096,N_5566);
nor U7804 (N_7804,N_5555,N_5586);
and U7805 (N_7805,N_7498,N_5124);
nand U7806 (N_7806,N_6807,N_6182);
xnor U7807 (N_7807,N_7167,N_5912);
xor U7808 (N_7808,N_5013,N_6453);
and U7809 (N_7809,N_7392,N_5898);
or U7810 (N_7810,N_5938,N_5500);
or U7811 (N_7811,N_7010,N_7485);
or U7812 (N_7812,N_5195,N_5130);
nor U7813 (N_7813,N_7256,N_5035);
nor U7814 (N_7814,N_5554,N_5158);
or U7815 (N_7815,N_5269,N_5854);
xor U7816 (N_7816,N_6928,N_5874);
or U7817 (N_7817,N_7362,N_7402);
or U7818 (N_7818,N_6728,N_6121);
nor U7819 (N_7819,N_6008,N_7023);
and U7820 (N_7820,N_6448,N_6652);
nand U7821 (N_7821,N_7171,N_5726);
xor U7822 (N_7822,N_6248,N_6804);
nor U7823 (N_7823,N_6048,N_7032);
and U7824 (N_7824,N_6629,N_6427);
nand U7825 (N_7825,N_5087,N_7416);
xnor U7826 (N_7826,N_6122,N_5565);
nand U7827 (N_7827,N_6026,N_6093);
and U7828 (N_7828,N_5855,N_5483);
xor U7829 (N_7829,N_6209,N_5010);
and U7830 (N_7830,N_5024,N_5360);
or U7831 (N_7831,N_7115,N_5611);
and U7832 (N_7832,N_6341,N_5864);
and U7833 (N_7833,N_6704,N_5118);
nor U7834 (N_7834,N_6937,N_6158);
nand U7835 (N_7835,N_7144,N_5562);
and U7836 (N_7836,N_5983,N_7350);
nand U7837 (N_7837,N_6472,N_6197);
or U7838 (N_7838,N_7103,N_5987);
xnor U7839 (N_7839,N_5408,N_6675);
nor U7840 (N_7840,N_6337,N_5139);
and U7841 (N_7841,N_5099,N_6224);
or U7842 (N_7842,N_6332,N_6892);
nand U7843 (N_7843,N_5941,N_5949);
nor U7844 (N_7844,N_5147,N_6029);
nand U7845 (N_7845,N_5409,N_5759);
nand U7846 (N_7846,N_5354,N_7321);
nor U7847 (N_7847,N_5250,N_5315);
or U7848 (N_7848,N_5844,N_7168);
nand U7849 (N_7849,N_6371,N_5007);
nand U7850 (N_7850,N_6721,N_6115);
and U7851 (N_7851,N_6363,N_6021);
or U7852 (N_7852,N_5438,N_7069);
xnor U7853 (N_7853,N_6795,N_5278);
nand U7854 (N_7854,N_5017,N_7216);
or U7855 (N_7855,N_5108,N_5849);
or U7856 (N_7856,N_5532,N_5032);
nand U7857 (N_7857,N_5080,N_6528);
and U7858 (N_7858,N_7273,N_5990);
nor U7859 (N_7859,N_6594,N_5004);
nand U7860 (N_7860,N_6083,N_5590);
nor U7861 (N_7861,N_5452,N_7211);
or U7862 (N_7862,N_6854,N_7465);
or U7863 (N_7863,N_6441,N_6734);
nand U7864 (N_7864,N_7294,N_6473);
and U7865 (N_7865,N_7005,N_7433);
nand U7866 (N_7866,N_6791,N_6031);
and U7867 (N_7867,N_6975,N_6737);
xor U7868 (N_7868,N_6656,N_7029);
nor U7869 (N_7869,N_7499,N_6309);
nand U7870 (N_7870,N_7460,N_7108);
or U7871 (N_7871,N_5971,N_6064);
or U7872 (N_7872,N_6603,N_5933);
and U7873 (N_7873,N_7043,N_7430);
nand U7874 (N_7874,N_7089,N_5782);
nor U7875 (N_7875,N_6387,N_7277);
or U7876 (N_7876,N_6503,N_5963);
nor U7877 (N_7877,N_6266,N_5385);
nand U7878 (N_7878,N_6112,N_7189);
or U7879 (N_7879,N_5243,N_6681);
and U7880 (N_7880,N_5902,N_6481);
xnor U7881 (N_7881,N_5685,N_6072);
xnor U7882 (N_7882,N_6518,N_6794);
and U7883 (N_7883,N_6869,N_5897);
or U7884 (N_7884,N_6340,N_5580);
xor U7885 (N_7885,N_5001,N_6313);
xnor U7886 (N_7886,N_6783,N_7347);
xor U7887 (N_7887,N_5915,N_5876);
and U7888 (N_7888,N_5071,N_6231);
xor U7889 (N_7889,N_6291,N_6577);
xor U7890 (N_7890,N_6553,N_5896);
xnor U7891 (N_7891,N_7431,N_7052);
nand U7892 (N_7892,N_5045,N_5123);
xor U7893 (N_7893,N_7325,N_7364);
or U7894 (N_7894,N_7450,N_5750);
nand U7895 (N_7895,N_7147,N_6169);
nor U7896 (N_7896,N_6138,N_5997);
and U7897 (N_7897,N_7051,N_5816);
or U7898 (N_7898,N_7367,N_5976);
nand U7899 (N_7899,N_5460,N_7312);
xor U7900 (N_7900,N_6490,N_6954);
nor U7901 (N_7901,N_5811,N_6500);
or U7902 (N_7902,N_6049,N_5392);
xor U7903 (N_7903,N_7082,N_6089);
nor U7904 (N_7904,N_5563,N_5216);
and U7905 (N_7905,N_7117,N_5937);
xor U7906 (N_7906,N_7487,N_6078);
nand U7907 (N_7907,N_6331,N_5349);
or U7908 (N_7908,N_6251,N_7400);
and U7909 (N_7909,N_5683,N_5711);
or U7910 (N_7910,N_6868,N_6285);
xor U7911 (N_7911,N_6776,N_7393);
nor U7912 (N_7912,N_6077,N_6646);
nand U7913 (N_7913,N_6099,N_5469);
and U7914 (N_7914,N_5325,N_5199);
nand U7915 (N_7915,N_5110,N_5223);
nor U7916 (N_7916,N_5649,N_7463);
nand U7917 (N_7917,N_7275,N_7233);
nand U7918 (N_7918,N_5253,N_5684);
xor U7919 (N_7919,N_7131,N_7220);
nand U7920 (N_7920,N_5066,N_6510);
and U7921 (N_7921,N_6921,N_6349);
nor U7922 (N_7922,N_7129,N_5197);
or U7923 (N_7923,N_6446,N_6678);
and U7924 (N_7924,N_5089,N_5129);
nor U7925 (N_7925,N_5747,N_6406);
or U7926 (N_7926,N_5461,N_5964);
and U7927 (N_7927,N_5394,N_6644);
nor U7928 (N_7928,N_5817,N_5196);
or U7929 (N_7929,N_5444,N_7435);
and U7930 (N_7930,N_6302,N_6017);
nand U7931 (N_7931,N_7109,N_6237);
nor U7932 (N_7932,N_5183,N_5036);
nor U7933 (N_7933,N_6960,N_7496);
or U7934 (N_7934,N_5485,N_6367);
nand U7935 (N_7935,N_5805,N_5655);
nand U7936 (N_7936,N_5852,N_7271);
and U7937 (N_7937,N_7002,N_5700);
and U7938 (N_7938,N_5029,N_5107);
nand U7939 (N_7939,N_7418,N_5551);
nor U7940 (N_7940,N_7170,N_6219);
and U7941 (N_7941,N_5247,N_5455);
nor U7942 (N_7942,N_6400,N_5982);
xor U7943 (N_7943,N_7353,N_6775);
nand U7944 (N_7944,N_5479,N_5263);
and U7945 (N_7945,N_5281,N_5831);
and U7946 (N_7946,N_6966,N_6998);
nand U7947 (N_7947,N_6465,N_7165);
xor U7948 (N_7948,N_6211,N_6929);
and U7949 (N_7949,N_6058,N_5397);
nor U7950 (N_7950,N_7083,N_5384);
nand U7951 (N_7951,N_5330,N_6707);
nor U7952 (N_7952,N_5731,N_6144);
nor U7953 (N_7953,N_7130,N_6994);
and U7954 (N_7954,N_5346,N_5406);
or U7955 (N_7955,N_5421,N_6556);
xor U7956 (N_7956,N_5464,N_5820);
nand U7957 (N_7957,N_5046,N_6041);
xor U7958 (N_7958,N_5174,N_5788);
nor U7959 (N_7959,N_6514,N_5350);
nand U7960 (N_7960,N_5310,N_6735);
nor U7961 (N_7961,N_6160,N_5680);
nor U7962 (N_7962,N_5420,N_6007);
xor U7963 (N_7963,N_6608,N_5168);
xor U7964 (N_7964,N_6307,N_7314);
or U7965 (N_7965,N_6139,N_7469);
xnor U7966 (N_7966,N_7007,N_5648);
and U7967 (N_7967,N_7067,N_6595);
nor U7968 (N_7968,N_5641,N_5610);
nand U7969 (N_7969,N_6106,N_7221);
nor U7970 (N_7970,N_7341,N_6022);
or U7971 (N_7971,N_5238,N_5673);
nor U7972 (N_7972,N_5252,N_5373);
or U7973 (N_7973,N_5800,N_7479);
nor U7974 (N_7974,N_5529,N_5053);
xor U7975 (N_7975,N_6718,N_5146);
nand U7976 (N_7976,N_5513,N_6054);
nor U7977 (N_7977,N_6784,N_6283);
or U7978 (N_7978,N_6230,N_5501);
nor U7979 (N_7979,N_5881,N_5132);
nand U7980 (N_7980,N_6452,N_5913);
nand U7981 (N_7981,N_6124,N_6389);
or U7982 (N_7982,N_5458,N_6085);
or U7983 (N_7983,N_6660,N_5671);
and U7984 (N_7984,N_7145,N_5120);
xor U7985 (N_7985,N_5169,N_5502);
nand U7986 (N_7986,N_6599,N_6541);
or U7987 (N_7987,N_6564,N_6606);
or U7988 (N_7988,N_5402,N_7120);
and U7989 (N_7989,N_5211,N_6091);
xnor U7990 (N_7990,N_5583,N_6864);
or U7991 (N_7991,N_6559,N_7457);
xnor U7992 (N_7992,N_5114,N_6486);
and U7993 (N_7993,N_5939,N_6290);
xnor U7994 (N_7994,N_5192,N_5732);
or U7995 (N_7995,N_5069,N_6961);
or U7996 (N_7996,N_6748,N_6110);
nor U7997 (N_7997,N_5134,N_5388);
xor U7998 (N_7998,N_6586,N_5465);
nor U7999 (N_7999,N_6709,N_5467);
and U8000 (N_8000,N_7057,N_6732);
nor U8001 (N_8001,N_6593,N_5792);
and U8002 (N_8002,N_6246,N_6947);
nand U8003 (N_8003,N_5363,N_7412);
nand U8004 (N_8004,N_5623,N_6671);
and U8005 (N_8005,N_5189,N_5742);
or U8006 (N_8006,N_6275,N_6812);
or U8007 (N_8007,N_5423,N_7408);
and U8008 (N_8008,N_5257,N_6778);
nor U8009 (N_8009,N_5128,N_6635);
or U8010 (N_8010,N_6565,N_6945);
or U8011 (N_8011,N_6645,N_7244);
or U8012 (N_8012,N_6033,N_5761);
xnor U8013 (N_8013,N_7063,N_7285);
and U8014 (N_8014,N_6798,N_7322);
and U8015 (N_8015,N_5975,N_7199);
nand U8016 (N_8016,N_6896,N_6262);
or U8017 (N_8017,N_5492,N_6053);
nor U8018 (N_8018,N_5443,N_6782);
and U8019 (N_8019,N_6557,N_5416);
xor U8020 (N_8020,N_5028,N_6700);
nand U8021 (N_8021,N_7296,N_6757);
and U8022 (N_8022,N_7053,N_6162);
nor U8023 (N_8023,N_6739,N_5633);
xnor U8024 (N_8024,N_7035,N_5210);
and U8025 (N_8025,N_5220,N_6897);
nor U8026 (N_8026,N_6423,N_6187);
and U8027 (N_8027,N_6123,N_5135);
nand U8028 (N_8028,N_7310,N_7114);
xnor U8029 (N_8029,N_5861,N_6421);
nand U8030 (N_8030,N_6601,N_6705);
nor U8031 (N_8031,N_7468,N_6096);
nor U8032 (N_8032,N_6045,N_5321);
and U8033 (N_8033,N_7116,N_6261);
or U8034 (N_8034,N_7332,N_6082);
xnor U8035 (N_8035,N_7012,N_6746);
nor U8036 (N_8036,N_5505,N_5914);
nor U8037 (N_8037,N_6926,N_6201);
nand U8038 (N_8038,N_5967,N_5558);
or U8039 (N_8039,N_6633,N_6189);
nand U8040 (N_8040,N_6025,N_6352);
xor U8041 (N_8041,N_6862,N_7177);
or U8042 (N_8042,N_5020,N_5067);
nand U8043 (N_8043,N_6663,N_6217);
and U8044 (N_8044,N_7014,N_7045);
xor U8045 (N_8045,N_5815,N_6647);
and U8046 (N_8046,N_5661,N_7071);
xor U8047 (N_8047,N_7218,N_5859);
or U8048 (N_8048,N_7421,N_6322);
nor U8049 (N_8049,N_6643,N_6909);
nor U8050 (N_8050,N_6519,N_5701);
xor U8051 (N_8051,N_5822,N_6154);
or U8052 (N_8052,N_6758,N_6888);
nand U8053 (N_8053,N_5287,N_6276);
nor U8054 (N_8054,N_5105,N_5206);
xor U8055 (N_8055,N_6374,N_6725);
or U8056 (N_8056,N_7403,N_5585);
nor U8057 (N_8057,N_6274,N_6860);
and U8058 (N_8058,N_7309,N_5539);
nand U8059 (N_8059,N_7381,N_6000);
or U8060 (N_8060,N_5286,N_6944);
or U8061 (N_8061,N_6579,N_6324);
nand U8062 (N_8062,N_6165,N_5618);
and U8063 (N_8063,N_6544,N_5818);
and U8064 (N_8064,N_5524,N_5885);
nand U8065 (N_8065,N_7405,N_6971);
nand U8066 (N_8066,N_5926,N_5704);
or U8067 (N_8067,N_5922,N_5104);
xnor U8068 (N_8068,N_7272,N_6113);
and U8069 (N_8069,N_7484,N_5918);
nand U8070 (N_8070,N_6227,N_7148);
and U8071 (N_8071,N_6417,N_5910);
and U8072 (N_8072,N_5375,N_6640);
or U8073 (N_8073,N_5825,N_6609);
nor U8074 (N_8074,N_6268,N_5791);
and U8075 (N_8075,N_6885,N_6895);
nand U8076 (N_8076,N_6570,N_6523);
nor U8077 (N_8077,N_5845,N_6526);
or U8078 (N_8078,N_5871,N_6199);
nor U8079 (N_8079,N_6623,N_5550);
and U8080 (N_8080,N_5802,N_5369);
or U8081 (N_8081,N_6143,N_7331);
xnor U8082 (N_8082,N_5378,N_7414);
nor U8083 (N_8083,N_7128,N_5407);
xnor U8084 (N_8084,N_6808,N_6370);
nand U8085 (N_8085,N_6245,N_5453);
xnor U8086 (N_8086,N_6009,N_5323);
and U8087 (N_8087,N_5778,N_6898);
nor U8088 (N_8088,N_6284,N_6981);
or U8089 (N_8089,N_5651,N_5647);
xor U8090 (N_8090,N_6153,N_5265);
xor U8091 (N_8091,N_6555,N_5653);
or U8092 (N_8092,N_7081,N_5725);
xnor U8093 (N_8093,N_6685,N_5674);
and U8094 (N_8094,N_7249,N_5893);
xnor U8095 (N_8095,N_7138,N_5514);
nand U8096 (N_8096,N_5117,N_5952);
xor U8097 (N_8097,N_6456,N_7388);
xor U8098 (N_8098,N_7352,N_7232);
or U8099 (N_8099,N_5929,N_5961);
xnor U8100 (N_8100,N_7006,N_6213);
nand U8101 (N_8101,N_6745,N_6702);
nand U8102 (N_8102,N_5541,N_5064);
and U8103 (N_8103,N_5528,N_5904);
nand U8104 (N_8104,N_6381,N_6080);
nand U8105 (N_8105,N_6826,N_6989);
or U8106 (N_8106,N_5398,N_7348);
nand U8107 (N_8107,N_5578,N_6908);
nor U8108 (N_8108,N_6538,N_6350);
nor U8109 (N_8109,N_6787,N_7274);
nor U8110 (N_8110,N_6815,N_7084);
nand U8111 (N_8111,N_6793,N_6339);
nand U8112 (N_8112,N_6974,N_6891);
nor U8113 (N_8113,N_5970,N_5518);
or U8114 (N_8114,N_6827,N_6889);
xnor U8115 (N_8115,N_6962,N_6818);
or U8116 (N_8116,N_7235,N_6533);
or U8117 (N_8117,N_6344,N_5285);
or U8118 (N_8118,N_6602,N_6176);
xnor U8119 (N_8119,N_5182,N_5361);
nor U8120 (N_8120,N_5448,N_6755);
nand U8121 (N_8121,N_6354,N_7305);
nor U8122 (N_8122,N_5367,N_6930);
nand U8123 (N_8123,N_6843,N_6409);
xnor U8124 (N_8124,N_7062,N_6697);
xnor U8125 (N_8125,N_7191,N_5993);
nor U8126 (N_8126,N_5016,N_6272);
xor U8127 (N_8127,N_7186,N_7385);
nor U8128 (N_8128,N_6415,N_6764);
or U8129 (N_8129,N_5098,N_5763);
nor U8130 (N_8130,N_6487,N_6051);
or U8131 (N_8131,N_6391,N_5927);
and U8132 (N_8132,N_5022,N_5712);
nand U8133 (N_8133,N_6877,N_6844);
xor U8134 (N_8134,N_6028,N_7236);
or U8135 (N_8135,N_5774,N_5115);
and U8136 (N_8136,N_6306,N_6694);
xnor U8137 (N_8137,N_5031,N_5968);
nand U8138 (N_8138,N_5355,N_6979);
nor U8139 (N_8139,N_5306,N_7125);
nand U8140 (N_8140,N_7009,N_6780);
or U8141 (N_8141,N_6856,N_5051);
xor U8142 (N_8142,N_5921,N_7486);
or U8143 (N_8143,N_6693,N_6484);
xnor U8144 (N_8144,N_5950,N_6607);
nor U8145 (N_8145,N_6545,N_6696);
nand U8146 (N_8146,N_5877,N_5217);
xor U8147 (N_8147,N_5535,N_5379);
xnor U8148 (N_8148,N_5224,N_6592);
xor U8149 (N_8149,N_6024,N_6939);
nand U8150 (N_8150,N_5426,N_6907);
or U8151 (N_8151,N_6717,N_6109);
or U8152 (N_8152,N_6995,N_6600);
xnor U8153 (N_8153,N_6398,N_6507);
or U8154 (N_8154,N_5256,N_5439);
nand U8155 (N_8155,N_6087,N_7132);
xor U8156 (N_8156,N_5944,N_7284);
xor U8157 (N_8157,N_5290,N_7230);
or U8158 (N_8158,N_6461,N_5254);
nor U8159 (N_8159,N_5440,N_5446);
xnor U8160 (N_8160,N_5312,N_5919);
xnor U8161 (N_8161,N_5714,N_5718);
or U8162 (N_8162,N_7087,N_6015);
nand U8163 (N_8163,N_5205,N_6569);
nor U8164 (N_8164,N_5411,N_7252);
nand U8165 (N_8165,N_5697,N_7384);
and U8166 (N_8166,N_7047,N_6010);
nor U8167 (N_8167,N_5481,N_5417);
xnor U8168 (N_8168,N_7241,N_7178);
nand U8169 (N_8169,N_6140,N_6550);
nor U8170 (N_8170,N_5170,N_5995);
nand U8171 (N_8171,N_5634,N_5846);
nand U8172 (N_8172,N_7127,N_6621);
nand U8173 (N_8173,N_6299,N_5632);
nor U8174 (N_8174,N_5272,N_5644);
nor U8175 (N_8175,N_6175,N_5342);
and U8176 (N_8176,N_6801,N_5989);
and U8177 (N_8177,N_5784,N_6317);
or U8178 (N_8178,N_6865,N_5380);
nor U8179 (N_8179,N_5100,N_5659);
or U8180 (N_8180,N_5412,N_6477);
xor U8181 (N_8181,N_6408,N_6388);
and U8182 (N_8182,N_6790,N_5277);
xor U8183 (N_8183,N_7432,N_6019);
nor U8184 (N_8184,N_5282,N_6591);
or U8185 (N_8185,N_5738,N_5592);
and U8186 (N_8186,N_5642,N_6412);
or U8187 (N_8187,N_5002,N_6380);
xnor U8188 (N_8188,N_6204,N_5672);
or U8189 (N_8189,N_5145,N_6133);
nor U8190 (N_8190,N_7439,N_7300);
or U8191 (N_8191,N_6902,N_6676);
and U8192 (N_8192,N_6321,N_5602);
xnor U8193 (N_8193,N_6571,N_7197);
or U8194 (N_8194,N_5042,N_5239);
nand U8195 (N_8195,N_5204,N_7354);
or U8196 (N_8196,N_6137,N_5386);
nor U8197 (N_8197,N_6667,N_5433);
and U8198 (N_8198,N_6933,N_5978);
nand U8199 (N_8199,N_5588,N_5297);
or U8200 (N_8200,N_5041,N_7041);
xnor U8201 (N_8201,N_7360,N_5823);
and U8202 (N_8202,N_6260,N_6418);
and U8203 (N_8203,N_6214,N_5977);
xnor U8204 (N_8204,N_6578,N_5546);
nand U8205 (N_8205,N_6442,N_5954);
or U8206 (N_8206,N_5548,N_5043);
xor U8207 (N_8207,N_7030,N_5499);
or U8208 (N_8208,N_5057,N_6476);
nor U8209 (N_8209,N_6358,N_6919);
nand U8210 (N_8210,N_6617,N_5543);
xor U8211 (N_8211,N_5765,N_6708);
xnor U8212 (N_8212,N_6348,N_6743);
or U8213 (N_8213,N_5515,N_5000);
and U8214 (N_8214,N_7494,N_5974);
or U8215 (N_8215,N_5911,N_6111);
and U8216 (N_8216,N_7456,N_6242);
and U8217 (N_8217,N_5657,N_5601);
xor U8218 (N_8218,N_5735,N_7202);
nor U8219 (N_8219,N_6711,N_5640);
xnor U8220 (N_8220,N_6469,N_6839);
and U8221 (N_8221,N_7424,N_6055);
or U8222 (N_8222,N_6378,N_6886);
or U8223 (N_8223,N_6480,N_6414);
nand U8224 (N_8224,N_5471,N_6539);
or U8225 (N_8225,N_5084,N_7245);
and U8226 (N_8226,N_6552,N_5625);
nor U8227 (N_8227,N_6073,N_6524);
and U8228 (N_8228,N_6014,N_6451);
xor U8229 (N_8229,N_5251,N_7268);
nor U8230 (N_8230,N_5812,N_6345);
xnor U8231 (N_8231,N_6634,N_6670);
nand U8232 (N_8232,N_6714,N_6867);
nor U8233 (N_8233,N_5382,N_5596);
or U8234 (N_8234,N_6881,N_7215);
and U8235 (N_8235,N_6831,N_5338);
and U8236 (N_8236,N_7075,N_5370);
or U8237 (N_8237,N_6188,N_5643);
xor U8238 (N_8238,N_6873,N_6572);
or U8239 (N_8239,N_7453,N_6649);
xor U8240 (N_8240,N_5533,N_5092);
or U8241 (N_8241,N_5273,N_6090);
or U8242 (N_8242,N_7124,N_5670);
and U8243 (N_8243,N_5015,N_7160);
xnor U8244 (N_8244,N_6653,N_6287);
or U8245 (N_8245,N_7420,N_6392);
nand U8246 (N_8246,N_7336,N_6004);
and U8247 (N_8247,N_6426,N_5076);
xor U8248 (N_8248,N_6252,N_7302);
xnor U8249 (N_8249,N_6614,N_5545);
nor U8250 (N_8250,N_7207,N_7182);
and U8251 (N_8251,N_7126,N_5014);
or U8252 (N_8252,N_7454,N_7327);
nand U8253 (N_8253,N_5645,N_5101);
and U8254 (N_8254,N_5715,N_5445);
nor U8255 (N_8255,N_6292,N_6916);
nor U8256 (N_8256,N_7458,N_6431);
or U8257 (N_8257,N_5781,N_7401);
or U8258 (N_8258,N_6910,N_5757);
xnor U8259 (N_8259,N_6806,N_7436);
nand U8260 (N_8260,N_5600,N_6876);
and U8261 (N_8261,N_7061,N_5577);
nand U8262 (N_8262,N_5389,N_6970);
nand U8263 (N_8263,N_5810,N_5698);
nor U8264 (N_8264,N_7413,N_7205);
nor U8265 (N_8265,N_5279,N_6482);
and U8266 (N_8266,N_7104,N_7210);
nand U8267 (N_8267,N_5973,N_6568);
nor U8268 (N_8268,N_5605,N_5335);
or U8269 (N_8269,N_5719,N_5793);
nand U8270 (N_8270,N_7151,N_5584);
or U8271 (N_8271,N_7292,N_6604);
and U8272 (N_8272,N_7093,N_6951);
nand U8273 (N_8273,N_5517,N_6852);
xor U8274 (N_8274,N_7459,N_5493);
nor U8275 (N_8275,N_6279,N_5424);
xor U8276 (N_8276,N_6803,N_5027);
and U8277 (N_8277,N_7175,N_5112);
xor U8278 (N_8278,N_6766,N_6731);
nor U8279 (N_8279,N_5474,N_5255);
nor U8280 (N_8280,N_7406,N_5786);
nand U8281 (N_8281,N_7471,N_5126);
nor U8282 (N_8282,N_7119,N_6874);
and U8283 (N_8283,N_6377,N_5821);
nor U8284 (N_8284,N_5767,N_5716);
nand U8285 (N_8285,N_6183,N_6105);
nand U8286 (N_8286,N_6509,N_6563);
nand U8287 (N_8287,N_5225,N_5894);
and U8288 (N_8288,N_7169,N_6792);
nor U8289 (N_8289,N_6899,N_5222);
xor U8290 (N_8290,N_7181,N_5058);
or U8291 (N_8291,N_5730,N_7427);
and U8292 (N_8292,N_5151,N_6301);
nor U8293 (N_8293,N_7192,N_5052);
xor U8294 (N_8294,N_7204,N_6624);
nand U8295 (N_8295,N_6134,N_7092);
nor U8296 (N_8296,N_5237,N_7445);
and U8297 (N_8297,N_7162,N_5059);
nor U8298 (N_8298,N_5228,N_7377);
and U8299 (N_8299,N_7366,N_7229);
nand U8300 (N_8300,N_7133,N_7096);
nand U8301 (N_8301,N_6913,N_7365);
nand U8302 (N_8302,N_7154,N_6575);
nor U8303 (N_8303,N_7356,N_5746);
nor U8304 (N_8304,N_6501,N_6304);
and U8305 (N_8305,N_7368,N_6173);
nor U8306 (N_8306,N_5457,N_7449);
or U8307 (N_8307,N_5525,N_7166);
nand U8308 (N_8308,N_6706,N_5531);
or U8309 (N_8309,N_6434,N_5106);
nand U8310 (N_8310,N_5740,N_6547);
nor U8311 (N_8311,N_6765,N_5873);
nand U8312 (N_8312,N_6872,N_7279);
nor U8313 (N_8313,N_6742,N_5696);
or U8314 (N_8314,N_7438,N_6940);
or U8315 (N_8315,N_5055,N_7340);
nor U8316 (N_8316,N_6314,N_5739);
and U8317 (N_8317,N_5547,N_7200);
xnor U8318 (N_8318,N_6511,N_5054);
xnor U8319 (N_8319,N_6984,N_7054);
and U8320 (N_8320,N_5116,N_7328);
xor U8321 (N_8321,N_5133,N_6741);
and U8322 (N_8322,N_5998,N_5957);
and U8323 (N_8323,N_6439,N_5149);
nor U8324 (N_8324,N_6294,N_5432);
nand U8325 (N_8325,N_6836,N_5160);
and U8326 (N_8326,N_6050,N_5347);
nand U8327 (N_8327,N_6359,N_6239);
or U8328 (N_8328,N_5796,N_7095);
nand U8329 (N_8329,N_7078,N_6403);
xnor U8330 (N_8330,N_5587,N_6543);
and U8331 (N_8331,N_5232,N_6657);
nor U8332 (N_8332,N_6824,N_6334);
nand U8333 (N_8333,N_6619,N_6081);
and U8334 (N_8334,N_7497,N_5303);
or U8335 (N_8335,N_7404,N_6620);
nor U8336 (N_8336,N_6829,N_7157);
nor U8337 (N_8337,N_7183,N_6425);
nand U8338 (N_8338,N_6847,N_6342);
nor U8339 (N_8339,N_6532,N_7156);
nand U8340 (N_8340,N_7446,N_5418);
or U8341 (N_8341,N_5540,N_6834);
nand U8342 (N_8342,N_5850,N_7193);
xnor U8343 (N_8343,N_6177,N_6148);
nor U8344 (N_8344,N_5624,N_6069);
nor U8345 (N_8345,N_6394,N_5526);
xnor U8346 (N_8346,N_6032,N_5372);
and U8347 (N_8347,N_5662,N_5311);
xor U8348 (N_8348,N_6638,N_7247);
and U8349 (N_8349,N_5637,N_7226);
xnor U8350 (N_8350,N_5833,N_5400);
and U8351 (N_8351,N_6016,N_7374);
and U8352 (N_8352,N_6682,N_7050);
nand U8353 (N_8353,N_7180,N_5184);
nor U8354 (N_8354,N_7248,N_7134);
xor U8355 (N_8355,N_5571,N_5776);
or U8356 (N_8356,N_6628,N_5227);
and U8357 (N_8357,N_5536,N_7448);
or U8358 (N_8358,N_6084,N_5077);
or U8359 (N_8359,N_6828,N_5865);
and U8360 (N_8360,N_6683,N_5889);
nor U8361 (N_8361,N_5737,N_5072);
and U8362 (N_8362,N_6355,N_6298);
nor U8363 (N_8363,N_5906,N_5519);
and U8364 (N_8364,N_6393,N_6132);
and U8365 (N_8365,N_5607,N_7337);
xor U8366 (N_8366,N_6904,N_5359);
nand U8367 (N_8367,N_5085,N_6215);
nor U8368 (N_8368,N_6485,N_7301);
xnor U8369 (N_8369,N_6222,N_5992);
xor U8370 (N_8370,N_6992,N_6825);
xor U8371 (N_8371,N_5708,N_7112);
xor U8372 (N_8372,N_7137,N_6920);
nand U8373 (N_8373,N_6811,N_6228);
xor U8374 (N_8374,N_5187,N_5468);
and U8375 (N_8375,N_6796,N_6991);
nand U8376 (N_8376,N_6554,N_7099);
nor U8377 (N_8377,N_7378,N_5959);
nand U8378 (N_8378,N_7163,N_5475);
or U8379 (N_8379,N_7351,N_6719);
nand U8380 (N_8380,N_6866,N_7477);
nor U8381 (N_8381,N_6770,N_7065);
nand U8382 (N_8382,N_6531,N_5834);
nor U8383 (N_8383,N_6492,N_7482);
xnor U8384 (N_8384,N_5713,N_5396);
and U8385 (N_8385,N_7106,N_6464);
or U8386 (N_8386,N_5159,N_6376);
and U8387 (N_8387,N_6052,N_6821);
xor U8388 (N_8388,N_6333,N_5218);
or U8389 (N_8389,N_5436,N_7239);
nor U8390 (N_8390,N_6566,N_7222);
xor U8391 (N_8391,N_5604,N_6774);
xnor U8392 (N_8392,N_5163,N_6880);
or U8393 (N_8393,N_5062,N_6720);
nor U8394 (N_8394,N_6560,N_6495);
nor U8395 (N_8395,N_5125,N_6233);
or U8396 (N_8396,N_5065,N_5851);
or U8397 (N_8397,N_5860,N_6234);
xnor U8398 (N_8398,N_6159,N_5773);
or U8399 (N_8399,N_5878,N_5650);
xnor U8400 (N_8400,N_6305,N_6444);
nand U8401 (N_8401,N_5291,N_6191);
nand U8402 (N_8402,N_7209,N_5795);
xnor U8403 (N_8403,N_7371,N_6335);
or U8404 (N_8404,N_7434,N_7060);
and U8405 (N_8405,N_5161,N_6271);
nand U8406 (N_8406,N_5390,N_5925);
and U8407 (N_8407,N_5429,N_5371);
xor U8408 (N_8408,N_5523,N_7311);
nor U8409 (N_8409,N_5798,N_6042);
nor U8410 (N_8410,N_6100,N_6263);
xnor U8411 (N_8411,N_5728,N_5832);
or U8412 (N_8412,N_6863,N_6756);
nor U8413 (N_8413,N_6561,N_6699);
nand U8414 (N_8414,N_7338,N_5137);
nand U8415 (N_8415,N_7031,N_6273);
nand U8416 (N_8416,N_5095,N_6654);
nand U8417 (N_8417,N_5466,N_6713);
nand U8418 (N_8418,N_7011,N_6396);
nand U8419 (N_8419,N_5207,N_5266);
xor U8420 (N_8420,N_6905,N_7475);
or U8421 (N_8421,N_7058,N_6343);
nand U8422 (N_8422,N_6736,N_5658);
and U8423 (N_8423,N_6917,N_6505);
or U8424 (N_8424,N_6558,N_6208);
and U8425 (N_8425,N_5393,N_5049);
nand U8426 (N_8426,N_6762,N_7097);
or U8427 (N_8427,N_6366,N_5768);
or U8428 (N_8428,N_5576,N_5749);
xnor U8429 (N_8429,N_6130,N_5141);
nand U8430 (N_8430,N_6356,N_6968);
or U8431 (N_8431,N_6729,N_6255);
or U8432 (N_8432,N_5934,N_7409);
or U8433 (N_8433,N_6927,N_5276);
xnor U8434 (N_8434,N_6664,N_5264);
or U8435 (N_8435,N_6062,N_7044);
nand U8436 (N_8436,N_5866,N_5905);
nor U8437 (N_8437,N_7101,N_5801);
nand U8438 (N_8438,N_6911,N_5706);
or U8439 (N_8439,N_5679,N_6046);
or U8440 (N_8440,N_7225,N_5900);
nor U8441 (N_8441,N_7326,N_5304);
nand U8442 (N_8442,N_5579,N_5245);
and U8443 (N_8443,N_6308,N_5488);
nand U8444 (N_8444,N_5827,N_5862);
xnor U8445 (N_8445,N_7425,N_5198);
nand U8446 (N_8446,N_6235,N_7122);
nor U8447 (N_8447,N_6958,N_5144);
nor U8448 (N_8448,N_7489,N_6357);
and U8449 (N_8449,N_6295,N_5909);
and U8450 (N_8450,N_6890,N_5879);
and U8451 (N_8451,N_7203,N_6965);
nor U8452 (N_8452,N_6771,N_5556);
nor U8453 (N_8453,N_6651,N_5510);
nor U8454 (N_8454,N_5676,N_6135);
and U8455 (N_8455,N_5319,N_7159);
nor U8456 (N_8456,N_5589,N_5268);
and U8457 (N_8457,N_5294,N_5758);
xnor U8458 (N_8458,N_5068,N_5431);
and U8459 (N_8459,N_6622,N_7040);
xnor U8460 (N_8460,N_5808,N_6987);
nor U8461 (N_8461,N_6672,N_7228);
and U8462 (N_8462,N_5480,N_5470);
nor U8463 (N_8463,N_6712,N_6070);
nand U8464 (N_8464,N_6264,N_6636);
or U8465 (N_8465,N_5283,N_6680);
nand U8466 (N_8466,N_6320,N_7266);
nand U8467 (N_8467,N_5259,N_6449);
or U8468 (N_8468,N_5403,N_6198);
xor U8469 (N_8469,N_6404,N_5039);
or U8470 (N_8470,N_6236,N_6726);
nor U8471 (N_8471,N_6797,N_5018);
nand U8472 (N_8472,N_6156,N_6369);
nor U8473 (N_8473,N_7260,N_5743);
nor U8474 (N_8474,N_6068,N_6990);
or U8475 (N_8475,N_6326,N_5615);
nand U8476 (N_8476,N_6458,N_5314);
nor U8477 (N_8477,N_5924,N_6061);
and U8478 (N_8478,N_5770,N_6611);
and U8479 (N_8479,N_7333,N_7334);
and U8480 (N_8480,N_5230,N_6980);
xnor U8481 (N_8481,N_6499,N_6819);
and U8482 (N_8482,N_5581,N_5603);
or U8483 (N_8483,N_5887,N_5487);
nor U8484 (N_8484,N_7462,N_6859);
xor U8485 (N_8485,N_5405,N_6938);
or U8486 (N_8486,N_5414,N_5178);
or U8487 (N_8487,N_7343,N_5186);
nand U8488 (N_8488,N_5381,N_6497);
and U8489 (N_8489,N_5103,N_6535);
nand U8490 (N_8490,N_7330,N_6724);
nor U8491 (N_8491,N_5428,N_7142);
xnor U8492 (N_8492,N_5534,N_5764);
and U8493 (N_8493,N_6094,N_6328);
xnor U8494 (N_8494,N_5486,N_5595);
or U8495 (N_8495,N_5516,N_7278);
xnor U8496 (N_8496,N_7086,N_5456);
and U8497 (N_8497,N_6946,N_6445);
and U8498 (N_8498,N_6420,N_6063);
nor U8499 (N_8499,N_6967,N_7411);
nor U8500 (N_8500,N_5521,N_7223);
and U8501 (N_8501,N_6626,N_5619);
and U8502 (N_8502,N_5613,N_6759);
xnor U8503 (N_8503,N_7102,N_6193);
nand U8504 (N_8504,N_5686,N_5235);
or U8505 (N_8505,N_7370,N_6047);
xor U8506 (N_8506,N_7212,N_5437);
nand U8507 (N_8507,N_6542,N_7072);
and U8508 (N_8508,N_5508,N_6435);
and U8509 (N_8509,N_6386,N_5327);
nand U8510 (N_8510,N_5270,N_5463);
and U8511 (N_8511,N_6769,N_5916);
nand U8512 (N_8512,N_7472,N_6221);
nand U8513 (N_8513,N_7022,N_7161);
xnor U8514 (N_8514,N_6474,N_6186);
or U8515 (N_8515,N_5756,N_6581);
xnor U8516 (N_8516,N_6303,N_6478);
nand U8517 (N_8517,N_6164,N_6368);
nor U8518 (N_8518,N_6364,N_6879);
xor U8519 (N_8519,N_5616,N_7121);
nand U8520 (N_8520,N_6044,N_6223);
or U8521 (N_8521,N_7025,N_5867);
nor U8522 (N_8522,N_5050,N_5012);
or U8523 (N_8523,N_6871,N_7422);
and U8524 (N_8524,N_5023,N_7290);
xnor U8525 (N_8525,N_6875,N_5061);
and U8526 (N_8526,N_5790,N_5088);
and U8527 (N_8527,N_6752,N_5048);
nand U8528 (N_8528,N_6618,N_6596);
xnor U8529 (N_8529,N_6104,N_5037);
nor U8530 (N_8530,N_7036,N_7231);
and U8531 (N_8531,N_6925,N_7480);
and U8532 (N_8532,N_7055,N_6703);
or U8533 (N_8533,N_6470,N_5172);
or U8534 (N_8534,N_5164,N_5336);
xnor U8535 (N_8535,N_5520,N_6763);
nor U8536 (N_8536,N_6407,N_5119);
and U8537 (N_8537,N_5442,N_7335);
and U8538 (N_8538,N_5138,N_5842);
xor U8539 (N_8539,N_7455,N_5040);
xnor U8540 (N_8540,N_7323,N_5958);
xnor U8541 (N_8541,N_6459,N_5621);
and U8542 (N_8542,N_7024,N_6277);
nand U8543 (N_8543,N_5664,N_5947);
nand U8544 (N_8544,N_5005,N_7265);
nor U8545 (N_8545,N_6166,N_5352);
and U8546 (N_8546,N_6075,N_5593);
or U8547 (N_8547,N_5213,N_5840);
nor U8548 (N_8548,N_5011,N_5171);
or U8549 (N_8549,N_7110,N_5721);
nand U8550 (N_8550,N_6203,N_5391);
xnor U8551 (N_8551,N_7208,N_7415);
nand U8552 (N_8552,N_5813,N_6128);
and U8553 (N_8553,N_6878,N_5705);
or U8554 (N_8554,N_6630,N_5094);
nor U8555 (N_8555,N_5351,N_6012);
nor U8556 (N_8556,N_6832,N_7493);
xor U8557 (N_8557,N_6360,N_6610);
nand U8558 (N_8558,N_6043,N_5113);
and U8559 (N_8559,N_6786,N_7001);
nor U8560 (N_8560,N_6817,N_7091);
xnor U8561 (N_8561,N_6316,N_7020);
xor U8562 (N_8562,N_6329,N_6816);
and U8563 (N_8563,N_6512,N_5190);
nand U8564 (N_8564,N_5262,N_5140);
nand U8565 (N_8565,N_7243,N_6498);
nor U8566 (N_8566,N_5594,N_6210);
and U8567 (N_8567,N_6297,N_5620);
xnor U8568 (N_8568,N_7033,N_5365);
or U8569 (N_8569,N_7190,N_7076);
xnor U8570 (N_8570,N_5333,N_5884);
xor U8571 (N_8571,N_5870,N_5527);
nand U8572 (N_8572,N_6650,N_6781);
xor U8573 (N_8573,N_7490,N_7135);
or U8574 (N_8574,N_6241,N_5830);
nor U8575 (N_8575,N_5056,N_7282);
nor U8576 (N_8576,N_6454,N_6338);
and U8577 (N_8577,N_6846,N_6805);
xnor U8578 (N_8578,N_6883,N_6810);
nor U8579 (N_8579,N_5188,N_5872);
nand U8580 (N_8580,N_5552,N_7291);
xor U8581 (N_8581,N_5783,N_6286);
and U8582 (N_8582,N_5785,N_5777);
or U8583 (N_8583,N_6034,N_5476);
xor U8584 (N_8584,N_6244,N_5194);
or U8585 (N_8585,N_7298,N_5891);
and U8586 (N_8586,N_5886,N_6433);
and U8587 (N_8587,N_5969,N_7070);
or U8588 (N_8588,N_6351,N_5980);
nor U8589 (N_8589,N_7238,N_6698);
nand U8590 (N_8590,N_5399,N_5839);
nand U8591 (N_8591,N_6020,N_6506);
or U8592 (N_8592,N_5271,N_7094);
xnor U8593 (N_8593,N_6943,N_6079);
nand U8594 (N_8594,N_5561,N_6969);
or U8595 (N_8595,N_5131,N_7253);
nand U8596 (N_8596,N_6789,N_6141);
nor U8597 (N_8597,N_5965,N_6679);
and U8598 (N_8598,N_6613,N_5923);
and U8599 (N_8599,N_7004,N_6585);
nor U8600 (N_8600,N_6661,N_6648);
xnor U8601 (N_8601,N_5951,N_7066);
nand U8602 (N_8602,N_5025,N_5544);
nand U8603 (N_8603,N_6108,N_6517);
xor U8604 (N_8604,N_5240,N_6972);
xnor U8605 (N_8605,N_6216,N_7474);
nor U8606 (N_8606,N_5720,N_5345);
and U8607 (N_8607,N_5383,N_6361);
nand U8608 (N_8608,N_6447,N_5191);
nand U8609 (N_8609,N_6278,N_7187);
nand U8610 (N_8610,N_5229,N_6845);
and U8611 (N_8611,N_5991,N_5744);
and U8612 (N_8612,N_6522,N_6226);
and U8613 (N_8613,N_5337,N_5289);
and U8614 (N_8614,N_5339,N_5609);
and U8615 (N_8615,N_7358,N_6095);
nor U8616 (N_8616,N_6460,N_6430);
nand U8617 (N_8617,N_6253,N_6964);
nor U8618 (N_8618,N_5702,N_5154);
nor U8619 (N_8619,N_6894,N_6692);
nor U8620 (N_8620,N_5091,N_7155);
and U8621 (N_8621,N_7059,N_6179);
nand U8622 (N_8622,N_7317,N_6530);
nand U8623 (N_8623,N_6744,N_5694);
and U8624 (N_8624,N_6747,N_6315);
or U8625 (N_8625,N_5366,N_7379);
xor U8626 (N_8626,N_7259,N_6120);
nand U8627 (N_8627,N_6674,N_6318);
xnor U8628 (N_8628,N_5591,N_5143);
nand U8629 (N_8629,N_5344,N_7410);
or U8630 (N_8630,N_6117,N_5682);
xnor U8631 (N_8631,N_5936,N_5249);
xnor U8632 (N_8632,N_5296,N_7437);
or U8633 (N_8633,N_5986,N_5324);
nor U8634 (N_8634,N_5215,N_5267);
or U8635 (N_8635,N_5331,N_7270);
xnor U8636 (N_8636,N_5462,N_6172);
nand U8637 (N_8637,N_6462,N_6382);
xnor U8638 (N_8638,N_5309,N_5847);
xnor U8639 (N_8639,N_5652,N_6155);
nand U8640 (N_8640,N_5722,N_6059);
xor U8641 (N_8641,N_5530,N_5122);
nand U8642 (N_8642,N_5559,N_7153);
and U8643 (N_8643,N_6118,N_6870);
nor U8644 (N_8644,N_5419,N_5755);
and U8645 (N_8645,N_7073,N_7491);
nand U8646 (N_8646,N_6529,N_5447);
and U8647 (N_8647,N_6065,N_7018);
or U8648 (N_8648,N_6149,N_5313);
nand U8649 (N_8649,N_5638,N_5246);
xor U8650 (N_8650,N_6730,N_5489);
and U8651 (N_8651,N_6496,N_5569);
nand U8652 (N_8652,N_6086,N_6802);
and U8653 (N_8653,N_5156,N_5295);
and U8654 (N_8654,N_6688,N_6733);
nor U8655 (N_8655,N_7176,N_6437);
and U8656 (N_8656,N_6390,N_6820);
nand U8657 (N_8657,N_6101,N_5401);
nor U8658 (N_8658,N_5430,N_7098);
nor U8659 (N_8659,N_6936,N_6701);
xor U8660 (N_8660,N_7423,N_7201);
xor U8661 (N_8661,N_5364,N_6194);
xnor U8662 (N_8662,N_6383,N_7306);
or U8663 (N_8663,N_5357,N_5454);
and U8664 (N_8664,N_5078,N_6402);
nand U8665 (N_8665,N_7276,N_7339);
nand U8666 (N_8666,N_7451,N_5075);
nor U8667 (N_8667,N_5646,N_5136);
nor U8668 (N_8668,N_7261,N_6168);
xor U8669 (N_8669,N_6710,N_5274);
or U8670 (N_8670,N_5966,N_5940);
nand U8671 (N_8671,N_5063,N_6655);
xor U8672 (N_8672,N_6948,N_5165);
or U8673 (N_8673,N_6536,N_5111);
or U8674 (N_8674,N_6192,N_5226);
xor U8675 (N_8675,N_7391,N_6288);
nor U8676 (N_8676,N_7313,N_5838);
or U8677 (N_8677,N_5693,N_5490);
nand U8678 (N_8678,N_5300,N_6232);
xnor U8679 (N_8679,N_5814,N_7150);
xnor U8680 (N_8680,N_6850,N_6373);
or U8681 (N_8681,N_6161,N_6695);
xnor U8682 (N_8682,N_7149,N_7056);
or U8683 (N_8683,N_5996,N_5903);
nand U8684 (N_8684,N_6687,N_5484);
xnor U8685 (N_8685,N_6983,N_6669);
nand U8686 (N_8686,N_5234,N_7038);
or U8687 (N_8687,N_7376,N_5931);
xnor U8688 (N_8688,N_5280,N_5824);
or U8689 (N_8689,N_5856,N_6311);
xor U8690 (N_8690,N_6534,N_5575);
and U8691 (N_8691,N_6327,N_6822);
xor U8692 (N_8692,N_7293,N_5828);
nor U8693 (N_8693,N_7398,N_7179);
and U8694 (N_8694,N_6857,N_6150);
nand U8695 (N_8695,N_6582,N_7447);
nand U8696 (N_8696,N_5752,N_5288);
or U8697 (N_8697,N_6384,N_6483);
and U8698 (N_8698,N_6668,N_7195);
nor U8699 (N_8699,N_7008,N_5882);
nor U8700 (N_8700,N_6146,N_5745);
nor U8701 (N_8701,N_7077,N_5019);
or U8702 (N_8702,N_7297,N_5677);
or U8703 (N_8703,N_7281,N_5512);
nor U8704 (N_8704,N_5574,N_5496);
nand U8705 (N_8705,N_6103,N_6833);
nand U8706 (N_8706,N_6422,N_7113);
nand U8707 (N_8707,N_5074,N_5185);
and U8708 (N_8708,N_6074,N_5668);
nor U8709 (N_8709,N_6107,N_6985);
and U8710 (N_8710,N_5751,N_6901);
nand U8711 (N_8711,N_5086,N_5928);
xor U8712 (N_8712,N_6855,N_6659);
nand U8713 (N_8713,N_5780,N_6395);
nor U8714 (N_8714,N_5599,N_7000);
nor U8715 (N_8715,N_5166,N_7188);
nor U8716 (N_8716,N_7164,N_7361);
nand U8717 (N_8717,N_6145,N_6988);
and U8718 (N_8718,N_6243,N_5880);
nor U8719 (N_8719,N_6114,N_6479);
and U8720 (N_8720,N_7280,N_6362);
nand U8721 (N_8721,N_6751,N_7015);
xor U8722 (N_8722,N_6935,N_6229);
nand U8723 (N_8723,N_7464,N_6323);
and U8724 (N_8724,N_6632,N_6220);
nor U8725 (N_8725,N_5317,N_5568);
xor U8726 (N_8726,N_5472,N_7027);
xnor U8727 (N_8727,N_5690,N_5495);
nor U8728 (N_8728,N_6574,N_6170);
and U8729 (N_8729,N_5377,N_6399);
or U8730 (N_8730,N_7046,N_5395);
nor U8731 (N_8731,N_6760,N_5340);
or U8732 (N_8732,N_6397,N_5943);
or U8733 (N_8733,N_6280,N_5953);
nor U8734 (N_8734,N_7003,N_5503);
xor U8735 (N_8735,N_7039,N_5179);
xnor U8736 (N_8736,N_5636,N_6293);
nor U8737 (N_8737,N_6567,N_5033);
or U8738 (N_8738,N_5248,N_5358);
nand U8739 (N_8739,N_7152,N_6615);
and U8740 (N_8740,N_7394,N_6858);
nand U8741 (N_8741,N_7452,N_7318);
nor U8742 (N_8742,N_6800,N_7407);
or U8743 (N_8743,N_5946,N_5729);
nand U8744 (N_8744,N_7251,N_6673);
nand U8745 (N_8745,N_5660,N_6023);
xnor U8746 (N_8746,N_6440,N_6516);
nand U8747 (N_8747,N_6932,N_7442);
and U8748 (N_8748,N_6999,N_5060);
and U8749 (N_8749,N_5899,N_5626);
and U8750 (N_8750,N_7279,N_5342);
or U8751 (N_8751,N_7483,N_6395);
nand U8752 (N_8752,N_5493,N_6130);
or U8753 (N_8753,N_5918,N_7013);
nor U8754 (N_8754,N_5820,N_7392);
nor U8755 (N_8755,N_6008,N_7357);
xor U8756 (N_8756,N_6969,N_5690);
nor U8757 (N_8757,N_5739,N_5616);
xnor U8758 (N_8758,N_5853,N_6324);
xor U8759 (N_8759,N_6059,N_7421);
or U8760 (N_8760,N_7337,N_5658);
or U8761 (N_8761,N_6571,N_5054);
nand U8762 (N_8762,N_7418,N_5684);
nor U8763 (N_8763,N_7037,N_6692);
nand U8764 (N_8764,N_5628,N_6553);
or U8765 (N_8765,N_5771,N_5512);
nand U8766 (N_8766,N_7071,N_5413);
and U8767 (N_8767,N_5176,N_6901);
or U8768 (N_8768,N_6790,N_5048);
and U8769 (N_8769,N_6339,N_5931);
and U8770 (N_8770,N_5107,N_5178);
or U8771 (N_8771,N_5022,N_5784);
nor U8772 (N_8772,N_5630,N_5526);
and U8773 (N_8773,N_5105,N_5842);
nand U8774 (N_8774,N_6929,N_7290);
xor U8775 (N_8775,N_5485,N_6198);
nor U8776 (N_8776,N_7427,N_7098);
or U8777 (N_8777,N_6259,N_6780);
or U8778 (N_8778,N_6357,N_6249);
xor U8779 (N_8779,N_6629,N_6164);
nand U8780 (N_8780,N_5722,N_5349);
and U8781 (N_8781,N_5261,N_6150);
xnor U8782 (N_8782,N_6716,N_6754);
xnor U8783 (N_8783,N_6091,N_6456);
and U8784 (N_8784,N_5802,N_5943);
or U8785 (N_8785,N_5711,N_6540);
and U8786 (N_8786,N_6736,N_7493);
nand U8787 (N_8787,N_7059,N_7054);
nor U8788 (N_8788,N_5714,N_5737);
nor U8789 (N_8789,N_5464,N_6321);
or U8790 (N_8790,N_6196,N_5694);
xnor U8791 (N_8791,N_6712,N_5403);
and U8792 (N_8792,N_6619,N_6318);
and U8793 (N_8793,N_5041,N_7191);
nand U8794 (N_8794,N_6429,N_5120);
xnor U8795 (N_8795,N_5665,N_5045);
or U8796 (N_8796,N_6442,N_7052);
and U8797 (N_8797,N_6284,N_6411);
nor U8798 (N_8798,N_7241,N_6237);
and U8799 (N_8799,N_7390,N_6340);
or U8800 (N_8800,N_5856,N_6524);
or U8801 (N_8801,N_5881,N_6196);
nand U8802 (N_8802,N_5230,N_6794);
or U8803 (N_8803,N_5246,N_6065);
nor U8804 (N_8804,N_6470,N_5180);
nand U8805 (N_8805,N_5557,N_5519);
nand U8806 (N_8806,N_6841,N_5118);
or U8807 (N_8807,N_6129,N_5905);
xnor U8808 (N_8808,N_5700,N_6252);
and U8809 (N_8809,N_6249,N_6290);
xor U8810 (N_8810,N_7350,N_6622);
and U8811 (N_8811,N_6315,N_6742);
or U8812 (N_8812,N_6763,N_5284);
nand U8813 (N_8813,N_6193,N_5249);
or U8814 (N_8814,N_5021,N_5436);
nor U8815 (N_8815,N_7418,N_6331);
nor U8816 (N_8816,N_6522,N_6799);
nor U8817 (N_8817,N_7425,N_5398);
nor U8818 (N_8818,N_6254,N_6753);
nand U8819 (N_8819,N_6271,N_6953);
nand U8820 (N_8820,N_6688,N_5423);
nor U8821 (N_8821,N_5920,N_7262);
and U8822 (N_8822,N_5041,N_6872);
nand U8823 (N_8823,N_5053,N_6351);
or U8824 (N_8824,N_7103,N_5693);
xor U8825 (N_8825,N_6068,N_7331);
nor U8826 (N_8826,N_5486,N_7343);
or U8827 (N_8827,N_5027,N_7380);
nand U8828 (N_8828,N_5781,N_5129);
xnor U8829 (N_8829,N_6012,N_6371);
nor U8830 (N_8830,N_7257,N_7403);
or U8831 (N_8831,N_5450,N_7459);
nand U8832 (N_8832,N_6829,N_6756);
nor U8833 (N_8833,N_5935,N_5852);
xnor U8834 (N_8834,N_6569,N_5732);
and U8835 (N_8835,N_6056,N_7397);
or U8836 (N_8836,N_7372,N_5786);
or U8837 (N_8837,N_7026,N_5176);
and U8838 (N_8838,N_5247,N_7479);
nor U8839 (N_8839,N_5371,N_5792);
and U8840 (N_8840,N_5175,N_6183);
nor U8841 (N_8841,N_5133,N_5597);
nand U8842 (N_8842,N_5981,N_6028);
nand U8843 (N_8843,N_5541,N_5326);
and U8844 (N_8844,N_5438,N_7247);
and U8845 (N_8845,N_7378,N_5654);
nor U8846 (N_8846,N_5685,N_6352);
xnor U8847 (N_8847,N_7474,N_5580);
and U8848 (N_8848,N_7164,N_7431);
nand U8849 (N_8849,N_5648,N_5416);
nor U8850 (N_8850,N_6227,N_6647);
and U8851 (N_8851,N_7458,N_6080);
xnor U8852 (N_8852,N_6838,N_6065);
nand U8853 (N_8853,N_7172,N_6850);
nand U8854 (N_8854,N_6120,N_6060);
and U8855 (N_8855,N_6976,N_5781);
nand U8856 (N_8856,N_5190,N_6063);
and U8857 (N_8857,N_5840,N_6671);
xnor U8858 (N_8858,N_6184,N_7316);
or U8859 (N_8859,N_6426,N_5732);
and U8860 (N_8860,N_5256,N_6827);
or U8861 (N_8861,N_7272,N_7044);
and U8862 (N_8862,N_6060,N_6555);
nor U8863 (N_8863,N_6622,N_6303);
nor U8864 (N_8864,N_6957,N_6290);
nand U8865 (N_8865,N_5292,N_6903);
nand U8866 (N_8866,N_7003,N_5249);
xnor U8867 (N_8867,N_7317,N_7214);
xnor U8868 (N_8868,N_7160,N_5295);
and U8869 (N_8869,N_6020,N_5672);
and U8870 (N_8870,N_6153,N_7288);
and U8871 (N_8871,N_6909,N_7221);
xor U8872 (N_8872,N_6496,N_6792);
nand U8873 (N_8873,N_6635,N_5735);
xnor U8874 (N_8874,N_7060,N_6765);
nand U8875 (N_8875,N_7218,N_6269);
xnor U8876 (N_8876,N_6932,N_5489);
nand U8877 (N_8877,N_6849,N_7208);
and U8878 (N_8878,N_6043,N_5448);
and U8879 (N_8879,N_6304,N_6063);
and U8880 (N_8880,N_6860,N_6487);
or U8881 (N_8881,N_5808,N_6720);
xnor U8882 (N_8882,N_7363,N_6848);
nand U8883 (N_8883,N_5749,N_6143);
nor U8884 (N_8884,N_7092,N_5512);
xnor U8885 (N_8885,N_6785,N_5197);
or U8886 (N_8886,N_7016,N_5967);
nand U8887 (N_8887,N_6464,N_6107);
and U8888 (N_8888,N_7113,N_6545);
nand U8889 (N_8889,N_7494,N_5024);
and U8890 (N_8890,N_7306,N_5735);
and U8891 (N_8891,N_6653,N_7071);
and U8892 (N_8892,N_5105,N_6791);
nor U8893 (N_8893,N_6152,N_7234);
xor U8894 (N_8894,N_6006,N_5486);
or U8895 (N_8895,N_5651,N_5281);
nor U8896 (N_8896,N_5229,N_5496);
xor U8897 (N_8897,N_6511,N_6487);
nor U8898 (N_8898,N_7240,N_7297);
nand U8899 (N_8899,N_5181,N_5312);
xor U8900 (N_8900,N_7241,N_5800);
and U8901 (N_8901,N_7408,N_6582);
or U8902 (N_8902,N_7032,N_6219);
and U8903 (N_8903,N_7266,N_5801);
nand U8904 (N_8904,N_5963,N_5085);
nand U8905 (N_8905,N_6606,N_5091);
xor U8906 (N_8906,N_6546,N_6179);
nor U8907 (N_8907,N_7418,N_5063);
xnor U8908 (N_8908,N_5658,N_6524);
nand U8909 (N_8909,N_5868,N_6622);
nor U8910 (N_8910,N_5601,N_7279);
nand U8911 (N_8911,N_6099,N_5219);
or U8912 (N_8912,N_6432,N_5838);
or U8913 (N_8913,N_5962,N_7239);
nor U8914 (N_8914,N_5703,N_6913);
and U8915 (N_8915,N_6153,N_7266);
or U8916 (N_8916,N_5189,N_7365);
and U8917 (N_8917,N_5629,N_5835);
nor U8918 (N_8918,N_6661,N_5533);
or U8919 (N_8919,N_5103,N_6710);
or U8920 (N_8920,N_6756,N_6923);
and U8921 (N_8921,N_5471,N_5127);
nor U8922 (N_8922,N_7083,N_5081);
nand U8923 (N_8923,N_6811,N_5931);
xnor U8924 (N_8924,N_6475,N_5291);
or U8925 (N_8925,N_5716,N_5699);
xnor U8926 (N_8926,N_5500,N_5533);
xnor U8927 (N_8927,N_6787,N_6623);
xor U8928 (N_8928,N_7453,N_6672);
or U8929 (N_8929,N_6133,N_7419);
or U8930 (N_8930,N_5374,N_5731);
nand U8931 (N_8931,N_5794,N_5525);
or U8932 (N_8932,N_7316,N_6867);
nor U8933 (N_8933,N_6975,N_7040);
nand U8934 (N_8934,N_6570,N_5957);
nand U8935 (N_8935,N_5776,N_5499);
and U8936 (N_8936,N_5112,N_6381);
nand U8937 (N_8937,N_6987,N_6805);
nand U8938 (N_8938,N_6862,N_5217);
and U8939 (N_8939,N_6575,N_6693);
or U8940 (N_8940,N_6059,N_5949);
xor U8941 (N_8941,N_6066,N_6454);
and U8942 (N_8942,N_5473,N_5094);
or U8943 (N_8943,N_5665,N_5915);
xor U8944 (N_8944,N_5175,N_6000);
xnor U8945 (N_8945,N_5255,N_6974);
nand U8946 (N_8946,N_5991,N_6094);
and U8947 (N_8947,N_5401,N_7092);
and U8948 (N_8948,N_5967,N_5093);
nand U8949 (N_8949,N_6664,N_7432);
nand U8950 (N_8950,N_7113,N_5831);
nor U8951 (N_8951,N_6951,N_5289);
and U8952 (N_8952,N_6077,N_7491);
xnor U8953 (N_8953,N_5896,N_5916);
xnor U8954 (N_8954,N_5956,N_6297);
nor U8955 (N_8955,N_6676,N_6117);
nor U8956 (N_8956,N_6701,N_5544);
or U8957 (N_8957,N_5482,N_7363);
nor U8958 (N_8958,N_7301,N_7380);
nand U8959 (N_8959,N_5658,N_7228);
or U8960 (N_8960,N_7253,N_7133);
nor U8961 (N_8961,N_6920,N_7395);
nor U8962 (N_8962,N_6411,N_5897);
xnor U8963 (N_8963,N_5997,N_7113);
and U8964 (N_8964,N_6300,N_6997);
and U8965 (N_8965,N_7286,N_5669);
nor U8966 (N_8966,N_6994,N_5733);
nor U8967 (N_8967,N_6892,N_7365);
nand U8968 (N_8968,N_7222,N_7228);
or U8969 (N_8969,N_6783,N_6576);
and U8970 (N_8970,N_5353,N_6110);
xor U8971 (N_8971,N_5465,N_5843);
nor U8972 (N_8972,N_6921,N_6634);
and U8973 (N_8973,N_5241,N_5091);
xor U8974 (N_8974,N_6085,N_5977);
and U8975 (N_8975,N_5426,N_6037);
xnor U8976 (N_8976,N_5449,N_6863);
nor U8977 (N_8977,N_5939,N_5148);
or U8978 (N_8978,N_7458,N_5761);
nand U8979 (N_8979,N_5950,N_6673);
xnor U8980 (N_8980,N_7418,N_5415);
or U8981 (N_8981,N_7400,N_6626);
xnor U8982 (N_8982,N_5038,N_7391);
nor U8983 (N_8983,N_5209,N_7102);
and U8984 (N_8984,N_7117,N_6740);
or U8985 (N_8985,N_6867,N_7052);
nor U8986 (N_8986,N_7373,N_6014);
nor U8987 (N_8987,N_5456,N_5446);
and U8988 (N_8988,N_5489,N_5527);
nor U8989 (N_8989,N_7333,N_6209);
and U8990 (N_8990,N_6492,N_7110);
and U8991 (N_8991,N_5453,N_6577);
or U8992 (N_8992,N_5664,N_6034);
nor U8993 (N_8993,N_6245,N_5097);
nand U8994 (N_8994,N_5256,N_7383);
and U8995 (N_8995,N_7169,N_6705);
xnor U8996 (N_8996,N_6375,N_5522);
xnor U8997 (N_8997,N_6361,N_6201);
nand U8998 (N_8998,N_5374,N_6116);
xnor U8999 (N_8999,N_5446,N_5465);
nor U9000 (N_9000,N_5225,N_7409);
xnor U9001 (N_9001,N_5603,N_5124);
nor U9002 (N_9002,N_7099,N_6771);
or U9003 (N_9003,N_6110,N_7443);
and U9004 (N_9004,N_5577,N_5859);
or U9005 (N_9005,N_5621,N_6599);
or U9006 (N_9006,N_5582,N_5775);
and U9007 (N_9007,N_7073,N_5578);
or U9008 (N_9008,N_5103,N_6382);
nor U9009 (N_9009,N_6559,N_6788);
and U9010 (N_9010,N_7283,N_6076);
and U9011 (N_9011,N_5102,N_5181);
nor U9012 (N_9012,N_6261,N_5728);
nor U9013 (N_9013,N_6241,N_6637);
and U9014 (N_9014,N_6665,N_6209);
and U9015 (N_9015,N_6816,N_6984);
nand U9016 (N_9016,N_6038,N_6789);
nand U9017 (N_9017,N_7325,N_5179);
xor U9018 (N_9018,N_7049,N_5797);
and U9019 (N_9019,N_5766,N_6762);
xor U9020 (N_9020,N_7154,N_5194);
or U9021 (N_9021,N_5109,N_6431);
or U9022 (N_9022,N_5398,N_6918);
xor U9023 (N_9023,N_6848,N_5225);
nor U9024 (N_9024,N_5965,N_7208);
nand U9025 (N_9025,N_6495,N_6930);
and U9026 (N_9026,N_6551,N_7335);
nor U9027 (N_9027,N_5987,N_6615);
nor U9028 (N_9028,N_7069,N_6832);
nor U9029 (N_9029,N_5222,N_6368);
and U9030 (N_9030,N_5277,N_6981);
or U9031 (N_9031,N_5143,N_6049);
or U9032 (N_9032,N_5144,N_6387);
or U9033 (N_9033,N_5414,N_6014);
and U9034 (N_9034,N_7250,N_6513);
nor U9035 (N_9035,N_6978,N_7431);
nor U9036 (N_9036,N_6628,N_5704);
and U9037 (N_9037,N_5495,N_5766);
nor U9038 (N_9038,N_7045,N_7131);
nor U9039 (N_9039,N_6718,N_5295);
nand U9040 (N_9040,N_7142,N_5394);
nand U9041 (N_9041,N_7390,N_6215);
nor U9042 (N_9042,N_6470,N_5615);
nor U9043 (N_9043,N_5073,N_7072);
nor U9044 (N_9044,N_5658,N_6941);
and U9045 (N_9045,N_6876,N_6745);
or U9046 (N_9046,N_5163,N_6854);
nand U9047 (N_9047,N_6366,N_5778);
xor U9048 (N_9048,N_5085,N_6376);
nand U9049 (N_9049,N_6172,N_5108);
xor U9050 (N_9050,N_5866,N_5302);
nor U9051 (N_9051,N_7155,N_6010);
xnor U9052 (N_9052,N_6125,N_5132);
or U9053 (N_9053,N_7419,N_7278);
nand U9054 (N_9054,N_6965,N_5008);
nand U9055 (N_9055,N_6846,N_5822);
and U9056 (N_9056,N_5711,N_5544);
nor U9057 (N_9057,N_6151,N_6019);
and U9058 (N_9058,N_5483,N_6884);
and U9059 (N_9059,N_6596,N_6722);
xor U9060 (N_9060,N_5056,N_6762);
nor U9061 (N_9061,N_5359,N_6684);
xor U9062 (N_9062,N_5606,N_6031);
and U9063 (N_9063,N_6884,N_5027);
xnor U9064 (N_9064,N_6285,N_6227);
nand U9065 (N_9065,N_7035,N_5809);
and U9066 (N_9066,N_6955,N_7487);
nand U9067 (N_9067,N_6376,N_5185);
nand U9068 (N_9068,N_5267,N_7082);
nor U9069 (N_9069,N_5118,N_5739);
nand U9070 (N_9070,N_5735,N_6127);
nor U9071 (N_9071,N_6216,N_7336);
or U9072 (N_9072,N_6189,N_7060);
nor U9073 (N_9073,N_6555,N_6855);
or U9074 (N_9074,N_6062,N_5795);
xnor U9075 (N_9075,N_6100,N_5158);
or U9076 (N_9076,N_5060,N_5572);
xor U9077 (N_9077,N_6794,N_6189);
or U9078 (N_9078,N_5116,N_6970);
or U9079 (N_9079,N_7008,N_5278);
and U9080 (N_9080,N_6778,N_5331);
xor U9081 (N_9081,N_6413,N_6708);
xor U9082 (N_9082,N_7444,N_6609);
or U9083 (N_9083,N_6281,N_6333);
xnor U9084 (N_9084,N_5308,N_7269);
xnor U9085 (N_9085,N_7263,N_5153);
xor U9086 (N_9086,N_6699,N_5910);
xnor U9087 (N_9087,N_7122,N_6338);
or U9088 (N_9088,N_6950,N_6665);
nand U9089 (N_9089,N_7454,N_6904);
nor U9090 (N_9090,N_5674,N_6222);
and U9091 (N_9091,N_5011,N_5378);
xor U9092 (N_9092,N_6108,N_5883);
and U9093 (N_9093,N_5388,N_6854);
nor U9094 (N_9094,N_5192,N_6231);
nor U9095 (N_9095,N_6096,N_6979);
or U9096 (N_9096,N_5674,N_6932);
xor U9097 (N_9097,N_6606,N_6020);
nand U9098 (N_9098,N_6100,N_6565);
nor U9099 (N_9099,N_6837,N_5494);
nor U9100 (N_9100,N_5032,N_5658);
and U9101 (N_9101,N_6883,N_5387);
nand U9102 (N_9102,N_5154,N_5727);
nand U9103 (N_9103,N_5953,N_6232);
nor U9104 (N_9104,N_6898,N_7037);
nand U9105 (N_9105,N_7484,N_6966);
nand U9106 (N_9106,N_6775,N_6939);
or U9107 (N_9107,N_6539,N_5495);
xnor U9108 (N_9108,N_7086,N_7037);
or U9109 (N_9109,N_5470,N_6547);
nand U9110 (N_9110,N_5489,N_7044);
nand U9111 (N_9111,N_6022,N_7250);
and U9112 (N_9112,N_6182,N_6927);
or U9113 (N_9113,N_7242,N_6120);
or U9114 (N_9114,N_6974,N_7430);
xnor U9115 (N_9115,N_5671,N_5274);
xnor U9116 (N_9116,N_7357,N_7438);
and U9117 (N_9117,N_5684,N_7194);
xnor U9118 (N_9118,N_7480,N_7199);
xnor U9119 (N_9119,N_6500,N_5211);
nor U9120 (N_9120,N_7059,N_7044);
and U9121 (N_9121,N_6337,N_6752);
or U9122 (N_9122,N_5628,N_6993);
or U9123 (N_9123,N_5164,N_6534);
and U9124 (N_9124,N_5226,N_6568);
and U9125 (N_9125,N_7396,N_5640);
nor U9126 (N_9126,N_6683,N_6097);
and U9127 (N_9127,N_5887,N_6521);
nand U9128 (N_9128,N_5524,N_5948);
xnor U9129 (N_9129,N_5826,N_5910);
xnor U9130 (N_9130,N_5405,N_6414);
and U9131 (N_9131,N_5880,N_6630);
or U9132 (N_9132,N_6407,N_6251);
xor U9133 (N_9133,N_6148,N_5568);
or U9134 (N_9134,N_5751,N_6111);
or U9135 (N_9135,N_6569,N_6116);
nor U9136 (N_9136,N_6756,N_5920);
xor U9137 (N_9137,N_5372,N_6704);
nand U9138 (N_9138,N_7297,N_5887);
nor U9139 (N_9139,N_7069,N_6548);
nand U9140 (N_9140,N_6718,N_7059);
nand U9141 (N_9141,N_5735,N_5836);
nor U9142 (N_9142,N_6705,N_6479);
nor U9143 (N_9143,N_5784,N_5858);
xor U9144 (N_9144,N_5387,N_7293);
xor U9145 (N_9145,N_6536,N_5065);
xnor U9146 (N_9146,N_6214,N_7134);
or U9147 (N_9147,N_5720,N_6297);
nand U9148 (N_9148,N_6105,N_6745);
xor U9149 (N_9149,N_7005,N_5984);
and U9150 (N_9150,N_6501,N_7159);
xnor U9151 (N_9151,N_5822,N_6483);
xnor U9152 (N_9152,N_6445,N_5857);
nor U9153 (N_9153,N_6126,N_6792);
and U9154 (N_9154,N_5089,N_6478);
nor U9155 (N_9155,N_5152,N_7018);
nor U9156 (N_9156,N_5599,N_7347);
nor U9157 (N_9157,N_5361,N_6841);
and U9158 (N_9158,N_6321,N_6634);
or U9159 (N_9159,N_7227,N_7392);
xor U9160 (N_9160,N_6867,N_5542);
xor U9161 (N_9161,N_6273,N_6894);
xor U9162 (N_9162,N_7261,N_6156);
nor U9163 (N_9163,N_5876,N_6081);
and U9164 (N_9164,N_6723,N_6257);
and U9165 (N_9165,N_5870,N_6143);
nor U9166 (N_9166,N_6564,N_6180);
or U9167 (N_9167,N_6616,N_6344);
xor U9168 (N_9168,N_5973,N_6566);
and U9169 (N_9169,N_5300,N_6170);
xor U9170 (N_9170,N_6508,N_5443);
nand U9171 (N_9171,N_6117,N_6957);
nor U9172 (N_9172,N_7244,N_6871);
nand U9173 (N_9173,N_6607,N_5414);
nor U9174 (N_9174,N_6272,N_6689);
or U9175 (N_9175,N_5644,N_5433);
or U9176 (N_9176,N_6840,N_5956);
or U9177 (N_9177,N_5555,N_5193);
and U9178 (N_9178,N_5474,N_5882);
and U9179 (N_9179,N_6430,N_5193);
or U9180 (N_9180,N_6962,N_6360);
and U9181 (N_9181,N_7335,N_5729);
nor U9182 (N_9182,N_6389,N_6331);
nor U9183 (N_9183,N_6527,N_6128);
or U9184 (N_9184,N_6024,N_6094);
xor U9185 (N_9185,N_6143,N_7367);
or U9186 (N_9186,N_5081,N_5874);
nor U9187 (N_9187,N_6443,N_5648);
or U9188 (N_9188,N_5191,N_5017);
nor U9189 (N_9189,N_6616,N_6812);
and U9190 (N_9190,N_5420,N_6966);
and U9191 (N_9191,N_5599,N_6107);
and U9192 (N_9192,N_6204,N_5818);
xnor U9193 (N_9193,N_6980,N_6855);
or U9194 (N_9194,N_5644,N_6940);
nor U9195 (N_9195,N_7134,N_7060);
nand U9196 (N_9196,N_6850,N_7482);
nand U9197 (N_9197,N_5756,N_6413);
and U9198 (N_9198,N_5013,N_6520);
or U9199 (N_9199,N_5910,N_6797);
nand U9200 (N_9200,N_7328,N_6359);
and U9201 (N_9201,N_5739,N_5982);
nor U9202 (N_9202,N_6939,N_6845);
or U9203 (N_9203,N_5889,N_7356);
and U9204 (N_9204,N_5441,N_7202);
nand U9205 (N_9205,N_7067,N_5960);
or U9206 (N_9206,N_6904,N_5191);
nand U9207 (N_9207,N_5360,N_5908);
nand U9208 (N_9208,N_5721,N_7077);
and U9209 (N_9209,N_6650,N_7320);
or U9210 (N_9210,N_5784,N_5744);
and U9211 (N_9211,N_7335,N_5523);
xnor U9212 (N_9212,N_5475,N_6910);
nor U9213 (N_9213,N_5462,N_6766);
xor U9214 (N_9214,N_6546,N_7044);
and U9215 (N_9215,N_6576,N_6085);
or U9216 (N_9216,N_6146,N_6360);
xnor U9217 (N_9217,N_6844,N_7455);
or U9218 (N_9218,N_6957,N_6433);
xnor U9219 (N_9219,N_5653,N_6816);
and U9220 (N_9220,N_6942,N_6027);
xor U9221 (N_9221,N_5458,N_6269);
and U9222 (N_9222,N_6055,N_6470);
nand U9223 (N_9223,N_6711,N_5549);
nand U9224 (N_9224,N_6954,N_6183);
xnor U9225 (N_9225,N_7307,N_6715);
and U9226 (N_9226,N_5054,N_6580);
or U9227 (N_9227,N_5000,N_7229);
xor U9228 (N_9228,N_6766,N_6528);
xor U9229 (N_9229,N_6275,N_6907);
and U9230 (N_9230,N_6236,N_6648);
nor U9231 (N_9231,N_6386,N_6012);
nand U9232 (N_9232,N_6393,N_5081);
nand U9233 (N_9233,N_6444,N_6666);
nand U9234 (N_9234,N_6768,N_6348);
or U9235 (N_9235,N_6388,N_6161);
xnor U9236 (N_9236,N_5845,N_5837);
nand U9237 (N_9237,N_7013,N_7370);
or U9238 (N_9238,N_5662,N_6073);
xnor U9239 (N_9239,N_5175,N_7324);
nor U9240 (N_9240,N_6496,N_6666);
or U9241 (N_9241,N_5151,N_5647);
xnor U9242 (N_9242,N_5640,N_6022);
nor U9243 (N_9243,N_6824,N_5385);
or U9244 (N_9244,N_5209,N_5784);
or U9245 (N_9245,N_5307,N_6564);
nor U9246 (N_9246,N_6162,N_5365);
xnor U9247 (N_9247,N_5035,N_6636);
nor U9248 (N_9248,N_5226,N_5572);
nand U9249 (N_9249,N_7462,N_6434);
xnor U9250 (N_9250,N_5488,N_7367);
xor U9251 (N_9251,N_7239,N_7338);
or U9252 (N_9252,N_7358,N_7090);
or U9253 (N_9253,N_6101,N_7034);
nor U9254 (N_9254,N_7185,N_7385);
nand U9255 (N_9255,N_6402,N_5517);
nor U9256 (N_9256,N_5521,N_6095);
nor U9257 (N_9257,N_5448,N_5930);
or U9258 (N_9258,N_5047,N_5945);
nor U9259 (N_9259,N_7327,N_5873);
xor U9260 (N_9260,N_6076,N_6615);
and U9261 (N_9261,N_6589,N_6368);
or U9262 (N_9262,N_5283,N_6362);
and U9263 (N_9263,N_5319,N_5963);
nor U9264 (N_9264,N_6510,N_5258);
and U9265 (N_9265,N_5174,N_6324);
or U9266 (N_9266,N_7479,N_6576);
nor U9267 (N_9267,N_5438,N_7252);
and U9268 (N_9268,N_5142,N_6638);
nor U9269 (N_9269,N_7400,N_5575);
nand U9270 (N_9270,N_6601,N_7450);
or U9271 (N_9271,N_5676,N_6907);
or U9272 (N_9272,N_7191,N_6391);
xor U9273 (N_9273,N_5679,N_7311);
xnor U9274 (N_9274,N_5886,N_7037);
or U9275 (N_9275,N_6742,N_6836);
xnor U9276 (N_9276,N_6814,N_6459);
nand U9277 (N_9277,N_6486,N_5235);
and U9278 (N_9278,N_7237,N_5914);
and U9279 (N_9279,N_7311,N_7131);
xnor U9280 (N_9280,N_6456,N_5203);
nor U9281 (N_9281,N_6946,N_5915);
or U9282 (N_9282,N_6891,N_6161);
xor U9283 (N_9283,N_6516,N_6169);
xnor U9284 (N_9284,N_7030,N_7036);
xor U9285 (N_9285,N_5740,N_5366);
nand U9286 (N_9286,N_5884,N_5120);
nand U9287 (N_9287,N_5241,N_5259);
xor U9288 (N_9288,N_6459,N_5900);
and U9289 (N_9289,N_6055,N_7069);
nand U9290 (N_9290,N_6302,N_6224);
xor U9291 (N_9291,N_6881,N_7487);
nor U9292 (N_9292,N_5167,N_5481);
xor U9293 (N_9293,N_5745,N_5148);
or U9294 (N_9294,N_5464,N_7029);
xnor U9295 (N_9295,N_6672,N_6352);
xnor U9296 (N_9296,N_6522,N_5671);
xor U9297 (N_9297,N_5093,N_7312);
and U9298 (N_9298,N_5999,N_6657);
and U9299 (N_9299,N_7072,N_5130);
nand U9300 (N_9300,N_5949,N_5050);
nand U9301 (N_9301,N_7194,N_6648);
nand U9302 (N_9302,N_5222,N_5930);
xor U9303 (N_9303,N_5105,N_5188);
nor U9304 (N_9304,N_5445,N_6100);
nand U9305 (N_9305,N_5670,N_6842);
xor U9306 (N_9306,N_7178,N_6310);
and U9307 (N_9307,N_5408,N_6727);
and U9308 (N_9308,N_7235,N_5370);
xor U9309 (N_9309,N_6339,N_6047);
nand U9310 (N_9310,N_6818,N_5767);
nand U9311 (N_9311,N_6269,N_5097);
nor U9312 (N_9312,N_5107,N_5540);
or U9313 (N_9313,N_7113,N_5315);
nand U9314 (N_9314,N_7176,N_5211);
nor U9315 (N_9315,N_7089,N_5354);
xor U9316 (N_9316,N_6169,N_7460);
xor U9317 (N_9317,N_6107,N_7016);
nand U9318 (N_9318,N_5485,N_6575);
and U9319 (N_9319,N_5828,N_6908);
nor U9320 (N_9320,N_5563,N_7103);
xnor U9321 (N_9321,N_5209,N_5822);
and U9322 (N_9322,N_7335,N_6743);
xnor U9323 (N_9323,N_5723,N_6769);
xor U9324 (N_9324,N_5453,N_6324);
or U9325 (N_9325,N_5504,N_5195);
nand U9326 (N_9326,N_6212,N_6236);
or U9327 (N_9327,N_5999,N_6501);
xor U9328 (N_9328,N_5924,N_6008);
or U9329 (N_9329,N_7333,N_5381);
or U9330 (N_9330,N_6788,N_5921);
and U9331 (N_9331,N_7171,N_5896);
nor U9332 (N_9332,N_7219,N_5744);
xnor U9333 (N_9333,N_5599,N_7257);
or U9334 (N_9334,N_5297,N_6071);
nor U9335 (N_9335,N_5751,N_7370);
or U9336 (N_9336,N_7251,N_5932);
nand U9337 (N_9337,N_7298,N_6691);
and U9338 (N_9338,N_6525,N_6840);
and U9339 (N_9339,N_5447,N_6536);
nor U9340 (N_9340,N_5043,N_5865);
nor U9341 (N_9341,N_6398,N_7229);
xnor U9342 (N_9342,N_6293,N_6080);
nor U9343 (N_9343,N_6498,N_6289);
or U9344 (N_9344,N_6427,N_7464);
and U9345 (N_9345,N_6113,N_5976);
nor U9346 (N_9346,N_5028,N_7017);
or U9347 (N_9347,N_6575,N_6046);
nor U9348 (N_9348,N_6036,N_5556);
and U9349 (N_9349,N_7490,N_5197);
nor U9350 (N_9350,N_5840,N_5952);
nor U9351 (N_9351,N_5089,N_5709);
xor U9352 (N_9352,N_7100,N_5435);
nor U9353 (N_9353,N_6410,N_5826);
nand U9354 (N_9354,N_5456,N_6055);
xnor U9355 (N_9355,N_6453,N_7116);
nand U9356 (N_9356,N_5958,N_7232);
nor U9357 (N_9357,N_5920,N_5439);
xor U9358 (N_9358,N_6420,N_5815);
nor U9359 (N_9359,N_5293,N_5747);
nor U9360 (N_9360,N_6914,N_6312);
and U9361 (N_9361,N_6512,N_7315);
or U9362 (N_9362,N_5388,N_5023);
nand U9363 (N_9363,N_6957,N_5584);
and U9364 (N_9364,N_5420,N_5785);
xor U9365 (N_9365,N_7016,N_7205);
nand U9366 (N_9366,N_7119,N_6718);
nor U9367 (N_9367,N_5195,N_6646);
nand U9368 (N_9368,N_6234,N_5205);
nand U9369 (N_9369,N_6393,N_6483);
xor U9370 (N_9370,N_7179,N_6941);
nand U9371 (N_9371,N_6468,N_7259);
and U9372 (N_9372,N_5739,N_7120);
or U9373 (N_9373,N_7311,N_6892);
nand U9374 (N_9374,N_5775,N_5456);
nor U9375 (N_9375,N_7350,N_6904);
nand U9376 (N_9376,N_6204,N_6208);
nand U9377 (N_9377,N_5612,N_7176);
and U9378 (N_9378,N_6378,N_7011);
xnor U9379 (N_9379,N_5967,N_6611);
and U9380 (N_9380,N_7030,N_7315);
and U9381 (N_9381,N_6819,N_5102);
xnor U9382 (N_9382,N_6518,N_6587);
nand U9383 (N_9383,N_6805,N_5730);
nand U9384 (N_9384,N_6922,N_5362);
or U9385 (N_9385,N_6309,N_5119);
nand U9386 (N_9386,N_5629,N_6300);
nand U9387 (N_9387,N_6604,N_6582);
and U9388 (N_9388,N_7364,N_7310);
and U9389 (N_9389,N_7083,N_5161);
nand U9390 (N_9390,N_5495,N_5610);
nand U9391 (N_9391,N_7272,N_5896);
nand U9392 (N_9392,N_5713,N_7196);
nor U9393 (N_9393,N_5550,N_5612);
nand U9394 (N_9394,N_7107,N_6200);
nand U9395 (N_9395,N_5613,N_5521);
nand U9396 (N_9396,N_6709,N_5983);
or U9397 (N_9397,N_7275,N_7077);
nand U9398 (N_9398,N_7211,N_5747);
and U9399 (N_9399,N_6694,N_7238);
nor U9400 (N_9400,N_5782,N_5311);
and U9401 (N_9401,N_5141,N_7113);
nand U9402 (N_9402,N_7274,N_5221);
and U9403 (N_9403,N_6101,N_6337);
nand U9404 (N_9404,N_6735,N_7426);
nand U9405 (N_9405,N_7491,N_5306);
nor U9406 (N_9406,N_5945,N_6424);
and U9407 (N_9407,N_5905,N_6060);
xnor U9408 (N_9408,N_6997,N_6361);
nor U9409 (N_9409,N_5269,N_5665);
nor U9410 (N_9410,N_5939,N_5070);
nor U9411 (N_9411,N_5387,N_6052);
xnor U9412 (N_9412,N_6914,N_6832);
and U9413 (N_9413,N_7180,N_5393);
nor U9414 (N_9414,N_7278,N_5795);
xnor U9415 (N_9415,N_5270,N_6163);
and U9416 (N_9416,N_5389,N_6719);
xor U9417 (N_9417,N_6306,N_7488);
nand U9418 (N_9418,N_5208,N_6196);
nor U9419 (N_9419,N_6062,N_6952);
nand U9420 (N_9420,N_6314,N_5680);
and U9421 (N_9421,N_5658,N_5229);
nand U9422 (N_9422,N_6710,N_6645);
and U9423 (N_9423,N_5333,N_6450);
xor U9424 (N_9424,N_7150,N_7486);
and U9425 (N_9425,N_7259,N_5185);
nor U9426 (N_9426,N_7415,N_5931);
nand U9427 (N_9427,N_5396,N_5716);
nor U9428 (N_9428,N_6084,N_6127);
nand U9429 (N_9429,N_5315,N_7104);
xnor U9430 (N_9430,N_7444,N_5040);
and U9431 (N_9431,N_6545,N_7228);
and U9432 (N_9432,N_6210,N_6121);
and U9433 (N_9433,N_5624,N_5547);
and U9434 (N_9434,N_5101,N_5344);
or U9435 (N_9435,N_5311,N_6534);
xor U9436 (N_9436,N_6946,N_5081);
or U9437 (N_9437,N_5949,N_7165);
nor U9438 (N_9438,N_6752,N_6336);
and U9439 (N_9439,N_6970,N_5818);
nand U9440 (N_9440,N_6751,N_6168);
nor U9441 (N_9441,N_5594,N_5571);
or U9442 (N_9442,N_6605,N_6781);
nor U9443 (N_9443,N_5836,N_6195);
nand U9444 (N_9444,N_6482,N_5594);
and U9445 (N_9445,N_6928,N_7255);
nor U9446 (N_9446,N_7208,N_6820);
nand U9447 (N_9447,N_5537,N_6794);
and U9448 (N_9448,N_6447,N_6689);
xnor U9449 (N_9449,N_6709,N_6330);
and U9450 (N_9450,N_5721,N_7252);
xnor U9451 (N_9451,N_7114,N_6118);
xor U9452 (N_9452,N_6511,N_6003);
nand U9453 (N_9453,N_6898,N_6969);
nand U9454 (N_9454,N_6226,N_6142);
or U9455 (N_9455,N_6409,N_6433);
and U9456 (N_9456,N_6732,N_6805);
nor U9457 (N_9457,N_5562,N_6474);
nor U9458 (N_9458,N_5618,N_5229);
nor U9459 (N_9459,N_5067,N_6748);
xnor U9460 (N_9460,N_5727,N_5092);
nand U9461 (N_9461,N_6412,N_5994);
or U9462 (N_9462,N_6883,N_7271);
nor U9463 (N_9463,N_6060,N_6490);
nand U9464 (N_9464,N_5239,N_6353);
nand U9465 (N_9465,N_7242,N_5870);
and U9466 (N_9466,N_7012,N_6156);
nor U9467 (N_9467,N_5702,N_5254);
nand U9468 (N_9468,N_6986,N_5099);
nand U9469 (N_9469,N_7465,N_7299);
xnor U9470 (N_9470,N_7045,N_6030);
xnor U9471 (N_9471,N_6363,N_5242);
xor U9472 (N_9472,N_5528,N_5757);
nor U9473 (N_9473,N_7325,N_7433);
and U9474 (N_9474,N_5452,N_6664);
nand U9475 (N_9475,N_5145,N_5084);
nor U9476 (N_9476,N_7184,N_7280);
xnor U9477 (N_9477,N_6287,N_6255);
nor U9478 (N_9478,N_6972,N_5549);
or U9479 (N_9479,N_5608,N_6380);
and U9480 (N_9480,N_7055,N_5078);
and U9481 (N_9481,N_5116,N_5479);
nand U9482 (N_9482,N_5702,N_6200);
xor U9483 (N_9483,N_6973,N_5982);
or U9484 (N_9484,N_5475,N_6090);
nor U9485 (N_9485,N_6609,N_6565);
xor U9486 (N_9486,N_6281,N_5897);
xnor U9487 (N_9487,N_5766,N_5137);
xor U9488 (N_9488,N_6272,N_5099);
nand U9489 (N_9489,N_5271,N_6280);
xor U9490 (N_9490,N_5215,N_6017);
nand U9491 (N_9491,N_6950,N_7375);
nand U9492 (N_9492,N_7475,N_6016);
and U9493 (N_9493,N_7129,N_5627);
nand U9494 (N_9494,N_5644,N_7220);
nand U9495 (N_9495,N_5186,N_5806);
nor U9496 (N_9496,N_6602,N_7294);
and U9497 (N_9497,N_5164,N_7339);
nor U9498 (N_9498,N_6833,N_5653);
nor U9499 (N_9499,N_5585,N_6607);
or U9500 (N_9500,N_5015,N_5664);
or U9501 (N_9501,N_6301,N_7179);
nor U9502 (N_9502,N_7107,N_6935);
xnor U9503 (N_9503,N_5350,N_5417);
xnor U9504 (N_9504,N_7140,N_5231);
and U9505 (N_9505,N_6787,N_7142);
nand U9506 (N_9506,N_5758,N_6239);
xnor U9507 (N_9507,N_6400,N_5990);
nor U9508 (N_9508,N_5431,N_6006);
xor U9509 (N_9509,N_5998,N_5228);
xor U9510 (N_9510,N_6183,N_5375);
xnor U9511 (N_9511,N_5156,N_6984);
nor U9512 (N_9512,N_6536,N_5233);
or U9513 (N_9513,N_6493,N_6244);
or U9514 (N_9514,N_6709,N_5253);
nand U9515 (N_9515,N_6009,N_7047);
nand U9516 (N_9516,N_6559,N_7090);
or U9517 (N_9517,N_5883,N_5613);
nand U9518 (N_9518,N_5844,N_6593);
or U9519 (N_9519,N_6624,N_5350);
nand U9520 (N_9520,N_6240,N_5445);
nand U9521 (N_9521,N_6764,N_5307);
nor U9522 (N_9522,N_7430,N_7115);
xnor U9523 (N_9523,N_7392,N_5822);
xnor U9524 (N_9524,N_6404,N_6839);
nor U9525 (N_9525,N_7017,N_7009);
xor U9526 (N_9526,N_7207,N_6912);
nand U9527 (N_9527,N_6785,N_7291);
nor U9528 (N_9528,N_6838,N_6140);
xnor U9529 (N_9529,N_7495,N_5465);
nor U9530 (N_9530,N_5128,N_6350);
nor U9531 (N_9531,N_5398,N_5391);
and U9532 (N_9532,N_5670,N_6506);
nor U9533 (N_9533,N_6188,N_5368);
xor U9534 (N_9534,N_7021,N_6503);
or U9535 (N_9535,N_6461,N_5575);
nand U9536 (N_9536,N_7489,N_5964);
and U9537 (N_9537,N_6038,N_7389);
xor U9538 (N_9538,N_5161,N_6001);
xnor U9539 (N_9539,N_6934,N_5954);
or U9540 (N_9540,N_5116,N_6494);
nand U9541 (N_9541,N_6450,N_7468);
nor U9542 (N_9542,N_5497,N_5303);
or U9543 (N_9543,N_6266,N_7215);
or U9544 (N_9544,N_7004,N_5005);
or U9545 (N_9545,N_5021,N_7222);
nor U9546 (N_9546,N_6205,N_6135);
or U9547 (N_9547,N_5243,N_5011);
nand U9548 (N_9548,N_5815,N_7337);
xnor U9549 (N_9549,N_6740,N_5637);
or U9550 (N_9550,N_5115,N_6764);
or U9551 (N_9551,N_5923,N_5399);
or U9552 (N_9552,N_5904,N_6888);
nand U9553 (N_9553,N_6090,N_7134);
nand U9554 (N_9554,N_5214,N_6825);
nor U9555 (N_9555,N_5444,N_6598);
xor U9556 (N_9556,N_6016,N_5518);
or U9557 (N_9557,N_5146,N_5625);
nor U9558 (N_9558,N_6877,N_5778);
xor U9559 (N_9559,N_7192,N_6653);
and U9560 (N_9560,N_6355,N_5527);
nor U9561 (N_9561,N_5965,N_6132);
or U9562 (N_9562,N_6223,N_7061);
nor U9563 (N_9563,N_6174,N_7272);
nand U9564 (N_9564,N_5677,N_5998);
or U9565 (N_9565,N_6418,N_6624);
nand U9566 (N_9566,N_5783,N_6995);
and U9567 (N_9567,N_6469,N_7446);
nand U9568 (N_9568,N_6762,N_5221);
nor U9569 (N_9569,N_6909,N_7063);
nand U9570 (N_9570,N_6317,N_6021);
and U9571 (N_9571,N_7058,N_6734);
nor U9572 (N_9572,N_6764,N_6270);
nand U9573 (N_9573,N_5187,N_7457);
xnor U9574 (N_9574,N_5886,N_6580);
or U9575 (N_9575,N_5287,N_5626);
or U9576 (N_9576,N_5962,N_5197);
nor U9577 (N_9577,N_6013,N_6618);
or U9578 (N_9578,N_5435,N_6868);
nand U9579 (N_9579,N_5906,N_6671);
xor U9580 (N_9580,N_7032,N_6743);
xor U9581 (N_9581,N_6005,N_5694);
xor U9582 (N_9582,N_5788,N_5880);
xnor U9583 (N_9583,N_6531,N_6965);
nor U9584 (N_9584,N_6628,N_6888);
nor U9585 (N_9585,N_5437,N_6658);
xor U9586 (N_9586,N_6688,N_6831);
or U9587 (N_9587,N_5450,N_6913);
nor U9588 (N_9588,N_7134,N_5834);
nand U9589 (N_9589,N_7181,N_6877);
and U9590 (N_9590,N_6522,N_5845);
nand U9591 (N_9591,N_6376,N_6808);
nand U9592 (N_9592,N_5631,N_5484);
nor U9593 (N_9593,N_6710,N_6096);
xnor U9594 (N_9594,N_7385,N_5620);
nor U9595 (N_9595,N_6143,N_5176);
or U9596 (N_9596,N_6435,N_5438);
nand U9597 (N_9597,N_7262,N_6697);
or U9598 (N_9598,N_6178,N_7247);
or U9599 (N_9599,N_7152,N_6464);
nor U9600 (N_9600,N_5043,N_6435);
nor U9601 (N_9601,N_7373,N_5450);
xnor U9602 (N_9602,N_6034,N_5242);
nand U9603 (N_9603,N_6367,N_6621);
and U9604 (N_9604,N_6274,N_6156);
nor U9605 (N_9605,N_5741,N_5071);
or U9606 (N_9606,N_6121,N_5810);
nor U9607 (N_9607,N_6138,N_6854);
nor U9608 (N_9608,N_5919,N_5772);
or U9609 (N_9609,N_7383,N_6407);
or U9610 (N_9610,N_5580,N_5830);
or U9611 (N_9611,N_7143,N_6020);
xnor U9612 (N_9612,N_5387,N_5587);
nand U9613 (N_9613,N_5609,N_5064);
xor U9614 (N_9614,N_5487,N_5562);
xor U9615 (N_9615,N_6060,N_5973);
nor U9616 (N_9616,N_6579,N_6420);
nand U9617 (N_9617,N_6760,N_7167);
and U9618 (N_9618,N_5542,N_7197);
or U9619 (N_9619,N_5191,N_5788);
xnor U9620 (N_9620,N_5552,N_5008);
and U9621 (N_9621,N_5506,N_5980);
xnor U9622 (N_9622,N_5448,N_5001);
or U9623 (N_9623,N_5446,N_7368);
nand U9624 (N_9624,N_5925,N_7064);
or U9625 (N_9625,N_6936,N_6866);
nor U9626 (N_9626,N_7238,N_6669);
nand U9627 (N_9627,N_5960,N_5354);
nand U9628 (N_9628,N_6955,N_6342);
nand U9629 (N_9629,N_5634,N_6363);
and U9630 (N_9630,N_6504,N_5245);
and U9631 (N_9631,N_5798,N_7161);
xnor U9632 (N_9632,N_6003,N_7097);
nand U9633 (N_9633,N_7176,N_6721);
nor U9634 (N_9634,N_5010,N_6283);
nand U9635 (N_9635,N_5876,N_6468);
or U9636 (N_9636,N_7042,N_7394);
nor U9637 (N_9637,N_6701,N_6661);
and U9638 (N_9638,N_6617,N_5690);
nand U9639 (N_9639,N_5908,N_7404);
nor U9640 (N_9640,N_5219,N_6234);
and U9641 (N_9641,N_5067,N_7352);
xnor U9642 (N_9642,N_7212,N_6242);
nand U9643 (N_9643,N_6342,N_5446);
and U9644 (N_9644,N_7062,N_5111);
xnor U9645 (N_9645,N_5053,N_6090);
nor U9646 (N_9646,N_6694,N_5126);
xor U9647 (N_9647,N_5995,N_5671);
nor U9648 (N_9648,N_5551,N_7429);
xnor U9649 (N_9649,N_5584,N_5175);
nand U9650 (N_9650,N_5565,N_7291);
nand U9651 (N_9651,N_6779,N_7438);
and U9652 (N_9652,N_6641,N_6071);
xnor U9653 (N_9653,N_6384,N_6555);
or U9654 (N_9654,N_6847,N_7215);
nand U9655 (N_9655,N_5471,N_5087);
xor U9656 (N_9656,N_6942,N_7002);
xor U9657 (N_9657,N_5551,N_6118);
and U9658 (N_9658,N_6228,N_6756);
or U9659 (N_9659,N_6161,N_6362);
nand U9660 (N_9660,N_7485,N_7358);
nor U9661 (N_9661,N_6749,N_5197);
or U9662 (N_9662,N_6097,N_5344);
and U9663 (N_9663,N_6425,N_6330);
and U9664 (N_9664,N_7213,N_6163);
xor U9665 (N_9665,N_6962,N_5457);
xnor U9666 (N_9666,N_6960,N_5733);
xnor U9667 (N_9667,N_7336,N_7098);
nand U9668 (N_9668,N_6569,N_5193);
nand U9669 (N_9669,N_6924,N_7075);
xnor U9670 (N_9670,N_6000,N_7096);
and U9671 (N_9671,N_6584,N_6884);
nor U9672 (N_9672,N_7277,N_6585);
nand U9673 (N_9673,N_7334,N_6818);
nand U9674 (N_9674,N_6366,N_6126);
nor U9675 (N_9675,N_5939,N_6573);
or U9676 (N_9676,N_5361,N_7290);
nand U9677 (N_9677,N_6589,N_5035);
nand U9678 (N_9678,N_5251,N_6958);
and U9679 (N_9679,N_6490,N_6307);
xor U9680 (N_9680,N_7328,N_6642);
and U9681 (N_9681,N_5007,N_5953);
or U9682 (N_9682,N_7363,N_7209);
or U9683 (N_9683,N_6068,N_5907);
xor U9684 (N_9684,N_7029,N_6215);
or U9685 (N_9685,N_6098,N_6132);
or U9686 (N_9686,N_6238,N_5503);
or U9687 (N_9687,N_7112,N_7265);
nand U9688 (N_9688,N_5859,N_7337);
nor U9689 (N_9689,N_5290,N_5352);
nor U9690 (N_9690,N_6962,N_6349);
or U9691 (N_9691,N_5377,N_6663);
nand U9692 (N_9692,N_5510,N_5439);
nand U9693 (N_9693,N_5306,N_7056);
nand U9694 (N_9694,N_7297,N_6440);
xor U9695 (N_9695,N_6515,N_5953);
or U9696 (N_9696,N_6277,N_5106);
or U9697 (N_9697,N_5648,N_5115);
nor U9698 (N_9698,N_5887,N_7125);
or U9699 (N_9699,N_6016,N_5228);
and U9700 (N_9700,N_6763,N_6974);
or U9701 (N_9701,N_7376,N_5925);
or U9702 (N_9702,N_6427,N_6223);
or U9703 (N_9703,N_5838,N_6067);
xor U9704 (N_9704,N_5063,N_6875);
xor U9705 (N_9705,N_5404,N_6735);
and U9706 (N_9706,N_7463,N_6906);
and U9707 (N_9707,N_6511,N_5338);
or U9708 (N_9708,N_7360,N_5372);
nand U9709 (N_9709,N_6555,N_6251);
and U9710 (N_9710,N_6586,N_5903);
nor U9711 (N_9711,N_5781,N_5972);
xor U9712 (N_9712,N_6098,N_5415);
nor U9713 (N_9713,N_5484,N_7236);
nor U9714 (N_9714,N_5235,N_6934);
xor U9715 (N_9715,N_7238,N_7090);
nor U9716 (N_9716,N_7225,N_6636);
xor U9717 (N_9717,N_5238,N_6631);
or U9718 (N_9718,N_5209,N_7162);
nor U9719 (N_9719,N_6773,N_5036);
and U9720 (N_9720,N_7460,N_5652);
nor U9721 (N_9721,N_7359,N_5833);
nor U9722 (N_9722,N_6844,N_6895);
xnor U9723 (N_9723,N_7164,N_5806);
nor U9724 (N_9724,N_5879,N_5228);
or U9725 (N_9725,N_7496,N_6759);
nor U9726 (N_9726,N_5203,N_6482);
or U9727 (N_9727,N_5398,N_7154);
or U9728 (N_9728,N_6533,N_7335);
xnor U9729 (N_9729,N_6653,N_6448);
nand U9730 (N_9730,N_6661,N_7013);
and U9731 (N_9731,N_7330,N_6121);
or U9732 (N_9732,N_5227,N_5262);
xnor U9733 (N_9733,N_5099,N_7281);
or U9734 (N_9734,N_6821,N_7116);
xor U9735 (N_9735,N_5402,N_7379);
and U9736 (N_9736,N_5751,N_6153);
nor U9737 (N_9737,N_6370,N_6890);
nand U9738 (N_9738,N_5513,N_6399);
nand U9739 (N_9739,N_6758,N_6873);
and U9740 (N_9740,N_7358,N_7119);
nand U9741 (N_9741,N_6052,N_7216);
nand U9742 (N_9742,N_6823,N_7369);
xnor U9743 (N_9743,N_5785,N_7024);
and U9744 (N_9744,N_6704,N_6670);
nand U9745 (N_9745,N_5263,N_5587);
xor U9746 (N_9746,N_5824,N_6594);
nor U9747 (N_9747,N_7192,N_6565);
or U9748 (N_9748,N_5409,N_6507);
or U9749 (N_9749,N_6666,N_5335);
or U9750 (N_9750,N_7207,N_5429);
and U9751 (N_9751,N_5504,N_5619);
and U9752 (N_9752,N_6754,N_5570);
and U9753 (N_9753,N_6556,N_5481);
and U9754 (N_9754,N_6236,N_6744);
nor U9755 (N_9755,N_6466,N_5056);
xor U9756 (N_9756,N_6479,N_7049);
xor U9757 (N_9757,N_5140,N_7491);
nor U9758 (N_9758,N_6215,N_7496);
and U9759 (N_9759,N_5197,N_5752);
xnor U9760 (N_9760,N_5217,N_6561);
nand U9761 (N_9761,N_6955,N_6833);
and U9762 (N_9762,N_6470,N_6034);
nand U9763 (N_9763,N_6681,N_5334);
or U9764 (N_9764,N_7342,N_6339);
nand U9765 (N_9765,N_7275,N_6600);
nand U9766 (N_9766,N_7131,N_7367);
xnor U9767 (N_9767,N_5719,N_5819);
xnor U9768 (N_9768,N_5470,N_6679);
nand U9769 (N_9769,N_5416,N_7101);
or U9770 (N_9770,N_6477,N_7263);
and U9771 (N_9771,N_6449,N_6871);
xor U9772 (N_9772,N_6464,N_5261);
nor U9773 (N_9773,N_6036,N_6464);
and U9774 (N_9774,N_5974,N_5782);
or U9775 (N_9775,N_5394,N_7159);
xnor U9776 (N_9776,N_5202,N_7232);
nand U9777 (N_9777,N_6200,N_6603);
or U9778 (N_9778,N_5506,N_6388);
nor U9779 (N_9779,N_7491,N_7435);
nor U9780 (N_9780,N_7106,N_5321);
nor U9781 (N_9781,N_6373,N_5152);
nand U9782 (N_9782,N_6219,N_7410);
and U9783 (N_9783,N_6573,N_5191);
xor U9784 (N_9784,N_5721,N_7133);
and U9785 (N_9785,N_6486,N_7282);
or U9786 (N_9786,N_7395,N_6144);
xor U9787 (N_9787,N_5665,N_7398);
xor U9788 (N_9788,N_6115,N_6928);
xnor U9789 (N_9789,N_5581,N_6862);
or U9790 (N_9790,N_7009,N_5040);
xor U9791 (N_9791,N_5997,N_7352);
or U9792 (N_9792,N_5701,N_5636);
or U9793 (N_9793,N_6784,N_6937);
or U9794 (N_9794,N_5851,N_6128);
nor U9795 (N_9795,N_6555,N_5096);
xnor U9796 (N_9796,N_5772,N_6676);
nor U9797 (N_9797,N_5532,N_7435);
nor U9798 (N_9798,N_6724,N_5299);
xnor U9799 (N_9799,N_7117,N_7198);
nor U9800 (N_9800,N_6937,N_6603);
or U9801 (N_9801,N_6684,N_6016);
or U9802 (N_9802,N_7258,N_5077);
or U9803 (N_9803,N_5608,N_6104);
and U9804 (N_9804,N_5651,N_5835);
nand U9805 (N_9805,N_5081,N_5881);
or U9806 (N_9806,N_5604,N_7448);
nand U9807 (N_9807,N_6130,N_5041);
or U9808 (N_9808,N_6336,N_7488);
nand U9809 (N_9809,N_5198,N_6550);
xnor U9810 (N_9810,N_6221,N_5014);
nor U9811 (N_9811,N_6751,N_7100);
nor U9812 (N_9812,N_6590,N_6834);
and U9813 (N_9813,N_7049,N_5148);
nor U9814 (N_9814,N_6818,N_6804);
or U9815 (N_9815,N_6548,N_6052);
nand U9816 (N_9816,N_7165,N_5194);
nand U9817 (N_9817,N_5870,N_6433);
nand U9818 (N_9818,N_6215,N_5559);
nand U9819 (N_9819,N_7041,N_6281);
and U9820 (N_9820,N_5860,N_6299);
and U9821 (N_9821,N_5913,N_5312);
nand U9822 (N_9822,N_6448,N_6020);
nor U9823 (N_9823,N_5860,N_7144);
and U9824 (N_9824,N_6668,N_5834);
and U9825 (N_9825,N_6050,N_7319);
nor U9826 (N_9826,N_7485,N_5245);
xnor U9827 (N_9827,N_5621,N_5970);
xnor U9828 (N_9828,N_5715,N_7129);
or U9829 (N_9829,N_5289,N_6103);
and U9830 (N_9830,N_5710,N_7310);
or U9831 (N_9831,N_6881,N_6630);
nor U9832 (N_9832,N_7091,N_6409);
xor U9833 (N_9833,N_5127,N_6461);
xor U9834 (N_9834,N_5187,N_5397);
or U9835 (N_9835,N_5754,N_6603);
nand U9836 (N_9836,N_5203,N_6242);
xnor U9837 (N_9837,N_7118,N_5478);
xor U9838 (N_9838,N_5056,N_6721);
nor U9839 (N_9839,N_6206,N_5771);
nand U9840 (N_9840,N_7185,N_6480);
and U9841 (N_9841,N_6253,N_6361);
nor U9842 (N_9842,N_6730,N_5607);
or U9843 (N_9843,N_7457,N_7078);
xnor U9844 (N_9844,N_6572,N_5917);
or U9845 (N_9845,N_6172,N_6873);
nor U9846 (N_9846,N_5658,N_6882);
or U9847 (N_9847,N_7219,N_5002);
nor U9848 (N_9848,N_5024,N_5902);
nand U9849 (N_9849,N_5215,N_6086);
nor U9850 (N_9850,N_7286,N_5783);
xnor U9851 (N_9851,N_5133,N_5810);
nor U9852 (N_9852,N_7054,N_7300);
xor U9853 (N_9853,N_6956,N_5951);
nor U9854 (N_9854,N_5838,N_7143);
and U9855 (N_9855,N_5019,N_6551);
or U9856 (N_9856,N_5389,N_5593);
and U9857 (N_9857,N_6018,N_6589);
and U9858 (N_9858,N_5742,N_5360);
xor U9859 (N_9859,N_5315,N_6601);
xnor U9860 (N_9860,N_5241,N_6313);
xnor U9861 (N_9861,N_5948,N_6646);
nor U9862 (N_9862,N_6381,N_7090);
or U9863 (N_9863,N_6806,N_7397);
nor U9864 (N_9864,N_6507,N_6617);
nor U9865 (N_9865,N_6786,N_6077);
or U9866 (N_9866,N_5227,N_6037);
and U9867 (N_9867,N_7041,N_7077);
xnor U9868 (N_9868,N_7425,N_6532);
and U9869 (N_9869,N_5903,N_5569);
or U9870 (N_9870,N_6708,N_5266);
and U9871 (N_9871,N_6341,N_5847);
nor U9872 (N_9872,N_7403,N_5371);
nor U9873 (N_9873,N_7258,N_6248);
or U9874 (N_9874,N_6413,N_7064);
nand U9875 (N_9875,N_7056,N_7152);
nand U9876 (N_9876,N_6968,N_5422);
xor U9877 (N_9877,N_6959,N_7360);
nor U9878 (N_9878,N_7060,N_5098);
or U9879 (N_9879,N_7068,N_6695);
or U9880 (N_9880,N_6328,N_5772);
nand U9881 (N_9881,N_6161,N_6409);
and U9882 (N_9882,N_5805,N_6536);
xnor U9883 (N_9883,N_5841,N_5911);
xnor U9884 (N_9884,N_5102,N_6312);
nand U9885 (N_9885,N_5424,N_6448);
xor U9886 (N_9886,N_5988,N_6343);
or U9887 (N_9887,N_6333,N_5616);
nor U9888 (N_9888,N_6040,N_5341);
nand U9889 (N_9889,N_6880,N_5715);
nand U9890 (N_9890,N_5306,N_7163);
nand U9891 (N_9891,N_6285,N_6842);
xor U9892 (N_9892,N_6170,N_5130);
nor U9893 (N_9893,N_5270,N_7463);
xor U9894 (N_9894,N_5886,N_6017);
nand U9895 (N_9895,N_6578,N_7406);
or U9896 (N_9896,N_5758,N_7248);
nor U9897 (N_9897,N_6213,N_5467);
and U9898 (N_9898,N_5922,N_6995);
nor U9899 (N_9899,N_5158,N_7163);
or U9900 (N_9900,N_6378,N_5136);
and U9901 (N_9901,N_6996,N_6621);
nand U9902 (N_9902,N_6939,N_7424);
nor U9903 (N_9903,N_5878,N_5626);
nor U9904 (N_9904,N_5771,N_5672);
or U9905 (N_9905,N_7490,N_5163);
xor U9906 (N_9906,N_7120,N_6949);
nor U9907 (N_9907,N_5650,N_6740);
nand U9908 (N_9908,N_5281,N_5478);
nor U9909 (N_9909,N_5760,N_7279);
xor U9910 (N_9910,N_6775,N_6428);
nor U9911 (N_9911,N_7111,N_5477);
nor U9912 (N_9912,N_5526,N_6211);
or U9913 (N_9913,N_7464,N_5002);
or U9914 (N_9914,N_5368,N_7031);
nand U9915 (N_9915,N_6294,N_5812);
nor U9916 (N_9916,N_6167,N_6544);
xor U9917 (N_9917,N_5029,N_7248);
or U9918 (N_9918,N_7010,N_5414);
and U9919 (N_9919,N_7121,N_5245);
xor U9920 (N_9920,N_6949,N_6818);
nor U9921 (N_9921,N_6599,N_5853);
or U9922 (N_9922,N_6349,N_7090);
and U9923 (N_9923,N_5563,N_7426);
nand U9924 (N_9924,N_5150,N_6695);
or U9925 (N_9925,N_5851,N_6892);
nand U9926 (N_9926,N_6242,N_5778);
nand U9927 (N_9927,N_6666,N_6808);
and U9928 (N_9928,N_5674,N_5531);
xnor U9929 (N_9929,N_5366,N_5075);
and U9930 (N_9930,N_6458,N_5739);
nor U9931 (N_9931,N_6392,N_5624);
or U9932 (N_9932,N_6375,N_5949);
nand U9933 (N_9933,N_6535,N_6184);
xor U9934 (N_9934,N_7013,N_6576);
nor U9935 (N_9935,N_5752,N_5248);
or U9936 (N_9936,N_6627,N_5513);
or U9937 (N_9937,N_5171,N_7164);
nand U9938 (N_9938,N_5870,N_6019);
and U9939 (N_9939,N_5301,N_5422);
or U9940 (N_9940,N_7251,N_5689);
nand U9941 (N_9941,N_5563,N_5513);
and U9942 (N_9942,N_6262,N_5871);
nor U9943 (N_9943,N_5796,N_6974);
nor U9944 (N_9944,N_5682,N_6425);
nand U9945 (N_9945,N_6030,N_5959);
nor U9946 (N_9946,N_5569,N_5271);
or U9947 (N_9947,N_5032,N_5357);
and U9948 (N_9948,N_5845,N_5414);
or U9949 (N_9949,N_6461,N_6871);
xnor U9950 (N_9950,N_5267,N_6670);
nor U9951 (N_9951,N_6334,N_5940);
and U9952 (N_9952,N_5880,N_6051);
nor U9953 (N_9953,N_5646,N_5494);
xnor U9954 (N_9954,N_5413,N_5703);
and U9955 (N_9955,N_7166,N_6306);
or U9956 (N_9956,N_6176,N_5284);
and U9957 (N_9957,N_7079,N_6506);
or U9958 (N_9958,N_6672,N_5532);
xor U9959 (N_9959,N_6323,N_6000);
nor U9960 (N_9960,N_7342,N_5180);
or U9961 (N_9961,N_6254,N_5296);
nand U9962 (N_9962,N_7244,N_7321);
xor U9963 (N_9963,N_6797,N_6589);
or U9964 (N_9964,N_5370,N_6259);
and U9965 (N_9965,N_6410,N_6777);
nand U9966 (N_9966,N_5067,N_7194);
or U9967 (N_9967,N_6942,N_6620);
nor U9968 (N_9968,N_6008,N_6518);
or U9969 (N_9969,N_5630,N_6944);
nand U9970 (N_9970,N_6885,N_5529);
nand U9971 (N_9971,N_6615,N_5500);
xnor U9972 (N_9972,N_6894,N_6081);
nor U9973 (N_9973,N_5270,N_7123);
xnor U9974 (N_9974,N_6300,N_6807);
and U9975 (N_9975,N_6795,N_6185);
and U9976 (N_9976,N_6407,N_7127);
nor U9977 (N_9977,N_7317,N_6813);
nand U9978 (N_9978,N_5960,N_5958);
nand U9979 (N_9979,N_7396,N_7371);
xor U9980 (N_9980,N_6378,N_5831);
xor U9981 (N_9981,N_6001,N_5366);
nand U9982 (N_9982,N_5166,N_5340);
and U9983 (N_9983,N_5718,N_6615);
xnor U9984 (N_9984,N_6831,N_6860);
nor U9985 (N_9985,N_5388,N_7332);
nor U9986 (N_9986,N_5833,N_5274);
and U9987 (N_9987,N_5811,N_6675);
xnor U9988 (N_9988,N_6576,N_6800);
xnor U9989 (N_9989,N_6426,N_7148);
and U9990 (N_9990,N_6139,N_6256);
xor U9991 (N_9991,N_7204,N_7103);
nor U9992 (N_9992,N_5328,N_6851);
xor U9993 (N_9993,N_7274,N_6292);
or U9994 (N_9994,N_7007,N_6406);
nor U9995 (N_9995,N_5021,N_6171);
nand U9996 (N_9996,N_6028,N_7044);
and U9997 (N_9997,N_6488,N_5530);
nand U9998 (N_9998,N_6630,N_6875);
or U9999 (N_9999,N_6874,N_5757);
and U10000 (N_10000,N_7859,N_9952);
or U10001 (N_10001,N_8394,N_9716);
nand U10002 (N_10002,N_7599,N_8629);
and U10003 (N_10003,N_9332,N_7724);
and U10004 (N_10004,N_7586,N_9596);
nand U10005 (N_10005,N_8578,N_9469);
xnor U10006 (N_10006,N_9497,N_8801);
or U10007 (N_10007,N_9437,N_8609);
or U10008 (N_10008,N_8999,N_9205);
or U10009 (N_10009,N_8740,N_7884);
nand U10010 (N_10010,N_7720,N_9159);
xor U10011 (N_10011,N_9589,N_7940);
nor U10012 (N_10012,N_8527,N_7662);
xnor U10013 (N_10013,N_9034,N_8473);
xnor U10014 (N_10014,N_8724,N_9068);
nor U10015 (N_10015,N_8431,N_9454);
xnor U10016 (N_10016,N_8677,N_7556);
nor U10017 (N_10017,N_8734,N_8448);
xor U10018 (N_10018,N_8576,N_9173);
or U10019 (N_10019,N_7627,N_7637);
nand U10020 (N_10020,N_9770,N_8455);
and U10021 (N_10021,N_8514,N_9496);
nor U10022 (N_10022,N_8602,N_8841);
or U10023 (N_10023,N_9305,N_9664);
xor U10024 (N_10024,N_8275,N_7995);
nor U10025 (N_10025,N_8018,N_7527);
nand U10026 (N_10026,N_9398,N_7520);
and U10027 (N_10027,N_8726,N_7957);
xor U10028 (N_10028,N_9624,N_9553);
xnor U10029 (N_10029,N_7779,N_8004);
xor U10030 (N_10030,N_7998,N_8761);
and U10031 (N_10031,N_8513,N_7747);
nand U10032 (N_10032,N_8402,N_9477);
xnor U10033 (N_10033,N_7781,N_7893);
or U10034 (N_10034,N_9765,N_9319);
xnor U10035 (N_10035,N_8154,N_7846);
nor U10036 (N_10036,N_8057,N_7948);
nor U10037 (N_10037,N_9775,N_9285);
nor U10038 (N_10038,N_9550,N_9012);
and U10039 (N_10039,N_9405,N_9588);
xor U10040 (N_10040,N_8763,N_8650);
and U10041 (N_10041,N_7541,N_7792);
nand U10042 (N_10042,N_9923,N_9857);
nor U10043 (N_10043,N_8096,N_7544);
nand U10044 (N_10044,N_9853,N_9823);
xnor U10045 (N_10045,N_8550,N_9184);
xor U10046 (N_10046,N_7934,N_8203);
xor U10047 (N_10047,N_8745,N_9888);
nand U10048 (N_10048,N_8844,N_9449);
and U10049 (N_10049,N_8707,N_8399);
nor U10050 (N_10050,N_9875,N_8437);
and U10051 (N_10051,N_9687,N_8387);
xnor U10052 (N_10052,N_8189,N_9583);
and U10053 (N_10053,N_8069,N_8517);
and U10054 (N_10054,N_9599,N_8406);
nand U10055 (N_10055,N_8133,N_8416);
xor U10056 (N_10056,N_9413,N_9925);
xor U10057 (N_10057,N_9994,N_9507);
and U10058 (N_10058,N_9468,N_7980);
xor U10059 (N_10059,N_8738,N_7587);
xor U10060 (N_10060,N_8414,N_8151);
xor U10061 (N_10061,N_8666,N_7689);
xor U10062 (N_10062,N_8451,N_9234);
nor U10063 (N_10063,N_9555,N_8026);
or U10064 (N_10064,N_7947,N_9804);
nand U10065 (N_10065,N_8815,N_7744);
nand U10066 (N_10066,N_7964,N_9799);
and U10067 (N_10067,N_8869,N_8560);
nor U10068 (N_10068,N_9979,N_8405);
and U10069 (N_10069,N_9341,N_9658);
nor U10070 (N_10070,N_7699,N_9115);
nor U10071 (N_10071,N_8935,N_8281);
or U10072 (N_10072,N_8000,N_8045);
nor U10073 (N_10073,N_8652,N_7959);
xnor U10074 (N_10074,N_9248,N_9053);
nor U10075 (N_10075,N_8078,N_8334);
or U10076 (N_10076,N_9648,N_8598);
and U10077 (N_10077,N_9443,N_8593);
nand U10078 (N_10078,N_8226,N_8600);
nor U10079 (N_10079,N_9239,N_8306);
or U10080 (N_10080,N_8065,N_8201);
nand U10081 (N_10081,N_7543,N_9220);
nor U10082 (N_10082,N_9554,N_8885);
nor U10083 (N_10083,N_8723,N_8524);
xor U10084 (N_10084,N_7723,N_8349);
or U10085 (N_10085,N_8710,N_9995);
or U10086 (N_10086,N_9734,N_7547);
nor U10087 (N_10087,N_9386,N_8345);
nor U10088 (N_10088,N_9841,N_8950);
nor U10089 (N_10089,N_9439,N_9794);
nor U10090 (N_10090,N_8274,N_7821);
and U10091 (N_10091,N_8411,N_7869);
and U10092 (N_10092,N_9755,N_8456);
xnor U10093 (N_10093,N_9038,N_8188);
or U10094 (N_10094,N_7665,N_9943);
xor U10095 (N_10095,N_9800,N_9733);
and U10096 (N_10096,N_8419,N_7932);
nor U10097 (N_10097,N_8941,N_7755);
nand U10098 (N_10098,N_9087,N_9339);
nor U10099 (N_10099,N_8436,N_8897);
and U10100 (N_10100,N_8244,N_9647);
nand U10101 (N_10101,N_8906,N_9263);
nor U10102 (N_10102,N_7643,N_9783);
xor U10103 (N_10103,N_9269,N_8596);
and U10104 (N_10104,N_8486,N_8376);
and U10105 (N_10105,N_9201,N_9340);
nor U10106 (N_10106,N_7786,N_7745);
nor U10107 (N_10107,N_8725,N_9662);
and U10108 (N_10108,N_9430,N_8315);
and U10109 (N_10109,N_9296,N_7944);
and U10110 (N_10110,N_9819,N_9007);
or U10111 (N_10111,N_9880,N_8110);
nand U10112 (N_10112,N_8926,N_7954);
and U10113 (N_10113,N_8965,N_9577);
and U10114 (N_10114,N_9098,N_8466);
xnor U10115 (N_10115,N_9621,N_8227);
nand U10116 (N_10116,N_9187,N_7560);
nor U10117 (N_10117,N_8880,N_7892);
nor U10118 (N_10118,N_9851,N_9354);
or U10119 (N_10119,N_7610,N_8491);
nor U10120 (N_10120,N_8239,N_9899);
nand U10121 (N_10121,N_8417,N_7653);
nor U10122 (N_10122,N_9470,N_8049);
or U10123 (N_10123,N_7870,N_8266);
nor U10124 (N_10124,N_8832,N_8344);
nor U10125 (N_10125,N_9283,N_8637);
or U10126 (N_10126,N_9627,N_9180);
nand U10127 (N_10127,N_8521,N_9459);
nor U10128 (N_10128,N_9362,N_9512);
or U10129 (N_10129,N_7507,N_9645);
or U10130 (N_10130,N_9135,N_8862);
xor U10131 (N_10131,N_8833,N_7806);
and U10132 (N_10132,N_7851,N_8016);
nor U10133 (N_10133,N_8930,N_9750);
or U10134 (N_10134,N_8787,N_9069);
or U10135 (N_10135,N_7624,N_8317);
nand U10136 (N_10136,N_8352,N_8307);
xnor U10137 (N_10137,N_7914,N_9077);
or U10138 (N_10138,N_9407,N_8704);
nor U10139 (N_10139,N_9921,N_8050);
nor U10140 (N_10140,N_8805,N_8942);
xnor U10141 (N_10141,N_9877,N_8728);
or U10142 (N_10142,N_8509,N_9969);
xnor U10143 (N_10143,N_8933,N_7801);
or U10144 (N_10144,N_9030,N_9297);
nand U10145 (N_10145,N_9705,N_8720);
and U10146 (N_10146,N_7608,N_8401);
and U10147 (N_10147,N_8665,N_9910);
xnor U10148 (N_10148,N_9552,N_8490);
nor U10149 (N_10149,N_8631,N_8443);
or U10150 (N_10150,N_8138,N_9196);
nand U10151 (N_10151,N_8791,N_9856);
or U10152 (N_10152,N_9421,N_9420);
or U10153 (N_10153,N_8536,N_7925);
and U10154 (N_10154,N_9935,N_9282);
nand U10155 (N_10155,N_9915,N_9380);
and U10156 (N_10156,N_7926,N_9186);
nand U10157 (N_10157,N_8530,N_8085);
or U10158 (N_10158,N_9118,N_8870);
xor U10159 (N_10159,N_9383,N_8161);
xor U10160 (N_10160,N_8464,N_8316);
nand U10161 (N_10161,N_8015,N_7579);
or U10162 (N_10162,N_9440,N_7636);
and U10163 (N_10163,N_9571,N_8569);
nor U10164 (N_10164,N_7928,N_8440);
xor U10165 (N_10165,N_9475,N_7886);
nand U10166 (N_10166,N_8916,N_9243);
or U10167 (N_10167,N_9491,N_7858);
and U10168 (N_10168,N_9618,N_9753);
and U10169 (N_10169,N_8852,N_8785);
nand U10170 (N_10170,N_7555,N_8231);
and U10171 (N_10171,N_9541,N_8857);
nor U10172 (N_10172,N_7885,N_9219);
nor U10173 (N_10173,N_8714,N_8322);
and U10174 (N_10174,N_8978,N_9999);
nand U10175 (N_10175,N_8716,N_8117);
nand U10176 (N_10176,N_8743,N_8675);
nor U10177 (N_10177,N_7728,N_8071);
or U10178 (N_10178,N_9972,N_9036);
nor U10179 (N_10179,N_9050,N_9978);
or U10180 (N_10180,N_7970,N_8195);
or U10181 (N_10181,N_8100,N_8846);
and U10182 (N_10182,N_7890,N_8503);
and U10183 (N_10183,N_9818,N_7647);
xnor U10184 (N_10184,N_9873,N_9633);
or U10185 (N_10185,N_9229,N_8892);
or U10186 (N_10186,N_9182,N_9506);
nand U10187 (N_10187,N_7984,N_9820);
nor U10188 (N_10188,N_9350,N_8347);
and U10189 (N_10189,N_7502,N_9892);
nand U10190 (N_10190,N_8175,N_7950);
xor U10191 (N_10191,N_9048,N_9883);
or U10192 (N_10192,N_8953,N_9501);
xnor U10193 (N_10193,N_9458,N_8485);
xnor U10194 (N_10194,N_9065,N_7688);
and U10195 (N_10195,N_9612,N_8337);
or U10196 (N_10196,N_8848,N_8077);
or U10197 (N_10197,N_9763,N_8945);
and U10198 (N_10198,N_8789,N_9456);
nand U10199 (N_10199,N_9587,N_7684);
and U10200 (N_10200,N_9836,N_8487);
and U10201 (N_10201,N_9432,N_7816);
nor U10202 (N_10202,N_9756,N_9997);
xnor U10203 (N_10203,N_8441,N_9345);
nand U10204 (N_10204,N_9408,N_9441);
and U10205 (N_10205,N_7788,N_9230);
nor U10206 (N_10206,N_8328,N_9232);
xor U10207 (N_10207,N_7711,N_7670);
xnor U10208 (N_10208,N_8254,N_8624);
and U10209 (N_10209,N_9902,N_9516);
or U10210 (N_10210,N_9642,N_7550);
xor U10211 (N_10211,N_8033,N_8397);
xor U10212 (N_10212,N_9998,N_9970);
and U10213 (N_10213,N_8169,N_9293);
xor U10214 (N_10214,N_8878,N_8899);
and U10215 (N_10215,N_7762,N_7820);
or U10216 (N_10216,N_9575,N_7659);
xnor U10217 (N_10217,N_8364,N_8649);
or U10218 (N_10218,N_8072,N_9211);
xnor U10219 (N_10219,N_8236,N_7585);
and U10220 (N_10220,N_9886,N_9780);
nor U10221 (N_10221,N_7805,N_8558);
or U10222 (N_10222,N_9813,N_9832);
nor U10223 (N_10223,N_9370,N_8034);
or U10224 (N_10224,N_9120,N_9758);
and U10225 (N_10225,N_9369,N_8752);
or U10226 (N_10226,N_9809,N_8181);
nor U10227 (N_10227,N_8240,N_7509);
and U10228 (N_10228,N_8238,N_8835);
xnor U10229 (N_10229,N_8084,N_8967);
or U10230 (N_10230,N_8127,N_9948);
nor U10231 (N_10231,N_9063,N_9467);
and U10232 (N_10232,N_8540,N_7853);
nand U10233 (N_10233,N_8186,N_9425);
or U10234 (N_10234,N_9958,N_8482);
nand U10235 (N_10235,N_9485,N_9314);
nor U10236 (N_10236,N_8934,N_9940);
or U10237 (N_10237,N_9917,N_8288);
xor U10238 (N_10238,N_8863,N_7833);
or U10239 (N_10239,N_9592,N_9391);
xor U10240 (N_10240,N_8040,N_9066);
and U10241 (N_10241,N_8037,N_9130);
nand U10242 (N_10242,N_7522,N_9827);
nand U10243 (N_10243,N_8125,N_8960);
nor U10244 (N_10244,N_9200,N_8770);
nand U10245 (N_10245,N_8054,N_9580);
nor U10246 (N_10246,N_9572,N_9812);
nor U10247 (N_10247,N_8961,N_9073);
xnor U10248 (N_10248,N_8122,N_9271);
xor U10249 (N_10249,N_9895,N_8512);
nand U10250 (N_10250,N_9792,N_8375);
nand U10251 (N_10251,N_7798,N_9942);
and U10252 (N_10252,N_8528,N_8171);
nor U10253 (N_10253,N_9183,N_9158);
nor U10254 (N_10254,N_8882,N_8116);
nor U10255 (N_10255,N_8006,N_8447);
nand U10256 (N_10256,N_7810,N_8595);
and U10257 (N_10257,N_8747,N_9304);
or U10258 (N_10258,N_9643,N_8165);
or U10259 (N_10259,N_8476,N_9249);
nor U10260 (N_10260,N_9896,N_9395);
nor U10261 (N_10261,N_7867,N_8147);
nand U10262 (N_10262,N_9690,N_8717);
nor U10263 (N_10263,N_8971,N_9672);
nor U10264 (N_10264,N_9737,N_7584);
and U10265 (N_10265,N_7681,N_8939);
nand U10266 (N_10266,N_8075,N_9493);
or U10267 (N_10267,N_9387,N_8366);
nor U10268 (N_10268,N_9424,N_7749);
nand U10269 (N_10269,N_8928,N_9075);
nand U10270 (N_10270,N_7633,N_7825);
and U10271 (N_10271,N_8706,N_8479);
nor U10272 (N_10272,N_8190,N_9093);
xnor U10273 (N_10273,N_8124,N_8561);
xnor U10274 (N_10274,N_8287,N_8118);
or U10275 (N_10275,N_9517,N_9535);
and U10276 (N_10276,N_8036,N_7878);
and U10277 (N_10277,N_8383,N_8759);
and U10278 (N_10278,N_8470,N_7648);
nor U10279 (N_10279,N_9450,N_8721);
nand U10280 (N_10280,N_7743,N_8319);
or U10281 (N_10281,N_7604,N_7561);
or U10282 (N_10282,N_7603,N_8424);
and U10283 (N_10283,N_8299,N_9963);
or U10284 (N_10284,N_7905,N_8699);
or U10285 (N_10285,N_8691,N_9004);
xnor U10286 (N_10286,N_9021,N_8647);
nor U10287 (N_10287,N_7916,N_8619);
xnor U10288 (N_10288,N_8948,N_9966);
nand U10289 (N_10289,N_8554,N_9035);
nand U10290 (N_10290,N_8768,N_7528);
and U10291 (N_10291,N_8333,N_9540);
nor U10292 (N_10292,N_8886,N_9730);
and U10293 (N_10293,N_9971,N_7739);
and U10294 (N_10294,N_7683,N_8879);
and U10295 (N_10295,N_8086,N_8755);
and U10296 (N_10296,N_7622,N_8727);
or U10297 (N_10297,N_9164,N_9166);
and U10298 (N_10298,N_7758,N_9129);
and U10299 (N_10299,N_8904,N_9404);
xnor U10300 (N_10300,N_7746,N_8061);
or U10301 (N_10301,N_8143,N_8263);
nor U10302 (N_10302,N_7500,N_8860);
or U10303 (N_10303,N_9289,N_8611);
nand U10304 (N_10304,N_9774,N_8659);
and U10305 (N_10305,N_8991,N_9167);
and U10306 (N_10306,N_7646,N_9381);
and U10307 (N_10307,N_8010,N_9336);
nand U10308 (N_10308,N_7795,N_9353);
or U10309 (N_10309,N_8856,N_8267);
nand U10310 (N_10310,N_8362,N_8280);
or U10311 (N_10311,N_8947,N_8449);
nand U10312 (N_10312,N_7857,N_7975);
xnor U10313 (N_10313,N_8702,N_9652);
nand U10314 (N_10314,N_7730,N_8774);
or U10315 (N_10315,N_8380,N_8511);
nor U10316 (N_10316,N_9584,N_8183);
nor U10317 (N_10317,N_8048,N_9711);
nand U10318 (N_10318,N_8258,N_9106);
and U10319 (N_10319,N_9586,N_9208);
nor U10320 (N_10320,N_9616,N_9879);
xor U10321 (N_10321,N_8821,N_8620);
and U10322 (N_10322,N_9446,N_8750);
nor U10323 (N_10323,N_7524,N_9505);
nand U10324 (N_10324,N_9975,N_9835);
and U10325 (N_10325,N_7922,N_7673);
or U10326 (N_10326,N_9842,N_9529);
nand U10327 (N_10327,N_8070,N_7834);
xnor U10328 (N_10328,N_9157,N_7563);
nor U10329 (N_10329,N_9613,N_8655);
nor U10330 (N_10330,N_7876,N_7967);
xor U10331 (N_10331,N_8887,N_9742);
or U10332 (N_10332,N_9677,N_9573);
or U10333 (N_10333,N_9214,N_8888);
nor U10334 (N_10334,N_7668,N_8775);
nand U10335 (N_10335,N_8229,N_9257);
and U10336 (N_10336,N_8444,N_9266);
nand U10337 (N_10337,N_9151,N_7824);
nand U10338 (N_10338,N_8241,N_7952);
xnor U10339 (N_10339,N_7750,N_8588);
and U10340 (N_10340,N_8243,N_9791);
and U10341 (N_10341,N_8784,N_9761);
nor U10342 (N_10342,N_9356,N_8095);
xor U10343 (N_10343,N_8901,N_8518);
or U10344 (N_10344,N_9258,N_8654);
or U10345 (N_10345,N_8042,N_8270);
and U10346 (N_10346,N_8359,N_9374);
nand U10347 (N_10347,N_8608,N_8673);
nand U10348 (N_10348,N_9005,N_9168);
or U10349 (N_10349,N_8415,N_8022);
xnor U10350 (N_10350,N_8722,N_8292);
or U10351 (N_10351,N_9010,N_9451);
or U10352 (N_10352,N_7906,N_8798);
and U10353 (N_10353,N_9124,N_8674);
and U10354 (N_10354,N_8741,N_7521);
xnor U10355 (N_10355,N_8246,N_8357);
nand U10356 (N_10356,N_8024,N_8693);
xor U10357 (N_10357,N_9489,N_8148);
and U10358 (N_10358,N_8515,N_7797);
and U10359 (N_10359,N_9872,N_9884);
nand U10360 (N_10360,N_8696,N_9309);
nor U10361 (N_10361,N_7686,N_9704);
xor U10362 (N_10362,N_9922,N_8166);
xnor U10363 (N_10363,N_9864,N_9984);
xnor U10364 (N_10364,N_9900,N_8995);
or U10365 (N_10365,N_9307,N_9498);
nand U10366 (N_10366,N_9788,N_9927);
nand U10367 (N_10367,N_7879,N_7613);
nand U10368 (N_10368,N_8635,N_7791);
nor U10369 (N_10369,N_9294,N_8421);
nand U10370 (N_10370,N_9524,N_8094);
xnor U10371 (N_10371,N_7794,N_8458);
xor U10372 (N_10372,N_9490,N_8480);
nor U10373 (N_10373,N_7590,N_8874);
nand U10374 (N_10374,N_9431,N_8410);
and U10375 (N_10375,N_8336,N_8404);
nor U10376 (N_10376,N_9122,N_9909);
nand U10377 (N_10377,N_9455,N_8200);
or U10378 (N_10378,N_9822,N_9171);
and U10379 (N_10379,N_8210,N_9946);
and U10380 (N_10380,N_8477,N_9646);
xnor U10381 (N_10381,N_8597,N_9310);
nand U10382 (N_10382,N_9938,N_8773);
nor U10383 (N_10383,N_8905,N_9981);
xnor U10384 (N_10384,N_8046,N_8329);
or U10385 (N_10385,N_9810,N_9131);
xor U10386 (N_10386,N_7883,N_8379);
and U10387 (N_10387,N_7815,N_9242);
nand U10388 (N_10388,N_8261,N_9422);
and U10389 (N_10389,N_8311,N_8194);
nor U10390 (N_10390,N_8756,N_9673);
xnor U10391 (N_10391,N_8925,N_9492);
xnor U10392 (N_10392,N_7796,N_9176);
nor U10393 (N_10393,N_8163,N_7865);
xnor U10394 (N_10394,N_8144,N_9047);
xor U10395 (N_10395,N_8790,N_8370);
and U10396 (N_10396,N_7992,N_9863);
xnor U10397 (N_10397,N_9654,N_8562);
and U10398 (N_10398,N_8221,N_7930);
xor U10399 (N_10399,N_9153,N_8374);
nand U10400 (N_10400,N_8247,N_8445);
or U10401 (N_10401,N_8736,N_7768);
nor U10402 (N_10402,N_9144,N_8234);
or U10403 (N_10403,N_8272,N_9785);
nand U10404 (N_10404,N_8807,N_9630);
or U10405 (N_10405,N_8868,N_9907);
and U10406 (N_10406,N_9790,N_7595);
nor U10407 (N_10407,N_8082,N_9148);
or U10408 (N_10408,N_9465,N_9328);
xnor U10409 (N_10409,N_8780,N_9960);
and U10410 (N_10410,N_9416,N_8850);
xnor U10411 (N_10411,N_8295,N_8943);
or U10412 (N_10412,N_8853,N_9090);
nand U10413 (N_10413,N_7920,N_7903);
nand U10414 (N_10414,N_7511,N_9499);
nor U10415 (N_10415,N_8742,N_7630);
xor U10416 (N_10416,N_8842,N_7625);
nor U10417 (N_10417,N_9409,N_7623);
or U10418 (N_10418,N_7960,N_9928);
or U10419 (N_10419,N_7671,N_7679);
nand U10420 (N_10420,N_8475,N_8718);
nor U10421 (N_10421,N_8660,N_9060);
nor U10422 (N_10422,N_9136,N_9312);
nor U10423 (N_10423,N_8946,N_9276);
nor U10424 (N_10424,N_9908,N_9565);
nand U10425 (N_10425,N_8697,N_9635);
or U10426 (N_10426,N_8400,N_8936);
nor U10427 (N_10427,N_8708,N_7504);
xor U10428 (N_10428,N_9762,N_8974);
xnor U10429 (N_10429,N_8427,N_8712);
xor U10430 (N_10430,N_7598,N_8881);
nand U10431 (N_10431,N_9562,N_9728);
nor U10432 (N_10432,N_9548,N_8912);
and U10433 (N_10433,N_7657,N_7533);
nand U10434 (N_10434,N_7628,N_8864);
nand U10435 (N_10435,N_8921,N_9134);
xor U10436 (N_10436,N_9582,N_7571);
and U10437 (N_10437,N_9264,N_9318);
xor U10438 (N_10438,N_9435,N_9474);
xor U10439 (N_10439,N_8029,N_8390);
xor U10440 (N_10440,N_7582,N_7828);
nor U10441 (N_10441,N_7654,N_9306);
and U10442 (N_10442,N_8845,N_8730);
xor U10443 (N_10443,N_9194,N_8360);
nor U10444 (N_10444,N_8523,N_7530);
xor U10445 (N_10445,N_8378,N_7937);
nand U10446 (N_10446,N_9121,N_9325);
nor U10447 (N_10447,N_8438,N_8889);
nor U10448 (N_10448,N_8915,N_9016);
or U10449 (N_10449,N_9125,N_9525);
or U10450 (N_10450,N_7596,N_7725);
or U10451 (N_10451,N_8672,N_9190);
xnor U10452 (N_10452,N_7951,N_9392);
nand U10453 (N_10453,N_9061,N_9521);
xor U10454 (N_10454,N_7936,N_9494);
nand U10455 (N_10455,N_8814,N_7921);
or U10456 (N_10456,N_9600,N_7753);
nand U10457 (N_10457,N_8684,N_7800);
or U10458 (N_10458,N_7569,N_9811);
nor U10459 (N_10459,N_9605,N_8613);
or U10460 (N_10460,N_8732,N_8796);
nand U10461 (N_10461,N_7852,N_8840);
nand U10462 (N_10462,N_8688,N_9629);
and U10463 (N_10463,N_8279,N_7880);
or U10464 (N_10464,N_9384,N_7696);
or U10465 (N_10465,N_8262,N_7501);
nand U10466 (N_10466,N_7844,N_9719);
and U10467 (N_10467,N_9920,N_8937);
and U10468 (N_10468,N_9657,N_7819);
xnor U10469 (N_10469,N_9078,N_9533);
xor U10470 (N_10470,N_8951,N_7776);
nand U10471 (N_10471,N_8529,N_8642);
xor U10472 (N_10472,N_8011,N_9233);
nor U10473 (N_10473,N_8146,N_8396);
xnor U10474 (N_10474,N_7901,N_8102);
nand U10475 (N_10475,N_7616,N_9667);
nand U10476 (N_10476,N_7705,N_7714);
nor U10477 (N_10477,N_9848,N_8500);
nand U10478 (N_10478,N_8825,N_8531);
and U10479 (N_10479,N_7703,N_8450);
nor U10480 (N_10480,N_8079,N_7915);
or U10481 (N_10481,N_9127,N_8520);
nand U10482 (N_10482,N_8758,N_9520);
and U10483 (N_10483,N_7551,N_9712);
nand U10484 (N_10484,N_9931,N_8172);
nor U10485 (N_10485,N_9227,N_7977);
and U10486 (N_10486,N_9924,N_9816);
or U10487 (N_10487,N_8501,N_9829);
and U10488 (N_10488,N_8395,N_9001);
xor U10489 (N_10489,N_9551,N_9286);
xor U10490 (N_10490,N_8664,N_8574);
nor U10491 (N_10491,N_9866,N_9675);
nand U10492 (N_10492,N_9595,N_9632);
nor U10493 (N_10493,N_7829,N_8504);
or U10494 (N_10494,N_8129,N_9887);
or U10495 (N_10495,N_8197,N_9890);
and U10496 (N_10496,N_8170,N_9941);
nand U10497 (N_10497,N_9393,N_9385);
nor U10498 (N_10498,N_9365,N_8859);
nand U10499 (N_10499,N_8800,N_9768);
and U10500 (N_10500,N_7897,N_7956);
or U10501 (N_10501,N_8662,N_8788);
nand U10502 (N_10502,N_9323,N_7618);
nand U10503 (N_10503,N_9260,N_7854);
and U10504 (N_10504,N_9538,N_9270);
xnor U10505 (N_10505,N_8325,N_8762);
or U10506 (N_10506,N_8676,N_8312);
or U10507 (N_10507,N_7842,N_7990);
and U10508 (N_10508,N_9561,N_9226);
nand U10509 (N_10509,N_9837,N_9504);
nand U10510 (N_10510,N_8591,N_8668);
or U10511 (N_10511,N_9102,N_9008);
nor U10512 (N_10512,N_9532,N_8273);
and U10513 (N_10513,N_8291,N_7756);
nand U10514 (N_10514,N_8997,N_7687);
xnor U10515 (N_10515,N_7606,N_9590);
xnor U10516 (N_10516,N_8626,N_9961);
or U10517 (N_10517,N_8812,N_8871);
and U10518 (N_10518,N_9212,N_9070);
xnor U10519 (N_10519,N_9937,N_7949);
nand U10520 (N_10520,N_8982,N_9250);
and U10521 (N_10521,N_7525,N_7775);
xor U10522 (N_10522,N_8572,N_7841);
nand U10523 (N_10523,N_8968,N_9874);
and U10524 (N_10524,N_8373,N_8969);
nand U10525 (N_10525,N_9959,N_8074);
nor U10526 (N_10526,N_9714,N_9055);
nand U10527 (N_10527,N_7935,N_8764);
or U10528 (N_10528,N_7660,N_8222);
nor U10529 (N_10529,N_8407,N_8638);
or U10530 (N_10530,N_9777,N_9707);
nand U10531 (N_10531,N_9481,N_8152);
or U10532 (N_10532,N_8484,N_7708);
nand U10533 (N_10533,N_8496,N_8284);
nand U10534 (N_10534,N_9359,N_8028);
nor U10535 (N_10535,N_8403,N_9252);
nand U10536 (N_10536,N_9338,N_7987);
nor U10537 (N_10537,N_9738,N_8692);
xor U10538 (N_10538,N_8985,N_9321);
or U10539 (N_10539,N_9795,N_7827);
nand U10540 (N_10540,N_9019,N_8786);
or U10541 (N_10541,N_9881,N_9607);
nor U10542 (N_10542,N_7685,N_9549);
nor U10543 (N_10543,N_8923,N_8130);
and U10544 (N_10544,N_8468,N_8657);
or U10545 (N_10545,N_8533,N_7706);
and U10546 (N_10546,N_8408,N_7721);
nand U10547 (N_10547,N_8683,N_7537);
xnor U10548 (N_10548,N_8179,N_9147);
xor U10549 (N_10549,N_8648,N_8549);
and U10550 (N_10550,N_9615,N_9058);
nand U10551 (N_10551,N_9585,N_8149);
nand U10552 (N_10552,N_7933,N_8382);
nor U10553 (N_10553,N_8565,N_9085);
and U10554 (N_10554,N_8245,N_8766);
nor U10555 (N_10555,N_8389,N_9360);
nor U10556 (N_10556,N_8829,N_7514);
or U10557 (N_10557,N_9870,N_9119);
nor U10558 (N_10558,N_8123,N_7731);
or U10559 (N_10559,N_8104,N_8196);
nand U10560 (N_10560,N_9028,N_8461);
and U10561 (N_10561,N_8367,N_9668);
nor U10562 (N_10562,N_8615,N_8205);
nor U10563 (N_10563,N_9317,N_8811);
and U10564 (N_10564,N_9379,N_9782);
or U10565 (N_10565,N_8783,N_9401);
or U10566 (N_10566,N_8884,N_9876);
and U10567 (N_10567,N_8137,N_8409);
or U10568 (N_10568,N_9982,N_9089);
or U10569 (N_10569,N_9530,N_9145);
or U10570 (N_10570,N_9913,N_9821);
and U10571 (N_10571,N_8224,N_8571);
or U10572 (N_10572,N_9105,N_9236);
and U10573 (N_10573,N_9546,N_9026);
or U10574 (N_10574,N_9757,N_7873);
nor U10575 (N_10575,N_7759,N_8293);
nor U10576 (N_10576,N_8837,N_8237);
nand U10577 (N_10577,N_8686,N_7574);
and U10578 (N_10578,N_8636,N_8681);
or U10579 (N_10579,N_8641,N_7568);
and U10580 (N_10580,N_7583,N_8749);
xnor U10581 (N_10581,N_8019,N_9142);
nand U10582 (N_10582,N_9235,N_8035);
nand U10583 (N_10583,N_8142,N_9406);
xnor U10584 (N_10584,N_8314,N_7912);
xnor U10585 (N_10585,N_8256,N_7766);
nor U10586 (N_10586,N_9348,N_9378);
nor U10587 (N_10587,N_8970,N_8507);
and U10588 (N_10588,N_7682,N_8510);
nor U10589 (N_10589,N_9709,N_8502);
or U10590 (N_10590,N_9445,N_9859);
and U10591 (N_10591,N_9476,N_7946);
xor U10592 (N_10592,N_7757,N_8338);
or U10593 (N_10593,N_7727,N_9778);
nand U10594 (N_10594,N_8393,N_8268);
nand U10595 (N_10595,N_9347,N_8767);
xnor U10596 (N_10596,N_9839,N_9679);
nand U10597 (N_10597,N_8585,N_8700);
nor U10598 (N_10598,N_8021,N_7512);
or U10599 (N_10599,N_8182,N_7771);
or U10600 (N_10600,N_9311,N_8087);
nand U10601 (N_10601,N_8908,N_8709);
nor U10602 (N_10602,N_8191,N_7580);
or U10603 (N_10603,N_9661,N_8746);
xor U10604 (N_10604,N_7534,N_9508);
xnor U10605 (N_10605,N_8855,N_8494);
nand U10606 (N_10606,N_8134,N_8873);
and U10607 (N_10607,N_8983,N_7763);
xor U10608 (N_10608,N_7812,N_8174);
xor U10609 (N_10609,N_9603,N_8080);
nand U10610 (N_10610,N_8979,N_7955);
or U10611 (N_10611,N_9715,N_9536);
nand U10612 (N_10612,N_8363,N_9898);
and U10613 (N_10613,N_7991,N_7862);
and U10614 (N_10614,N_9361,N_9651);
xnor U10615 (N_10615,N_8633,N_9082);
nor U10616 (N_10616,N_8605,N_8795);
nand U10617 (N_10617,N_9267,N_9056);
xnor U10618 (N_10618,N_8044,N_8119);
or U10619 (N_10619,N_9364,N_8304);
and U10620 (N_10620,N_7986,N_9865);
xnor U10621 (N_10621,N_9172,N_9199);
and U10622 (N_10622,N_9617,N_9926);
xnor U10623 (N_10623,N_7545,N_8289);
or U10624 (N_10624,N_7564,N_8964);
xnor U10625 (N_10625,N_9693,N_7864);
or U10626 (N_10626,N_7900,N_8973);
or U10627 (N_10627,N_7848,N_7860);
xor U10628 (N_10628,N_8032,N_9040);
or U10629 (N_10629,N_7650,N_7953);
or U10630 (N_10630,N_7738,N_7516);
and U10631 (N_10631,N_8679,N_8867);
xor U10632 (N_10632,N_7894,N_8039);
and U10633 (N_10633,N_7742,N_9608);
or U10634 (N_10634,N_9696,N_8290);
xor U10635 (N_10635,N_8285,N_8506);
nand U10636 (N_10636,N_9483,N_7832);
nand U10637 (N_10637,N_8067,N_9203);
nand U10638 (N_10638,N_9817,N_8038);
or U10639 (N_10639,N_8875,N_7802);
nor U10640 (N_10640,N_9101,N_9116);
xor U10641 (N_10641,N_8914,N_9204);
or U10642 (N_10642,N_7874,N_7799);
xor U10643 (N_10643,N_8340,N_7523);
xnor U10644 (N_10644,N_9241,N_9748);
and U10645 (N_10645,N_9224,N_8300);
and U10646 (N_10646,N_7994,N_7716);
nand U10647 (N_10647,N_8202,N_9198);
or U10648 (N_10648,N_8385,N_7830);
or U10649 (N_10649,N_9814,N_9951);
nand U10650 (N_10650,N_7715,N_8264);
xor U10651 (N_10651,N_9861,N_8233);
nor U10652 (N_10652,N_8809,N_9175);
nor U10653 (N_10653,N_7818,N_8701);
nor U10654 (N_10654,N_9185,N_9251);
or U10655 (N_10655,N_8330,N_8353);
or U10656 (N_10656,N_9891,N_8326);
or U10657 (N_10657,N_9487,N_9313);
and U10658 (N_10658,N_9188,N_9046);
nand U10659 (N_10659,N_9831,N_7678);
xnor U10660 (N_10660,N_7863,N_7929);
xor U10661 (N_10661,N_8185,N_8669);
nor U10662 (N_10662,N_9570,N_8567);
xor U10663 (N_10663,N_8656,N_9330);
nor U10664 (N_10664,N_7765,N_7552);
nor U10665 (N_10665,N_8136,N_7943);
and U10666 (N_10666,N_9691,N_9457);
nand U10667 (N_10667,N_9274,N_8135);
nand U10668 (N_10668,N_8932,N_7764);
and U10669 (N_10669,N_8794,N_7602);
nor U10670 (N_10670,N_8131,N_7917);
or U10671 (N_10671,N_9682,N_7576);
nor U10672 (N_10672,N_9161,N_9210);
nor U10673 (N_10673,N_9735,N_8141);
nor U10674 (N_10674,N_9844,N_9281);
xnor U10675 (N_10675,N_9802,N_7734);
xnor U10676 (N_10676,N_7924,N_9287);
or U10677 (N_10677,N_7666,N_9072);
or U10678 (N_10678,N_8228,N_7588);
and U10679 (N_10679,N_9964,N_8425);
and U10680 (N_10680,N_7611,N_8980);
and U10681 (N_10681,N_8109,N_8838);
nand U10682 (N_10682,N_7554,N_9429);
nand U10683 (N_10683,N_8580,N_9051);
nor U10684 (N_10684,N_9713,N_9784);
nand U10685 (N_10685,N_9747,N_7770);
xnor U10686 (N_10686,N_7619,N_9149);
or U10687 (N_10687,N_9003,N_9945);
nor U10688 (N_10688,N_8545,N_9803);
nor U10689 (N_10689,N_8765,N_9302);
and U10690 (N_10690,N_7549,N_8516);
nor U10691 (N_10691,N_8097,N_8027);
xor U10692 (N_10692,N_7993,N_8834);
nand U10693 (N_10693,N_9358,N_8640);
xnor U10694 (N_10694,N_8248,N_8827);
and U10695 (N_10695,N_7909,N_8952);
nor U10696 (N_10696,N_8296,N_9014);
nand U10697 (N_10697,N_9606,N_9154);
nor U10698 (N_10698,N_8418,N_9746);
or U10699 (N_10699,N_8658,N_8121);
nor U10700 (N_10700,N_9195,N_8434);
nor U10701 (N_10701,N_8303,N_8625);
and U10702 (N_10702,N_8826,N_8180);
nand U10703 (N_10703,N_9095,N_9155);
nand U10704 (N_10704,N_9333,N_9464);
nor U10705 (N_10705,N_8014,N_7713);
xnor U10706 (N_10706,N_7913,N_9619);
nor U10707 (N_10707,N_9108,N_7877);
and U10708 (N_10708,N_9566,N_7601);
and U10709 (N_10709,N_9545,N_8754);
or U10710 (N_10710,N_9284,N_8577);
nor U10711 (N_10711,N_8017,N_7789);
or U10712 (N_10712,N_9372,N_9976);
nor U10713 (N_10713,N_9526,N_9394);
nand U10714 (N_10714,N_9472,N_8924);
xnor U10715 (N_10715,N_8031,N_7767);
and U10716 (N_10716,N_9918,N_9833);
and U10717 (N_10717,N_9634,N_8478);
nand U10718 (N_10718,N_9514,N_8843);
nor U10719 (N_10719,N_9703,N_7782);
or U10720 (N_10720,N_7888,N_9097);
and U10721 (N_10721,N_8140,N_9557);
nor U10722 (N_10722,N_7620,N_9732);
nand U10723 (N_10723,N_7761,N_9885);
and U10724 (N_10724,N_8792,N_9178);
nand U10725 (N_10725,N_9620,N_8715);
or U10726 (N_10726,N_8160,N_8007);
nand U10727 (N_10727,N_8977,N_9855);
nand U10728 (N_10728,N_8062,N_8064);
xor U10729 (N_10729,N_7640,N_7594);
and U10730 (N_10730,N_8368,N_9983);
nor U10731 (N_10731,N_9100,N_9977);
or U10732 (N_10732,N_8108,N_9547);
or U10733 (N_10733,N_8214,N_9444);
xor U10734 (N_10734,N_8323,N_9346);
and U10735 (N_10735,N_9787,N_9564);
or U10736 (N_10736,N_8092,N_9137);
nand U10737 (N_10737,N_8454,N_7839);
xor U10738 (N_10738,N_8877,N_9563);
nand U10739 (N_10739,N_9906,N_9141);
or U10740 (N_10740,N_8731,N_7667);
or U10741 (N_10741,N_9871,N_9598);
xnor U10742 (N_10742,N_9080,N_9766);
xor U10743 (N_10743,N_7996,N_8929);
and U10744 (N_10744,N_7923,N_7822);
and U10745 (N_10745,N_9860,N_8098);
xnor U10746 (N_10746,N_9759,N_7503);
or U10747 (N_10747,N_9006,N_8564);
nor U10748 (N_10748,N_8639,N_8217);
nor U10749 (N_10749,N_9045,N_8259);
xor U10750 (N_10750,N_9559,N_8614);
or U10751 (N_10751,N_7732,N_8249);
nand U10752 (N_10752,N_9191,N_7754);
nor U10753 (N_10753,N_7872,N_9807);
or U10754 (N_10754,N_8623,N_9858);
and U10755 (N_10755,N_9366,N_9622);
and U10756 (N_10756,N_8566,N_9044);
nor U10757 (N_10757,N_9382,N_8327);
xor U10758 (N_10758,N_8320,N_9544);
nand U10759 (N_10759,N_9843,N_8607);
nand U10760 (N_10760,N_8808,N_8828);
and U10761 (N_10761,N_8208,N_9152);
nand U10762 (N_10762,N_9478,N_7803);
nand U10763 (N_10763,N_8497,N_7612);
xor U10764 (N_10764,N_8276,N_9576);
and U10765 (N_10765,N_8653,N_7697);
nand U10766 (N_10766,N_8063,N_8621);
and U10767 (N_10767,N_7726,N_7572);
xor U10768 (N_10768,N_8093,N_9801);
nor U10769 (N_10769,N_7515,N_7656);
xnor U10770 (N_10770,N_9460,N_8159);
or U10771 (N_10771,N_7589,N_7540);
nor U10772 (N_10772,N_7733,N_8301);
xnor U10773 (N_10773,N_8645,N_7985);
xnor U10774 (N_10774,N_9179,N_8310);
and U10775 (N_10775,N_7592,N_8184);
and U10776 (N_10776,N_9601,N_7973);
or U10777 (N_10777,N_8917,N_9417);
xor U10778 (N_10778,N_8575,N_8976);
and U10779 (N_10779,N_7965,N_8113);
and U10780 (N_10780,N_8209,N_9660);
nor U10781 (N_10781,N_9238,N_8579);
and U10782 (N_10782,N_8526,N_8592);
xnor U10783 (N_10783,N_8628,N_8355);
nand U10784 (N_10784,N_8115,N_9025);
or U10785 (N_10785,N_8341,N_9944);
xor U10786 (N_10786,N_9965,N_9772);
nor U10787 (N_10787,N_9139,N_9000);
nor U10788 (N_10788,N_7621,N_8430);
and U10789 (N_10789,N_8963,N_8990);
or U10790 (N_10790,N_9683,N_8553);
or U10791 (N_10791,N_7600,N_9912);
nand U10792 (N_10792,N_9953,N_9295);
nor U10793 (N_10793,N_7783,N_8023);
nor U10794 (N_10794,N_9723,N_7680);
nand U10795 (N_10795,N_9695,N_8043);
nand U10796 (N_10796,N_9447,N_9240);
nor U10797 (N_10797,N_9626,N_9434);
nand U10798 (N_10798,N_7908,N_9639);
or U10799 (N_10799,N_8126,N_7969);
nand U10800 (N_10800,N_9727,N_7649);
and U10801 (N_10801,N_9031,N_9140);
nand U10802 (N_10802,N_7529,N_9308);
xnor U10803 (N_10803,N_8493,N_9411);
nor U10804 (N_10804,N_7780,N_7809);
nor U10805 (N_10805,N_8954,N_8803);
and U10806 (N_10806,N_9169,N_9736);
xor U10807 (N_10807,N_8522,N_8002);
and U10808 (N_10808,N_8959,N_8918);
or U10809 (N_10809,N_8435,N_9769);
nor U10810 (N_10810,N_7942,N_9609);
nand U10811 (N_10811,N_8206,N_9581);
and U10812 (N_10812,N_7505,N_9290);
and U10813 (N_10813,N_9022,N_9974);
nor U10814 (N_10814,N_8739,N_8058);
nor U10815 (N_10815,N_9020,N_7823);
or U10816 (N_10816,N_7945,N_7814);
xor U10817 (N_10817,N_9752,N_8106);
nor U10818 (N_10818,N_7850,N_7736);
or U10819 (N_10819,N_8429,N_8155);
and U10820 (N_10820,N_7553,N_8150);
and U10821 (N_10821,N_9027,N_8594);
nor U10822 (N_10822,N_7773,N_9373);
xnor U10823 (N_10823,N_7694,N_8599);
xor U10824 (N_10824,N_7607,N_7691);
nor U10825 (N_10825,N_8498,N_9949);
xnor U10826 (N_10826,N_8955,N_8519);
nor U10827 (N_10827,N_8911,N_9064);
xor U10828 (N_10828,N_7866,N_8958);
and U10829 (N_10829,N_7614,N_9694);
and U10830 (N_10830,N_9659,N_8286);
or U10831 (N_10831,N_7676,N_9329);
nand U10832 (N_10832,N_7966,N_7695);
xor U10833 (N_10833,N_8525,N_9237);
or U10834 (N_10834,N_9088,N_8537);
and U10835 (N_10835,N_9623,N_8685);
or U10836 (N_10836,N_7609,N_9515);
nor U10837 (N_10837,N_7831,N_9604);
nor U10838 (N_10838,N_8278,N_8861);
xor U10839 (N_10839,N_7626,N_8091);
nand U10840 (N_10840,N_8173,N_8053);
or U10841 (N_10841,N_7517,N_8548);
or U10842 (N_10842,N_8839,N_8059);
xnor U10843 (N_10843,N_9665,N_8682);
or U10844 (N_10844,N_9265,N_8847);
and U10845 (N_10845,N_9676,N_9128);
or U10846 (N_10846,N_7868,N_9701);
or U10847 (N_10847,N_9897,N_9717);
xnor U10848 (N_10848,N_8318,N_9315);
xor U10849 (N_10849,N_9656,N_9262);
or U10850 (N_10850,N_9987,N_8351);
xor U10851 (N_10851,N_9352,N_8177);
xnor U10852 (N_10852,N_9878,N_8145);
and U10853 (N_10853,N_9402,N_8713);
or U10854 (N_10854,N_7661,N_9862);
xnor U10855 (N_10855,N_8158,N_7875);
nand U10856 (N_10856,N_9729,N_7634);
nor U10857 (N_10857,N_7717,N_8089);
and U10858 (N_10858,N_7939,N_9032);
xor U10859 (N_10859,N_7826,N_8198);
or U10860 (N_10860,N_9223,N_8810);
nand U10861 (N_10861,N_7729,N_8678);
xnor U10862 (N_10862,N_9543,N_8446);
nor U10863 (N_10863,N_7690,N_8283);
nor U10864 (N_10864,N_8413,N_8153);
nor U10865 (N_10865,N_9698,N_8371);
or U10866 (N_10866,N_8213,N_9640);
and U10867 (N_10867,N_9914,N_8819);
and U10868 (N_10868,N_9278,N_9002);
xor U10869 (N_10869,N_9396,N_8573);
and U10870 (N_10870,N_9018,N_8112);
xnor U10871 (N_10871,N_7813,N_8223);
and U10872 (N_10872,N_8543,N_8559);
and U10873 (N_10873,N_8698,N_9511);
nor U10874 (N_10874,N_9650,N_8893);
nor U10875 (N_10875,N_9697,N_9796);
nor U10876 (N_10876,N_9114,N_8589);
nand U10877 (N_10877,N_9261,N_9202);
or U10878 (N_10878,N_9869,N_8465);
nor U10879 (N_10879,N_8128,N_9218);
and U10880 (N_10880,N_7644,N_9706);
or U10881 (N_10881,N_9009,N_9112);
xor U10882 (N_10882,N_8508,N_9893);
nor U10883 (N_10883,N_9503,N_8910);
nand U10884 (N_10884,N_7849,N_9789);
nand U10885 (N_10885,N_8907,N_8705);
xor U10886 (N_10886,N_8586,N_7597);
nor U10887 (N_10887,N_7658,N_9666);
and U10888 (N_10888,N_9092,N_7740);
xor U10889 (N_10889,N_8120,N_7968);
nand U10890 (N_10890,N_9739,N_7719);
and U10891 (N_10891,N_7790,N_9955);
nor U10892 (N_10892,N_8627,N_7712);
nand U10893 (N_10893,N_9275,N_8361);
and U10894 (N_10894,N_8294,N_9649);
and U10895 (N_10895,N_7881,N_8342);
nand U10896 (N_10896,N_8469,N_9111);
and U10897 (N_10897,N_8492,N_8544);
nor U10898 (N_10898,N_9423,N_9641);
xor U10899 (N_10899,N_7843,N_8836);
and U10900 (N_10900,N_9628,N_8902);
or U10901 (N_10901,N_7835,N_9929);
nand U10902 (N_10902,N_9644,N_7793);
or U10903 (N_10903,N_9932,N_8687);
nor U10904 (N_10904,N_8957,N_9574);
xnor U10905 (N_10905,N_9852,N_7807);
nand U10906 (N_10906,N_8737,N_9399);
or U10907 (N_10907,N_7591,N_9638);
and U10908 (N_10908,N_9245,N_8806);
or U10909 (N_10909,N_8212,N_8132);
or U10910 (N_10910,N_9388,N_8606);
xnor U10911 (N_10911,N_7652,N_9480);
nor U10912 (N_10912,N_7664,N_9334);
nor U10913 (N_10913,N_8412,N_9357);
nor U10914 (N_10914,N_7506,N_9988);
and U10915 (N_10915,N_7855,N_8225);
or U10916 (N_10916,N_9950,N_7976);
xor U10917 (N_10917,N_8634,N_7907);
nor U10918 (N_10918,N_8391,N_9527);
nor U10919 (N_10919,N_9718,N_9322);
and U10920 (N_10920,N_7811,N_9671);
nor U10921 (N_10921,N_9259,N_9542);
nor U10922 (N_10922,N_8903,N_8622);
nor U10923 (N_10923,N_7669,N_8644);
or U10924 (N_10924,N_9255,N_9107);
nor U10925 (N_10925,N_9798,N_8442);
nor U10926 (N_10926,N_9568,N_8354);
nor U10927 (N_10927,N_8047,N_9327);
and U10928 (N_10928,N_8081,N_8073);
nor U10929 (N_10929,N_8392,N_9303);
and U10930 (N_10930,N_8711,N_9916);
xor U10931 (N_10931,N_8782,N_9519);
or U10932 (N_10932,N_8277,N_8433);
xnor U10933 (N_10933,N_8269,N_8949);
nor U10934 (N_10934,N_9962,N_8984);
nand U10935 (N_10935,N_8219,N_8428);
nor U10936 (N_10936,N_8927,N_9996);
and U10937 (N_10937,N_7981,N_8818);
nor U10938 (N_10938,N_8076,N_7577);
or U10939 (N_10939,N_8055,N_9057);
nand U10940 (N_10940,N_9049,N_9680);
nand U10941 (N_10941,N_9463,N_8372);
nor U10942 (N_10942,N_7889,N_9461);
xnor U10943 (N_10943,N_8432,N_8996);
nor U10944 (N_10944,N_9724,N_8218);
nor U10945 (N_10945,N_8667,N_9781);
xnor U10946 (N_10946,N_8913,N_9578);
nand U10947 (N_10947,N_8020,N_9017);
nand U10948 (N_10948,N_9418,N_8308);
or U10949 (N_10949,N_8557,N_8547);
and U10950 (N_10950,N_8008,N_9367);
nand U10951 (N_10951,N_9793,N_9523);
or U10952 (N_10952,N_9299,N_8799);
or U10953 (N_10953,N_7882,N_8255);
or U10954 (N_10954,N_8193,N_9611);
and U10955 (N_10955,N_9500,N_8694);
nand U10956 (N_10956,N_9749,N_9246);
nand U10957 (N_10957,N_9117,N_7902);
and U10958 (N_10958,N_7837,N_8066);
nand U10959 (N_10959,N_8735,N_8824);
xor U10960 (N_10960,N_7931,N_8895);
nor U10961 (N_10961,N_7531,N_9170);
nand U10962 (N_10962,N_7751,N_7508);
nand U10963 (N_10963,N_8568,N_8876);
nor U10964 (N_10964,N_9674,N_7999);
xor U10965 (N_10965,N_8604,N_9669);
or U10966 (N_10966,N_9614,N_9113);
nand U10967 (N_10967,N_9231,N_9288);
and U10968 (N_10968,N_9991,N_8365);
or U10969 (N_10969,N_9268,N_9433);
xnor U10970 (N_10970,N_8822,N_8797);
and U10971 (N_10971,N_9375,N_9631);
or U10972 (N_10972,N_9688,N_9160);
nand U10973 (N_10973,N_8757,N_9126);
nand U10974 (N_10974,N_9882,N_9156);
xnor U10975 (N_10975,N_8781,N_9109);
nor U10976 (N_10976,N_8332,N_9104);
xnor U10977 (N_10977,N_7847,N_8896);
nand U10978 (N_10978,N_9254,N_7989);
or U10979 (N_10979,N_8335,N_9150);
or U10980 (N_10980,N_9956,N_8539);
xnor U10981 (N_10981,N_7631,N_8041);
and U10982 (N_10982,N_9351,N_9071);
nor U10983 (N_10983,N_9277,N_8729);
or U10984 (N_10984,N_8643,N_8538);
xnor U10985 (N_10985,N_9023,N_7557);
nand U10986 (N_10986,N_8162,N_8384);
xnor U10987 (N_10987,N_7651,N_7704);
nor U10988 (N_10988,N_9655,N_9039);
nand U10989 (N_10989,N_7861,N_8211);
nor U10990 (N_10990,N_9670,N_8851);
or U10991 (N_10991,N_8753,N_8854);
xor U10992 (N_10992,N_9298,N_7777);
xnor U10993 (N_10993,N_9189,N_8013);
or U10994 (N_10994,N_7593,N_7918);
nor U10995 (N_10995,N_7978,N_8009);
or U10996 (N_10996,N_9725,N_8298);
or U10997 (N_10997,N_9934,N_9933);
nor U10998 (N_10998,N_9518,N_8956);
xnor U10999 (N_10999,N_8056,N_8025);
xor U11000 (N_11000,N_9967,N_8398);
xor U11001 (N_11001,N_9337,N_9024);
nor U11002 (N_11002,N_7919,N_8369);
nand U11003 (N_11003,N_7938,N_9681);
or U11004 (N_11004,N_7895,N_9412);
xor U11005 (N_11005,N_8164,N_9637);
xor U11006 (N_11006,N_8618,N_7538);
or U11007 (N_11007,N_9939,N_8891);
nand U11008 (N_11008,N_8830,N_7693);
and U11009 (N_11009,N_7674,N_7752);
xor U11010 (N_11010,N_9905,N_7566);
or U11011 (N_11011,N_9834,N_9488);
nand U11012 (N_11012,N_8003,N_8088);
or U11013 (N_11013,N_9625,N_7760);
xor U11014 (N_11014,N_9436,N_8872);
xnor U11015 (N_11015,N_7548,N_8823);
or U11016 (N_11016,N_9692,N_8103);
nand U11017 (N_11017,N_8474,N_7941);
or U11018 (N_11018,N_9054,N_8343);
nand U11019 (N_11019,N_9452,N_9062);
nand U11020 (N_11020,N_9708,N_8751);
xnor U11021 (N_11021,N_9806,N_8663);
nor U11022 (N_11022,N_9850,N_9165);
xor U11023 (N_11023,N_9610,N_8988);
nor U11024 (N_11024,N_8253,N_9653);
nor U11025 (N_11025,N_8695,N_7558);
xnor U11026 (N_11026,N_8998,N_8931);
nand U11027 (N_11027,N_9059,N_8313);
and U11028 (N_11028,N_8883,N_8242);
nand U11029 (N_11029,N_7808,N_8563);
and U11030 (N_11030,N_8235,N_8981);
and U11031 (N_11031,N_7891,N_8068);
xor U11032 (N_11032,N_9684,N_8358);
nand U11033 (N_11033,N_7961,N_9292);
nand U11034 (N_11034,N_9947,N_9110);
xnor U11035 (N_11035,N_8422,N_9225);
and U11036 (N_11036,N_9174,N_9221);
and U11037 (N_11037,N_8505,N_9349);
and U11038 (N_11038,N_8250,N_9754);
nor U11039 (N_11039,N_8321,N_8381);
or U11040 (N_11040,N_7972,N_7979);
xnor U11041 (N_11041,N_9414,N_8099);
xor U11042 (N_11042,N_9331,N_9904);
or U11043 (N_11043,N_9919,N_9528);
nor U11044 (N_11044,N_7562,N_9390);
xor U11045 (N_11045,N_9539,N_7963);
nor U11046 (N_11046,N_7638,N_8890);
nand U11047 (N_11047,N_7510,N_9291);
xnor U11048 (N_11048,N_7787,N_7642);
or U11049 (N_11049,N_8297,N_9556);
nand U11050 (N_11050,N_8052,N_7710);
or U11051 (N_11051,N_8938,N_9720);
xor U11052 (N_11052,N_7741,N_8817);
nor U11053 (N_11053,N_9052,N_8167);
nand U11054 (N_11054,N_8820,N_9847);
or U11055 (N_11055,N_9815,N_8651);
nor U11056 (N_11056,N_8471,N_7675);
nor U11057 (N_11057,N_9700,N_9567);
nand U11058 (N_11058,N_8989,N_9479);
nand U11059 (N_11059,N_7856,N_8646);
and U11060 (N_11060,N_7535,N_7709);
nand U11061 (N_11061,N_9721,N_9426);
and U11062 (N_11062,N_8617,N_7542);
nor U11063 (N_11063,N_9840,N_9247);
nor U11064 (N_11064,N_7575,N_8230);
nand U11065 (N_11065,N_9099,N_9094);
nand U11066 (N_11066,N_8051,N_7513);
nor U11067 (N_11067,N_8587,N_9828);
nor U11068 (N_11068,N_7573,N_9192);
nor U11069 (N_11069,N_9037,N_9419);
xor U11070 (N_11070,N_9011,N_9805);
or U11071 (N_11071,N_9228,N_8216);
nand U11072 (N_11072,N_8452,N_9043);
nand U11073 (N_11073,N_8680,N_9132);
and U11074 (N_11074,N_8542,N_8541);
or U11075 (N_11075,N_9534,N_9280);
and U11076 (N_11076,N_9741,N_8778);
or U11077 (N_11077,N_9797,N_9537);
or U11078 (N_11078,N_9764,N_9731);
nand U11079 (N_11079,N_9980,N_7581);
xor U11080 (N_11080,N_9371,N_9397);
xor U11081 (N_11081,N_7629,N_8083);
or U11082 (N_11082,N_8802,N_9824);
nor U11083 (N_11083,N_9745,N_8251);
nand U11084 (N_11084,N_7817,N_9096);
nor U11085 (N_11085,N_9678,N_8388);
nor U11086 (N_11086,N_9076,N_9699);
xor U11087 (N_11087,N_7836,N_9986);
nand U11088 (N_11088,N_7570,N_7737);
nor U11089 (N_11089,N_9256,N_8975);
or U11090 (N_11090,N_9569,N_8793);
nor U11091 (N_11091,N_9636,N_9103);
xor U11092 (N_11092,N_8779,N_8260);
nand U11093 (N_11093,N_7536,N_9213);
xor U11094 (N_11094,N_9854,N_7997);
xnor U11095 (N_11095,N_9990,N_9825);
nor U11096 (N_11096,N_8944,N_9992);
nor U11097 (N_11097,N_8499,N_9486);
or U11098 (N_11098,N_8690,N_9400);
or U11099 (N_11099,N_7701,N_8760);
and U11100 (N_11100,N_8462,N_7748);
or U11101 (N_11101,N_8590,N_8101);
xnor U11102 (N_11102,N_9903,N_9597);
nand U11103 (N_11103,N_9448,N_9502);
xnor U11104 (N_11104,N_9041,N_7605);
nor U11105 (N_11105,N_9663,N_8972);
or U11106 (N_11106,N_9957,N_7700);
nor U11107 (N_11107,N_8467,N_8986);
or U11108 (N_11108,N_9473,N_7784);
xnor U11109 (N_11109,N_9326,N_7838);
or U11110 (N_11110,N_9133,N_9702);
or U11111 (N_11111,N_9826,N_7565);
xnor U11112 (N_11112,N_9686,N_8661);
or U11113 (N_11113,N_9042,N_8426);
nor U11114 (N_11114,N_9067,N_8772);
nor U11115 (N_11115,N_9029,N_7707);
xor U11116 (N_11116,N_8546,N_7840);
nor U11117 (N_11117,N_8168,N_7718);
nand U11118 (N_11118,N_9301,N_9593);
or U11119 (N_11119,N_8030,N_8987);
or U11120 (N_11120,N_8204,N_9138);
nand U11121 (N_11121,N_9901,N_7539);
nand U11122 (N_11122,N_9760,N_9377);
xnor U11123 (N_11123,N_8339,N_8894);
nor U11124 (N_11124,N_8816,N_7911);
and U11125 (N_11125,N_7546,N_9344);
xnor U11126 (N_11126,N_9084,N_8187);
or U11127 (N_11127,N_7702,N_7971);
and U11128 (N_11128,N_8282,N_7632);
nand U11129 (N_11129,N_9722,N_8582);
and U11130 (N_11130,N_7526,N_8215);
and U11131 (N_11131,N_8265,N_8463);
or U11132 (N_11132,N_7958,N_8488);
nand U11133 (N_11133,N_9368,N_7672);
nor U11134 (N_11134,N_9453,N_9363);
nand U11135 (N_11135,N_8616,N_9244);
nand U11136 (N_11136,N_9355,N_9197);
nor U11137 (N_11137,N_8670,N_7532);
nand U11138 (N_11138,N_7698,N_8900);
nand U11139 (N_11139,N_8744,N_7774);
nor U11140 (N_11140,N_8178,N_8107);
nor U11141 (N_11141,N_9689,N_8992);
and U11142 (N_11142,N_9808,N_7617);
nand U11143 (N_11143,N_9143,N_9091);
xnor U11144 (N_11144,N_9316,N_9602);
and U11145 (N_11145,N_8966,N_9074);
xnor U11146 (N_11146,N_9846,N_8551);
nor U11147 (N_11147,N_9206,N_7567);
xnor U11148 (N_11148,N_9989,N_8689);
nand U11149 (N_11149,N_9685,N_8583);
nand U11150 (N_11150,N_9771,N_8377);
or U11151 (N_11151,N_8555,N_7639);
xnor U11152 (N_11152,N_8199,N_9272);
or U11153 (N_11153,N_8331,N_7655);
nor U11154 (N_11154,N_8472,N_8495);
nor U11155 (N_11155,N_9081,N_8612);
and U11156 (N_11156,N_9320,N_8324);
xnor U11157 (N_11157,N_8457,N_9083);
nor U11158 (N_11158,N_9215,N_9579);
xor U11159 (N_11159,N_8271,N_9415);
or U11160 (N_11160,N_7778,N_8192);
or U11161 (N_11161,N_8534,N_9751);
nor U11162 (N_11162,N_9335,N_8804);
or U11163 (N_11163,N_9773,N_8005);
nand U11164 (N_11164,N_7692,N_9300);
xor U11165 (N_11165,N_9954,N_8630);
or U11166 (N_11166,N_7635,N_9482);
xnor U11167 (N_11167,N_8176,N_9845);
nand U11168 (N_11168,N_9410,N_9594);
or U11169 (N_11169,N_7887,N_9222);
nand U11170 (N_11170,N_8603,N_9462);
nand U11171 (N_11171,N_9779,N_8813);
xor U11172 (N_11172,N_8962,N_8632);
or U11173 (N_11173,N_8671,N_7772);
nor U11174 (N_11174,N_9442,N_8532);
nand U11175 (N_11175,N_8535,N_8420);
or U11176 (N_11176,N_7910,N_9740);
nand U11177 (N_11177,N_7785,N_9471);
nor U11178 (N_11178,N_7804,N_9033);
or U11179 (N_11179,N_9531,N_8866);
nor U11180 (N_11180,N_9744,N_8570);
or U11181 (N_11181,N_8252,N_7677);
xnor U11182 (N_11182,N_7927,N_9993);
and U11183 (N_11183,N_7518,N_8157);
and U11184 (N_11184,N_8232,N_9510);
nand U11185 (N_11185,N_9376,N_9849);
or U11186 (N_11186,N_9162,N_9123);
or U11187 (N_11187,N_8439,N_8257);
and U11188 (N_11188,N_8610,N_8849);
nand U11189 (N_11189,N_9273,N_8090);
xnor U11190 (N_11190,N_9985,N_8156);
xnor U11191 (N_11191,N_9181,N_9776);
nor U11192 (N_11192,N_9013,N_9343);
or U11193 (N_11193,N_9743,N_7845);
or U11194 (N_11194,N_8114,N_8601);
or U11195 (N_11195,N_8584,N_8581);
nor U11196 (N_11196,N_9786,N_7983);
nor U11197 (N_11197,N_8919,N_7641);
nor U11198 (N_11198,N_8207,N_7898);
nor U11199 (N_11199,N_7722,N_9438);
nor U11200 (N_11200,N_7871,N_8139);
and U11201 (N_11201,N_8305,N_9868);
or U11202 (N_11202,N_8556,N_7578);
xor U11203 (N_11203,N_7982,N_8719);
xnor U11204 (N_11204,N_9867,N_7974);
nor U11205 (N_11205,N_9560,N_8940);
nand U11206 (N_11206,N_9495,N_8831);
nand U11207 (N_11207,N_8356,N_8922);
nand U11208 (N_11208,N_9209,N_7899);
or U11209 (N_11209,N_8858,N_8993);
or U11210 (N_11210,N_8348,N_9509);
xor U11211 (N_11211,N_8309,N_8769);
nor U11212 (N_11212,N_8386,N_8771);
nand U11213 (N_11213,N_9936,N_8898);
or U11214 (N_11214,N_9403,N_8459);
xnor U11215 (N_11215,N_8346,N_7663);
and U11216 (N_11216,N_9015,N_9163);
xor U11217 (N_11217,N_8777,N_9324);
nor U11218 (N_11218,N_8001,N_9558);
nand U11219 (N_11219,N_9726,N_9930);
nor U11220 (N_11220,N_9484,N_9894);
or U11221 (N_11221,N_8220,N_9911);
or U11222 (N_11222,N_9591,N_9767);
xor U11223 (N_11223,N_7615,N_8865);
or U11224 (N_11224,N_9079,N_8350);
and U11225 (N_11225,N_7896,N_9710);
or U11226 (N_11226,N_9146,N_9513);
and U11227 (N_11227,N_9389,N_9342);
and U11228 (N_11228,N_8105,N_7904);
nand U11229 (N_11229,N_9216,N_8481);
nor U11230 (N_11230,N_7645,N_8483);
nand U11231 (N_11231,N_8733,N_9973);
or U11232 (N_11232,N_9086,N_7519);
xor U11233 (N_11233,N_9207,N_9522);
xor U11234 (N_11234,N_8060,N_8703);
nand U11235 (N_11235,N_7962,N_8302);
nor U11236 (N_11236,N_7988,N_7769);
nand U11237 (N_11237,N_9279,N_8460);
or U11238 (N_11238,N_9889,N_8994);
nand U11239 (N_11239,N_8453,N_8423);
or U11240 (N_11240,N_9830,N_9177);
xor U11241 (N_11241,N_9466,N_9193);
and U11242 (N_11242,N_9427,N_9217);
and U11243 (N_11243,N_9428,N_9968);
nor U11244 (N_11244,N_7559,N_8776);
nor U11245 (N_11245,N_9253,N_8920);
or U11246 (N_11246,N_8012,N_8748);
or U11247 (N_11247,N_8552,N_8909);
nand U11248 (N_11248,N_8111,N_8489);
or U11249 (N_11249,N_9838,N_7735);
or U11250 (N_11250,N_9729,N_9636);
or U11251 (N_11251,N_9030,N_9897);
xnor U11252 (N_11252,N_9803,N_9551);
nor U11253 (N_11253,N_8640,N_7756);
xnor U11254 (N_11254,N_8792,N_8510);
and U11255 (N_11255,N_8782,N_8001);
nor U11256 (N_11256,N_8686,N_9681);
nand U11257 (N_11257,N_9603,N_9918);
xor U11258 (N_11258,N_9583,N_7552);
xnor U11259 (N_11259,N_9909,N_9980);
and U11260 (N_11260,N_8400,N_8326);
and U11261 (N_11261,N_9733,N_9475);
or U11262 (N_11262,N_7737,N_7947);
and U11263 (N_11263,N_8579,N_7845);
nor U11264 (N_11264,N_8965,N_7786);
and U11265 (N_11265,N_8395,N_9804);
or U11266 (N_11266,N_9945,N_7736);
and U11267 (N_11267,N_7542,N_7802);
nor U11268 (N_11268,N_7571,N_9493);
nor U11269 (N_11269,N_8434,N_8178);
nand U11270 (N_11270,N_9764,N_9904);
nand U11271 (N_11271,N_9647,N_7511);
xor U11272 (N_11272,N_9342,N_8808);
and U11273 (N_11273,N_9903,N_8079);
nand U11274 (N_11274,N_7625,N_8583);
nor U11275 (N_11275,N_9806,N_7799);
nor U11276 (N_11276,N_8011,N_8013);
and U11277 (N_11277,N_9290,N_8654);
nand U11278 (N_11278,N_9945,N_9236);
xor U11279 (N_11279,N_9406,N_9045);
nand U11280 (N_11280,N_9231,N_8407);
nand U11281 (N_11281,N_8300,N_8735);
xnor U11282 (N_11282,N_8416,N_7867);
nor U11283 (N_11283,N_8196,N_8293);
xor U11284 (N_11284,N_9061,N_8449);
xnor U11285 (N_11285,N_7960,N_7544);
nand U11286 (N_11286,N_9745,N_9514);
nand U11287 (N_11287,N_9156,N_8756);
or U11288 (N_11288,N_8226,N_8374);
xor U11289 (N_11289,N_7607,N_8033);
nor U11290 (N_11290,N_9068,N_8266);
nor U11291 (N_11291,N_9360,N_8363);
or U11292 (N_11292,N_7712,N_9256);
nand U11293 (N_11293,N_9480,N_9785);
and U11294 (N_11294,N_8916,N_8566);
or U11295 (N_11295,N_8276,N_9228);
nand U11296 (N_11296,N_8420,N_8021);
nor U11297 (N_11297,N_8719,N_9655);
or U11298 (N_11298,N_9091,N_9881);
xnor U11299 (N_11299,N_8878,N_8315);
or U11300 (N_11300,N_7538,N_8809);
or U11301 (N_11301,N_8200,N_9704);
nor U11302 (N_11302,N_9939,N_9424);
or U11303 (N_11303,N_9288,N_8391);
and U11304 (N_11304,N_8068,N_8372);
or U11305 (N_11305,N_8523,N_8159);
or U11306 (N_11306,N_9855,N_8898);
or U11307 (N_11307,N_9925,N_8969);
xnor U11308 (N_11308,N_8732,N_9599);
nor U11309 (N_11309,N_8489,N_8281);
nand U11310 (N_11310,N_9198,N_9426);
nor U11311 (N_11311,N_8606,N_9310);
or U11312 (N_11312,N_9146,N_7628);
nor U11313 (N_11313,N_7604,N_9200);
or U11314 (N_11314,N_9637,N_9078);
nand U11315 (N_11315,N_8875,N_9155);
or U11316 (N_11316,N_9200,N_7733);
or U11317 (N_11317,N_9021,N_8749);
nor U11318 (N_11318,N_9940,N_8263);
or U11319 (N_11319,N_7750,N_9318);
or U11320 (N_11320,N_9918,N_8665);
or U11321 (N_11321,N_9943,N_8901);
and U11322 (N_11322,N_9192,N_9664);
and U11323 (N_11323,N_9452,N_8736);
xor U11324 (N_11324,N_9081,N_9643);
xnor U11325 (N_11325,N_8913,N_8395);
nand U11326 (N_11326,N_9859,N_7564);
xor U11327 (N_11327,N_8052,N_7622);
or U11328 (N_11328,N_9467,N_9654);
nor U11329 (N_11329,N_8847,N_8560);
nand U11330 (N_11330,N_9830,N_7712);
xnor U11331 (N_11331,N_8982,N_9468);
or U11332 (N_11332,N_9576,N_8195);
nor U11333 (N_11333,N_8754,N_8626);
and U11334 (N_11334,N_8802,N_9545);
xnor U11335 (N_11335,N_9665,N_9734);
nand U11336 (N_11336,N_8974,N_8164);
and U11337 (N_11337,N_9386,N_8756);
nor U11338 (N_11338,N_7715,N_8712);
nand U11339 (N_11339,N_9415,N_9128);
and U11340 (N_11340,N_7677,N_9744);
nor U11341 (N_11341,N_8942,N_9884);
or U11342 (N_11342,N_9150,N_7980);
xnor U11343 (N_11343,N_7720,N_8011);
nor U11344 (N_11344,N_8611,N_8262);
nand U11345 (N_11345,N_9232,N_8701);
nor U11346 (N_11346,N_7584,N_8481);
xor U11347 (N_11347,N_7509,N_9734);
nand U11348 (N_11348,N_9128,N_9409);
nand U11349 (N_11349,N_8294,N_8536);
and U11350 (N_11350,N_9227,N_8567);
nor U11351 (N_11351,N_9171,N_9979);
nor U11352 (N_11352,N_8099,N_9811);
or U11353 (N_11353,N_9713,N_9531);
and U11354 (N_11354,N_7907,N_8994);
nor U11355 (N_11355,N_8697,N_8750);
xnor U11356 (N_11356,N_8117,N_9426);
or U11357 (N_11357,N_7976,N_9807);
nor U11358 (N_11358,N_7960,N_8945);
and U11359 (N_11359,N_7793,N_9413);
or U11360 (N_11360,N_9824,N_8781);
xor U11361 (N_11361,N_7856,N_8690);
or U11362 (N_11362,N_9820,N_9717);
or U11363 (N_11363,N_8418,N_9754);
xnor U11364 (N_11364,N_7957,N_7597);
nand U11365 (N_11365,N_8120,N_8658);
nand U11366 (N_11366,N_7746,N_8646);
and U11367 (N_11367,N_9953,N_8212);
or U11368 (N_11368,N_9701,N_7980);
and U11369 (N_11369,N_8798,N_9260);
and U11370 (N_11370,N_8735,N_8463);
xnor U11371 (N_11371,N_9421,N_9149);
or U11372 (N_11372,N_9542,N_9912);
nand U11373 (N_11373,N_7572,N_8889);
nor U11374 (N_11374,N_9807,N_9562);
or U11375 (N_11375,N_8442,N_9820);
nor U11376 (N_11376,N_8803,N_8057);
nor U11377 (N_11377,N_7745,N_9324);
and U11378 (N_11378,N_9856,N_8360);
nand U11379 (N_11379,N_8720,N_9944);
xnor U11380 (N_11380,N_9054,N_9338);
xnor U11381 (N_11381,N_9766,N_8695);
xor U11382 (N_11382,N_9876,N_8719);
or U11383 (N_11383,N_9027,N_9675);
nor U11384 (N_11384,N_8558,N_9242);
nand U11385 (N_11385,N_9882,N_8921);
nor U11386 (N_11386,N_8077,N_8584);
nor U11387 (N_11387,N_8584,N_9420);
or U11388 (N_11388,N_8462,N_9949);
and U11389 (N_11389,N_9738,N_9706);
nor U11390 (N_11390,N_8685,N_8084);
nand U11391 (N_11391,N_8654,N_7786);
xor U11392 (N_11392,N_9069,N_8897);
xnor U11393 (N_11393,N_8142,N_9772);
nor U11394 (N_11394,N_9276,N_7562);
and U11395 (N_11395,N_7746,N_9318);
nor U11396 (N_11396,N_9722,N_7915);
and U11397 (N_11397,N_9974,N_8662);
nand U11398 (N_11398,N_8710,N_9168);
nand U11399 (N_11399,N_9362,N_9250);
or U11400 (N_11400,N_7997,N_8417);
nor U11401 (N_11401,N_9665,N_8573);
nor U11402 (N_11402,N_9402,N_8432);
and U11403 (N_11403,N_9920,N_8719);
nand U11404 (N_11404,N_8966,N_9490);
and U11405 (N_11405,N_9379,N_7578);
or U11406 (N_11406,N_8612,N_8216);
or U11407 (N_11407,N_9458,N_9298);
nor U11408 (N_11408,N_9900,N_7804);
xor U11409 (N_11409,N_9104,N_8339);
and U11410 (N_11410,N_8326,N_9990);
and U11411 (N_11411,N_9953,N_9253);
and U11412 (N_11412,N_8027,N_9483);
or U11413 (N_11413,N_8780,N_8753);
nor U11414 (N_11414,N_7545,N_8399);
nand U11415 (N_11415,N_8534,N_7866);
nor U11416 (N_11416,N_9052,N_7866);
or U11417 (N_11417,N_8636,N_7675);
nand U11418 (N_11418,N_7861,N_9663);
nor U11419 (N_11419,N_9457,N_7787);
and U11420 (N_11420,N_8328,N_8896);
and U11421 (N_11421,N_8869,N_8024);
xor U11422 (N_11422,N_7812,N_7529);
and U11423 (N_11423,N_8251,N_8096);
and U11424 (N_11424,N_9507,N_8605);
and U11425 (N_11425,N_8983,N_8813);
xor U11426 (N_11426,N_7709,N_7995);
or U11427 (N_11427,N_9497,N_8096);
xnor U11428 (N_11428,N_7893,N_9099);
xor U11429 (N_11429,N_9377,N_7714);
nor U11430 (N_11430,N_9805,N_8626);
nand U11431 (N_11431,N_9981,N_9214);
nor U11432 (N_11432,N_9971,N_8225);
nor U11433 (N_11433,N_8028,N_9305);
or U11434 (N_11434,N_8216,N_7888);
xnor U11435 (N_11435,N_9468,N_9162);
or U11436 (N_11436,N_7728,N_9110);
nand U11437 (N_11437,N_8249,N_9405);
nor U11438 (N_11438,N_9773,N_9920);
xor U11439 (N_11439,N_8953,N_9429);
nor U11440 (N_11440,N_9912,N_9046);
xor U11441 (N_11441,N_8164,N_9766);
and U11442 (N_11442,N_9732,N_9831);
or U11443 (N_11443,N_9449,N_8477);
xor U11444 (N_11444,N_9445,N_8553);
nor U11445 (N_11445,N_8717,N_9227);
xor U11446 (N_11446,N_8411,N_7784);
nor U11447 (N_11447,N_7896,N_8174);
nand U11448 (N_11448,N_7834,N_8524);
nand U11449 (N_11449,N_9698,N_9618);
or U11450 (N_11450,N_8561,N_7981);
nor U11451 (N_11451,N_9778,N_9531);
xnor U11452 (N_11452,N_7872,N_8145);
or U11453 (N_11453,N_8146,N_7646);
or U11454 (N_11454,N_7535,N_7821);
nand U11455 (N_11455,N_9179,N_9424);
nor U11456 (N_11456,N_7503,N_8484);
xnor U11457 (N_11457,N_8436,N_7765);
nor U11458 (N_11458,N_9381,N_7955);
and U11459 (N_11459,N_9159,N_8252);
xnor U11460 (N_11460,N_9064,N_9176);
and U11461 (N_11461,N_9309,N_8441);
nor U11462 (N_11462,N_8646,N_8846);
xnor U11463 (N_11463,N_9744,N_9885);
nor U11464 (N_11464,N_9207,N_7731);
nor U11465 (N_11465,N_9269,N_9573);
nand U11466 (N_11466,N_8955,N_9926);
and U11467 (N_11467,N_8389,N_9365);
or U11468 (N_11468,N_8309,N_8465);
or U11469 (N_11469,N_9737,N_8694);
nand U11470 (N_11470,N_8843,N_9354);
xnor U11471 (N_11471,N_9037,N_8884);
or U11472 (N_11472,N_8340,N_7759);
nand U11473 (N_11473,N_8228,N_9054);
or U11474 (N_11474,N_9496,N_9661);
xor U11475 (N_11475,N_7736,N_9311);
and U11476 (N_11476,N_9205,N_9167);
or U11477 (N_11477,N_8668,N_7653);
and U11478 (N_11478,N_9430,N_9771);
nor U11479 (N_11479,N_8924,N_8076);
nor U11480 (N_11480,N_8690,N_7799);
and U11481 (N_11481,N_8475,N_8764);
xnor U11482 (N_11482,N_9080,N_7540);
and U11483 (N_11483,N_7936,N_8513);
xor U11484 (N_11484,N_8639,N_9493);
nand U11485 (N_11485,N_7913,N_8702);
and U11486 (N_11486,N_9169,N_9945);
nand U11487 (N_11487,N_8261,N_9552);
nor U11488 (N_11488,N_9709,N_9474);
nand U11489 (N_11489,N_8196,N_8789);
nand U11490 (N_11490,N_8052,N_9970);
nor U11491 (N_11491,N_8102,N_9564);
or U11492 (N_11492,N_7929,N_9959);
and U11493 (N_11493,N_9645,N_8498);
nand U11494 (N_11494,N_9615,N_9931);
nor U11495 (N_11495,N_9651,N_9329);
or U11496 (N_11496,N_8623,N_9435);
nand U11497 (N_11497,N_8414,N_7814);
or U11498 (N_11498,N_8655,N_7986);
xnor U11499 (N_11499,N_9198,N_9048);
nor U11500 (N_11500,N_9193,N_7879);
or U11501 (N_11501,N_8780,N_9224);
or U11502 (N_11502,N_9699,N_9206);
nor U11503 (N_11503,N_7571,N_8648);
nand U11504 (N_11504,N_9833,N_7694);
nand U11505 (N_11505,N_8803,N_9383);
nor U11506 (N_11506,N_8540,N_8682);
nand U11507 (N_11507,N_8274,N_7854);
or U11508 (N_11508,N_8104,N_8578);
nand U11509 (N_11509,N_8046,N_7921);
and U11510 (N_11510,N_7519,N_7728);
and U11511 (N_11511,N_9162,N_7840);
xor U11512 (N_11512,N_7960,N_8244);
xor U11513 (N_11513,N_9715,N_9721);
or U11514 (N_11514,N_9654,N_8382);
nand U11515 (N_11515,N_8985,N_9644);
nor U11516 (N_11516,N_7846,N_7694);
xor U11517 (N_11517,N_8764,N_9790);
and U11518 (N_11518,N_9415,N_8452);
nand U11519 (N_11519,N_9486,N_9057);
nand U11520 (N_11520,N_9895,N_8144);
or U11521 (N_11521,N_9915,N_9591);
and U11522 (N_11522,N_9697,N_9936);
nand U11523 (N_11523,N_9103,N_7975);
nand U11524 (N_11524,N_8184,N_9842);
nand U11525 (N_11525,N_9236,N_8087);
nor U11526 (N_11526,N_7919,N_8619);
nand U11527 (N_11527,N_9990,N_8501);
xor U11528 (N_11528,N_8373,N_8231);
and U11529 (N_11529,N_8924,N_9399);
and U11530 (N_11530,N_8050,N_8430);
or U11531 (N_11531,N_8259,N_7944);
or U11532 (N_11532,N_9638,N_8592);
and U11533 (N_11533,N_7897,N_7570);
nor U11534 (N_11534,N_7871,N_8177);
or U11535 (N_11535,N_8338,N_9213);
xnor U11536 (N_11536,N_9011,N_8375);
and U11537 (N_11537,N_8608,N_9529);
xnor U11538 (N_11538,N_9979,N_7948);
and U11539 (N_11539,N_9409,N_7673);
nor U11540 (N_11540,N_9079,N_9834);
and U11541 (N_11541,N_9354,N_7552);
and U11542 (N_11542,N_9156,N_7917);
and U11543 (N_11543,N_9611,N_9686);
and U11544 (N_11544,N_8327,N_9685);
nand U11545 (N_11545,N_8663,N_7786);
or U11546 (N_11546,N_7834,N_8079);
xor U11547 (N_11547,N_8343,N_7890);
xor U11548 (N_11548,N_7818,N_8480);
nor U11549 (N_11549,N_9297,N_9634);
xor U11550 (N_11550,N_8796,N_8221);
or U11551 (N_11551,N_9135,N_9632);
nor U11552 (N_11552,N_7679,N_8785);
xor U11553 (N_11553,N_8127,N_9535);
xnor U11554 (N_11554,N_9645,N_8912);
nand U11555 (N_11555,N_8107,N_8893);
and U11556 (N_11556,N_9524,N_9642);
and U11557 (N_11557,N_8660,N_8890);
xnor U11558 (N_11558,N_8091,N_8239);
or U11559 (N_11559,N_7621,N_9375);
nand U11560 (N_11560,N_8142,N_9147);
nand U11561 (N_11561,N_8404,N_7666);
or U11562 (N_11562,N_8094,N_9041);
nor U11563 (N_11563,N_8091,N_9069);
and U11564 (N_11564,N_7760,N_9165);
xnor U11565 (N_11565,N_9856,N_9133);
and U11566 (N_11566,N_9604,N_8557);
nor U11567 (N_11567,N_9688,N_8857);
nand U11568 (N_11568,N_8634,N_7729);
nor U11569 (N_11569,N_7694,N_7650);
nor U11570 (N_11570,N_8501,N_7957);
nand U11571 (N_11571,N_8033,N_8799);
nand U11572 (N_11572,N_7671,N_9665);
nand U11573 (N_11573,N_9079,N_9951);
or U11574 (N_11574,N_9160,N_8069);
nor U11575 (N_11575,N_7606,N_9756);
or U11576 (N_11576,N_9038,N_9326);
or U11577 (N_11577,N_9513,N_8112);
or U11578 (N_11578,N_8615,N_8827);
xnor U11579 (N_11579,N_9446,N_7847);
and U11580 (N_11580,N_9085,N_8861);
and U11581 (N_11581,N_7525,N_7532);
and U11582 (N_11582,N_8252,N_7619);
and U11583 (N_11583,N_8047,N_8443);
xor U11584 (N_11584,N_8982,N_8357);
or U11585 (N_11585,N_9489,N_7534);
nor U11586 (N_11586,N_8079,N_9184);
nor U11587 (N_11587,N_9372,N_8645);
nand U11588 (N_11588,N_9871,N_8291);
xnor U11589 (N_11589,N_9163,N_7891);
xnor U11590 (N_11590,N_9291,N_8156);
xor U11591 (N_11591,N_8421,N_9233);
nor U11592 (N_11592,N_9403,N_7971);
and U11593 (N_11593,N_9844,N_9532);
nand U11594 (N_11594,N_8255,N_9205);
xor U11595 (N_11595,N_9583,N_8924);
nor U11596 (N_11596,N_7666,N_9516);
or U11597 (N_11597,N_7578,N_7995);
nand U11598 (N_11598,N_7705,N_7911);
nand U11599 (N_11599,N_8808,N_9639);
nor U11600 (N_11600,N_8788,N_7759);
or U11601 (N_11601,N_8084,N_9028);
xnor U11602 (N_11602,N_7725,N_9321);
nand U11603 (N_11603,N_8152,N_8510);
or U11604 (N_11604,N_9518,N_8971);
nor U11605 (N_11605,N_8806,N_8368);
nand U11606 (N_11606,N_9804,N_8510);
nand U11607 (N_11607,N_8909,N_7653);
nor U11608 (N_11608,N_7724,N_7520);
or U11609 (N_11609,N_9922,N_9198);
xor U11610 (N_11610,N_7698,N_8583);
nand U11611 (N_11611,N_7840,N_9909);
and U11612 (N_11612,N_8310,N_7979);
xor U11613 (N_11613,N_9696,N_9669);
and U11614 (N_11614,N_9982,N_8475);
xnor U11615 (N_11615,N_9297,N_7688);
nand U11616 (N_11616,N_9389,N_9904);
xor U11617 (N_11617,N_9698,N_9208);
or U11618 (N_11618,N_7736,N_8663);
or U11619 (N_11619,N_9698,N_9892);
or U11620 (N_11620,N_7943,N_8703);
or U11621 (N_11621,N_7898,N_7537);
nor U11622 (N_11622,N_9224,N_9358);
and U11623 (N_11623,N_9525,N_9798);
nand U11624 (N_11624,N_8125,N_8211);
and U11625 (N_11625,N_9341,N_7904);
xor U11626 (N_11626,N_9897,N_7689);
nand U11627 (N_11627,N_9011,N_8111);
xor U11628 (N_11628,N_8429,N_8763);
and U11629 (N_11629,N_9027,N_8783);
and U11630 (N_11630,N_9306,N_9702);
nand U11631 (N_11631,N_8969,N_8595);
nand U11632 (N_11632,N_9952,N_7893);
xor U11633 (N_11633,N_8826,N_9788);
nor U11634 (N_11634,N_8771,N_9220);
xor U11635 (N_11635,N_9565,N_7854);
and U11636 (N_11636,N_7770,N_9945);
or U11637 (N_11637,N_8622,N_9719);
nand U11638 (N_11638,N_9545,N_8521);
or U11639 (N_11639,N_9654,N_8241);
and U11640 (N_11640,N_8753,N_8757);
nand U11641 (N_11641,N_8579,N_7748);
and U11642 (N_11642,N_9131,N_8927);
nand U11643 (N_11643,N_8809,N_9903);
nand U11644 (N_11644,N_7875,N_7764);
nand U11645 (N_11645,N_8913,N_8381);
xnor U11646 (N_11646,N_9480,N_9969);
xor U11647 (N_11647,N_8004,N_8086);
xnor U11648 (N_11648,N_9495,N_8651);
xor U11649 (N_11649,N_8231,N_8701);
and U11650 (N_11650,N_8517,N_9585);
or U11651 (N_11651,N_9360,N_8731);
nand U11652 (N_11652,N_8139,N_8880);
or U11653 (N_11653,N_8511,N_8976);
and U11654 (N_11654,N_8146,N_8051);
or U11655 (N_11655,N_9079,N_9798);
xnor U11656 (N_11656,N_8705,N_9389);
or U11657 (N_11657,N_7673,N_8856);
xor U11658 (N_11658,N_8973,N_9933);
nand U11659 (N_11659,N_8962,N_8344);
xnor U11660 (N_11660,N_8127,N_7701);
xor U11661 (N_11661,N_9633,N_7517);
xor U11662 (N_11662,N_8089,N_7706);
nor U11663 (N_11663,N_9313,N_8468);
or U11664 (N_11664,N_9245,N_7790);
and U11665 (N_11665,N_7921,N_9283);
nand U11666 (N_11666,N_9248,N_8406);
nand U11667 (N_11667,N_9287,N_8389);
or U11668 (N_11668,N_9082,N_8156);
nand U11669 (N_11669,N_9185,N_8625);
or U11670 (N_11670,N_8537,N_9467);
xnor U11671 (N_11671,N_8511,N_9076);
xnor U11672 (N_11672,N_9481,N_9179);
xnor U11673 (N_11673,N_8085,N_8089);
or U11674 (N_11674,N_8246,N_9099);
nand U11675 (N_11675,N_7954,N_8229);
xor U11676 (N_11676,N_9420,N_9587);
and U11677 (N_11677,N_9901,N_9208);
and U11678 (N_11678,N_7945,N_9521);
and U11679 (N_11679,N_8941,N_8176);
xnor U11680 (N_11680,N_9251,N_8436);
nand U11681 (N_11681,N_8382,N_7603);
nor U11682 (N_11682,N_9252,N_8012);
xor U11683 (N_11683,N_7999,N_8778);
nand U11684 (N_11684,N_8364,N_8391);
or U11685 (N_11685,N_8926,N_9282);
nor U11686 (N_11686,N_8591,N_9328);
xor U11687 (N_11687,N_8096,N_8402);
nand U11688 (N_11688,N_9256,N_9852);
or U11689 (N_11689,N_8422,N_8077);
nand U11690 (N_11690,N_9550,N_8831);
or U11691 (N_11691,N_8223,N_9590);
nand U11692 (N_11692,N_8148,N_8759);
or U11693 (N_11693,N_7941,N_8713);
nor U11694 (N_11694,N_8133,N_9442);
nor U11695 (N_11695,N_9168,N_8072);
or U11696 (N_11696,N_8707,N_8481);
nor U11697 (N_11697,N_8935,N_8844);
xor U11698 (N_11698,N_9925,N_8538);
xnor U11699 (N_11699,N_7668,N_8526);
xor U11700 (N_11700,N_8903,N_9079);
or U11701 (N_11701,N_9719,N_8666);
or U11702 (N_11702,N_9046,N_7644);
xnor U11703 (N_11703,N_8336,N_9254);
or U11704 (N_11704,N_7998,N_9880);
nand U11705 (N_11705,N_8822,N_9544);
or U11706 (N_11706,N_9999,N_9022);
nor U11707 (N_11707,N_8604,N_8755);
nor U11708 (N_11708,N_8696,N_8305);
or U11709 (N_11709,N_9622,N_9520);
nor U11710 (N_11710,N_9371,N_7763);
and U11711 (N_11711,N_9292,N_8402);
nand U11712 (N_11712,N_8516,N_8519);
or U11713 (N_11713,N_9989,N_9142);
nand U11714 (N_11714,N_9818,N_8827);
nand U11715 (N_11715,N_8356,N_8322);
xnor U11716 (N_11716,N_9972,N_9142);
nor U11717 (N_11717,N_7993,N_9935);
or U11718 (N_11718,N_9773,N_9972);
nor U11719 (N_11719,N_8040,N_8809);
xnor U11720 (N_11720,N_9551,N_7594);
or U11721 (N_11721,N_7741,N_9297);
and U11722 (N_11722,N_8015,N_7597);
and U11723 (N_11723,N_7783,N_7690);
nor U11724 (N_11724,N_9135,N_9330);
nor U11725 (N_11725,N_7753,N_8028);
nand U11726 (N_11726,N_9607,N_8136);
xnor U11727 (N_11727,N_9821,N_8530);
or U11728 (N_11728,N_7510,N_8110);
and U11729 (N_11729,N_7940,N_9163);
and U11730 (N_11730,N_8671,N_9108);
nor U11731 (N_11731,N_7623,N_8245);
nand U11732 (N_11732,N_8547,N_8066);
nor U11733 (N_11733,N_8471,N_8498);
nor U11734 (N_11734,N_8588,N_7735);
and U11735 (N_11735,N_7959,N_8065);
or U11736 (N_11736,N_9396,N_8270);
and U11737 (N_11737,N_8145,N_8752);
xnor U11738 (N_11738,N_8939,N_8492);
nor U11739 (N_11739,N_7686,N_9027);
nor U11740 (N_11740,N_9594,N_7685);
xnor U11741 (N_11741,N_8296,N_9513);
or U11742 (N_11742,N_7550,N_8838);
xnor U11743 (N_11743,N_8811,N_8363);
xor U11744 (N_11744,N_8659,N_8692);
nand U11745 (N_11745,N_9235,N_9625);
xnor U11746 (N_11746,N_8843,N_7648);
xor U11747 (N_11747,N_8314,N_9589);
and U11748 (N_11748,N_7755,N_9461);
and U11749 (N_11749,N_8671,N_9555);
nand U11750 (N_11750,N_8456,N_7774);
nand U11751 (N_11751,N_7946,N_8727);
nand U11752 (N_11752,N_8585,N_9598);
or U11753 (N_11753,N_9669,N_8431);
nor U11754 (N_11754,N_8271,N_8763);
nand U11755 (N_11755,N_8896,N_8726);
nor U11756 (N_11756,N_8561,N_7720);
and U11757 (N_11757,N_9659,N_9690);
nor U11758 (N_11758,N_8254,N_8073);
or U11759 (N_11759,N_9313,N_8025);
and U11760 (N_11760,N_9290,N_7757);
nand U11761 (N_11761,N_7963,N_9991);
xor U11762 (N_11762,N_9512,N_9710);
nand U11763 (N_11763,N_8762,N_9403);
xnor U11764 (N_11764,N_8298,N_7652);
and U11765 (N_11765,N_8062,N_9011);
and U11766 (N_11766,N_8209,N_8559);
or U11767 (N_11767,N_8721,N_8649);
nor U11768 (N_11768,N_8941,N_9936);
xor U11769 (N_11769,N_9838,N_8333);
xnor U11770 (N_11770,N_7644,N_7797);
nor U11771 (N_11771,N_8545,N_9490);
and U11772 (N_11772,N_9450,N_7612);
nor U11773 (N_11773,N_9914,N_8257);
or U11774 (N_11774,N_8181,N_8978);
and U11775 (N_11775,N_9227,N_8954);
nor U11776 (N_11776,N_9543,N_8400);
and U11777 (N_11777,N_8651,N_9977);
nand U11778 (N_11778,N_8147,N_8085);
nand U11779 (N_11779,N_8662,N_9114);
nor U11780 (N_11780,N_8116,N_8585);
nand U11781 (N_11781,N_9088,N_8807);
xnor U11782 (N_11782,N_8696,N_8809);
nor U11783 (N_11783,N_9059,N_8178);
or U11784 (N_11784,N_9214,N_9548);
xor U11785 (N_11785,N_9260,N_9038);
nor U11786 (N_11786,N_8544,N_9779);
and U11787 (N_11787,N_7660,N_9284);
xnor U11788 (N_11788,N_9547,N_8783);
and U11789 (N_11789,N_8826,N_9398);
nand U11790 (N_11790,N_8381,N_8498);
nand U11791 (N_11791,N_8525,N_8605);
nand U11792 (N_11792,N_9246,N_7759);
and U11793 (N_11793,N_9740,N_8721);
and U11794 (N_11794,N_9689,N_8525);
and U11795 (N_11795,N_7647,N_8218);
nand U11796 (N_11796,N_9482,N_7906);
and U11797 (N_11797,N_7502,N_8815);
nand U11798 (N_11798,N_8362,N_7940);
nand U11799 (N_11799,N_9255,N_7780);
xnor U11800 (N_11800,N_9915,N_8778);
nor U11801 (N_11801,N_7611,N_9320);
nor U11802 (N_11802,N_9179,N_9125);
or U11803 (N_11803,N_9682,N_8648);
and U11804 (N_11804,N_9054,N_8530);
nor U11805 (N_11805,N_8932,N_8315);
nor U11806 (N_11806,N_8655,N_9112);
nand U11807 (N_11807,N_9239,N_7662);
xnor U11808 (N_11808,N_9447,N_7641);
xnor U11809 (N_11809,N_8503,N_7579);
nor U11810 (N_11810,N_7927,N_9458);
or U11811 (N_11811,N_9113,N_7746);
xnor U11812 (N_11812,N_8671,N_9944);
nand U11813 (N_11813,N_9556,N_9456);
or U11814 (N_11814,N_9105,N_8342);
and U11815 (N_11815,N_7607,N_8441);
and U11816 (N_11816,N_7940,N_7702);
xor U11817 (N_11817,N_9356,N_8437);
or U11818 (N_11818,N_9328,N_8794);
nand U11819 (N_11819,N_7864,N_7580);
or U11820 (N_11820,N_8945,N_8088);
xor U11821 (N_11821,N_8140,N_7948);
and U11822 (N_11822,N_7687,N_9615);
and U11823 (N_11823,N_7687,N_9207);
nand U11824 (N_11824,N_8605,N_9070);
and U11825 (N_11825,N_9241,N_9036);
and U11826 (N_11826,N_8474,N_8036);
nand U11827 (N_11827,N_8927,N_7703);
or U11828 (N_11828,N_9752,N_8844);
nor U11829 (N_11829,N_9567,N_8532);
or U11830 (N_11830,N_7709,N_8613);
nor U11831 (N_11831,N_8740,N_7540);
or U11832 (N_11832,N_8140,N_8506);
xor U11833 (N_11833,N_8645,N_8303);
xnor U11834 (N_11834,N_8909,N_9721);
nor U11835 (N_11835,N_7960,N_9349);
nand U11836 (N_11836,N_8208,N_9052);
or U11837 (N_11837,N_9528,N_9699);
or U11838 (N_11838,N_9453,N_8502);
xnor U11839 (N_11839,N_8890,N_9556);
xor U11840 (N_11840,N_7686,N_7694);
xnor U11841 (N_11841,N_8077,N_7598);
or U11842 (N_11842,N_8903,N_8890);
and U11843 (N_11843,N_9225,N_7524);
and U11844 (N_11844,N_8456,N_7745);
or U11845 (N_11845,N_8172,N_8214);
or U11846 (N_11846,N_7663,N_8789);
xnor U11847 (N_11847,N_9723,N_9882);
or U11848 (N_11848,N_8386,N_8068);
xor U11849 (N_11849,N_9366,N_9027);
nor U11850 (N_11850,N_8718,N_8266);
nor U11851 (N_11851,N_9164,N_7949);
nor U11852 (N_11852,N_7971,N_9018);
xnor U11853 (N_11853,N_9583,N_8974);
and U11854 (N_11854,N_9418,N_9760);
nand U11855 (N_11855,N_9749,N_9614);
xor U11856 (N_11856,N_7787,N_8052);
or U11857 (N_11857,N_9008,N_8539);
nand U11858 (N_11858,N_9963,N_9857);
and U11859 (N_11859,N_7878,N_7969);
xnor U11860 (N_11860,N_9329,N_8616);
or U11861 (N_11861,N_9044,N_7861);
and U11862 (N_11862,N_9619,N_9424);
nand U11863 (N_11863,N_9083,N_7774);
or U11864 (N_11864,N_7950,N_9854);
or U11865 (N_11865,N_9962,N_7855);
xnor U11866 (N_11866,N_8383,N_8143);
and U11867 (N_11867,N_7511,N_9643);
nor U11868 (N_11868,N_7982,N_9615);
and U11869 (N_11869,N_8581,N_8155);
nor U11870 (N_11870,N_9487,N_8815);
nand U11871 (N_11871,N_8802,N_8704);
and U11872 (N_11872,N_8868,N_7917);
or U11873 (N_11873,N_7857,N_9919);
nand U11874 (N_11874,N_7591,N_7680);
or U11875 (N_11875,N_8639,N_9637);
nand U11876 (N_11876,N_8554,N_8107);
xnor U11877 (N_11877,N_9425,N_8255);
nor U11878 (N_11878,N_8572,N_7604);
or U11879 (N_11879,N_7997,N_7698);
or U11880 (N_11880,N_9960,N_9905);
and U11881 (N_11881,N_9002,N_8620);
xor U11882 (N_11882,N_7974,N_9641);
xor U11883 (N_11883,N_9110,N_9842);
and U11884 (N_11884,N_7590,N_9034);
or U11885 (N_11885,N_7500,N_8990);
nand U11886 (N_11886,N_8705,N_8722);
nand U11887 (N_11887,N_8941,N_9337);
xnor U11888 (N_11888,N_9293,N_8229);
or U11889 (N_11889,N_9577,N_7811);
nand U11890 (N_11890,N_9470,N_9947);
nor U11891 (N_11891,N_9799,N_9419);
and U11892 (N_11892,N_9881,N_9681);
or U11893 (N_11893,N_9059,N_8445);
and U11894 (N_11894,N_7880,N_9219);
or U11895 (N_11895,N_8592,N_8220);
and U11896 (N_11896,N_9421,N_8386);
nand U11897 (N_11897,N_7677,N_8911);
and U11898 (N_11898,N_7975,N_8980);
xor U11899 (N_11899,N_7522,N_9664);
xor U11900 (N_11900,N_9705,N_9072);
nor U11901 (N_11901,N_9108,N_8150);
or U11902 (N_11902,N_7918,N_9057);
nor U11903 (N_11903,N_8199,N_9247);
and U11904 (N_11904,N_7680,N_9158);
nor U11905 (N_11905,N_8996,N_8939);
and U11906 (N_11906,N_7983,N_8742);
or U11907 (N_11907,N_8906,N_9308);
nor U11908 (N_11908,N_7816,N_8580);
nor U11909 (N_11909,N_9994,N_9490);
nand U11910 (N_11910,N_8073,N_9553);
nand U11911 (N_11911,N_7985,N_7606);
xnor U11912 (N_11912,N_9623,N_9588);
xnor U11913 (N_11913,N_9955,N_8151);
and U11914 (N_11914,N_8173,N_8981);
and U11915 (N_11915,N_9722,N_9863);
nand U11916 (N_11916,N_8093,N_8434);
and U11917 (N_11917,N_7567,N_7981);
xnor U11918 (N_11918,N_7762,N_9161);
or U11919 (N_11919,N_9022,N_7660);
nand U11920 (N_11920,N_8822,N_8315);
nand U11921 (N_11921,N_9943,N_9243);
xnor U11922 (N_11922,N_9170,N_9032);
and U11923 (N_11923,N_9859,N_9308);
xnor U11924 (N_11924,N_7506,N_7808);
xnor U11925 (N_11925,N_9144,N_7850);
xor U11926 (N_11926,N_8429,N_9431);
and U11927 (N_11927,N_8873,N_9980);
or U11928 (N_11928,N_8231,N_7673);
xnor U11929 (N_11929,N_7927,N_7648);
and U11930 (N_11930,N_9554,N_8076);
xor U11931 (N_11931,N_7792,N_9688);
xnor U11932 (N_11932,N_9650,N_7662);
or U11933 (N_11933,N_8754,N_8230);
nand U11934 (N_11934,N_7974,N_8617);
nand U11935 (N_11935,N_8699,N_8221);
nand U11936 (N_11936,N_8237,N_7684);
xor U11937 (N_11937,N_7985,N_9376);
nor U11938 (N_11938,N_7723,N_8531);
xnor U11939 (N_11939,N_9161,N_7957);
and U11940 (N_11940,N_9031,N_9695);
nor U11941 (N_11941,N_9396,N_9637);
xnor U11942 (N_11942,N_8796,N_8797);
xnor U11943 (N_11943,N_8389,N_8807);
nand U11944 (N_11944,N_8953,N_7508);
and U11945 (N_11945,N_9756,N_9601);
and U11946 (N_11946,N_9554,N_9548);
xnor U11947 (N_11947,N_8105,N_8715);
nor U11948 (N_11948,N_8853,N_8406);
xnor U11949 (N_11949,N_7625,N_9550);
and U11950 (N_11950,N_8935,N_8307);
xnor U11951 (N_11951,N_7839,N_9092);
nand U11952 (N_11952,N_7515,N_7521);
and U11953 (N_11953,N_8966,N_7561);
nand U11954 (N_11954,N_8348,N_8061);
and U11955 (N_11955,N_8924,N_9988);
or U11956 (N_11956,N_8393,N_8689);
or U11957 (N_11957,N_8258,N_8463);
or U11958 (N_11958,N_9590,N_8822);
or U11959 (N_11959,N_9932,N_7942);
nand U11960 (N_11960,N_7602,N_7840);
nand U11961 (N_11961,N_7735,N_8940);
xnor U11962 (N_11962,N_9493,N_7543);
and U11963 (N_11963,N_9915,N_9240);
nor U11964 (N_11964,N_9869,N_9051);
nand U11965 (N_11965,N_7826,N_7698);
nor U11966 (N_11966,N_8912,N_8169);
nand U11967 (N_11967,N_7926,N_9396);
or U11968 (N_11968,N_9655,N_9221);
or U11969 (N_11969,N_8652,N_8168);
xor U11970 (N_11970,N_9957,N_9608);
xnor U11971 (N_11971,N_8186,N_9199);
or U11972 (N_11972,N_9226,N_8616);
xor U11973 (N_11973,N_7841,N_8922);
nand U11974 (N_11974,N_8878,N_8641);
xor U11975 (N_11975,N_8876,N_9063);
nor U11976 (N_11976,N_9563,N_7691);
nand U11977 (N_11977,N_7998,N_8686);
and U11978 (N_11978,N_8463,N_8183);
xnor U11979 (N_11979,N_9030,N_8329);
nor U11980 (N_11980,N_8446,N_7968);
and U11981 (N_11981,N_7629,N_8525);
nor U11982 (N_11982,N_8982,N_9157);
or U11983 (N_11983,N_9400,N_8056);
nand U11984 (N_11984,N_8051,N_7960);
or U11985 (N_11985,N_7979,N_8458);
xnor U11986 (N_11986,N_8595,N_9821);
nand U11987 (N_11987,N_8348,N_9626);
nor U11988 (N_11988,N_7995,N_8090);
nand U11989 (N_11989,N_9132,N_7950);
and U11990 (N_11990,N_8610,N_7993);
nor U11991 (N_11991,N_8171,N_9305);
or U11992 (N_11992,N_8898,N_9922);
nand U11993 (N_11993,N_9624,N_9842);
or U11994 (N_11994,N_7983,N_8648);
or U11995 (N_11995,N_9906,N_9842);
nand U11996 (N_11996,N_8003,N_8167);
nor U11997 (N_11997,N_9402,N_7684);
xnor U11998 (N_11998,N_9834,N_8893);
nand U11999 (N_11999,N_7884,N_9304);
xnor U12000 (N_12000,N_9332,N_8825);
xnor U12001 (N_12001,N_9428,N_8192);
and U12002 (N_12002,N_8486,N_7544);
xnor U12003 (N_12003,N_8587,N_9961);
nor U12004 (N_12004,N_8740,N_9491);
and U12005 (N_12005,N_9089,N_7579);
xnor U12006 (N_12006,N_8330,N_8869);
and U12007 (N_12007,N_8790,N_9634);
nand U12008 (N_12008,N_9213,N_9489);
nand U12009 (N_12009,N_9347,N_9353);
xnor U12010 (N_12010,N_8263,N_9012);
and U12011 (N_12011,N_8103,N_8452);
nand U12012 (N_12012,N_7791,N_8460);
nor U12013 (N_12013,N_9096,N_8589);
and U12014 (N_12014,N_9147,N_8924);
or U12015 (N_12015,N_8602,N_8516);
or U12016 (N_12016,N_7558,N_8476);
or U12017 (N_12017,N_9810,N_9143);
or U12018 (N_12018,N_9068,N_7952);
nand U12019 (N_12019,N_7905,N_9571);
nor U12020 (N_12020,N_9510,N_9642);
nor U12021 (N_12021,N_9618,N_9719);
or U12022 (N_12022,N_7643,N_8874);
or U12023 (N_12023,N_8931,N_9380);
or U12024 (N_12024,N_9430,N_8591);
nand U12025 (N_12025,N_9859,N_9284);
nor U12026 (N_12026,N_7734,N_8801);
nand U12027 (N_12027,N_9105,N_7873);
nand U12028 (N_12028,N_8339,N_8590);
xor U12029 (N_12029,N_8095,N_8798);
or U12030 (N_12030,N_8887,N_9061);
nor U12031 (N_12031,N_8680,N_7985);
nand U12032 (N_12032,N_9539,N_9607);
nor U12033 (N_12033,N_9659,N_8327);
nor U12034 (N_12034,N_7630,N_8007);
nor U12035 (N_12035,N_8730,N_7969);
nand U12036 (N_12036,N_7528,N_9574);
or U12037 (N_12037,N_8756,N_7934);
nand U12038 (N_12038,N_7844,N_7592);
nor U12039 (N_12039,N_9144,N_9774);
nand U12040 (N_12040,N_7917,N_7628);
and U12041 (N_12041,N_8560,N_7586);
nand U12042 (N_12042,N_8405,N_8599);
and U12043 (N_12043,N_9141,N_9568);
nand U12044 (N_12044,N_9974,N_9598);
xor U12045 (N_12045,N_9326,N_7765);
nor U12046 (N_12046,N_8800,N_7734);
or U12047 (N_12047,N_8695,N_9797);
nand U12048 (N_12048,N_8345,N_9008);
or U12049 (N_12049,N_8010,N_7980);
and U12050 (N_12050,N_8290,N_8596);
nor U12051 (N_12051,N_8118,N_7642);
or U12052 (N_12052,N_9081,N_9281);
nand U12053 (N_12053,N_8163,N_7750);
and U12054 (N_12054,N_7699,N_9376);
and U12055 (N_12055,N_9714,N_7706);
xor U12056 (N_12056,N_7695,N_9862);
and U12057 (N_12057,N_9079,N_8557);
and U12058 (N_12058,N_9280,N_8212);
nor U12059 (N_12059,N_8064,N_8830);
and U12060 (N_12060,N_7555,N_9718);
nand U12061 (N_12061,N_9850,N_9223);
and U12062 (N_12062,N_8538,N_8794);
xor U12063 (N_12063,N_9972,N_7509);
and U12064 (N_12064,N_8347,N_7644);
nor U12065 (N_12065,N_9057,N_9566);
nand U12066 (N_12066,N_8910,N_7923);
or U12067 (N_12067,N_9487,N_9633);
or U12068 (N_12068,N_9749,N_9944);
or U12069 (N_12069,N_8083,N_8406);
nor U12070 (N_12070,N_9548,N_7593);
and U12071 (N_12071,N_9943,N_8813);
or U12072 (N_12072,N_7947,N_8815);
and U12073 (N_12073,N_8849,N_7728);
or U12074 (N_12074,N_9277,N_9752);
and U12075 (N_12075,N_9178,N_8939);
xnor U12076 (N_12076,N_9085,N_7871);
or U12077 (N_12077,N_9680,N_8442);
and U12078 (N_12078,N_7692,N_7987);
or U12079 (N_12079,N_8817,N_9738);
nor U12080 (N_12080,N_8957,N_8687);
and U12081 (N_12081,N_9128,N_8461);
xnor U12082 (N_12082,N_9407,N_9242);
and U12083 (N_12083,N_8382,N_8433);
and U12084 (N_12084,N_7866,N_8942);
and U12085 (N_12085,N_9904,N_8730);
or U12086 (N_12086,N_8587,N_9689);
and U12087 (N_12087,N_9837,N_8944);
and U12088 (N_12088,N_8733,N_8263);
nand U12089 (N_12089,N_7659,N_8999);
or U12090 (N_12090,N_7647,N_7506);
xnor U12091 (N_12091,N_7626,N_8059);
nand U12092 (N_12092,N_9840,N_9046);
nor U12093 (N_12093,N_7862,N_8343);
nand U12094 (N_12094,N_9181,N_8270);
and U12095 (N_12095,N_9147,N_7514);
nor U12096 (N_12096,N_9018,N_7958);
xor U12097 (N_12097,N_9958,N_7508);
or U12098 (N_12098,N_8991,N_9536);
or U12099 (N_12099,N_8086,N_8961);
nand U12100 (N_12100,N_9385,N_8182);
or U12101 (N_12101,N_8102,N_8801);
or U12102 (N_12102,N_8600,N_8739);
xnor U12103 (N_12103,N_9418,N_8294);
xor U12104 (N_12104,N_8434,N_8871);
nand U12105 (N_12105,N_8954,N_9439);
nand U12106 (N_12106,N_9543,N_8343);
or U12107 (N_12107,N_8825,N_8972);
nand U12108 (N_12108,N_9233,N_7681);
and U12109 (N_12109,N_9862,N_9003);
nor U12110 (N_12110,N_8708,N_8575);
nor U12111 (N_12111,N_8957,N_9072);
or U12112 (N_12112,N_7836,N_8944);
or U12113 (N_12113,N_9627,N_9517);
nor U12114 (N_12114,N_9399,N_7505);
xnor U12115 (N_12115,N_9629,N_7662);
and U12116 (N_12116,N_9218,N_9991);
nor U12117 (N_12117,N_8548,N_9187);
xnor U12118 (N_12118,N_9438,N_9822);
nor U12119 (N_12119,N_8430,N_9087);
and U12120 (N_12120,N_9038,N_8823);
or U12121 (N_12121,N_9881,N_8066);
or U12122 (N_12122,N_8353,N_9439);
or U12123 (N_12123,N_9682,N_9304);
nor U12124 (N_12124,N_8742,N_8321);
nand U12125 (N_12125,N_9489,N_9080);
nor U12126 (N_12126,N_9874,N_7550);
or U12127 (N_12127,N_7549,N_8789);
xnor U12128 (N_12128,N_7791,N_8041);
xor U12129 (N_12129,N_9406,N_7704);
xnor U12130 (N_12130,N_8441,N_9684);
or U12131 (N_12131,N_9215,N_7629);
xor U12132 (N_12132,N_7605,N_8095);
and U12133 (N_12133,N_8844,N_8144);
nand U12134 (N_12134,N_7827,N_7966);
and U12135 (N_12135,N_7973,N_7811);
xor U12136 (N_12136,N_9359,N_9833);
nor U12137 (N_12137,N_9713,N_8769);
and U12138 (N_12138,N_9530,N_7534);
xnor U12139 (N_12139,N_7675,N_8836);
xor U12140 (N_12140,N_9898,N_8422);
xnor U12141 (N_12141,N_7942,N_9170);
nor U12142 (N_12142,N_8436,N_9195);
nor U12143 (N_12143,N_9299,N_9666);
or U12144 (N_12144,N_9197,N_8050);
nor U12145 (N_12145,N_9024,N_9071);
and U12146 (N_12146,N_8327,N_8896);
xnor U12147 (N_12147,N_8397,N_7966);
nand U12148 (N_12148,N_9688,N_8441);
xor U12149 (N_12149,N_7529,N_9966);
or U12150 (N_12150,N_9461,N_9620);
xor U12151 (N_12151,N_8733,N_8122);
xor U12152 (N_12152,N_9026,N_8911);
nor U12153 (N_12153,N_9673,N_9348);
or U12154 (N_12154,N_9424,N_7503);
or U12155 (N_12155,N_7936,N_7847);
nand U12156 (N_12156,N_9575,N_7729);
nor U12157 (N_12157,N_8059,N_7744);
nand U12158 (N_12158,N_8057,N_8086);
nand U12159 (N_12159,N_9474,N_9772);
and U12160 (N_12160,N_9192,N_8223);
xor U12161 (N_12161,N_7949,N_7550);
nor U12162 (N_12162,N_9644,N_7651);
or U12163 (N_12163,N_9794,N_9211);
nor U12164 (N_12164,N_9815,N_9436);
or U12165 (N_12165,N_8148,N_7502);
nor U12166 (N_12166,N_8791,N_8540);
xnor U12167 (N_12167,N_8271,N_8330);
or U12168 (N_12168,N_7698,N_9632);
nor U12169 (N_12169,N_8405,N_8431);
or U12170 (N_12170,N_8096,N_9534);
and U12171 (N_12171,N_8943,N_9427);
nand U12172 (N_12172,N_7705,N_7755);
nor U12173 (N_12173,N_7756,N_8601);
nand U12174 (N_12174,N_8480,N_8470);
and U12175 (N_12175,N_8065,N_9334);
nor U12176 (N_12176,N_9277,N_7590);
xor U12177 (N_12177,N_8693,N_7828);
nor U12178 (N_12178,N_9532,N_9095);
and U12179 (N_12179,N_8378,N_8678);
nand U12180 (N_12180,N_8100,N_8038);
and U12181 (N_12181,N_9307,N_9343);
nor U12182 (N_12182,N_8573,N_9802);
xor U12183 (N_12183,N_8320,N_9381);
or U12184 (N_12184,N_8341,N_8799);
or U12185 (N_12185,N_7778,N_9307);
xnor U12186 (N_12186,N_8821,N_8867);
and U12187 (N_12187,N_7838,N_9545);
or U12188 (N_12188,N_8193,N_9114);
nand U12189 (N_12189,N_9370,N_9479);
or U12190 (N_12190,N_7556,N_7527);
xnor U12191 (N_12191,N_7993,N_9813);
and U12192 (N_12192,N_9771,N_8780);
or U12193 (N_12193,N_9345,N_8074);
and U12194 (N_12194,N_9759,N_8432);
nand U12195 (N_12195,N_9119,N_7579);
nor U12196 (N_12196,N_8013,N_8842);
and U12197 (N_12197,N_7797,N_8063);
and U12198 (N_12198,N_8849,N_8761);
nor U12199 (N_12199,N_8197,N_9592);
nor U12200 (N_12200,N_8323,N_9854);
xor U12201 (N_12201,N_7542,N_8785);
nor U12202 (N_12202,N_8364,N_9434);
nand U12203 (N_12203,N_9543,N_9232);
xor U12204 (N_12204,N_9536,N_8230);
xnor U12205 (N_12205,N_8437,N_9896);
nor U12206 (N_12206,N_9530,N_9162);
and U12207 (N_12207,N_9935,N_9383);
nor U12208 (N_12208,N_7890,N_8759);
or U12209 (N_12209,N_9359,N_8676);
xor U12210 (N_12210,N_9257,N_7847);
nor U12211 (N_12211,N_9353,N_9543);
nor U12212 (N_12212,N_8876,N_9578);
and U12213 (N_12213,N_7731,N_8335);
nor U12214 (N_12214,N_7829,N_7879);
nor U12215 (N_12215,N_7934,N_8857);
or U12216 (N_12216,N_8679,N_8929);
nand U12217 (N_12217,N_9841,N_9434);
nand U12218 (N_12218,N_8998,N_8953);
nand U12219 (N_12219,N_8744,N_8873);
nand U12220 (N_12220,N_8396,N_9174);
nor U12221 (N_12221,N_8586,N_7837);
xor U12222 (N_12222,N_8964,N_8773);
or U12223 (N_12223,N_7595,N_8914);
nor U12224 (N_12224,N_8843,N_7741);
nand U12225 (N_12225,N_7932,N_9660);
or U12226 (N_12226,N_9131,N_8046);
and U12227 (N_12227,N_8778,N_8783);
or U12228 (N_12228,N_9079,N_7900);
nand U12229 (N_12229,N_7951,N_7617);
nor U12230 (N_12230,N_7763,N_8916);
nand U12231 (N_12231,N_7727,N_7958);
and U12232 (N_12232,N_7919,N_9931);
and U12233 (N_12233,N_7792,N_8942);
nor U12234 (N_12234,N_8765,N_8207);
and U12235 (N_12235,N_9823,N_7600);
nor U12236 (N_12236,N_8254,N_8768);
nor U12237 (N_12237,N_9771,N_9867);
nor U12238 (N_12238,N_8698,N_7541);
and U12239 (N_12239,N_8225,N_8259);
nor U12240 (N_12240,N_9001,N_9132);
nor U12241 (N_12241,N_9972,N_8336);
or U12242 (N_12242,N_9319,N_9522);
nor U12243 (N_12243,N_8557,N_9178);
or U12244 (N_12244,N_7604,N_9809);
nand U12245 (N_12245,N_7945,N_7616);
and U12246 (N_12246,N_8848,N_8932);
or U12247 (N_12247,N_8290,N_9251);
nor U12248 (N_12248,N_9520,N_7681);
xor U12249 (N_12249,N_8984,N_9501);
or U12250 (N_12250,N_7882,N_9483);
xnor U12251 (N_12251,N_7684,N_8155);
or U12252 (N_12252,N_9471,N_8138);
or U12253 (N_12253,N_9871,N_8695);
xnor U12254 (N_12254,N_8237,N_8546);
nand U12255 (N_12255,N_9088,N_9739);
xnor U12256 (N_12256,N_8902,N_9228);
xor U12257 (N_12257,N_9809,N_7670);
xnor U12258 (N_12258,N_8337,N_8682);
nand U12259 (N_12259,N_9926,N_9510);
nand U12260 (N_12260,N_8923,N_7599);
xnor U12261 (N_12261,N_8389,N_9658);
or U12262 (N_12262,N_9524,N_8456);
or U12263 (N_12263,N_8740,N_8411);
and U12264 (N_12264,N_9451,N_8309);
and U12265 (N_12265,N_9909,N_7633);
nor U12266 (N_12266,N_8566,N_8111);
nor U12267 (N_12267,N_7526,N_9497);
or U12268 (N_12268,N_8962,N_9419);
nand U12269 (N_12269,N_8720,N_8828);
xnor U12270 (N_12270,N_7964,N_9013);
xnor U12271 (N_12271,N_9162,N_8533);
nor U12272 (N_12272,N_8555,N_9588);
nand U12273 (N_12273,N_8500,N_8223);
nand U12274 (N_12274,N_7589,N_9085);
and U12275 (N_12275,N_9882,N_8030);
nor U12276 (N_12276,N_8517,N_9752);
xnor U12277 (N_12277,N_8762,N_7865);
nor U12278 (N_12278,N_9771,N_9200);
and U12279 (N_12279,N_8974,N_9411);
and U12280 (N_12280,N_8939,N_9532);
and U12281 (N_12281,N_8898,N_8756);
and U12282 (N_12282,N_7983,N_9173);
or U12283 (N_12283,N_9435,N_9232);
nand U12284 (N_12284,N_9558,N_8520);
and U12285 (N_12285,N_9539,N_9651);
and U12286 (N_12286,N_8437,N_9042);
or U12287 (N_12287,N_8668,N_8630);
or U12288 (N_12288,N_8827,N_8637);
or U12289 (N_12289,N_8568,N_7879);
and U12290 (N_12290,N_9287,N_9194);
nor U12291 (N_12291,N_9148,N_9800);
xnor U12292 (N_12292,N_7622,N_9165);
or U12293 (N_12293,N_8887,N_7694);
and U12294 (N_12294,N_8498,N_9975);
xnor U12295 (N_12295,N_8685,N_9963);
nor U12296 (N_12296,N_8709,N_8358);
nor U12297 (N_12297,N_8872,N_8609);
xnor U12298 (N_12298,N_8397,N_8664);
and U12299 (N_12299,N_8242,N_9801);
nand U12300 (N_12300,N_8454,N_9651);
and U12301 (N_12301,N_8158,N_8580);
nand U12302 (N_12302,N_9546,N_9448);
and U12303 (N_12303,N_9695,N_9421);
nor U12304 (N_12304,N_9097,N_8549);
or U12305 (N_12305,N_8569,N_8735);
xor U12306 (N_12306,N_9595,N_9435);
nand U12307 (N_12307,N_8945,N_8504);
nor U12308 (N_12308,N_8709,N_9142);
or U12309 (N_12309,N_9114,N_9556);
and U12310 (N_12310,N_9981,N_7802);
xnor U12311 (N_12311,N_8053,N_9930);
or U12312 (N_12312,N_8601,N_9790);
and U12313 (N_12313,N_8094,N_9419);
nand U12314 (N_12314,N_9346,N_9378);
or U12315 (N_12315,N_8477,N_9159);
xnor U12316 (N_12316,N_7561,N_7887);
nor U12317 (N_12317,N_9006,N_9387);
nand U12318 (N_12318,N_8289,N_9844);
or U12319 (N_12319,N_7732,N_8556);
xor U12320 (N_12320,N_8502,N_7795);
and U12321 (N_12321,N_9860,N_9313);
and U12322 (N_12322,N_9179,N_9339);
or U12323 (N_12323,N_9787,N_9595);
or U12324 (N_12324,N_7502,N_8293);
nor U12325 (N_12325,N_7584,N_8549);
nand U12326 (N_12326,N_8170,N_7626);
and U12327 (N_12327,N_9245,N_9380);
nor U12328 (N_12328,N_8363,N_8746);
xor U12329 (N_12329,N_9916,N_7959);
or U12330 (N_12330,N_8076,N_9618);
nand U12331 (N_12331,N_8682,N_8882);
nand U12332 (N_12332,N_9214,N_8263);
and U12333 (N_12333,N_7632,N_8876);
nand U12334 (N_12334,N_8032,N_9053);
or U12335 (N_12335,N_9512,N_8968);
xnor U12336 (N_12336,N_9308,N_9004);
or U12337 (N_12337,N_8403,N_7775);
nor U12338 (N_12338,N_9761,N_9855);
or U12339 (N_12339,N_8952,N_9166);
xor U12340 (N_12340,N_9733,N_8949);
nor U12341 (N_12341,N_9167,N_7783);
xnor U12342 (N_12342,N_8926,N_9614);
xnor U12343 (N_12343,N_9050,N_9923);
or U12344 (N_12344,N_7662,N_8429);
or U12345 (N_12345,N_8020,N_9094);
and U12346 (N_12346,N_7708,N_8286);
and U12347 (N_12347,N_8469,N_9712);
xor U12348 (N_12348,N_9021,N_9136);
or U12349 (N_12349,N_7663,N_7566);
and U12350 (N_12350,N_9870,N_9383);
and U12351 (N_12351,N_7863,N_7645);
xnor U12352 (N_12352,N_8744,N_9038);
xnor U12353 (N_12353,N_9948,N_8971);
xnor U12354 (N_12354,N_9553,N_8204);
nor U12355 (N_12355,N_8481,N_8499);
or U12356 (N_12356,N_8356,N_9915);
nand U12357 (N_12357,N_9600,N_8477);
nor U12358 (N_12358,N_9644,N_8334);
nand U12359 (N_12359,N_9304,N_9875);
nor U12360 (N_12360,N_9121,N_7872);
xor U12361 (N_12361,N_9490,N_8566);
xor U12362 (N_12362,N_9364,N_7545);
or U12363 (N_12363,N_9192,N_7508);
or U12364 (N_12364,N_7830,N_9155);
xor U12365 (N_12365,N_7731,N_8542);
xor U12366 (N_12366,N_8273,N_7589);
nor U12367 (N_12367,N_8075,N_8112);
and U12368 (N_12368,N_9670,N_8877);
or U12369 (N_12369,N_9401,N_9817);
nor U12370 (N_12370,N_8041,N_7659);
and U12371 (N_12371,N_9962,N_9254);
and U12372 (N_12372,N_8575,N_8600);
nor U12373 (N_12373,N_7598,N_8287);
or U12374 (N_12374,N_9371,N_9058);
or U12375 (N_12375,N_7710,N_9225);
nand U12376 (N_12376,N_7988,N_8453);
nor U12377 (N_12377,N_8010,N_9657);
or U12378 (N_12378,N_8317,N_8429);
nand U12379 (N_12379,N_9603,N_9859);
xnor U12380 (N_12380,N_9678,N_7592);
or U12381 (N_12381,N_9277,N_9493);
and U12382 (N_12382,N_9242,N_8631);
nand U12383 (N_12383,N_8513,N_9223);
nor U12384 (N_12384,N_9048,N_7860);
or U12385 (N_12385,N_9372,N_7557);
or U12386 (N_12386,N_9969,N_7587);
nand U12387 (N_12387,N_9425,N_8359);
and U12388 (N_12388,N_8769,N_9046);
nand U12389 (N_12389,N_8311,N_9256);
nor U12390 (N_12390,N_9671,N_7652);
nor U12391 (N_12391,N_8072,N_8096);
or U12392 (N_12392,N_9377,N_8526);
xnor U12393 (N_12393,N_8515,N_9327);
xor U12394 (N_12394,N_9478,N_9297);
and U12395 (N_12395,N_7942,N_7604);
nand U12396 (N_12396,N_9926,N_8704);
nand U12397 (N_12397,N_8831,N_9389);
nor U12398 (N_12398,N_8548,N_9448);
nor U12399 (N_12399,N_9616,N_9271);
and U12400 (N_12400,N_8786,N_8980);
nand U12401 (N_12401,N_9217,N_7612);
or U12402 (N_12402,N_7574,N_9819);
or U12403 (N_12403,N_8832,N_8799);
nor U12404 (N_12404,N_9223,N_9069);
xor U12405 (N_12405,N_8627,N_9531);
or U12406 (N_12406,N_8527,N_8854);
or U12407 (N_12407,N_7602,N_9915);
and U12408 (N_12408,N_7572,N_8238);
nand U12409 (N_12409,N_8064,N_9506);
and U12410 (N_12410,N_8356,N_8865);
or U12411 (N_12411,N_9673,N_9145);
and U12412 (N_12412,N_9937,N_9914);
and U12413 (N_12413,N_8410,N_9646);
xnor U12414 (N_12414,N_7619,N_9571);
nor U12415 (N_12415,N_8431,N_8847);
and U12416 (N_12416,N_8830,N_7576);
xnor U12417 (N_12417,N_9069,N_8904);
xnor U12418 (N_12418,N_8479,N_9205);
xor U12419 (N_12419,N_9350,N_8344);
and U12420 (N_12420,N_9101,N_8406);
nor U12421 (N_12421,N_9096,N_8635);
and U12422 (N_12422,N_7756,N_8988);
nand U12423 (N_12423,N_9767,N_8860);
xor U12424 (N_12424,N_7902,N_9549);
or U12425 (N_12425,N_8658,N_8063);
nand U12426 (N_12426,N_9789,N_7694);
and U12427 (N_12427,N_7574,N_7803);
nand U12428 (N_12428,N_7684,N_8832);
or U12429 (N_12429,N_8490,N_9519);
and U12430 (N_12430,N_8130,N_7717);
nand U12431 (N_12431,N_8524,N_8415);
and U12432 (N_12432,N_9279,N_8019);
nor U12433 (N_12433,N_9939,N_9761);
nand U12434 (N_12434,N_8444,N_8423);
and U12435 (N_12435,N_9966,N_9027);
or U12436 (N_12436,N_8797,N_9339);
nand U12437 (N_12437,N_9266,N_8855);
or U12438 (N_12438,N_8156,N_8758);
nand U12439 (N_12439,N_7537,N_9753);
or U12440 (N_12440,N_8355,N_8637);
or U12441 (N_12441,N_8217,N_7722);
nand U12442 (N_12442,N_9830,N_9228);
nor U12443 (N_12443,N_9035,N_9960);
xnor U12444 (N_12444,N_9478,N_7726);
or U12445 (N_12445,N_9203,N_8127);
xor U12446 (N_12446,N_8945,N_8458);
and U12447 (N_12447,N_7838,N_8656);
or U12448 (N_12448,N_7779,N_8741);
and U12449 (N_12449,N_9528,N_8326);
xnor U12450 (N_12450,N_9228,N_8911);
nor U12451 (N_12451,N_8960,N_9707);
xor U12452 (N_12452,N_8004,N_8473);
or U12453 (N_12453,N_8535,N_8283);
nor U12454 (N_12454,N_9310,N_8278);
xor U12455 (N_12455,N_8027,N_9645);
or U12456 (N_12456,N_8707,N_8422);
nand U12457 (N_12457,N_9297,N_8458);
xor U12458 (N_12458,N_9580,N_7853);
and U12459 (N_12459,N_8807,N_9082);
or U12460 (N_12460,N_7510,N_8582);
and U12461 (N_12461,N_8622,N_9841);
nand U12462 (N_12462,N_7906,N_8934);
and U12463 (N_12463,N_8745,N_7901);
and U12464 (N_12464,N_8701,N_9785);
nand U12465 (N_12465,N_9013,N_7615);
xnor U12466 (N_12466,N_7679,N_9417);
xnor U12467 (N_12467,N_9611,N_8304);
and U12468 (N_12468,N_9916,N_8915);
nor U12469 (N_12469,N_8698,N_8116);
xor U12470 (N_12470,N_8814,N_8553);
and U12471 (N_12471,N_9696,N_8542);
xor U12472 (N_12472,N_9641,N_8003);
nand U12473 (N_12473,N_8252,N_7682);
nand U12474 (N_12474,N_8884,N_9818);
nor U12475 (N_12475,N_9556,N_9480);
and U12476 (N_12476,N_9746,N_8379);
or U12477 (N_12477,N_8119,N_9486);
nand U12478 (N_12478,N_8076,N_9200);
xnor U12479 (N_12479,N_8001,N_7531);
or U12480 (N_12480,N_7729,N_8578);
nand U12481 (N_12481,N_8548,N_9318);
nor U12482 (N_12482,N_9839,N_9102);
nor U12483 (N_12483,N_7513,N_9122);
and U12484 (N_12484,N_8004,N_7637);
and U12485 (N_12485,N_7555,N_8442);
and U12486 (N_12486,N_9025,N_9353);
nor U12487 (N_12487,N_8506,N_8609);
nand U12488 (N_12488,N_9149,N_7603);
or U12489 (N_12489,N_9661,N_8846);
nand U12490 (N_12490,N_9348,N_8662);
nand U12491 (N_12491,N_8753,N_9891);
xnor U12492 (N_12492,N_8913,N_9759);
or U12493 (N_12493,N_8736,N_7850);
nor U12494 (N_12494,N_9393,N_7541);
or U12495 (N_12495,N_9713,N_8793);
and U12496 (N_12496,N_8840,N_8479);
and U12497 (N_12497,N_8230,N_7819);
nor U12498 (N_12498,N_7813,N_7595);
and U12499 (N_12499,N_9478,N_9081);
nor U12500 (N_12500,N_11972,N_10538);
nor U12501 (N_12501,N_11047,N_10762);
xor U12502 (N_12502,N_11995,N_12279);
nand U12503 (N_12503,N_10872,N_11500);
xor U12504 (N_12504,N_10053,N_11631);
nand U12505 (N_12505,N_12121,N_10671);
or U12506 (N_12506,N_10967,N_12191);
and U12507 (N_12507,N_11542,N_10735);
nor U12508 (N_12508,N_10311,N_11054);
and U12509 (N_12509,N_11055,N_10086);
or U12510 (N_12510,N_10740,N_12293);
and U12511 (N_12511,N_11416,N_12143);
nor U12512 (N_12512,N_11557,N_10235);
nor U12513 (N_12513,N_12390,N_12125);
and U12514 (N_12514,N_12495,N_11398);
nand U12515 (N_12515,N_11588,N_11623);
or U12516 (N_12516,N_10632,N_11771);
nor U12517 (N_12517,N_11442,N_10726);
xor U12518 (N_12518,N_10320,N_12337);
xnor U12519 (N_12519,N_10244,N_11966);
xnor U12520 (N_12520,N_10029,N_10756);
xor U12521 (N_12521,N_10854,N_10763);
or U12522 (N_12522,N_11478,N_10817);
nand U12523 (N_12523,N_11074,N_11366);
nor U12524 (N_12524,N_11343,N_10189);
xnor U12525 (N_12525,N_12324,N_12194);
xor U12526 (N_12526,N_10602,N_11547);
xnor U12527 (N_12527,N_11855,N_10813);
and U12528 (N_12528,N_10048,N_12025);
or U12529 (N_12529,N_11341,N_10770);
or U12530 (N_12530,N_10623,N_10272);
xor U12531 (N_12531,N_11744,N_12227);
xnor U12532 (N_12532,N_11955,N_11549);
xor U12533 (N_12533,N_12375,N_10540);
or U12534 (N_12534,N_12126,N_11583);
nor U12535 (N_12535,N_11395,N_11419);
xnor U12536 (N_12536,N_11560,N_12344);
nor U12537 (N_12537,N_12475,N_11906);
and U12538 (N_12538,N_10665,N_12192);
or U12539 (N_12539,N_11913,N_11206);
nand U12540 (N_12540,N_10774,N_11863);
nor U12541 (N_12541,N_10258,N_10067);
or U12542 (N_12542,N_10675,N_10100);
nor U12543 (N_12543,N_12240,N_10928);
xnor U12544 (N_12544,N_11185,N_10388);
nand U12545 (N_12545,N_10986,N_12270);
nand U12546 (N_12546,N_11666,N_11065);
xor U12547 (N_12547,N_11192,N_12373);
nor U12548 (N_12548,N_11857,N_12338);
or U12549 (N_12549,N_10358,N_10240);
xor U12550 (N_12550,N_10641,N_12133);
nand U12551 (N_12551,N_11003,N_11522);
or U12552 (N_12552,N_11516,N_11014);
xor U12553 (N_12553,N_10597,N_10991);
and U12554 (N_12554,N_11632,N_11480);
nand U12555 (N_12555,N_10808,N_10246);
nand U12556 (N_12556,N_11933,N_10282);
nand U12557 (N_12557,N_11162,N_11705);
or U12558 (N_12558,N_12258,N_10378);
xor U12559 (N_12559,N_12439,N_12478);
nor U12560 (N_12560,N_11724,N_12265);
nor U12561 (N_12561,N_11902,N_11778);
xor U12562 (N_12562,N_10290,N_12347);
nor U12563 (N_12563,N_10230,N_12357);
nand U12564 (N_12564,N_11153,N_12307);
and U12565 (N_12565,N_12171,N_12459);
and U12566 (N_12566,N_12185,N_10911);
nand U12567 (N_12567,N_11172,N_12148);
nor U12568 (N_12568,N_11887,N_12306);
nor U12569 (N_12569,N_10487,N_11710);
nand U12570 (N_12570,N_11593,N_12209);
and U12571 (N_12571,N_10288,N_11506);
xnor U12572 (N_12572,N_10440,N_10899);
nor U12573 (N_12573,N_11550,N_11633);
nand U12574 (N_12574,N_10079,N_10070);
nand U12575 (N_12575,N_12158,N_10385);
xnor U12576 (N_12576,N_11757,N_12496);
or U12577 (N_12577,N_12303,N_12248);
nor U12578 (N_12578,N_12094,N_12323);
and U12579 (N_12579,N_10020,N_12470);
or U12580 (N_12580,N_11302,N_10741);
nor U12581 (N_12581,N_11152,N_10834);
and U12582 (N_12582,N_10448,N_10043);
or U12583 (N_12583,N_10044,N_12273);
nand U12584 (N_12584,N_11555,N_11002);
and U12585 (N_12585,N_11989,N_12421);
or U12586 (N_12586,N_12352,N_10289);
and U12587 (N_12587,N_11434,N_11931);
and U12588 (N_12588,N_11012,N_11754);
nand U12589 (N_12589,N_12297,N_10682);
and U12590 (N_12590,N_11649,N_11646);
or U12591 (N_12591,N_11218,N_10422);
or U12592 (N_12592,N_12413,N_11477);
xnor U12593 (N_12593,N_11561,N_11204);
nand U12594 (N_12594,N_10278,N_11051);
xnor U12595 (N_12595,N_12467,N_11774);
and U12596 (N_12596,N_10635,N_10200);
nand U12597 (N_12597,N_11504,N_10130);
and U12598 (N_12598,N_12316,N_10075);
nor U12599 (N_12599,N_11585,N_12354);
or U12600 (N_12600,N_11182,N_10861);
nor U12601 (N_12601,N_10150,N_11930);
or U12602 (N_12602,N_10201,N_11041);
xor U12603 (N_12603,N_11028,N_12198);
or U12604 (N_12604,N_12465,N_10430);
nand U12605 (N_12605,N_11075,N_11077);
nor U12606 (N_12606,N_11792,N_10192);
xnor U12607 (N_12607,N_12230,N_11865);
xor U12608 (N_12608,N_10112,N_11409);
nand U12609 (N_12609,N_12268,N_10927);
and U12610 (N_12610,N_11451,N_12489);
and U12611 (N_12611,N_12416,N_10934);
nand U12612 (N_12612,N_10653,N_11997);
nor U12613 (N_12613,N_11163,N_10082);
or U12614 (N_12614,N_12207,N_10620);
or U12615 (N_12615,N_11348,N_10081);
nor U12616 (N_12616,N_10280,N_10490);
and U12617 (N_12617,N_10248,N_10794);
xor U12618 (N_12618,N_10441,N_10666);
and U12619 (N_12619,N_10199,N_11001);
or U12620 (N_12620,N_11715,N_11134);
xor U12621 (N_12621,N_11030,N_12423);
or U12622 (N_12622,N_11203,N_12369);
or U12623 (N_12623,N_12221,N_10517);
or U12624 (N_12624,N_12320,N_12244);
nor U12625 (N_12625,N_11764,N_10639);
nor U12626 (N_12626,N_12104,N_10616);
xor U12627 (N_12627,N_10113,N_11685);
nand U12628 (N_12628,N_12041,N_12098);
nand U12629 (N_12629,N_12069,N_11293);
or U12630 (N_12630,N_11107,N_10019);
nor U12631 (N_12631,N_12417,N_11297);
or U12632 (N_12632,N_11460,N_10874);
and U12633 (N_12633,N_10603,N_10463);
xor U12634 (N_12634,N_11927,N_12267);
nor U12635 (N_12635,N_11546,N_11166);
nor U12636 (N_12636,N_10369,N_10454);
nand U12637 (N_12637,N_11637,N_12278);
nand U12638 (N_12638,N_12447,N_11136);
nor U12639 (N_12639,N_11604,N_12335);
nor U12640 (N_12640,N_11333,N_12301);
xnor U12641 (N_12641,N_11713,N_10224);
xnor U12642 (N_12642,N_10379,N_10807);
nand U12643 (N_12643,N_10955,N_12071);
nand U12644 (N_12644,N_10804,N_11895);
nand U12645 (N_12645,N_12407,N_10537);
and U12646 (N_12646,N_10532,N_12032);
nand U12647 (N_12647,N_11271,N_11843);
and U12648 (N_12648,N_11474,N_11468);
and U12649 (N_12649,N_12034,N_12432);
and U12650 (N_12650,N_11935,N_11740);
nor U12651 (N_12651,N_10847,N_12313);
and U12652 (N_12652,N_10042,N_11452);
nand U12653 (N_12653,N_10268,N_11575);
nor U12654 (N_12654,N_11952,N_11455);
nor U12655 (N_12655,N_11841,N_10174);
xor U12656 (N_12656,N_10466,N_11096);
or U12657 (N_12657,N_10459,N_12366);
xor U12658 (N_12658,N_10047,N_11237);
nand U12659 (N_12659,N_10000,N_11507);
nand U12660 (N_12660,N_10767,N_11563);
xor U12661 (N_12661,N_10974,N_10543);
xor U12662 (N_12662,N_11537,N_11839);
nand U12663 (N_12663,N_11183,N_10060);
nor U12664 (N_12664,N_12492,N_11362);
nor U12665 (N_12665,N_12113,N_10140);
nand U12666 (N_12666,N_10502,N_11878);
nor U12667 (N_12667,N_10723,N_11769);
nor U12668 (N_12668,N_11234,N_11834);
nor U12669 (N_12669,N_10030,N_11923);
nor U12670 (N_12670,N_10106,N_11804);
and U12671 (N_12671,N_10428,N_11675);
nand U12672 (N_12672,N_10349,N_12372);
nand U12673 (N_12673,N_12015,N_10315);
nand U12674 (N_12674,N_11365,N_11378);
and U12675 (N_12675,N_11728,N_12424);
or U12676 (N_12676,N_12280,N_11023);
and U12677 (N_12677,N_12111,N_10445);
nand U12678 (N_12678,N_12208,N_12181);
and U12679 (N_12679,N_12154,N_11700);
and U12680 (N_12680,N_11386,N_11674);
or U12681 (N_12681,N_11315,N_12136);
or U12682 (N_12682,N_10058,N_11978);
nand U12683 (N_12683,N_12242,N_10931);
nand U12684 (N_12684,N_11655,N_10800);
nand U12685 (N_12685,N_12277,N_11999);
nand U12686 (N_12686,N_10330,N_11198);
nand U12687 (N_12687,N_11737,N_10432);
nand U12688 (N_12688,N_11594,N_12341);
and U12689 (N_12689,N_12430,N_11007);
nand U12690 (N_12690,N_11161,N_12330);
xor U12691 (N_12691,N_11783,N_10568);
nand U12692 (N_12692,N_10015,N_11382);
nor U12693 (N_12693,N_10701,N_11412);
and U12694 (N_12694,N_11803,N_11064);
nand U12695 (N_12695,N_11200,N_10037);
nand U12696 (N_12696,N_11038,N_11309);
nor U12697 (N_12697,N_11929,N_11784);
and U12698 (N_12698,N_12093,N_10371);
or U12699 (N_12699,N_11829,N_12348);
and U12700 (N_12700,N_11485,N_12183);
nor U12701 (N_12701,N_10122,N_12095);
xnor U12702 (N_12702,N_11773,N_11566);
nand U12703 (N_12703,N_12151,N_11669);
xnor U12704 (N_12704,N_10582,N_11858);
nand U12705 (N_12705,N_10710,N_10750);
nand U12706 (N_12706,N_12252,N_10832);
or U12707 (N_12707,N_11105,N_10071);
nand U12708 (N_12708,N_12073,N_10564);
nand U12709 (N_12709,N_11894,N_10747);
and U12710 (N_12710,N_10470,N_10522);
xor U12711 (N_12711,N_12394,N_10998);
or U12712 (N_12712,N_11414,N_10354);
nor U12713 (N_12713,N_12395,N_10786);
nand U12714 (N_12714,N_11496,N_12130);
or U12715 (N_12715,N_11367,N_10152);
and U12716 (N_12716,N_12190,N_11712);
nand U12717 (N_12717,N_10527,N_12315);
nor U12718 (N_12718,N_11726,N_10018);
or U12719 (N_12719,N_11093,N_10728);
and U12720 (N_12720,N_10417,N_11187);
or U12721 (N_12721,N_12457,N_12122);
nand U12722 (N_12722,N_11687,N_10294);
or U12723 (N_12723,N_11558,N_10232);
and U12724 (N_12724,N_12441,N_10227);
xor U12725 (N_12725,N_11639,N_11866);
nor U12726 (N_12726,N_12055,N_10685);
or U12727 (N_12727,N_11891,N_11606);
or U12728 (N_12728,N_12234,N_11600);
or U12729 (N_12729,N_11595,N_10051);
nand U12730 (N_12730,N_11760,N_11938);
nor U12731 (N_12731,N_12051,N_11736);
xnor U12732 (N_12732,N_12440,N_11984);
nor U12733 (N_12733,N_10080,N_11100);
xor U12734 (N_12734,N_12172,N_10016);
nand U12735 (N_12735,N_11644,N_12396);
and U12736 (N_12736,N_11813,N_10118);
nor U12737 (N_12737,N_10326,N_11943);
xnor U12738 (N_12738,N_10924,N_11654);
or U12739 (N_12739,N_10922,N_10775);
nand U12740 (N_12740,N_12117,N_10863);
or U12741 (N_12741,N_10674,N_12139);
or U12742 (N_12742,N_12110,N_11659);
and U12743 (N_12743,N_12067,N_10707);
nor U12744 (N_12744,N_10376,N_10835);
nor U12745 (N_12745,N_10604,N_11679);
xor U12746 (N_12746,N_10598,N_10401);
nand U12747 (N_12747,N_12317,N_10894);
xnor U12748 (N_12748,N_10254,N_12219);
or U12749 (N_12749,N_10331,N_12291);
or U12750 (N_12750,N_11832,N_10884);
nor U12751 (N_12751,N_12493,N_10077);
nand U12752 (N_12752,N_11083,N_10695);
nand U12753 (N_12753,N_10117,N_11363);
nand U12754 (N_12754,N_11856,N_11559);
nand U12755 (N_12755,N_11324,N_10771);
nor U12756 (N_12756,N_10057,N_11120);
nor U12757 (N_12757,N_11073,N_10742);
nor U12758 (N_12758,N_11961,N_10933);
and U12759 (N_12759,N_11733,N_10852);
nor U12760 (N_12760,N_10626,N_10452);
nand U12761 (N_12761,N_10175,N_11782);
nor U12762 (N_12762,N_11720,N_10557);
or U12763 (N_12763,N_12384,N_11351);
and U12764 (N_12764,N_12134,N_10395);
nand U12765 (N_12765,N_12364,N_12068);
or U12766 (N_12766,N_10116,N_11266);
nand U12767 (N_12767,N_10091,N_12088);
or U12768 (N_12768,N_11610,N_11458);
or U12769 (N_12769,N_11758,N_10877);
nor U12770 (N_12770,N_10815,N_10782);
xor U12771 (N_12771,N_10381,N_11650);
nor U12772 (N_12772,N_11605,N_10929);
nor U12773 (N_12773,N_10049,N_10629);
and U12774 (N_12774,N_11181,N_11087);
xnor U12775 (N_12775,N_12005,N_10660);
xnor U12776 (N_12776,N_11115,N_11953);
nand U12777 (N_12777,N_11326,N_12434);
nor U12778 (N_12778,N_12004,N_10752);
nor U12779 (N_12779,N_10158,N_11838);
and U12780 (N_12780,N_10034,N_10054);
nor U12781 (N_12781,N_11336,N_10337);
or U12782 (N_12782,N_11979,N_12131);
and U12783 (N_12783,N_11624,N_12193);
nand U12784 (N_12784,N_10838,N_11323);
nand U12785 (N_12785,N_11421,N_10634);
nand U12786 (N_12786,N_10275,N_11168);
or U12787 (N_12787,N_11881,N_10627);
nand U12788 (N_12788,N_12188,N_12061);
xor U12789 (N_12789,N_10870,N_10344);
and U12790 (N_12790,N_11750,N_11454);
or U12791 (N_12791,N_11860,N_12075);
and U12792 (N_12792,N_11868,N_11069);
or U12793 (N_12793,N_10410,N_10920);
or U12794 (N_12794,N_10722,N_11143);
xnor U12795 (N_12795,N_11660,N_11084);
xnor U12796 (N_12796,N_12254,N_11034);
nand U12797 (N_12797,N_10413,N_10788);
nor U12798 (N_12798,N_11056,N_11031);
and U12799 (N_12799,N_11971,N_11411);
nor U12800 (N_12800,N_10370,N_11290);
xnor U12801 (N_12801,N_12035,N_11375);
nor U12802 (N_12802,N_10947,N_10718);
xor U12803 (N_12803,N_11657,N_10903);
xnor U12804 (N_12804,N_11908,N_11911);
xor U12805 (N_12805,N_12162,N_12445);
or U12806 (N_12806,N_11167,N_11948);
nor U12807 (N_12807,N_11548,N_10758);
nor U12808 (N_12808,N_10207,N_10485);
xor U12809 (N_12809,N_10969,N_10407);
and U12810 (N_12810,N_11368,N_10383);
or U12811 (N_12811,N_10738,N_10971);
nand U12812 (N_12812,N_11556,N_11922);
nor U12813 (N_12813,N_10438,N_10261);
nor U12814 (N_12814,N_11877,N_12000);
nand U12815 (N_12815,N_12246,N_11889);
xnor U12816 (N_12816,N_12002,N_12226);
and U12817 (N_12817,N_11830,N_11128);
nor U12818 (N_12818,N_11755,N_11518);
or U12819 (N_12819,N_11253,N_12247);
xor U12820 (N_12820,N_12468,N_11114);
and U12821 (N_12821,N_12175,N_11471);
and U12822 (N_12822,N_12250,N_11423);
xnor U12823 (N_12823,N_11864,N_11587);
or U12824 (N_12824,N_10943,N_10423);
nor U12825 (N_12825,N_12201,N_11207);
or U12826 (N_12826,N_12415,N_12054);
and U12827 (N_12827,N_11288,N_10185);
xor U12828 (N_12828,N_10721,N_11491);
nand U12829 (N_12829,N_10220,N_11042);
and U12830 (N_12830,N_10239,N_11890);
nand U12831 (N_12831,N_11872,N_10587);
xnor U12832 (N_12832,N_10589,N_12319);
nor U12833 (N_12833,N_10149,N_10109);
nand U12834 (N_12834,N_11123,N_10892);
and U12835 (N_12835,N_10216,N_10889);
or U12836 (N_12836,N_10827,N_10002);
xnor U12837 (N_12837,N_12135,N_10688);
or U12838 (N_12838,N_12355,N_10431);
nor U12839 (N_12839,N_10038,N_11811);
nor U12840 (N_12840,N_10901,N_10777);
nor U12841 (N_12841,N_11138,N_12107);
and U12842 (N_12842,N_12414,N_11974);
nor U12843 (N_12843,N_12129,N_10253);
nand U12844 (N_12844,N_10864,N_11818);
xor U12845 (N_12845,N_11707,N_10760);
or U12846 (N_12846,N_11800,N_11040);
xnor U12847 (N_12847,N_11260,N_11080);
and U12848 (N_12848,N_11230,N_10271);
or U12849 (N_12849,N_11325,N_11697);
xnor U12850 (N_12850,N_10702,N_11827);
nand U12851 (N_12851,N_11157,N_11987);
or U12852 (N_12852,N_10497,N_11968);
and U12853 (N_12853,N_10663,N_10733);
and U12854 (N_12854,N_12361,N_10706);
and U12855 (N_12855,N_11934,N_11239);
or U12856 (N_12856,N_11199,N_12286);
and U12857 (N_12857,N_12109,N_12228);
or U12858 (N_12858,N_12099,N_11453);
or U12859 (N_12859,N_12389,N_10757);
nor U12860 (N_12860,N_12036,N_10599);
nor U12861 (N_12861,N_11410,N_12149);
nand U12862 (N_12862,N_11656,N_10393);
and U12863 (N_12863,N_11721,N_11330);
and U12864 (N_12864,N_11063,N_10387);
nor U12865 (N_12865,N_10549,N_11033);
and U12866 (N_12866,N_12399,N_11553);
and U12867 (N_12867,N_10453,N_12127);
xnor U12868 (N_12868,N_11436,N_11472);
nor U12869 (N_12869,N_12266,N_11193);
nand U12870 (N_12870,N_10836,N_10995);
or U12871 (N_12871,N_10693,N_10961);
nor U12872 (N_12872,N_12038,N_11339);
and U12873 (N_12873,N_11910,N_11232);
nor U12874 (N_12874,N_11523,N_12308);
nand U12875 (N_12875,N_12174,N_12236);
xnor U12876 (N_12876,N_10176,N_11150);
nand U12877 (N_12877,N_11229,N_10050);
nand U12878 (N_12878,N_11861,N_10380);
or U12879 (N_12879,N_11291,N_10755);
and U12880 (N_12880,N_10567,N_10828);
nand U12881 (N_12881,N_10111,N_11772);
xnor U12882 (N_12882,N_11062,N_11994);
xor U12883 (N_12883,N_11739,N_12178);
nor U12884 (N_12884,N_10433,N_10559);
nor U12885 (N_12885,N_11567,N_10252);
nor U12886 (N_12886,N_10556,N_10196);
nor U12887 (N_12887,N_11884,N_12437);
and U12888 (N_12888,N_10759,N_10143);
and U12889 (N_12889,N_12435,N_11503);
or U12890 (N_12890,N_12145,N_11667);
or U12891 (N_12891,N_10643,N_11244);
and U12892 (N_12892,N_10979,N_12214);
and U12893 (N_12893,N_10435,N_12449);
nand U12894 (N_12894,N_12063,N_11327);
nand U12895 (N_12895,N_10263,N_11068);
nor U12896 (N_12896,N_10093,N_11964);
and U12897 (N_12897,N_11126,N_10411);
or U12898 (N_12898,N_11652,N_11638);
and U12899 (N_12899,N_11917,N_11456);
xor U12900 (N_12900,N_11924,N_12321);
or U12901 (N_12901,N_10753,N_10437);
and U12902 (N_12902,N_10744,N_11463);
nand U12903 (N_12903,N_11248,N_12391);
or U12904 (N_12904,N_10624,N_10180);
xnor U12905 (N_12905,N_10749,N_10679);
nor U12906 (N_12906,N_12412,N_11036);
and U12907 (N_12907,N_11440,N_10914);
nand U12908 (N_12908,N_11396,N_11225);
nor U12909 (N_12909,N_11734,N_11625);
xor U12910 (N_12910,N_10655,N_10724);
and U12911 (N_12911,N_11189,N_10913);
nor U12912 (N_12912,N_10205,N_10391);
nor U12913 (N_12913,N_11562,N_11190);
xor U12914 (N_12914,N_11196,N_11617);
nor U12915 (N_12915,N_10473,N_11982);
nor U12916 (N_12916,N_12382,N_12229);
nand U12917 (N_12917,N_12023,N_12065);
and U12918 (N_12918,N_11937,N_10853);
xnor U12919 (N_12919,N_10628,N_10831);
nor U12920 (N_12920,N_12084,N_10548);
or U12921 (N_12921,N_10965,N_10908);
nor U12922 (N_12922,N_10363,N_11949);
nand U12923 (N_12923,N_10193,N_11552);
nand U12924 (N_12924,N_12046,N_11766);
nand U12925 (N_12925,N_11429,N_11278);
or U12926 (N_12926,N_11591,N_10550);
and U12927 (N_12927,N_10519,N_11270);
and U12928 (N_12928,N_10382,N_11641);
and U12929 (N_12929,N_11526,N_11113);
nor U12930 (N_12930,N_10163,N_11347);
nand U12931 (N_12931,N_12272,N_11939);
xor U12932 (N_12932,N_10691,N_12351);
nor U12933 (N_12933,N_10825,N_11268);
or U12934 (N_12934,N_12251,N_12264);
or U12935 (N_12935,N_12360,N_12215);
nor U12936 (N_12936,N_10694,N_11110);
nand U12937 (N_12937,N_10493,N_12403);
and U12938 (N_12938,N_12336,N_10136);
xnor U12939 (N_12939,N_10021,N_11869);
xnor U12940 (N_12940,N_11301,N_11287);
nand U12941 (N_12941,N_10526,N_10650);
nor U12942 (N_12942,N_10234,N_12462);
nand U12943 (N_12943,N_10342,N_10449);
and U12944 (N_12944,N_12377,N_12011);
nor U12945 (N_12945,N_11169,N_11495);
and U12946 (N_12946,N_11517,N_10214);
nor U12947 (N_12947,N_11907,N_12097);
and U12948 (N_12948,N_11497,N_10966);
nand U12949 (N_12949,N_11532,N_11319);
or U12950 (N_12950,N_10241,N_12072);
and U12951 (N_12951,N_10824,N_10040);
nor U12952 (N_12952,N_11004,N_11767);
xor U12953 (N_12953,N_11180,N_11801);
or U12954 (N_12954,N_12045,N_11950);
or U12955 (N_12955,N_10439,N_12056);
nand U12956 (N_12956,N_11525,N_11662);
nor U12957 (N_12957,N_10229,N_11240);
and U12958 (N_12958,N_12472,N_11725);
xor U12959 (N_12959,N_10520,N_10313);
nor U12960 (N_12960,N_10510,N_11298);
nand U12961 (N_12961,N_10959,N_11570);
nand U12962 (N_12962,N_10094,N_10949);
nand U12963 (N_12963,N_11747,N_10173);
nand U12964 (N_12964,N_11275,N_11775);
xnor U12965 (N_12965,N_11130,N_10778);
xnor U12966 (N_12966,N_11027,N_12452);
xnor U12967 (N_12967,N_12367,N_11576);
and U12968 (N_12968,N_10651,N_11904);
or U12969 (N_12969,N_10687,N_12342);
nor U12970 (N_12970,N_11139,N_11751);
or U12971 (N_12971,N_10262,N_11620);
xnor U12972 (N_12972,N_10504,N_12076);
nor U12973 (N_12973,N_12257,N_10181);
or U12974 (N_12974,N_11228,N_11618);
nor U12975 (N_12975,N_11826,N_11371);
nor U12976 (N_12976,N_11885,N_11936);
and U12977 (N_12977,N_10713,N_11086);
nand U12978 (N_12978,N_12179,N_10322);
nor U12979 (N_12979,N_11462,N_11350);
nand U12980 (N_12980,N_11825,N_11101);
or U12981 (N_12981,N_11400,N_10638);
or U12982 (N_12982,N_11389,N_12461);
or U12983 (N_12983,N_11510,N_11777);
nor U12984 (N_12984,N_11888,N_11008);
and U12985 (N_12985,N_11787,N_12256);
nor U12986 (N_12986,N_12140,N_11158);
nor U12987 (N_12987,N_12189,N_10878);
nor U12988 (N_12988,N_10829,N_10987);
xnor U12989 (N_12989,N_10572,N_12410);
nand U12990 (N_12990,N_10225,N_12484);
nand U12991 (N_12991,N_10219,N_10101);
nor U12992 (N_12992,N_10684,N_10197);
nand U12993 (N_12993,N_12477,N_12294);
xnor U12994 (N_12994,N_10008,N_11520);
xnor U12995 (N_12995,N_11672,N_10301);
and U12996 (N_12996,N_11630,N_12120);
xor U12997 (N_12997,N_11572,N_11524);
nand U12998 (N_12998,N_11942,N_10221);
nor U12999 (N_12999,N_11046,N_12491);
nand U13000 (N_13000,N_10890,N_10056);
nor U13001 (N_13001,N_12379,N_11538);
nand U13002 (N_13002,N_10912,N_11693);
nor U13003 (N_13003,N_10714,N_12383);
or U13004 (N_13004,N_12261,N_11844);
nand U13005 (N_13005,N_10228,N_10999);
xnor U13006 (N_13006,N_10231,N_10170);
xnor U13007 (N_13007,N_11596,N_10575);
or U13008 (N_13008,N_11098,N_11407);
nand U13009 (N_13009,N_10489,N_10962);
and U13010 (N_13010,N_10508,N_12473);
nand U13011 (N_13011,N_10898,N_10474);
and U13012 (N_13012,N_11519,N_12304);
nor U13013 (N_13013,N_11692,N_12406);
nor U13014 (N_13014,N_12083,N_10468);
xnor U13015 (N_13015,N_10730,N_10590);
nor U13016 (N_13016,N_12499,N_12033);
nand U13017 (N_13017,N_10768,N_10881);
nor U13018 (N_13018,N_11197,N_11164);
or U13019 (N_13019,N_10946,N_12381);
nand U13020 (N_13020,N_11794,N_11816);
and U13021 (N_13021,N_10668,N_11636);
nor U13022 (N_13022,N_11089,N_12322);
or U13023 (N_13023,N_11338,N_12027);
nand U13024 (N_13024,N_10588,N_10343);
nand U13025 (N_13025,N_11094,N_11545);
nor U13026 (N_13026,N_11686,N_12216);
or U13027 (N_13027,N_10345,N_12276);
or U13028 (N_13028,N_10837,N_12048);
nor U13029 (N_13029,N_10285,N_12263);
nor U13030 (N_13030,N_12147,N_12150);
nand U13031 (N_13031,N_10412,N_11403);
xnor U13032 (N_13032,N_11815,N_12152);
and U13033 (N_13033,N_11284,N_11781);
or U13034 (N_13034,N_11727,N_11564);
or U13035 (N_13035,N_11765,N_11117);
or U13036 (N_13036,N_11808,N_10918);
xor U13037 (N_13037,N_11684,N_10062);
nand U13038 (N_13038,N_11109,N_10960);
nor U13039 (N_13039,N_10985,N_10776);
nor U13040 (N_13040,N_11645,N_10544);
nor U13041 (N_13041,N_10035,N_11621);
and U13042 (N_13042,N_10904,N_11973);
or U13043 (N_13043,N_11106,N_10236);
nor U13044 (N_13044,N_10636,N_10184);
xor U13045 (N_13045,N_11381,N_11321);
nor U13046 (N_13046,N_10260,N_12311);
nand U13047 (N_13047,N_11099,N_11482);
xor U13048 (N_13048,N_10584,N_10558);
and U13049 (N_13049,N_11354,N_10512);
and U13050 (N_13050,N_10484,N_10478);
nor U13051 (N_13051,N_11067,N_10507);
or U13052 (N_13052,N_10715,N_10367);
nand U13053 (N_13053,N_11776,N_10039);
and U13054 (N_13054,N_11292,N_10155);
or U13055 (N_13055,N_11958,N_11049);
and U13056 (N_13056,N_11489,N_11435);
xnor U13057 (N_13057,N_10950,N_12451);
or U13058 (N_13058,N_10129,N_12476);
xnor U13059 (N_13059,N_10296,N_10186);
nand U13060 (N_13060,N_10213,N_10909);
nor U13061 (N_13061,N_12062,N_10446);
and U13062 (N_13062,N_11282,N_11217);
xor U13063 (N_13063,N_11677,N_11616);
and U13064 (N_13064,N_11147,N_11241);
nand U13065 (N_13065,N_10795,N_10183);
and U13066 (N_13066,N_11254,N_12223);
and U13067 (N_13067,N_12044,N_10318);
nor U13068 (N_13068,N_10102,N_11789);
and U13069 (N_13069,N_12089,N_10885);
nor U13070 (N_13070,N_11688,N_11018);
xor U13071 (N_13071,N_10975,N_10862);
and U13072 (N_13072,N_12007,N_11141);
nor U13073 (N_13073,N_11060,N_10996);
nor U13074 (N_13074,N_12419,N_12274);
or U13075 (N_13075,N_10579,N_11356);
nand U13076 (N_13076,N_11357,N_10299);
or U13077 (N_13077,N_11928,N_10001);
nor U13078 (N_13078,N_12332,N_10123);
and U13079 (N_13079,N_11791,N_10156);
and U13080 (N_13080,N_10095,N_10547);
nand U13081 (N_13081,N_11222,N_11058);
nand U13082 (N_13082,N_10699,N_10577);
or U13083 (N_13083,N_11819,N_10511);
nor U13084 (N_13084,N_11464,N_11188);
nand U13085 (N_13085,N_10717,N_11457);
nor U13086 (N_13086,N_11151,N_12212);
or U13087 (N_13087,N_11511,N_10451);
or U13088 (N_13088,N_10810,N_10633);
and U13089 (N_13089,N_10866,N_11874);
xnor U13090 (N_13090,N_10727,N_11097);
or U13091 (N_13091,N_10953,N_10879);
nor U13092 (N_13092,N_11243,N_10456);
xnor U13093 (N_13093,N_10177,N_10954);
and U13094 (N_13094,N_11483,N_10206);
and U13095 (N_13095,N_11438,N_11037);
nor U13096 (N_13096,N_12019,N_10061);
nor U13097 (N_13097,N_11369,N_10818);
xnor U13098 (N_13098,N_12167,N_10600);
nand U13099 (N_13099,N_11738,N_12053);
or U13100 (N_13100,N_10135,N_11820);
nand U13101 (N_13101,N_12168,N_11171);
or U13102 (N_13102,N_10743,N_11536);
xnor U13103 (N_13103,N_11186,N_10471);
and U13104 (N_13104,N_11648,N_10963);
and U13105 (N_13105,N_11170,N_10637);
nand U13106 (N_13106,N_11148,N_11195);
and U13107 (N_13107,N_11897,N_10563);
nor U13108 (N_13108,N_11629,N_11568);
or U13109 (N_13109,N_12103,N_10372);
and U13110 (N_13110,N_10868,N_10578);
or U13111 (N_13111,N_10161,N_10033);
xnor U13112 (N_13112,N_10676,N_11899);
nor U13113 (N_13113,N_11599,N_12448);
and U13114 (N_13114,N_10848,N_11124);
nand U13115 (N_13115,N_11010,N_11609);
nor U13116 (N_13116,N_11372,N_10384);
nand U13117 (N_13117,N_11273,N_10797);
nor U13118 (N_13118,N_11780,N_10126);
xor U13119 (N_13119,N_10128,N_10151);
or U13120 (N_13120,N_11264,N_10843);
nor U13121 (N_13121,N_10705,N_10300);
or U13122 (N_13122,N_12018,N_10350);
nand U13123 (N_13123,N_12197,N_11173);
nor U13124 (N_13124,N_11571,N_12333);
nor U13125 (N_13125,N_11131,N_10068);
xor U13126 (N_13126,N_10286,N_10542);
and U13127 (N_13127,N_12105,N_12300);
nor U13128 (N_13128,N_11121,N_10277);
and U13129 (N_13129,N_10297,N_10509);
and U13130 (N_13130,N_10267,N_12282);
nand U13131 (N_13131,N_11481,N_10157);
xnor U13132 (N_13132,N_11534,N_11277);
and U13133 (N_13133,N_10210,N_12100);
xor U13134 (N_13134,N_10595,N_10686);
or U13135 (N_13135,N_10335,N_11242);
nor U13136 (N_13136,N_10087,N_11647);
nor U13137 (N_13137,N_11149,N_12494);
or U13138 (N_13138,N_11317,N_11331);
xnor U13139 (N_13139,N_10801,N_12312);
xnor U13140 (N_13140,N_10467,N_11824);
or U13141 (N_13141,N_11116,N_10159);
or U13142 (N_13142,N_12156,N_10883);
and U13143 (N_13143,N_12429,N_11274);
or U13144 (N_13144,N_11428,N_11263);
nor U13145 (N_13145,N_10506,N_11748);
and U13146 (N_13146,N_11388,N_10436);
or U13147 (N_13147,N_12444,N_11903);
nor U13148 (N_13148,N_10324,N_12123);
or U13149 (N_13149,N_10546,N_11332);
nand U13150 (N_13150,N_11052,N_12378);
nor U13151 (N_13151,N_10857,N_10245);
and U13152 (N_13152,N_11252,N_10841);
or U13153 (N_13153,N_12305,N_10359);
xor U13154 (N_13154,N_10614,N_11770);
nor U13155 (N_13155,N_12079,N_12021);
and U13156 (N_13156,N_11081,N_11340);
nand U13157 (N_13157,N_11871,N_10787);
and U13158 (N_13158,N_10392,N_11628);
nor U13159 (N_13159,N_10951,N_10799);
nand U13160 (N_13160,N_10725,N_10014);
and U13161 (N_13161,N_11699,N_11385);
xor U13162 (N_13162,N_11603,N_11059);
and U13163 (N_13163,N_10266,N_10066);
or U13164 (N_13164,N_10785,N_12340);
nor U13165 (N_13165,N_12186,N_10065);
and U13166 (N_13166,N_11634,N_10869);
nand U13167 (N_13167,N_11577,N_11092);
nand U13168 (N_13168,N_10119,N_10690);
or U13169 (N_13169,N_10569,N_10670);
or U13170 (N_13170,N_11790,N_10880);
nand U13171 (N_13171,N_10017,N_10190);
or U13172 (N_13172,N_10022,N_12288);
xor U13173 (N_13173,N_10916,N_12289);
and U13174 (N_13174,N_10978,N_12009);
and U13175 (N_13175,N_11539,N_11853);
xnor U13176 (N_13176,N_11255,N_12371);
xnor U13177 (N_13177,N_12411,N_11306);
nor U13178 (N_13178,N_11308,N_10539);
nor U13179 (N_13179,N_11342,N_12217);
xnor U13180 (N_13180,N_10360,N_10976);
or U13181 (N_13181,N_11683,N_11424);
nor U13182 (N_13182,N_10646,N_10925);
and U13183 (N_13183,N_11492,N_10408);
xor U13184 (N_13184,N_10993,N_10494);
or U13185 (N_13185,N_10399,N_10462);
and U13186 (N_13186,N_11286,N_11682);
nand U13187 (N_13187,N_11175,N_10131);
nor U13188 (N_13188,N_12404,N_11359);
xor U13189 (N_13189,N_11296,N_12165);
or U13190 (N_13190,N_12138,N_11473);
nand U13191 (N_13191,N_11883,N_11281);
nand U13192 (N_13192,N_12295,N_12334);
xnor U13193 (N_13193,N_10366,N_10442);
nand U13194 (N_13194,N_10896,N_10709);
and U13195 (N_13195,N_12281,N_10907);
xor U13196 (N_13196,N_10593,N_11391);
nand U13197 (N_13197,N_11963,N_10078);
and U13198 (N_13198,N_11445,N_11223);
and U13199 (N_13199,N_11810,N_10025);
and U13200 (N_13200,N_11219,N_10419);
xor U13201 (N_13201,N_10580,N_11394);
xor U13202 (N_13202,N_11802,N_10704);
nor U13203 (N_13203,N_11430,N_10496);
nand U13204 (N_13204,N_12350,N_11450);
nor U13205 (N_13205,N_10238,N_11211);
or U13206 (N_13206,N_11212,N_12058);
xor U13207 (N_13207,N_11954,N_11959);
nor U13208 (N_13208,N_10719,N_11017);
or U13209 (N_13209,N_12239,N_10011);
nand U13210 (N_13210,N_10720,N_11786);
or U13211 (N_13211,N_11635,N_12020);
xor U13212 (N_13212,N_10346,N_11285);
or U13213 (N_13213,N_11346,N_12255);
xor U13214 (N_13214,N_11898,N_11439);
xor U13215 (N_13215,N_10919,N_10525);
nor U13216 (N_13216,N_10731,N_10457);
or U13217 (N_13217,N_11312,N_11111);
nand U13218 (N_13218,N_12164,N_10850);
or U13219 (N_13219,N_10198,N_11714);
nor U13220 (N_13220,N_10012,N_12284);
and U13221 (N_13221,N_10644,N_10678);
nor U13222 (N_13222,N_12132,N_10373);
nand U13223 (N_13223,N_11508,N_11103);
or U13224 (N_13224,N_11016,N_11090);
and U13225 (N_13225,N_11718,N_10535);
nand U13226 (N_13226,N_10233,N_12141);
nand U13227 (N_13227,N_11812,N_12231);
and U13228 (N_13228,N_11976,N_10064);
and U13229 (N_13229,N_10652,N_10873);
nor U13230 (N_13230,N_10876,N_11867);
or U13231 (N_13231,N_11261,N_11900);
or U13232 (N_13232,N_11661,N_10167);
or U13233 (N_13233,N_12082,N_10662);
or U13234 (N_13234,N_11731,N_10317);
nor U13235 (N_13235,N_11956,N_11376);
and U13236 (N_13236,N_12184,N_10377);
and U13237 (N_13237,N_12485,N_10609);
nor U13238 (N_13238,N_11444,N_11512);
nor U13239 (N_13239,N_12353,N_12487);
nor U13240 (N_13240,N_12380,N_10171);
nor U13241 (N_13241,N_10226,N_12349);
or U13242 (N_13242,N_11806,N_12409);
nand U13243 (N_13243,N_10310,N_11749);
nor U13244 (N_13244,N_11479,N_11209);
xnor U13245 (N_13245,N_11102,N_11159);
and U13246 (N_13246,N_10781,N_10279);
nand U13247 (N_13247,N_12479,N_12339);
or U13248 (N_13248,N_11227,N_12454);
and U13249 (N_13249,N_10332,N_10606);
nor U13250 (N_13250,N_11798,N_10851);
and U13251 (N_13251,N_10138,N_12469);
nor U13252 (N_13252,N_12199,N_10307);
nor U13253 (N_13253,N_10055,N_11387);
nand U13254 (N_13254,N_11246,N_12157);
and U13255 (N_13255,N_11615,N_12057);
and U13256 (N_13256,N_11226,N_11651);
xnor U13257 (N_13257,N_11335,N_12066);
nand U13258 (N_13258,N_11044,N_11678);
or U13259 (N_13259,N_10611,N_12241);
nor U13260 (N_13260,N_11201,N_11852);
nand U13261 (N_13261,N_10247,N_10274);
and U13262 (N_13262,N_12249,N_11940);
and U13263 (N_13263,N_10647,N_10498);
nor U13264 (N_13264,N_12206,N_10553);
nor U13265 (N_13265,N_11009,N_10667);
and U13266 (N_13266,N_11238,N_12013);
or U13267 (N_13267,N_10340,N_11980);
nand U13268 (N_13268,N_12050,N_10023);
and U13269 (N_13269,N_12426,N_11882);
nor U13270 (N_13270,N_10179,N_10074);
or U13271 (N_13271,N_11601,N_11026);
xor U13272 (N_13272,N_10165,N_11875);
and U13273 (N_13273,N_10833,N_12159);
nor U13274 (N_13274,N_10141,N_10581);
nand U13275 (N_13275,N_11300,N_10669);
nand U13276 (N_13276,N_10594,N_11850);
or U13277 (N_13277,N_12302,N_10988);
nand U13278 (N_13278,N_11231,N_12106);
xor U13279 (N_13279,N_12052,N_11531);
or U13280 (N_13280,N_11413,N_10696);
and U13281 (N_13281,N_10739,N_11673);
or U13282 (N_13282,N_10982,N_11029);
nand U13283 (N_13283,N_11849,N_11879);
xor U13284 (N_13284,N_11095,N_12116);
nor U13285 (N_13285,N_12345,N_12220);
nand U13286 (N_13286,N_11614,N_11214);
nor U13287 (N_13287,N_11947,N_10906);
nand U13288 (N_13288,N_11919,N_10460);
and U13289 (N_13289,N_11494,N_10811);
nor U13290 (N_13290,N_10188,N_11598);
nor U13291 (N_13291,N_11814,N_11422);
xnor U13292 (N_13292,N_10917,N_12343);
nor U13293 (N_13293,N_11730,N_12374);
and U13294 (N_13294,N_10072,N_10745);
nand U13295 (N_13295,N_12195,N_10394);
or U13296 (N_13296,N_11797,N_11314);
nand U13297 (N_13297,N_10139,N_12271);
nand U13298 (N_13298,N_12235,N_12049);
nand U13299 (N_13299,N_12078,N_11048);
xor U13300 (N_13300,N_10374,N_11785);
xnor U13301 (N_13301,N_11502,N_10860);
nor U13302 (N_13302,N_10697,N_10640);
or U13303 (N_13303,N_10255,N_10024);
and U13304 (N_13304,N_10500,N_11475);
and U13305 (N_13305,N_12387,N_11466);
nor U13306 (N_13306,N_11643,N_12474);
or U13307 (N_13307,N_10154,N_10356);
or U13308 (N_13308,N_10191,N_12029);
xnor U13309 (N_13309,N_12443,N_11000);
xor U13310 (N_13310,N_10945,N_10327);
or U13311 (N_13311,N_10132,N_12428);
nand U13312 (N_13312,N_11912,N_11763);
nor U13313 (N_13313,N_10482,N_11461);
and U13314 (N_13314,N_10888,N_12446);
and U13315 (N_13315,N_10416,N_10166);
xor U13316 (N_13316,N_10491,N_11653);
xor U13317 (N_13317,N_10630,N_12385);
nor U13318 (N_13318,N_11515,N_10649);
or U13319 (N_13319,N_12040,N_10406);
or U13320 (N_13320,N_11265,N_11761);
and U13321 (N_13321,N_11280,N_10195);
nor U13322 (N_13322,N_10968,N_12450);
xnor U13323 (N_13323,N_10893,N_11091);
or U13324 (N_13324,N_10523,N_11951);
nor U13325 (N_13325,N_11486,N_12405);
nand U13326 (N_13326,N_12362,N_10144);
xor U13327 (N_13327,N_11528,N_11133);
or U13328 (N_13328,N_11578,N_10243);
xnor U13329 (N_13329,N_10364,N_11393);
or U13330 (N_13330,N_11799,N_10472);
or U13331 (N_13331,N_10842,N_12422);
nand U13332 (N_13332,N_10347,N_11156);
nor U13333 (N_13333,N_11809,N_11735);
nand U13334 (N_13334,N_10309,N_11752);
and U13335 (N_13335,N_10821,N_11390);
xor U13336 (N_13336,N_12318,N_12237);
xor U13337 (N_13337,N_11045,N_12031);
or U13338 (N_13338,N_10415,N_11756);
nor U13339 (N_13339,N_10479,N_10295);
nand U13340 (N_13340,N_11220,N_10041);
or U13341 (N_13341,N_11580,N_10672);
xnor U13342 (N_13342,N_11337,N_11493);
and U13343 (N_13343,N_10153,N_11716);
xnor U13344 (N_13344,N_11032,N_12269);
nand U13345 (N_13345,N_11746,N_11490);
nand U13346 (N_13346,N_10856,N_11914);
or U13347 (N_13347,N_10212,N_11836);
xor U13348 (N_13348,N_11194,N_10565);
and U13349 (N_13349,N_10846,N_11216);
or U13350 (N_13350,N_12456,N_11602);
and U13351 (N_13351,N_11127,N_10803);
and U13352 (N_13352,N_11425,N_12298);
or U13353 (N_13353,N_11135,N_10897);
and U13354 (N_13354,N_10751,N_11467);
xor U13355 (N_13355,N_11070,N_12030);
and U13356 (N_13356,N_11215,N_12086);
xnor U13357 (N_13357,N_11926,N_12327);
xor U13358 (N_13358,N_10513,N_12128);
nor U13359 (N_13359,N_11447,N_12166);
or U13360 (N_13360,N_12356,N_10536);
xor U13361 (N_13361,N_10657,N_10121);
and U13362 (N_13362,N_11025,N_10127);
or U13363 (N_13363,N_11380,N_10932);
or U13364 (N_13364,N_12299,N_10656);
nor U13365 (N_13365,N_10530,N_11729);
xnor U13366 (N_13366,N_11793,N_10566);
xor U13367 (N_13367,N_11676,N_11529);
and U13368 (N_13368,N_11753,N_10551);
and U13369 (N_13369,N_10302,N_11702);
nand U13370 (N_13370,N_12285,N_10560);
nor U13371 (N_13371,N_11607,N_10338);
nand U13372 (N_13372,N_10303,N_11155);
and U13373 (N_13373,N_10555,N_11142);
xor U13374 (N_13374,N_11344,N_12463);
xnor U13375 (N_13375,N_11488,N_10097);
nand U13376 (N_13376,N_11541,N_11967);
nand U13377 (N_13377,N_10926,N_10004);
or U13378 (N_13378,N_11915,N_10096);
nor U13379 (N_13379,N_10562,N_10867);
or U13380 (N_13380,N_12329,N_12370);
xor U13381 (N_13381,N_10554,N_10027);
or U13382 (N_13382,N_11072,N_10276);
xnor U13383 (N_13383,N_10396,N_11741);
and U13384 (N_13384,N_11840,N_10761);
xor U13385 (N_13385,N_11991,N_10443);
nor U13386 (N_13386,N_10291,N_12436);
xor U13387 (N_13387,N_10625,N_10796);
xnor U13388 (N_13388,N_10168,N_12014);
or U13389 (N_13389,N_11276,N_11544);
and U13390 (N_13390,N_10108,N_10242);
xnor U13391 (N_13391,N_11779,N_11392);
nor U13392 (N_13392,N_10826,N_12187);
xor U13393 (N_13393,N_12070,N_12153);
xor U13394 (N_13394,N_12408,N_11996);
and U13395 (N_13395,N_10169,N_12077);
nor U13396 (N_13396,N_11358,N_10404);
nand U13397 (N_13397,N_11892,N_11020);
xnor U13398 (N_13398,N_10939,N_11521);
xnor U13399 (N_13399,N_11316,N_10902);
xor U13400 (N_13400,N_11788,N_11210);
or U13401 (N_13401,N_11013,N_11993);
xnor U13402 (N_13402,N_11406,N_11144);
nor U13403 (N_13403,N_10887,N_10477);
nor U13404 (N_13404,N_11446,N_11842);
nor U13405 (N_13405,N_11082,N_10103);
or U13406 (N_13406,N_11379,N_10712);
nand U13407 (N_13407,N_11990,N_11104);
nor U13408 (N_13408,N_10716,N_10984);
and U13409 (N_13409,N_11259,N_11565);
nand U13410 (N_13410,N_10223,N_10973);
nand U13411 (N_13411,N_10085,N_10923);
and U13412 (N_13412,N_10314,N_11021);
xor U13413 (N_13413,N_10187,N_11859);
or U13414 (N_13414,N_12388,N_12096);
nand U13415 (N_13415,N_10125,N_10990);
xor U13416 (N_13416,N_11944,N_12458);
nand U13417 (N_13417,N_11663,N_12142);
or U13418 (N_13418,N_12398,N_11640);
xor U13419 (N_13419,N_12101,N_10026);
or U13420 (N_13420,N_12482,N_10514);
xor U13421 (N_13421,N_11619,N_10871);
or U13422 (N_13422,N_12498,N_10533);
or U13423 (N_13423,N_10561,N_11345);
or U13424 (N_13424,N_12196,N_10823);
or U13425 (N_13425,N_10009,N_11717);
and U13426 (N_13426,N_12001,N_10005);
nor U13427 (N_13427,N_10420,N_11509);
and U13428 (N_13428,N_10708,N_10414);
nand U13429 (N_13429,N_11665,N_12146);
nand U13430 (N_13430,N_10780,N_11449);
nand U13431 (N_13431,N_11310,N_11448);
or U13432 (N_13432,N_10980,N_10458);
nor U13433 (N_13433,N_10940,N_11817);
nand U13434 (N_13434,N_10596,N_11294);
xor U13435 (N_13435,N_12210,N_10052);
or U13436 (N_13436,N_10013,N_10773);
nor U13437 (N_13437,N_10455,N_10312);
nor U13438 (N_13438,N_10434,N_10092);
or U13439 (N_13439,N_12124,N_10293);
or U13440 (N_13440,N_10618,N_10400);
xnor U13441 (N_13441,N_10619,N_11122);
nand U13442 (N_13442,N_10849,N_10217);
nor U13443 (N_13443,N_11233,N_12085);
xnor U13444 (N_13444,N_10677,N_11311);
or U13445 (N_13445,N_10250,N_10469);
xnor U13446 (N_13446,N_10237,N_10270);
or U13447 (N_13447,N_11579,N_10505);
and U13448 (N_13448,N_10608,N_11476);
nor U13449 (N_13449,N_10390,N_11880);
nor U13450 (N_13450,N_11334,N_12425);
and U13451 (N_13451,N_10099,N_12224);
xnor U13452 (N_13452,N_10992,N_10427);
xor U13453 (N_13453,N_10336,N_10613);
and U13454 (N_13454,N_11703,N_12401);
or U13455 (N_13455,N_10793,N_11664);
and U13456 (N_13456,N_11328,N_10202);
xor U13457 (N_13457,N_12026,N_11893);
nor U13458 (N_13458,N_11251,N_10610);
and U13459 (N_13459,N_10886,N_12016);
nand U13460 (N_13460,N_11283,N_11066);
and U13461 (N_13461,N_10257,N_10910);
nor U13462 (N_13462,N_11235,N_11627);
nand U13463 (N_13463,N_10421,N_10700);
nor U13464 (N_13464,N_12039,N_11533);
and U13465 (N_13465,N_11112,N_11313);
and U13466 (N_13466,N_10115,N_10424);
xnor U13467 (N_13467,N_11586,N_10503);
and U13468 (N_13468,N_10145,N_12028);
or U13469 (N_13469,N_11043,N_11484);
nand U13470 (N_13470,N_11289,N_12243);
nand U13471 (N_13471,N_11823,N_11658);
xnor U13472 (N_13472,N_10323,N_12115);
and U13473 (N_13473,N_12177,N_10830);
and U13474 (N_13474,N_10772,N_10259);
or U13475 (N_13475,N_10944,N_10215);
and U13476 (N_13476,N_10134,N_12238);
xor U13477 (N_13477,N_12042,N_11581);
xor U13478 (N_13478,N_12471,N_10251);
xor U13479 (N_13479,N_11184,N_11795);
or U13480 (N_13480,N_11318,N_10805);
nand U13481 (N_13481,N_11965,N_11873);
or U13482 (N_13482,N_12119,N_11745);
xnor U13483 (N_13483,N_11932,N_10353);
and U13484 (N_13484,N_12245,N_10298);
nand U13485 (N_13485,N_10952,N_11851);
nand U13486 (N_13486,N_12427,N_11140);
xor U13487 (N_13487,N_11039,N_10090);
nor U13488 (N_13488,N_11373,N_12309);
and U13489 (N_13489,N_10612,N_10790);
or U13490 (N_13490,N_11807,N_11590);
and U13491 (N_13491,N_11833,N_10711);
nor U13492 (N_13492,N_12314,N_11946);
and U13493 (N_13493,N_10585,N_10819);
and U13494 (N_13494,N_11499,N_12402);
or U13495 (N_13495,N_10941,N_10882);
xor U13496 (N_13496,N_10789,N_10855);
nand U13497 (N_13497,N_10531,N_10178);
and U13498 (N_13498,N_12003,N_10264);
xnor U13499 (N_13499,N_12363,N_11909);
xor U13500 (N_13500,N_10895,N_11527);
nor U13501 (N_13501,N_11420,N_11837);
nand U13502 (N_13502,N_10956,N_10137);
nor U13503 (N_13503,N_11828,N_12225);
or U13504 (N_13504,N_10586,N_11015);
nor U13505 (N_13505,N_11945,N_11011);
xor U13506 (N_13506,N_11821,N_12213);
and U13507 (N_13507,N_10162,N_10105);
nor U13508 (N_13508,N_10792,N_11574);
or U13509 (N_13509,N_11920,N_12259);
nand U13510 (N_13510,N_10348,N_10283);
and U13511 (N_13511,N_12204,N_10281);
xor U13512 (N_13512,N_10765,N_11295);
or U13513 (N_13513,N_12310,N_10798);
xnor U13514 (N_13514,N_12160,N_12365);
and U13515 (N_13515,N_11024,N_11896);
xnor U13516 (N_13516,N_11706,N_11985);
nand U13517 (N_13517,N_10256,N_11405);
nand U13518 (N_13518,N_10110,N_10938);
xor U13519 (N_13519,N_10160,N_10534);
or U13520 (N_13520,N_11119,N_10203);
or U13521 (N_13521,N_11145,N_11969);
xnor U13522 (N_13522,N_10769,N_10045);
or U13523 (N_13523,N_12480,N_11256);
and U13524 (N_13524,N_11078,N_12006);
nor U13525 (N_13525,N_12368,N_11404);
xor U13526 (N_13526,N_11986,N_12253);
nand U13527 (N_13527,N_10107,N_11690);
or U13528 (N_13528,N_11925,N_10518);
xor U13529 (N_13529,N_10645,N_10692);
nor U13530 (N_13530,N_11681,N_10089);
xor U13531 (N_13531,N_10036,N_10994);
xor U13532 (N_13532,N_12087,N_11845);
nand U13533 (N_13533,N_11177,N_12074);
nor U13534 (N_13534,N_12438,N_12176);
and U13535 (N_13535,N_10501,N_12392);
nor U13536 (N_13536,N_10891,N_11918);
and U13537 (N_13537,N_10541,N_12022);
and U13538 (N_13538,N_10754,N_11320);
nor U13539 (N_13539,N_10461,N_11019);
xor U13540 (N_13540,N_10308,N_11723);
nor U13541 (N_13541,N_11304,N_12043);
nor U13542 (N_13542,N_11418,N_11431);
nand U13543 (N_13543,N_10591,N_10194);
or U13544 (N_13544,N_11543,N_11709);
nor U13545 (N_13545,N_12205,N_10736);
and U13546 (N_13546,N_10698,N_10822);
xor U13547 (N_13547,N_10573,N_10476);
nand U13548 (N_13548,N_12262,N_12064);
or U13549 (N_13549,N_10182,N_10069);
or U13550 (N_13550,N_12497,N_12481);
xor U13551 (N_13551,N_10859,N_11360);
nand U13552 (N_13552,N_10319,N_10204);
and U13553 (N_13553,N_10104,N_12060);
and U13554 (N_13554,N_11433,N_10007);
or U13555 (N_13555,N_11006,N_11355);
xor U13556 (N_13556,N_10265,N_11160);
nor U13557 (N_13557,N_10673,N_11437);
nor U13558 (N_13558,N_10642,N_10059);
xnor U13559 (N_13559,N_11998,N_11695);
or U13560 (N_13560,N_11165,N_10570);
or U13561 (N_13561,N_12108,N_10164);
and U13562 (N_13562,N_10287,N_11612);
or U13563 (N_13563,N_10583,N_11584);
xor U13564 (N_13564,N_11960,N_10935);
nor U13565 (N_13565,N_10398,N_10734);
nor U13566 (N_13566,N_11408,N_10905);
and U13567 (N_13567,N_12400,N_10405);
or U13568 (N_13568,N_11076,N_11221);
and U13569 (N_13569,N_11671,N_11822);
nand U13570 (N_13570,N_11698,N_11530);
nor U13571 (N_13571,N_12328,N_12180);
nand U13572 (N_13572,N_10003,N_10397);
xor U13573 (N_13573,N_10329,N_10146);
nand U13574 (N_13574,N_12326,N_11835);
xor U13575 (N_13575,N_11022,N_10972);
or U13576 (N_13576,N_11704,N_12170);
and U13577 (N_13577,N_12037,N_10444);
or U13578 (N_13578,N_10865,N_11514);
nor U13579 (N_13579,N_10631,N_10936);
xnor U13580 (N_13580,N_10839,N_10528);
nor U13581 (N_13581,N_11303,N_11962);
nor U13582 (N_13582,N_10820,N_11694);
nor U13583 (N_13583,N_12233,N_11768);
nand U13584 (N_13584,N_11129,N_10447);
nor U13585 (N_13585,N_10306,N_10208);
or U13586 (N_13586,N_10816,N_12092);
nand U13587 (N_13587,N_10814,N_11513);
xor U13588 (N_13588,N_10339,N_12008);
or U13589 (N_13589,N_12290,N_11329);
xor U13590 (N_13590,N_12325,N_12460);
nor U13591 (N_13591,N_11236,N_10031);
xor U13592 (N_13592,N_11178,N_10812);
nor U13593 (N_13593,N_11569,N_10601);
nand U13594 (N_13594,N_12486,N_11554);
nand U13595 (N_13595,N_10409,N_12203);
and U13596 (N_13596,N_10680,N_12287);
xor U13597 (N_13597,N_11249,N_10748);
or U13598 (N_13598,N_11981,N_10766);
nand U13599 (N_13599,N_11540,N_12386);
or U13600 (N_13600,N_12080,N_12182);
or U13601 (N_13601,N_11307,N_11551);
nand U13602 (N_13602,N_10746,N_10304);
and U13603 (N_13603,N_10622,N_11680);
xnor U13604 (N_13604,N_11642,N_10703);
nor U13605 (N_13605,N_10147,N_10486);
nor U13606 (N_13606,N_10098,N_12442);
or U13607 (N_13607,N_10269,N_11613);
nor U13608 (N_13608,N_11079,N_11154);
nor U13609 (N_13609,N_10088,N_12112);
nor U13610 (N_13610,N_10930,N_11916);
or U13611 (N_13611,N_11352,N_11759);
and U13612 (N_13612,N_12218,N_10032);
nand U13613 (N_13613,N_12397,N_12490);
and U13614 (N_13614,N_10218,N_11349);
nand U13615 (N_13615,N_11108,N_10341);
nand U13616 (N_13616,N_10571,N_10545);
xor U13617 (N_13617,N_11970,N_12118);
xor U13618 (N_13618,N_10076,N_12283);
xnor U13619 (N_13619,N_10316,N_12114);
nor U13620 (N_13620,N_10607,N_11870);
and U13621 (N_13621,N_12222,N_10426);
xor U13622 (N_13622,N_12483,N_11174);
xor U13623 (N_13623,N_11370,N_11053);
nor U13624 (N_13624,N_11213,N_10006);
xnor U13625 (N_13625,N_10475,N_11071);
nand U13626 (N_13626,N_10515,N_11258);
nand U13627 (N_13627,N_10333,N_12024);
and U13628 (N_13628,N_10209,N_11137);
xnor U13629 (N_13629,N_10942,N_10386);
xnor U13630 (N_13630,N_11762,N_11711);
nand U13631 (N_13631,N_10483,N_11443);
nor U13632 (N_13632,N_10664,N_10495);
and U13633 (N_13633,N_12163,N_11417);
or U13634 (N_13634,N_11732,N_10389);
xor U13635 (N_13635,N_10355,N_11377);
or U13636 (N_13636,N_11626,N_12047);
and U13637 (N_13637,N_12464,N_11941);
nor U13638 (N_13638,N_11267,N_10292);
xor U13639 (N_13639,N_12232,N_10499);
and U13640 (N_13640,N_10172,N_10784);
or U13641 (N_13641,N_11689,N_10970);
nor U13642 (N_13642,N_11088,N_11279);
and U13643 (N_13643,N_10592,N_10368);
and U13644 (N_13644,N_11592,N_11205);
nand U13645 (N_13645,N_11459,N_11383);
nand U13646 (N_13646,N_12393,N_11582);
nand U13647 (N_13647,N_12012,N_11118);
and U13648 (N_13648,N_11876,N_11691);
nor U13649 (N_13649,N_10621,N_11305);
nand U13650 (N_13650,N_11353,N_11469);
or U13651 (N_13651,N_12081,N_11505);
and U13652 (N_13652,N_10840,N_11125);
and U13653 (N_13653,N_11905,N_12200);
or U13654 (N_13654,N_11470,N_11401);
or U13655 (N_13655,N_10915,N_11670);
nand U13656 (N_13656,N_10010,N_10211);
and U13657 (N_13657,N_10681,N_10958);
xor U13658 (N_13658,N_10351,N_12144);
or U13659 (N_13659,N_11202,N_10222);
nand U13660 (N_13660,N_11061,N_12010);
or U13661 (N_13661,N_11245,N_10615);
nand U13662 (N_13662,N_12420,N_10481);
xnor U13663 (N_13663,N_11035,N_12418);
nor U13664 (N_13664,N_11465,N_11224);
xor U13665 (N_13665,N_10654,N_10809);
xnor U13666 (N_13666,N_11722,N_12358);
nand U13667 (N_13667,N_12292,N_12359);
or U13668 (N_13668,N_11299,N_11005);
nor U13669 (N_13669,N_10983,N_10875);
and U13670 (N_13670,N_11805,N_12453);
nor U13671 (N_13671,N_10921,N_11426);
xor U13672 (N_13672,N_12455,N_12161);
or U13673 (N_13673,N_11848,N_11501);
and U13674 (N_13674,N_10273,N_11250);
nand U13675 (N_13675,N_11847,N_11432);
or U13676 (N_13676,N_10576,N_11441);
or U13677 (N_13677,N_11696,N_11191);
nand U13678 (N_13678,N_10492,N_12202);
nand U13679 (N_13679,N_11498,N_10083);
and U13680 (N_13680,N_11622,N_11886);
or U13681 (N_13681,N_10063,N_10648);
nor U13682 (N_13682,N_11269,N_12169);
nand U13683 (N_13683,N_10997,N_10529);
nand U13684 (N_13684,N_12296,N_10806);
and U13685 (N_13685,N_12260,N_10661);
or U13686 (N_13686,N_10402,N_10516);
xnor U13687 (N_13687,N_12431,N_11668);
nor U13688 (N_13688,N_10732,N_10403);
xnor U13689 (N_13689,N_10142,N_10683);
or U13690 (N_13690,N_11057,N_12090);
or U13691 (N_13691,N_11988,N_11322);
xnor U13692 (N_13692,N_10844,N_10779);
and U13693 (N_13693,N_12376,N_10365);
nor U13694 (N_13694,N_11719,N_10352);
xor U13695 (N_13695,N_11957,N_12155);
nor U13696 (N_13696,N_10480,N_10845);
or U13697 (N_13697,N_12466,N_10729);
and U13698 (N_13698,N_12275,N_10948);
nor U13699 (N_13699,N_10305,N_10977);
nand U13700 (N_13700,N_11611,N_10046);
nor U13701 (N_13701,N_10488,N_10783);
nand U13702 (N_13702,N_10989,N_11975);
or U13703 (N_13703,N_10737,N_10937);
nor U13704 (N_13704,N_10957,N_11384);
xor U13705 (N_13705,N_10073,N_10284);
nand U13706 (N_13706,N_11608,N_11862);
nor U13707 (N_13707,N_11597,N_10964);
nor U13708 (N_13708,N_10084,N_10249);
nor U13709 (N_13709,N_10764,N_11179);
or U13710 (N_13710,N_10114,N_11247);
nor U13711 (N_13711,N_11983,N_11176);
nand U13712 (N_13712,N_12137,N_11402);
and U13713 (N_13713,N_10133,N_10464);
xnor U13714 (N_13714,N_10425,N_10124);
and U13715 (N_13715,N_10328,N_10981);
nor U13716 (N_13716,N_10321,N_11364);
or U13717 (N_13717,N_11992,N_11132);
and U13718 (N_13718,N_10418,N_10659);
nor U13719 (N_13719,N_12017,N_12102);
xor U13720 (N_13720,N_12173,N_11272);
nor U13721 (N_13721,N_11846,N_10362);
and U13722 (N_13722,N_11397,N_10605);
nand U13723 (N_13723,N_12059,N_10617);
and U13724 (N_13724,N_12331,N_11708);
and U13725 (N_13725,N_11901,N_11257);
and U13726 (N_13726,N_11146,N_12346);
xor U13727 (N_13727,N_10429,N_11701);
xor U13728 (N_13728,N_10658,N_12488);
nand U13729 (N_13729,N_11854,N_10858);
and U13730 (N_13730,N_11399,N_11427);
nand U13731 (N_13731,N_11050,N_11415);
xnor U13732 (N_13732,N_10689,N_11487);
or U13733 (N_13733,N_12433,N_10325);
and U13734 (N_13734,N_11743,N_10552);
xnor U13735 (N_13735,N_11361,N_10465);
xnor U13736 (N_13736,N_12091,N_10028);
nor U13737 (N_13737,N_10900,N_12211);
nand U13738 (N_13738,N_10148,N_10574);
nand U13739 (N_13739,N_10357,N_11374);
or U13740 (N_13740,N_11831,N_11208);
nand U13741 (N_13741,N_11085,N_10334);
nor U13742 (N_13742,N_10375,N_10450);
xor U13743 (N_13743,N_11262,N_10524);
nor U13744 (N_13744,N_10120,N_11921);
and U13745 (N_13745,N_10802,N_10361);
nand U13746 (N_13746,N_11742,N_11589);
xnor U13747 (N_13747,N_10521,N_11535);
nand U13748 (N_13748,N_11573,N_11796);
and U13749 (N_13749,N_10791,N_11977);
nand U13750 (N_13750,N_12059,N_10634);
nand U13751 (N_13751,N_12239,N_11776);
or U13752 (N_13752,N_11683,N_11182);
or U13753 (N_13753,N_10443,N_10038);
nor U13754 (N_13754,N_11263,N_11627);
xnor U13755 (N_13755,N_10392,N_11063);
or U13756 (N_13756,N_11160,N_11475);
xor U13757 (N_13757,N_11854,N_10014);
nor U13758 (N_13758,N_12095,N_10042);
nand U13759 (N_13759,N_11046,N_12448);
and U13760 (N_13760,N_11894,N_11124);
and U13761 (N_13761,N_10496,N_12309);
xnor U13762 (N_13762,N_11402,N_10422);
nor U13763 (N_13763,N_10183,N_12092);
nor U13764 (N_13764,N_10965,N_11397);
nand U13765 (N_13765,N_10798,N_11452);
or U13766 (N_13766,N_12045,N_12415);
nor U13767 (N_13767,N_11334,N_11678);
nor U13768 (N_13768,N_11184,N_10323);
nor U13769 (N_13769,N_11047,N_11333);
and U13770 (N_13770,N_12241,N_12486);
and U13771 (N_13771,N_12332,N_11836);
nor U13772 (N_13772,N_11084,N_11684);
and U13773 (N_13773,N_11720,N_12477);
nand U13774 (N_13774,N_10867,N_10335);
and U13775 (N_13775,N_12093,N_10574);
nand U13776 (N_13776,N_10343,N_10043);
xnor U13777 (N_13777,N_10502,N_11311);
and U13778 (N_13778,N_11302,N_10907);
nand U13779 (N_13779,N_11537,N_12375);
nand U13780 (N_13780,N_10290,N_11774);
xor U13781 (N_13781,N_11626,N_12404);
and U13782 (N_13782,N_10686,N_10458);
or U13783 (N_13783,N_12158,N_12032);
nand U13784 (N_13784,N_10860,N_12379);
and U13785 (N_13785,N_11460,N_11981);
nor U13786 (N_13786,N_10661,N_10551);
xor U13787 (N_13787,N_10955,N_10001);
or U13788 (N_13788,N_12299,N_12055);
nand U13789 (N_13789,N_11417,N_10518);
and U13790 (N_13790,N_11822,N_12273);
nor U13791 (N_13791,N_11117,N_10821);
nand U13792 (N_13792,N_10054,N_11075);
or U13793 (N_13793,N_11554,N_11837);
or U13794 (N_13794,N_10276,N_10743);
xnor U13795 (N_13795,N_11861,N_11916);
and U13796 (N_13796,N_11864,N_10513);
nor U13797 (N_13797,N_10714,N_11741);
nor U13798 (N_13798,N_10695,N_10918);
nand U13799 (N_13799,N_12063,N_10589);
or U13800 (N_13800,N_11354,N_11853);
or U13801 (N_13801,N_10676,N_11424);
or U13802 (N_13802,N_12282,N_10397);
nand U13803 (N_13803,N_11429,N_10120);
xnor U13804 (N_13804,N_12309,N_10718);
xor U13805 (N_13805,N_11679,N_10992);
or U13806 (N_13806,N_11227,N_11319);
nand U13807 (N_13807,N_11085,N_11859);
nor U13808 (N_13808,N_11078,N_12230);
xnor U13809 (N_13809,N_10854,N_10659);
nor U13810 (N_13810,N_12202,N_11439);
and U13811 (N_13811,N_11934,N_10764);
or U13812 (N_13812,N_10833,N_10474);
or U13813 (N_13813,N_10854,N_10866);
xor U13814 (N_13814,N_12494,N_11480);
nand U13815 (N_13815,N_11532,N_10915);
xnor U13816 (N_13816,N_12407,N_10797);
or U13817 (N_13817,N_10728,N_11675);
or U13818 (N_13818,N_11441,N_11223);
nand U13819 (N_13819,N_10984,N_11208);
or U13820 (N_13820,N_10773,N_11356);
or U13821 (N_13821,N_10298,N_10118);
nor U13822 (N_13822,N_10721,N_10565);
xnor U13823 (N_13823,N_10807,N_10244);
nand U13824 (N_13824,N_10107,N_10912);
and U13825 (N_13825,N_10299,N_10700);
xnor U13826 (N_13826,N_11539,N_11341);
or U13827 (N_13827,N_10765,N_12124);
or U13828 (N_13828,N_11026,N_11166);
xnor U13829 (N_13829,N_11678,N_10592);
nand U13830 (N_13830,N_10018,N_12145);
xnor U13831 (N_13831,N_12399,N_10526);
xor U13832 (N_13832,N_11818,N_11503);
nor U13833 (N_13833,N_12153,N_11031);
and U13834 (N_13834,N_12412,N_12444);
or U13835 (N_13835,N_10521,N_11912);
or U13836 (N_13836,N_11440,N_11926);
nor U13837 (N_13837,N_10462,N_11411);
and U13838 (N_13838,N_10859,N_10752);
nor U13839 (N_13839,N_11051,N_11243);
and U13840 (N_13840,N_10338,N_10238);
nor U13841 (N_13841,N_12121,N_11707);
nand U13842 (N_13842,N_10881,N_12262);
nand U13843 (N_13843,N_12454,N_11885);
and U13844 (N_13844,N_11367,N_11334);
nor U13845 (N_13845,N_10769,N_10503);
nor U13846 (N_13846,N_11933,N_10249);
nor U13847 (N_13847,N_11755,N_11314);
xnor U13848 (N_13848,N_10055,N_10367);
xnor U13849 (N_13849,N_11679,N_11814);
and U13850 (N_13850,N_12280,N_12324);
or U13851 (N_13851,N_10291,N_10376);
nand U13852 (N_13852,N_10593,N_11819);
xnor U13853 (N_13853,N_10534,N_12095);
xor U13854 (N_13854,N_11967,N_11889);
and U13855 (N_13855,N_10480,N_10848);
and U13856 (N_13856,N_12354,N_11032);
nor U13857 (N_13857,N_12106,N_10331);
xor U13858 (N_13858,N_11919,N_10267);
and U13859 (N_13859,N_11615,N_12378);
and U13860 (N_13860,N_10994,N_11689);
and U13861 (N_13861,N_10475,N_12064);
or U13862 (N_13862,N_12128,N_10927);
nor U13863 (N_13863,N_12385,N_10559);
or U13864 (N_13864,N_11772,N_11764);
or U13865 (N_13865,N_10471,N_10315);
xnor U13866 (N_13866,N_11187,N_10996);
nor U13867 (N_13867,N_10898,N_11095);
nor U13868 (N_13868,N_10648,N_10003);
nor U13869 (N_13869,N_10508,N_10294);
nand U13870 (N_13870,N_12208,N_10507);
nand U13871 (N_13871,N_12086,N_11634);
xor U13872 (N_13872,N_10737,N_12329);
nand U13873 (N_13873,N_11493,N_12081);
and U13874 (N_13874,N_11008,N_12046);
or U13875 (N_13875,N_10849,N_10597);
or U13876 (N_13876,N_11517,N_10245);
and U13877 (N_13877,N_11516,N_11826);
or U13878 (N_13878,N_10064,N_11802);
nor U13879 (N_13879,N_10980,N_10567);
and U13880 (N_13880,N_11778,N_11151);
and U13881 (N_13881,N_12026,N_10909);
xor U13882 (N_13882,N_10009,N_11032);
nor U13883 (N_13883,N_11938,N_12421);
nor U13884 (N_13884,N_10454,N_11756);
and U13885 (N_13885,N_12227,N_10123);
xor U13886 (N_13886,N_10471,N_12419);
nand U13887 (N_13887,N_11991,N_12167);
xor U13888 (N_13888,N_12340,N_12381);
and U13889 (N_13889,N_10810,N_11240);
and U13890 (N_13890,N_10288,N_11491);
xor U13891 (N_13891,N_10534,N_12498);
nor U13892 (N_13892,N_11707,N_10988);
nand U13893 (N_13893,N_10544,N_11871);
nor U13894 (N_13894,N_11773,N_10273);
or U13895 (N_13895,N_11956,N_11049);
nand U13896 (N_13896,N_10998,N_10773);
xnor U13897 (N_13897,N_10260,N_11811);
nor U13898 (N_13898,N_11223,N_11259);
or U13899 (N_13899,N_12296,N_11759);
xor U13900 (N_13900,N_11745,N_11110);
and U13901 (N_13901,N_11498,N_11926);
nand U13902 (N_13902,N_10692,N_12030);
or U13903 (N_13903,N_11839,N_10629);
nand U13904 (N_13904,N_11983,N_10769);
and U13905 (N_13905,N_11841,N_12323);
xor U13906 (N_13906,N_10196,N_10709);
xor U13907 (N_13907,N_11748,N_10664);
nor U13908 (N_13908,N_11573,N_10557);
xnor U13909 (N_13909,N_10795,N_12093);
xor U13910 (N_13910,N_12029,N_10535);
and U13911 (N_13911,N_11832,N_10910);
or U13912 (N_13912,N_11420,N_12312);
xnor U13913 (N_13913,N_11084,N_10497);
nor U13914 (N_13914,N_10484,N_12435);
xnor U13915 (N_13915,N_10058,N_11411);
or U13916 (N_13916,N_10872,N_10442);
nor U13917 (N_13917,N_10701,N_10847);
and U13918 (N_13918,N_11744,N_10245);
xnor U13919 (N_13919,N_10145,N_11614);
and U13920 (N_13920,N_11309,N_12157);
nand U13921 (N_13921,N_12329,N_11615);
nor U13922 (N_13922,N_11196,N_10287);
nand U13923 (N_13923,N_10484,N_10181);
xnor U13924 (N_13924,N_11520,N_11689);
xor U13925 (N_13925,N_11416,N_10591);
xnor U13926 (N_13926,N_11258,N_12160);
nor U13927 (N_13927,N_10820,N_11613);
nand U13928 (N_13928,N_12058,N_10075);
nand U13929 (N_13929,N_12394,N_11363);
xnor U13930 (N_13930,N_10560,N_10387);
nand U13931 (N_13931,N_11256,N_11854);
and U13932 (N_13932,N_11202,N_10903);
nand U13933 (N_13933,N_11711,N_10518);
nor U13934 (N_13934,N_12191,N_10265);
or U13935 (N_13935,N_11724,N_10470);
or U13936 (N_13936,N_10072,N_11566);
xor U13937 (N_13937,N_10911,N_11642);
nor U13938 (N_13938,N_11369,N_10658);
nand U13939 (N_13939,N_10822,N_12149);
nor U13940 (N_13940,N_10560,N_11642);
xnor U13941 (N_13941,N_12029,N_11908);
or U13942 (N_13942,N_11873,N_10736);
or U13943 (N_13943,N_11527,N_11640);
nor U13944 (N_13944,N_11419,N_10927);
nor U13945 (N_13945,N_10269,N_10486);
xor U13946 (N_13946,N_12008,N_10932);
xor U13947 (N_13947,N_12276,N_10578);
or U13948 (N_13948,N_10620,N_11084);
and U13949 (N_13949,N_10954,N_11060);
or U13950 (N_13950,N_10622,N_10795);
xor U13951 (N_13951,N_10992,N_11408);
nand U13952 (N_13952,N_10797,N_11962);
nor U13953 (N_13953,N_10772,N_10540);
xnor U13954 (N_13954,N_11443,N_10622);
nand U13955 (N_13955,N_11290,N_11189);
nor U13956 (N_13956,N_10872,N_11675);
nand U13957 (N_13957,N_11134,N_10317);
nor U13958 (N_13958,N_10521,N_12273);
and U13959 (N_13959,N_11542,N_10344);
nor U13960 (N_13960,N_11690,N_10925);
and U13961 (N_13961,N_11304,N_11997);
nor U13962 (N_13962,N_12229,N_12140);
xor U13963 (N_13963,N_12140,N_12103);
xor U13964 (N_13964,N_12241,N_10660);
and U13965 (N_13965,N_10815,N_10267);
nor U13966 (N_13966,N_11351,N_10320);
xor U13967 (N_13967,N_10662,N_10618);
nand U13968 (N_13968,N_11098,N_10177);
or U13969 (N_13969,N_11116,N_11000);
nor U13970 (N_13970,N_11137,N_12465);
nand U13971 (N_13971,N_10025,N_11996);
xor U13972 (N_13972,N_11496,N_11945);
xor U13973 (N_13973,N_10844,N_11696);
and U13974 (N_13974,N_11129,N_12223);
or U13975 (N_13975,N_11257,N_10744);
and U13976 (N_13976,N_11921,N_10195);
nand U13977 (N_13977,N_10296,N_10463);
nand U13978 (N_13978,N_10414,N_11644);
and U13979 (N_13979,N_11460,N_10242);
xnor U13980 (N_13980,N_12165,N_10218);
xor U13981 (N_13981,N_10516,N_11155);
and U13982 (N_13982,N_12106,N_10383);
nand U13983 (N_13983,N_12258,N_11838);
nand U13984 (N_13984,N_11589,N_10352);
nand U13985 (N_13985,N_12152,N_11450);
nor U13986 (N_13986,N_10180,N_10733);
or U13987 (N_13987,N_11568,N_11167);
nor U13988 (N_13988,N_11390,N_10187);
nand U13989 (N_13989,N_11851,N_11667);
and U13990 (N_13990,N_11196,N_12303);
and U13991 (N_13991,N_11755,N_12393);
or U13992 (N_13992,N_11036,N_12349);
nand U13993 (N_13993,N_10435,N_11634);
xnor U13994 (N_13994,N_11459,N_10578);
or U13995 (N_13995,N_11282,N_12249);
nor U13996 (N_13996,N_11781,N_11969);
nor U13997 (N_13997,N_12362,N_10528);
nor U13998 (N_13998,N_11962,N_11204);
or U13999 (N_13999,N_10596,N_10040);
nand U14000 (N_14000,N_10275,N_10746);
or U14001 (N_14001,N_12033,N_12104);
or U14002 (N_14002,N_11610,N_11367);
nor U14003 (N_14003,N_11804,N_10300);
and U14004 (N_14004,N_11826,N_12493);
or U14005 (N_14005,N_10579,N_11460);
and U14006 (N_14006,N_11064,N_10536);
xnor U14007 (N_14007,N_10993,N_11916);
and U14008 (N_14008,N_10272,N_11918);
xnor U14009 (N_14009,N_12157,N_12015);
or U14010 (N_14010,N_11829,N_10748);
nor U14011 (N_14011,N_12429,N_11469);
nor U14012 (N_14012,N_10708,N_11781);
and U14013 (N_14013,N_10428,N_10000);
xnor U14014 (N_14014,N_10198,N_10135);
and U14015 (N_14015,N_10103,N_10926);
or U14016 (N_14016,N_10173,N_11480);
nand U14017 (N_14017,N_11361,N_11122);
nand U14018 (N_14018,N_12488,N_10783);
or U14019 (N_14019,N_10468,N_11846);
or U14020 (N_14020,N_11190,N_11840);
and U14021 (N_14021,N_10818,N_12436);
and U14022 (N_14022,N_10650,N_12033);
nand U14023 (N_14023,N_10465,N_11769);
nor U14024 (N_14024,N_11946,N_11342);
nand U14025 (N_14025,N_11634,N_10438);
and U14026 (N_14026,N_11526,N_10402);
nor U14027 (N_14027,N_10738,N_11654);
and U14028 (N_14028,N_10730,N_10450);
xor U14029 (N_14029,N_12148,N_10002);
nand U14030 (N_14030,N_10649,N_11314);
xor U14031 (N_14031,N_10691,N_10586);
and U14032 (N_14032,N_11242,N_10971);
or U14033 (N_14033,N_10452,N_12181);
nand U14034 (N_14034,N_10687,N_12162);
xor U14035 (N_14035,N_10796,N_10907);
or U14036 (N_14036,N_11811,N_12320);
nor U14037 (N_14037,N_12403,N_10844);
and U14038 (N_14038,N_10726,N_11945);
nor U14039 (N_14039,N_12378,N_10800);
and U14040 (N_14040,N_10853,N_12200);
nand U14041 (N_14041,N_10495,N_10516);
or U14042 (N_14042,N_11408,N_11101);
xnor U14043 (N_14043,N_10083,N_10921);
and U14044 (N_14044,N_12451,N_11436);
xor U14045 (N_14045,N_11057,N_12044);
or U14046 (N_14046,N_10839,N_10665);
nand U14047 (N_14047,N_11842,N_11669);
and U14048 (N_14048,N_10203,N_11075);
and U14049 (N_14049,N_11898,N_10174);
nor U14050 (N_14050,N_10047,N_10586);
nor U14051 (N_14051,N_12399,N_11388);
or U14052 (N_14052,N_11065,N_10538);
or U14053 (N_14053,N_11934,N_11241);
or U14054 (N_14054,N_10574,N_10215);
nor U14055 (N_14055,N_10366,N_11821);
nand U14056 (N_14056,N_11965,N_11179);
nand U14057 (N_14057,N_12340,N_10352);
nand U14058 (N_14058,N_10808,N_11503);
xor U14059 (N_14059,N_12331,N_11872);
or U14060 (N_14060,N_10810,N_11423);
or U14061 (N_14061,N_12344,N_10007);
or U14062 (N_14062,N_12421,N_11622);
nand U14063 (N_14063,N_11856,N_12313);
xnor U14064 (N_14064,N_10525,N_10747);
xnor U14065 (N_14065,N_11607,N_12024);
or U14066 (N_14066,N_12250,N_12091);
nor U14067 (N_14067,N_10842,N_10193);
xnor U14068 (N_14068,N_11043,N_11077);
or U14069 (N_14069,N_10803,N_10804);
nand U14070 (N_14070,N_12420,N_12297);
nand U14071 (N_14071,N_11926,N_10350);
and U14072 (N_14072,N_11123,N_11457);
nand U14073 (N_14073,N_10325,N_11651);
and U14074 (N_14074,N_11297,N_11288);
nor U14075 (N_14075,N_10034,N_11445);
xnor U14076 (N_14076,N_10191,N_12139);
nor U14077 (N_14077,N_11066,N_11341);
nand U14078 (N_14078,N_11124,N_12170);
xnor U14079 (N_14079,N_10679,N_11056);
nor U14080 (N_14080,N_10538,N_10307);
nor U14081 (N_14081,N_12462,N_10952);
nand U14082 (N_14082,N_11740,N_11000);
or U14083 (N_14083,N_12487,N_11630);
nand U14084 (N_14084,N_10132,N_11704);
xnor U14085 (N_14085,N_12473,N_11498);
xor U14086 (N_14086,N_11406,N_12151);
or U14087 (N_14087,N_11121,N_10730);
nand U14088 (N_14088,N_12322,N_11723);
or U14089 (N_14089,N_12320,N_12111);
nor U14090 (N_14090,N_11816,N_12355);
nor U14091 (N_14091,N_12306,N_11680);
or U14092 (N_14092,N_11270,N_10330);
or U14093 (N_14093,N_11324,N_11548);
or U14094 (N_14094,N_12474,N_10039);
or U14095 (N_14095,N_11337,N_10965);
or U14096 (N_14096,N_10498,N_10038);
xor U14097 (N_14097,N_10517,N_12167);
nand U14098 (N_14098,N_10740,N_12201);
or U14099 (N_14099,N_11079,N_10760);
or U14100 (N_14100,N_12236,N_10270);
nor U14101 (N_14101,N_10753,N_11127);
nand U14102 (N_14102,N_10961,N_11231);
nand U14103 (N_14103,N_12146,N_10927);
and U14104 (N_14104,N_10416,N_10602);
nor U14105 (N_14105,N_10957,N_10392);
or U14106 (N_14106,N_12350,N_12190);
or U14107 (N_14107,N_11058,N_10256);
or U14108 (N_14108,N_12179,N_10095);
nand U14109 (N_14109,N_11434,N_11183);
or U14110 (N_14110,N_10884,N_10857);
and U14111 (N_14111,N_11696,N_11773);
nor U14112 (N_14112,N_10249,N_11686);
nor U14113 (N_14113,N_11190,N_11864);
nand U14114 (N_14114,N_10609,N_11632);
or U14115 (N_14115,N_11661,N_10414);
and U14116 (N_14116,N_10386,N_11498);
xnor U14117 (N_14117,N_12170,N_11678);
xnor U14118 (N_14118,N_12397,N_11219);
and U14119 (N_14119,N_12393,N_11314);
and U14120 (N_14120,N_10905,N_11879);
xnor U14121 (N_14121,N_10090,N_11926);
and U14122 (N_14122,N_11872,N_10906);
or U14123 (N_14123,N_10044,N_12283);
xor U14124 (N_14124,N_11885,N_11827);
xor U14125 (N_14125,N_11383,N_11613);
nor U14126 (N_14126,N_10147,N_12408);
nand U14127 (N_14127,N_11622,N_12371);
xnor U14128 (N_14128,N_12071,N_11118);
xnor U14129 (N_14129,N_11505,N_12239);
nor U14130 (N_14130,N_11896,N_10921);
and U14131 (N_14131,N_11614,N_12075);
xor U14132 (N_14132,N_11021,N_10001);
and U14133 (N_14133,N_12297,N_10293);
and U14134 (N_14134,N_10244,N_10262);
nand U14135 (N_14135,N_10986,N_12472);
nand U14136 (N_14136,N_12420,N_10278);
and U14137 (N_14137,N_10034,N_10206);
xor U14138 (N_14138,N_10864,N_10708);
nor U14139 (N_14139,N_10025,N_10655);
or U14140 (N_14140,N_12372,N_11816);
and U14141 (N_14141,N_10915,N_11254);
nor U14142 (N_14142,N_10785,N_10897);
or U14143 (N_14143,N_12100,N_10545);
nand U14144 (N_14144,N_10594,N_11949);
or U14145 (N_14145,N_11756,N_11256);
nand U14146 (N_14146,N_11308,N_11864);
nand U14147 (N_14147,N_11302,N_11866);
nand U14148 (N_14148,N_12253,N_10073);
nor U14149 (N_14149,N_12474,N_10686);
or U14150 (N_14150,N_12160,N_10912);
nand U14151 (N_14151,N_11263,N_11393);
nand U14152 (N_14152,N_11482,N_12462);
nor U14153 (N_14153,N_11034,N_10961);
and U14154 (N_14154,N_11708,N_11302);
nand U14155 (N_14155,N_11703,N_10863);
nor U14156 (N_14156,N_11144,N_10669);
nand U14157 (N_14157,N_10429,N_11919);
nand U14158 (N_14158,N_12352,N_11383);
xnor U14159 (N_14159,N_10773,N_11733);
nand U14160 (N_14160,N_11588,N_10349);
xnor U14161 (N_14161,N_10279,N_12443);
nor U14162 (N_14162,N_11272,N_12293);
xnor U14163 (N_14163,N_11659,N_11903);
nand U14164 (N_14164,N_12271,N_10644);
and U14165 (N_14165,N_10333,N_10393);
nor U14166 (N_14166,N_10874,N_11436);
xor U14167 (N_14167,N_12142,N_10032);
xor U14168 (N_14168,N_12300,N_11898);
nand U14169 (N_14169,N_11428,N_11467);
xnor U14170 (N_14170,N_12255,N_11751);
nand U14171 (N_14171,N_10174,N_10842);
or U14172 (N_14172,N_10193,N_11079);
and U14173 (N_14173,N_10773,N_12187);
or U14174 (N_14174,N_10302,N_10510);
xnor U14175 (N_14175,N_12178,N_11679);
or U14176 (N_14176,N_10961,N_10911);
or U14177 (N_14177,N_11342,N_12019);
nor U14178 (N_14178,N_10712,N_12495);
nor U14179 (N_14179,N_12361,N_11013);
xor U14180 (N_14180,N_12412,N_11534);
and U14181 (N_14181,N_10865,N_11618);
xnor U14182 (N_14182,N_10686,N_10596);
nor U14183 (N_14183,N_12396,N_12486);
nand U14184 (N_14184,N_10377,N_10667);
xnor U14185 (N_14185,N_10692,N_10475);
and U14186 (N_14186,N_12264,N_10174);
nor U14187 (N_14187,N_11202,N_11464);
and U14188 (N_14188,N_11369,N_10887);
nand U14189 (N_14189,N_11720,N_10314);
nor U14190 (N_14190,N_11741,N_12292);
nand U14191 (N_14191,N_10462,N_11583);
nand U14192 (N_14192,N_11349,N_11768);
and U14193 (N_14193,N_10414,N_11179);
and U14194 (N_14194,N_10204,N_10306);
and U14195 (N_14195,N_11819,N_11247);
and U14196 (N_14196,N_10429,N_11714);
nor U14197 (N_14197,N_10761,N_10007);
nand U14198 (N_14198,N_10100,N_12029);
xnor U14199 (N_14199,N_11417,N_11753);
nor U14200 (N_14200,N_11268,N_10733);
or U14201 (N_14201,N_10974,N_12007);
nor U14202 (N_14202,N_12330,N_12016);
and U14203 (N_14203,N_10528,N_10156);
nand U14204 (N_14204,N_11014,N_11126);
xor U14205 (N_14205,N_10571,N_10062);
xnor U14206 (N_14206,N_11248,N_10151);
xor U14207 (N_14207,N_11581,N_11774);
nand U14208 (N_14208,N_11068,N_10931);
and U14209 (N_14209,N_12444,N_11036);
nand U14210 (N_14210,N_11729,N_12192);
nor U14211 (N_14211,N_10900,N_11707);
and U14212 (N_14212,N_10789,N_11602);
nand U14213 (N_14213,N_10695,N_10184);
or U14214 (N_14214,N_11417,N_11253);
nor U14215 (N_14215,N_10688,N_10863);
nor U14216 (N_14216,N_11183,N_11036);
xnor U14217 (N_14217,N_11792,N_12019);
or U14218 (N_14218,N_10892,N_11337);
and U14219 (N_14219,N_10297,N_10630);
or U14220 (N_14220,N_10206,N_10155);
or U14221 (N_14221,N_11111,N_10658);
xor U14222 (N_14222,N_11275,N_12391);
or U14223 (N_14223,N_11898,N_11946);
nor U14224 (N_14224,N_12299,N_11282);
xor U14225 (N_14225,N_11137,N_12184);
nor U14226 (N_14226,N_12049,N_10348);
nor U14227 (N_14227,N_10705,N_10224);
and U14228 (N_14228,N_10575,N_10423);
nand U14229 (N_14229,N_11702,N_10447);
xnor U14230 (N_14230,N_11261,N_10809);
and U14231 (N_14231,N_12073,N_12156);
xnor U14232 (N_14232,N_10129,N_11745);
nand U14233 (N_14233,N_10562,N_11987);
nor U14234 (N_14234,N_11116,N_11827);
xor U14235 (N_14235,N_12054,N_11633);
nor U14236 (N_14236,N_11696,N_12497);
xnor U14237 (N_14237,N_10696,N_10796);
and U14238 (N_14238,N_12109,N_10174);
xnor U14239 (N_14239,N_12490,N_12365);
or U14240 (N_14240,N_11392,N_11410);
and U14241 (N_14241,N_12030,N_11482);
xor U14242 (N_14242,N_12130,N_10352);
and U14243 (N_14243,N_12325,N_11056);
nand U14244 (N_14244,N_11000,N_12415);
nor U14245 (N_14245,N_11062,N_12269);
or U14246 (N_14246,N_10310,N_12056);
xnor U14247 (N_14247,N_11359,N_11387);
xor U14248 (N_14248,N_10030,N_10885);
nand U14249 (N_14249,N_11252,N_10531);
nand U14250 (N_14250,N_11504,N_12362);
xor U14251 (N_14251,N_10061,N_10992);
or U14252 (N_14252,N_10559,N_11827);
nand U14253 (N_14253,N_11258,N_10027);
and U14254 (N_14254,N_11182,N_10220);
and U14255 (N_14255,N_10676,N_11219);
xnor U14256 (N_14256,N_11494,N_11073);
nor U14257 (N_14257,N_10151,N_11756);
nand U14258 (N_14258,N_10374,N_11208);
xnor U14259 (N_14259,N_10695,N_10613);
or U14260 (N_14260,N_10757,N_11529);
and U14261 (N_14261,N_10970,N_10536);
xnor U14262 (N_14262,N_12306,N_10340);
and U14263 (N_14263,N_11223,N_10784);
or U14264 (N_14264,N_11477,N_11800);
or U14265 (N_14265,N_10848,N_11632);
and U14266 (N_14266,N_12150,N_11311);
nand U14267 (N_14267,N_10038,N_11157);
or U14268 (N_14268,N_11433,N_10650);
nor U14269 (N_14269,N_11733,N_11392);
nor U14270 (N_14270,N_10023,N_11964);
xnor U14271 (N_14271,N_10122,N_10773);
nor U14272 (N_14272,N_12332,N_10569);
and U14273 (N_14273,N_11210,N_10333);
nand U14274 (N_14274,N_10984,N_11079);
and U14275 (N_14275,N_10764,N_10664);
or U14276 (N_14276,N_12116,N_11861);
and U14277 (N_14277,N_10445,N_10071);
xor U14278 (N_14278,N_11548,N_10826);
xnor U14279 (N_14279,N_10347,N_11230);
nand U14280 (N_14280,N_12059,N_12298);
nor U14281 (N_14281,N_12143,N_10189);
or U14282 (N_14282,N_10225,N_10652);
and U14283 (N_14283,N_11132,N_11009);
nor U14284 (N_14284,N_12066,N_10984);
xnor U14285 (N_14285,N_11719,N_12372);
xnor U14286 (N_14286,N_11196,N_10097);
xor U14287 (N_14287,N_11460,N_10392);
or U14288 (N_14288,N_10363,N_11984);
nand U14289 (N_14289,N_10581,N_11199);
nand U14290 (N_14290,N_11008,N_10481);
and U14291 (N_14291,N_11735,N_10927);
and U14292 (N_14292,N_10553,N_11858);
or U14293 (N_14293,N_10214,N_10990);
and U14294 (N_14294,N_10723,N_12449);
xor U14295 (N_14295,N_10059,N_10953);
or U14296 (N_14296,N_12307,N_10124);
xor U14297 (N_14297,N_11099,N_12085);
xor U14298 (N_14298,N_10267,N_12048);
xnor U14299 (N_14299,N_10177,N_10820);
xor U14300 (N_14300,N_12154,N_11050);
or U14301 (N_14301,N_10260,N_12480);
nor U14302 (N_14302,N_10535,N_11726);
or U14303 (N_14303,N_11479,N_12289);
nand U14304 (N_14304,N_12412,N_10837);
xnor U14305 (N_14305,N_10924,N_11791);
xor U14306 (N_14306,N_10143,N_12422);
xor U14307 (N_14307,N_10697,N_11110);
nand U14308 (N_14308,N_11764,N_11904);
or U14309 (N_14309,N_12340,N_10021);
nor U14310 (N_14310,N_12184,N_10875);
nor U14311 (N_14311,N_11794,N_10570);
and U14312 (N_14312,N_11982,N_10293);
nand U14313 (N_14313,N_10768,N_10337);
xor U14314 (N_14314,N_10374,N_12339);
nand U14315 (N_14315,N_12407,N_11861);
nor U14316 (N_14316,N_10908,N_11806);
or U14317 (N_14317,N_12402,N_11655);
xnor U14318 (N_14318,N_11095,N_11337);
nor U14319 (N_14319,N_11084,N_11978);
or U14320 (N_14320,N_11994,N_10367);
and U14321 (N_14321,N_12409,N_11950);
nand U14322 (N_14322,N_11768,N_10114);
and U14323 (N_14323,N_11715,N_12313);
nor U14324 (N_14324,N_11343,N_11666);
and U14325 (N_14325,N_11620,N_10879);
xnor U14326 (N_14326,N_10283,N_11256);
nor U14327 (N_14327,N_11994,N_11422);
nand U14328 (N_14328,N_10489,N_11552);
xnor U14329 (N_14329,N_11366,N_10572);
or U14330 (N_14330,N_11998,N_12254);
or U14331 (N_14331,N_12357,N_10742);
xnor U14332 (N_14332,N_11587,N_10288);
nor U14333 (N_14333,N_11215,N_11458);
or U14334 (N_14334,N_11183,N_12423);
nand U14335 (N_14335,N_12414,N_10835);
and U14336 (N_14336,N_12190,N_11551);
and U14337 (N_14337,N_10205,N_11727);
or U14338 (N_14338,N_11716,N_10253);
nand U14339 (N_14339,N_12189,N_10312);
or U14340 (N_14340,N_10406,N_11333);
or U14341 (N_14341,N_10475,N_10917);
xor U14342 (N_14342,N_11302,N_11907);
xor U14343 (N_14343,N_10760,N_10068);
and U14344 (N_14344,N_11435,N_11400);
or U14345 (N_14345,N_10127,N_10391);
xor U14346 (N_14346,N_10702,N_12236);
xor U14347 (N_14347,N_10710,N_10133);
or U14348 (N_14348,N_11599,N_11610);
nor U14349 (N_14349,N_10230,N_11502);
and U14350 (N_14350,N_10125,N_12128);
and U14351 (N_14351,N_11182,N_11035);
nor U14352 (N_14352,N_12490,N_11472);
nor U14353 (N_14353,N_12432,N_11736);
and U14354 (N_14354,N_10799,N_10691);
nor U14355 (N_14355,N_11608,N_12170);
nor U14356 (N_14356,N_12463,N_10098);
xnor U14357 (N_14357,N_10237,N_11858);
nor U14358 (N_14358,N_12442,N_12105);
nand U14359 (N_14359,N_12254,N_11693);
and U14360 (N_14360,N_12352,N_10329);
and U14361 (N_14361,N_11979,N_10092);
xnor U14362 (N_14362,N_12224,N_10881);
xnor U14363 (N_14363,N_12315,N_11117);
and U14364 (N_14364,N_10532,N_10016);
nand U14365 (N_14365,N_10296,N_11054);
and U14366 (N_14366,N_10481,N_11236);
nor U14367 (N_14367,N_10445,N_10531);
nor U14368 (N_14368,N_10879,N_12186);
nor U14369 (N_14369,N_11760,N_12180);
and U14370 (N_14370,N_12320,N_12323);
or U14371 (N_14371,N_11791,N_11696);
or U14372 (N_14372,N_11686,N_10561);
and U14373 (N_14373,N_11638,N_10368);
nor U14374 (N_14374,N_12466,N_12196);
xor U14375 (N_14375,N_11472,N_11223);
and U14376 (N_14376,N_10402,N_12267);
nor U14377 (N_14377,N_12379,N_12069);
nand U14378 (N_14378,N_11485,N_10733);
or U14379 (N_14379,N_12440,N_12097);
xor U14380 (N_14380,N_10892,N_11503);
nor U14381 (N_14381,N_10321,N_10089);
and U14382 (N_14382,N_11705,N_12110);
nor U14383 (N_14383,N_10004,N_11948);
xnor U14384 (N_14384,N_12215,N_10957);
and U14385 (N_14385,N_11208,N_10489);
or U14386 (N_14386,N_11925,N_11567);
xor U14387 (N_14387,N_11721,N_10875);
nor U14388 (N_14388,N_12464,N_11124);
or U14389 (N_14389,N_12201,N_11848);
or U14390 (N_14390,N_11468,N_10247);
xnor U14391 (N_14391,N_11281,N_11906);
nand U14392 (N_14392,N_10533,N_11337);
and U14393 (N_14393,N_11269,N_10690);
and U14394 (N_14394,N_11858,N_12319);
and U14395 (N_14395,N_11315,N_11303);
or U14396 (N_14396,N_11363,N_11792);
nand U14397 (N_14397,N_11367,N_11346);
and U14398 (N_14398,N_10889,N_10454);
or U14399 (N_14399,N_11388,N_11166);
nor U14400 (N_14400,N_11407,N_11667);
nand U14401 (N_14401,N_12097,N_10062);
xor U14402 (N_14402,N_10725,N_12027);
and U14403 (N_14403,N_11174,N_12093);
nand U14404 (N_14404,N_12280,N_10101);
xor U14405 (N_14405,N_11631,N_10721);
nand U14406 (N_14406,N_10859,N_12131);
xor U14407 (N_14407,N_10655,N_11702);
or U14408 (N_14408,N_11179,N_10118);
or U14409 (N_14409,N_10323,N_11515);
nor U14410 (N_14410,N_11490,N_11205);
or U14411 (N_14411,N_10595,N_11251);
nand U14412 (N_14412,N_11401,N_11365);
xor U14413 (N_14413,N_11910,N_10592);
and U14414 (N_14414,N_12125,N_11715);
nor U14415 (N_14415,N_11156,N_10601);
nor U14416 (N_14416,N_11841,N_10518);
and U14417 (N_14417,N_10285,N_12131);
nor U14418 (N_14418,N_10219,N_11203);
nand U14419 (N_14419,N_10784,N_11547);
or U14420 (N_14420,N_11334,N_12387);
and U14421 (N_14421,N_10597,N_10280);
nor U14422 (N_14422,N_12465,N_10958);
xnor U14423 (N_14423,N_10718,N_11220);
xnor U14424 (N_14424,N_10189,N_12306);
nor U14425 (N_14425,N_11987,N_11214);
or U14426 (N_14426,N_12466,N_10196);
nand U14427 (N_14427,N_11525,N_11762);
xor U14428 (N_14428,N_12169,N_12183);
xnor U14429 (N_14429,N_10523,N_11934);
xor U14430 (N_14430,N_10162,N_11883);
and U14431 (N_14431,N_12176,N_10148);
xor U14432 (N_14432,N_11308,N_10126);
xnor U14433 (N_14433,N_11613,N_12323);
xnor U14434 (N_14434,N_10582,N_11510);
nor U14435 (N_14435,N_12407,N_10269);
nor U14436 (N_14436,N_10663,N_10961);
xor U14437 (N_14437,N_11754,N_12417);
xor U14438 (N_14438,N_11610,N_12078);
nand U14439 (N_14439,N_11336,N_12388);
nor U14440 (N_14440,N_11814,N_11684);
nor U14441 (N_14441,N_11747,N_10110);
xor U14442 (N_14442,N_11437,N_10012);
or U14443 (N_14443,N_12327,N_12117);
nand U14444 (N_14444,N_11650,N_11901);
xnor U14445 (N_14445,N_12073,N_11972);
nor U14446 (N_14446,N_10160,N_10894);
xnor U14447 (N_14447,N_11532,N_10951);
nand U14448 (N_14448,N_11380,N_11779);
xnor U14449 (N_14449,N_10098,N_11853);
and U14450 (N_14450,N_10184,N_12391);
or U14451 (N_14451,N_10880,N_10179);
and U14452 (N_14452,N_11993,N_10736);
nand U14453 (N_14453,N_10179,N_12333);
nand U14454 (N_14454,N_11151,N_10345);
xnor U14455 (N_14455,N_10395,N_11410);
and U14456 (N_14456,N_11457,N_12081);
and U14457 (N_14457,N_10141,N_10246);
nor U14458 (N_14458,N_11151,N_10788);
nor U14459 (N_14459,N_10007,N_11736);
or U14460 (N_14460,N_10544,N_11343);
xor U14461 (N_14461,N_10303,N_10450);
xor U14462 (N_14462,N_10526,N_10804);
or U14463 (N_14463,N_11630,N_11971);
and U14464 (N_14464,N_10182,N_12029);
xnor U14465 (N_14465,N_12468,N_11978);
xor U14466 (N_14466,N_11717,N_10423);
or U14467 (N_14467,N_10006,N_10051);
xor U14468 (N_14468,N_11063,N_10717);
nor U14469 (N_14469,N_11397,N_10824);
xnor U14470 (N_14470,N_10693,N_12077);
xnor U14471 (N_14471,N_11405,N_11072);
nand U14472 (N_14472,N_10644,N_10044);
xnor U14473 (N_14473,N_12173,N_12092);
nor U14474 (N_14474,N_10118,N_12453);
nand U14475 (N_14475,N_11203,N_10916);
or U14476 (N_14476,N_12288,N_12009);
or U14477 (N_14477,N_11276,N_11148);
xnor U14478 (N_14478,N_12392,N_12189);
or U14479 (N_14479,N_10115,N_12203);
or U14480 (N_14480,N_11847,N_10702);
or U14481 (N_14481,N_11365,N_11292);
and U14482 (N_14482,N_10616,N_10725);
nand U14483 (N_14483,N_11298,N_11578);
or U14484 (N_14484,N_10424,N_11646);
xor U14485 (N_14485,N_10979,N_11863);
nor U14486 (N_14486,N_10597,N_10494);
nor U14487 (N_14487,N_12144,N_11645);
nand U14488 (N_14488,N_10087,N_10221);
nand U14489 (N_14489,N_11899,N_12055);
xor U14490 (N_14490,N_10283,N_11621);
and U14491 (N_14491,N_12008,N_11912);
nor U14492 (N_14492,N_10586,N_11345);
and U14493 (N_14493,N_11177,N_12324);
and U14494 (N_14494,N_10685,N_11402);
nor U14495 (N_14495,N_10191,N_11197);
xor U14496 (N_14496,N_10367,N_11570);
xor U14497 (N_14497,N_10845,N_12336);
nand U14498 (N_14498,N_11583,N_11961);
nand U14499 (N_14499,N_12291,N_10982);
or U14500 (N_14500,N_11178,N_11213);
xor U14501 (N_14501,N_11454,N_11600);
and U14502 (N_14502,N_10944,N_11190);
xnor U14503 (N_14503,N_10185,N_12410);
nor U14504 (N_14504,N_12450,N_11436);
xnor U14505 (N_14505,N_10149,N_10561);
nand U14506 (N_14506,N_12461,N_10384);
nor U14507 (N_14507,N_12006,N_11816);
nand U14508 (N_14508,N_11773,N_10411);
and U14509 (N_14509,N_10927,N_11623);
nor U14510 (N_14510,N_10823,N_12270);
xor U14511 (N_14511,N_11600,N_11280);
or U14512 (N_14512,N_10155,N_10736);
xnor U14513 (N_14513,N_12483,N_12476);
nor U14514 (N_14514,N_10732,N_11842);
xor U14515 (N_14515,N_10439,N_12459);
or U14516 (N_14516,N_10619,N_10314);
nor U14517 (N_14517,N_11030,N_11586);
nand U14518 (N_14518,N_11660,N_11589);
and U14519 (N_14519,N_11360,N_10372);
nor U14520 (N_14520,N_12274,N_10266);
nand U14521 (N_14521,N_10767,N_11773);
nor U14522 (N_14522,N_11397,N_12200);
and U14523 (N_14523,N_10817,N_10136);
xnor U14524 (N_14524,N_11756,N_11910);
or U14525 (N_14525,N_12103,N_11824);
nor U14526 (N_14526,N_11602,N_11442);
or U14527 (N_14527,N_11954,N_11144);
and U14528 (N_14528,N_10016,N_10761);
nor U14529 (N_14529,N_10879,N_11034);
nor U14530 (N_14530,N_11039,N_11941);
nor U14531 (N_14531,N_10174,N_11756);
or U14532 (N_14532,N_10824,N_12133);
nand U14533 (N_14533,N_10563,N_10195);
xor U14534 (N_14534,N_10268,N_10959);
nand U14535 (N_14535,N_11279,N_11139);
nand U14536 (N_14536,N_11841,N_11800);
xnor U14537 (N_14537,N_10692,N_11707);
or U14538 (N_14538,N_12220,N_11226);
nand U14539 (N_14539,N_10642,N_11659);
and U14540 (N_14540,N_10679,N_11439);
and U14541 (N_14541,N_10875,N_11377);
or U14542 (N_14542,N_11231,N_10317);
xnor U14543 (N_14543,N_10225,N_10399);
and U14544 (N_14544,N_11142,N_12288);
or U14545 (N_14545,N_10076,N_10004);
or U14546 (N_14546,N_10355,N_12152);
and U14547 (N_14547,N_10714,N_11596);
nand U14548 (N_14548,N_11331,N_10363);
and U14549 (N_14549,N_12453,N_11747);
and U14550 (N_14550,N_10272,N_10491);
nor U14551 (N_14551,N_10569,N_10566);
xnor U14552 (N_14552,N_10320,N_10086);
nand U14553 (N_14553,N_11892,N_11899);
or U14554 (N_14554,N_10109,N_12018);
nor U14555 (N_14555,N_10982,N_10307);
or U14556 (N_14556,N_11319,N_10613);
nor U14557 (N_14557,N_10038,N_10707);
xor U14558 (N_14558,N_11974,N_10291);
and U14559 (N_14559,N_10604,N_11763);
and U14560 (N_14560,N_12084,N_10509);
and U14561 (N_14561,N_12409,N_10422);
or U14562 (N_14562,N_10981,N_10396);
and U14563 (N_14563,N_12070,N_11982);
and U14564 (N_14564,N_11705,N_12353);
xor U14565 (N_14565,N_10173,N_12149);
and U14566 (N_14566,N_11339,N_12147);
xnor U14567 (N_14567,N_11141,N_12375);
nand U14568 (N_14568,N_12063,N_11922);
xor U14569 (N_14569,N_10811,N_12153);
nor U14570 (N_14570,N_10289,N_12333);
xnor U14571 (N_14571,N_10931,N_10662);
nor U14572 (N_14572,N_11877,N_11749);
and U14573 (N_14573,N_11507,N_11910);
nand U14574 (N_14574,N_12444,N_12334);
or U14575 (N_14575,N_11869,N_10607);
nand U14576 (N_14576,N_12312,N_11708);
or U14577 (N_14577,N_10193,N_12059);
nand U14578 (N_14578,N_11546,N_10685);
xor U14579 (N_14579,N_10006,N_10548);
or U14580 (N_14580,N_10666,N_10023);
nor U14581 (N_14581,N_10346,N_10187);
or U14582 (N_14582,N_11319,N_11674);
xor U14583 (N_14583,N_11296,N_11827);
nand U14584 (N_14584,N_11361,N_11845);
or U14585 (N_14585,N_10722,N_11808);
and U14586 (N_14586,N_10153,N_12057);
nand U14587 (N_14587,N_11324,N_12360);
xnor U14588 (N_14588,N_11955,N_10125);
xor U14589 (N_14589,N_11178,N_10748);
or U14590 (N_14590,N_12254,N_11007);
or U14591 (N_14591,N_11490,N_11458);
and U14592 (N_14592,N_11906,N_12212);
xnor U14593 (N_14593,N_12416,N_10913);
nand U14594 (N_14594,N_11328,N_12205);
or U14595 (N_14595,N_10000,N_10114);
nand U14596 (N_14596,N_11791,N_10713);
nor U14597 (N_14597,N_10318,N_10529);
or U14598 (N_14598,N_10165,N_12072);
nand U14599 (N_14599,N_10123,N_10712);
and U14600 (N_14600,N_10226,N_12158);
xnor U14601 (N_14601,N_10735,N_11760);
or U14602 (N_14602,N_10086,N_11808);
or U14603 (N_14603,N_11655,N_10125);
or U14604 (N_14604,N_10616,N_10527);
nand U14605 (N_14605,N_10488,N_11253);
and U14606 (N_14606,N_12209,N_10810);
nor U14607 (N_14607,N_12063,N_10405);
or U14608 (N_14608,N_12484,N_10385);
nor U14609 (N_14609,N_11759,N_10272);
or U14610 (N_14610,N_12424,N_11537);
nand U14611 (N_14611,N_10021,N_10504);
or U14612 (N_14612,N_10537,N_11107);
or U14613 (N_14613,N_10034,N_11951);
nand U14614 (N_14614,N_10525,N_10264);
nor U14615 (N_14615,N_12206,N_11300);
xnor U14616 (N_14616,N_11018,N_10606);
nor U14617 (N_14617,N_12018,N_12246);
nor U14618 (N_14618,N_11649,N_11761);
nand U14619 (N_14619,N_10257,N_10859);
xnor U14620 (N_14620,N_12400,N_12474);
and U14621 (N_14621,N_11499,N_11607);
xor U14622 (N_14622,N_11205,N_12320);
and U14623 (N_14623,N_10005,N_12289);
xnor U14624 (N_14624,N_10568,N_12378);
nor U14625 (N_14625,N_10524,N_11269);
nand U14626 (N_14626,N_12374,N_10846);
nand U14627 (N_14627,N_10395,N_10279);
and U14628 (N_14628,N_11183,N_10401);
xnor U14629 (N_14629,N_10776,N_10640);
nand U14630 (N_14630,N_12300,N_12463);
or U14631 (N_14631,N_12131,N_10110);
xnor U14632 (N_14632,N_12440,N_11926);
xor U14633 (N_14633,N_11832,N_12322);
or U14634 (N_14634,N_11822,N_10892);
or U14635 (N_14635,N_10300,N_11377);
nand U14636 (N_14636,N_10889,N_11349);
nand U14637 (N_14637,N_11980,N_11406);
nand U14638 (N_14638,N_11997,N_12181);
or U14639 (N_14639,N_10686,N_12366);
nand U14640 (N_14640,N_10607,N_10703);
and U14641 (N_14641,N_11984,N_12341);
nor U14642 (N_14642,N_12123,N_10729);
xnor U14643 (N_14643,N_10623,N_11769);
nor U14644 (N_14644,N_10246,N_11226);
nand U14645 (N_14645,N_11894,N_11901);
nand U14646 (N_14646,N_10415,N_12062);
nand U14647 (N_14647,N_12113,N_11306);
nand U14648 (N_14648,N_11415,N_10795);
xor U14649 (N_14649,N_10729,N_10885);
and U14650 (N_14650,N_10285,N_10604);
nor U14651 (N_14651,N_12130,N_10061);
or U14652 (N_14652,N_12299,N_10696);
xor U14653 (N_14653,N_11557,N_11907);
or U14654 (N_14654,N_11077,N_10256);
nand U14655 (N_14655,N_10278,N_12008);
xnor U14656 (N_14656,N_10145,N_10458);
or U14657 (N_14657,N_12223,N_10518);
nor U14658 (N_14658,N_10713,N_12330);
and U14659 (N_14659,N_10476,N_12474);
and U14660 (N_14660,N_10694,N_12305);
nor U14661 (N_14661,N_11445,N_11543);
nor U14662 (N_14662,N_10120,N_10812);
and U14663 (N_14663,N_10965,N_11159);
and U14664 (N_14664,N_12363,N_11875);
xnor U14665 (N_14665,N_10942,N_10169);
or U14666 (N_14666,N_12155,N_10768);
and U14667 (N_14667,N_11766,N_10987);
and U14668 (N_14668,N_12436,N_12168);
and U14669 (N_14669,N_10608,N_11315);
xor U14670 (N_14670,N_10932,N_11215);
or U14671 (N_14671,N_12147,N_10791);
nand U14672 (N_14672,N_10367,N_11731);
xnor U14673 (N_14673,N_11371,N_10691);
nor U14674 (N_14674,N_11627,N_12249);
xor U14675 (N_14675,N_10522,N_12452);
nor U14676 (N_14676,N_10172,N_10128);
xor U14677 (N_14677,N_11656,N_10719);
and U14678 (N_14678,N_10354,N_11276);
nor U14679 (N_14679,N_11604,N_11003);
nor U14680 (N_14680,N_11249,N_11969);
nand U14681 (N_14681,N_11034,N_10897);
xnor U14682 (N_14682,N_11751,N_11924);
and U14683 (N_14683,N_10862,N_10677);
xnor U14684 (N_14684,N_11624,N_12478);
and U14685 (N_14685,N_12057,N_12194);
nor U14686 (N_14686,N_12195,N_11737);
and U14687 (N_14687,N_11304,N_10871);
nand U14688 (N_14688,N_11722,N_10859);
xor U14689 (N_14689,N_11481,N_11287);
nand U14690 (N_14690,N_10644,N_10209);
and U14691 (N_14691,N_11090,N_10763);
xnor U14692 (N_14692,N_10541,N_10827);
nand U14693 (N_14693,N_10758,N_10132);
or U14694 (N_14694,N_10048,N_10424);
nor U14695 (N_14695,N_10448,N_11935);
or U14696 (N_14696,N_10924,N_11365);
nor U14697 (N_14697,N_10755,N_11300);
nand U14698 (N_14698,N_12213,N_12351);
nand U14699 (N_14699,N_12287,N_10985);
nor U14700 (N_14700,N_11293,N_12052);
nand U14701 (N_14701,N_11646,N_10882);
or U14702 (N_14702,N_11129,N_10985);
and U14703 (N_14703,N_11434,N_10424);
nand U14704 (N_14704,N_11748,N_11545);
nor U14705 (N_14705,N_12213,N_10999);
nand U14706 (N_14706,N_12185,N_10083);
and U14707 (N_14707,N_11077,N_11321);
nand U14708 (N_14708,N_10739,N_10247);
xor U14709 (N_14709,N_11297,N_11483);
or U14710 (N_14710,N_10782,N_11409);
and U14711 (N_14711,N_11103,N_10374);
and U14712 (N_14712,N_11053,N_10289);
or U14713 (N_14713,N_11206,N_10777);
nor U14714 (N_14714,N_12449,N_10657);
or U14715 (N_14715,N_10947,N_10488);
xor U14716 (N_14716,N_12135,N_11760);
nand U14717 (N_14717,N_10538,N_10587);
nand U14718 (N_14718,N_10580,N_10188);
nor U14719 (N_14719,N_10074,N_12197);
and U14720 (N_14720,N_12451,N_10615);
nand U14721 (N_14721,N_10569,N_11355);
and U14722 (N_14722,N_11777,N_12063);
and U14723 (N_14723,N_10104,N_11987);
nand U14724 (N_14724,N_11614,N_11398);
and U14725 (N_14725,N_11082,N_11591);
xor U14726 (N_14726,N_10279,N_10127);
nand U14727 (N_14727,N_10432,N_10018);
nand U14728 (N_14728,N_11611,N_10148);
or U14729 (N_14729,N_10587,N_11716);
nor U14730 (N_14730,N_10193,N_11548);
nor U14731 (N_14731,N_10989,N_11909);
xor U14732 (N_14732,N_11228,N_10539);
nand U14733 (N_14733,N_11711,N_10498);
xor U14734 (N_14734,N_11017,N_10420);
or U14735 (N_14735,N_10226,N_11553);
or U14736 (N_14736,N_10889,N_10562);
and U14737 (N_14737,N_11934,N_12021);
or U14738 (N_14738,N_12447,N_11348);
nand U14739 (N_14739,N_11593,N_10621);
xor U14740 (N_14740,N_11108,N_12320);
and U14741 (N_14741,N_11241,N_10126);
xnor U14742 (N_14742,N_11623,N_11781);
xnor U14743 (N_14743,N_12333,N_11413);
nor U14744 (N_14744,N_10348,N_12060);
xnor U14745 (N_14745,N_12170,N_10480);
or U14746 (N_14746,N_11174,N_11875);
and U14747 (N_14747,N_11615,N_10025);
nand U14748 (N_14748,N_11055,N_10495);
or U14749 (N_14749,N_10403,N_10020);
xnor U14750 (N_14750,N_11893,N_10548);
nand U14751 (N_14751,N_12460,N_11166);
nand U14752 (N_14752,N_11187,N_11796);
nor U14753 (N_14753,N_11143,N_10492);
xnor U14754 (N_14754,N_10732,N_10999);
and U14755 (N_14755,N_11403,N_11272);
or U14756 (N_14756,N_11438,N_11967);
and U14757 (N_14757,N_10449,N_12153);
or U14758 (N_14758,N_10312,N_12058);
and U14759 (N_14759,N_12035,N_10245);
nand U14760 (N_14760,N_10271,N_10516);
xor U14761 (N_14761,N_10022,N_12351);
nand U14762 (N_14762,N_10412,N_11825);
and U14763 (N_14763,N_11987,N_12092);
nand U14764 (N_14764,N_11599,N_12261);
nand U14765 (N_14765,N_11008,N_10517);
nor U14766 (N_14766,N_11379,N_12072);
or U14767 (N_14767,N_12445,N_12382);
nor U14768 (N_14768,N_10924,N_11872);
or U14769 (N_14769,N_11301,N_11475);
xor U14770 (N_14770,N_10266,N_10268);
xnor U14771 (N_14771,N_11072,N_11203);
or U14772 (N_14772,N_11881,N_11775);
nand U14773 (N_14773,N_11425,N_10911);
or U14774 (N_14774,N_10183,N_10073);
or U14775 (N_14775,N_10087,N_11324);
or U14776 (N_14776,N_11634,N_10530);
nor U14777 (N_14777,N_10377,N_10934);
or U14778 (N_14778,N_12244,N_10165);
nand U14779 (N_14779,N_12097,N_12327);
or U14780 (N_14780,N_10155,N_12080);
and U14781 (N_14781,N_11096,N_10508);
nand U14782 (N_14782,N_10275,N_10082);
nand U14783 (N_14783,N_11080,N_12428);
xnor U14784 (N_14784,N_12491,N_10773);
nor U14785 (N_14785,N_10226,N_10287);
xnor U14786 (N_14786,N_12320,N_11369);
and U14787 (N_14787,N_12206,N_12254);
and U14788 (N_14788,N_11784,N_11336);
nand U14789 (N_14789,N_11172,N_12444);
xor U14790 (N_14790,N_10914,N_12056);
nand U14791 (N_14791,N_10167,N_12056);
nor U14792 (N_14792,N_10416,N_11282);
or U14793 (N_14793,N_11696,N_10955);
xor U14794 (N_14794,N_11659,N_11363);
or U14795 (N_14795,N_10683,N_11775);
and U14796 (N_14796,N_10461,N_12126);
and U14797 (N_14797,N_11281,N_10727);
xnor U14798 (N_14798,N_11547,N_10530);
xnor U14799 (N_14799,N_11551,N_10020);
or U14800 (N_14800,N_11868,N_11981);
or U14801 (N_14801,N_10502,N_12228);
or U14802 (N_14802,N_12447,N_12288);
nand U14803 (N_14803,N_10159,N_10626);
or U14804 (N_14804,N_10944,N_10144);
or U14805 (N_14805,N_11755,N_11642);
and U14806 (N_14806,N_10485,N_11581);
xor U14807 (N_14807,N_11452,N_10309);
or U14808 (N_14808,N_11948,N_11787);
or U14809 (N_14809,N_11409,N_11972);
or U14810 (N_14810,N_10614,N_12146);
and U14811 (N_14811,N_10674,N_11115);
nor U14812 (N_14812,N_12201,N_11618);
nand U14813 (N_14813,N_10778,N_11724);
and U14814 (N_14814,N_11974,N_12344);
and U14815 (N_14815,N_10505,N_12044);
or U14816 (N_14816,N_11597,N_12178);
and U14817 (N_14817,N_10364,N_11729);
xnor U14818 (N_14818,N_10133,N_11972);
or U14819 (N_14819,N_10861,N_10337);
nand U14820 (N_14820,N_10334,N_10342);
or U14821 (N_14821,N_12167,N_12062);
xnor U14822 (N_14822,N_11475,N_10259);
or U14823 (N_14823,N_10705,N_10512);
nand U14824 (N_14824,N_12008,N_10694);
nand U14825 (N_14825,N_11074,N_11614);
and U14826 (N_14826,N_11526,N_10952);
or U14827 (N_14827,N_10314,N_10523);
nor U14828 (N_14828,N_12462,N_10388);
nor U14829 (N_14829,N_11069,N_11105);
nand U14830 (N_14830,N_11400,N_11084);
xnor U14831 (N_14831,N_12311,N_12136);
nor U14832 (N_14832,N_12057,N_11663);
and U14833 (N_14833,N_10918,N_12211);
or U14834 (N_14834,N_12065,N_11888);
xnor U14835 (N_14835,N_11475,N_10032);
nand U14836 (N_14836,N_11277,N_11610);
or U14837 (N_14837,N_11902,N_11436);
and U14838 (N_14838,N_10844,N_10323);
xnor U14839 (N_14839,N_11222,N_12205);
nand U14840 (N_14840,N_12457,N_10027);
nand U14841 (N_14841,N_12236,N_11437);
nand U14842 (N_14842,N_10563,N_11009);
xor U14843 (N_14843,N_10129,N_11447);
xnor U14844 (N_14844,N_11751,N_12161);
nand U14845 (N_14845,N_11164,N_10066);
or U14846 (N_14846,N_11333,N_10513);
and U14847 (N_14847,N_10286,N_11570);
nor U14848 (N_14848,N_11144,N_11189);
xnor U14849 (N_14849,N_11789,N_11130);
and U14850 (N_14850,N_11826,N_11163);
nor U14851 (N_14851,N_10736,N_12458);
nor U14852 (N_14852,N_11110,N_12424);
xnor U14853 (N_14853,N_11212,N_10003);
and U14854 (N_14854,N_12436,N_11962);
nor U14855 (N_14855,N_11213,N_10854);
nor U14856 (N_14856,N_11765,N_11071);
nor U14857 (N_14857,N_11921,N_11691);
or U14858 (N_14858,N_12206,N_10484);
nor U14859 (N_14859,N_10391,N_12370);
or U14860 (N_14860,N_11185,N_11145);
xnor U14861 (N_14861,N_10396,N_10519);
xor U14862 (N_14862,N_11261,N_10759);
or U14863 (N_14863,N_12047,N_11872);
or U14864 (N_14864,N_12435,N_10760);
and U14865 (N_14865,N_11028,N_10948);
nand U14866 (N_14866,N_12217,N_10072);
nor U14867 (N_14867,N_11324,N_11420);
nand U14868 (N_14868,N_11070,N_10430);
xor U14869 (N_14869,N_12447,N_11005);
nand U14870 (N_14870,N_12376,N_12437);
xnor U14871 (N_14871,N_11557,N_10371);
xnor U14872 (N_14872,N_12401,N_11767);
xor U14873 (N_14873,N_12172,N_10863);
nor U14874 (N_14874,N_10371,N_10156);
or U14875 (N_14875,N_11695,N_11411);
nor U14876 (N_14876,N_10741,N_10610);
xnor U14877 (N_14877,N_10921,N_11536);
and U14878 (N_14878,N_10709,N_10678);
or U14879 (N_14879,N_10287,N_10271);
and U14880 (N_14880,N_10573,N_11451);
and U14881 (N_14881,N_11708,N_12274);
xor U14882 (N_14882,N_12437,N_11434);
xnor U14883 (N_14883,N_11330,N_10015);
xnor U14884 (N_14884,N_11271,N_12447);
nand U14885 (N_14885,N_10974,N_10587);
nor U14886 (N_14886,N_12300,N_10400);
nand U14887 (N_14887,N_10381,N_10587);
or U14888 (N_14888,N_11082,N_12150);
nor U14889 (N_14889,N_11845,N_10931);
xor U14890 (N_14890,N_12466,N_11247);
xor U14891 (N_14891,N_12201,N_11884);
or U14892 (N_14892,N_10066,N_12118);
xor U14893 (N_14893,N_12277,N_11813);
xor U14894 (N_14894,N_10198,N_11998);
nor U14895 (N_14895,N_11809,N_12366);
nor U14896 (N_14896,N_11232,N_11100);
and U14897 (N_14897,N_10554,N_11746);
and U14898 (N_14898,N_12145,N_10550);
nor U14899 (N_14899,N_12450,N_11410);
or U14900 (N_14900,N_10719,N_11294);
or U14901 (N_14901,N_12483,N_12275);
nand U14902 (N_14902,N_11423,N_11241);
nand U14903 (N_14903,N_10516,N_11628);
xor U14904 (N_14904,N_12120,N_12189);
xor U14905 (N_14905,N_11171,N_10015);
or U14906 (N_14906,N_10217,N_10621);
or U14907 (N_14907,N_10748,N_10739);
and U14908 (N_14908,N_11327,N_11689);
xor U14909 (N_14909,N_11884,N_10097);
nand U14910 (N_14910,N_12430,N_10328);
and U14911 (N_14911,N_10044,N_11724);
nand U14912 (N_14912,N_10223,N_11932);
nor U14913 (N_14913,N_11846,N_10853);
and U14914 (N_14914,N_12092,N_12479);
or U14915 (N_14915,N_12075,N_10099);
nand U14916 (N_14916,N_11831,N_12218);
and U14917 (N_14917,N_10479,N_12387);
nor U14918 (N_14918,N_10144,N_12437);
and U14919 (N_14919,N_11637,N_10415);
and U14920 (N_14920,N_10361,N_12046);
xnor U14921 (N_14921,N_10152,N_10760);
nor U14922 (N_14922,N_11010,N_11242);
and U14923 (N_14923,N_11838,N_11208);
or U14924 (N_14924,N_10067,N_11124);
xnor U14925 (N_14925,N_11169,N_11642);
nand U14926 (N_14926,N_11140,N_10998);
xor U14927 (N_14927,N_10156,N_10612);
and U14928 (N_14928,N_10166,N_10341);
nand U14929 (N_14929,N_12406,N_11335);
and U14930 (N_14930,N_11452,N_10491);
or U14931 (N_14931,N_12015,N_11707);
nand U14932 (N_14932,N_12141,N_11688);
or U14933 (N_14933,N_11042,N_11768);
and U14934 (N_14934,N_11283,N_12402);
xor U14935 (N_14935,N_10376,N_11369);
xnor U14936 (N_14936,N_11407,N_11726);
nand U14937 (N_14937,N_12033,N_10258);
xor U14938 (N_14938,N_11300,N_10316);
xnor U14939 (N_14939,N_10077,N_11194);
and U14940 (N_14940,N_11179,N_10305);
and U14941 (N_14941,N_10594,N_11195);
and U14942 (N_14942,N_10488,N_11612);
and U14943 (N_14943,N_11187,N_11001);
xor U14944 (N_14944,N_10872,N_12158);
nand U14945 (N_14945,N_10930,N_12456);
nand U14946 (N_14946,N_10947,N_10994);
xor U14947 (N_14947,N_11201,N_11479);
xnor U14948 (N_14948,N_10256,N_10186);
nand U14949 (N_14949,N_11728,N_11687);
xnor U14950 (N_14950,N_11200,N_11305);
xnor U14951 (N_14951,N_12261,N_10823);
or U14952 (N_14952,N_11274,N_11089);
and U14953 (N_14953,N_11609,N_11672);
nand U14954 (N_14954,N_10404,N_10550);
xor U14955 (N_14955,N_10184,N_10262);
or U14956 (N_14956,N_10664,N_12251);
xnor U14957 (N_14957,N_10349,N_11798);
nor U14958 (N_14958,N_10539,N_12277);
and U14959 (N_14959,N_11522,N_10532);
nand U14960 (N_14960,N_12020,N_10800);
and U14961 (N_14961,N_12235,N_10794);
nor U14962 (N_14962,N_11918,N_11330);
and U14963 (N_14963,N_10690,N_10343);
and U14964 (N_14964,N_10208,N_11751);
and U14965 (N_14965,N_10259,N_11145);
and U14966 (N_14966,N_10483,N_10340);
and U14967 (N_14967,N_11140,N_10291);
and U14968 (N_14968,N_10850,N_10729);
nor U14969 (N_14969,N_10093,N_12207);
nor U14970 (N_14970,N_11411,N_11713);
or U14971 (N_14971,N_11417,N_10691);
nor U14972 (N_14972,N_11506,N_10755);
and U14973 (N_14973,N_11027,N_10804);
xor U14974 (N_14974,N_10109,N_11282);
and U14975 (N_14975,N_11122,N_12164);
nand U14976 (N_14976,N_10919,N_10550);
xor U14977 (N_14977,N_12341,N_11569);
xor U14978 (N_14978,N_11641,N_11272);
xor U14979 (N_14979,N_11990,N_10876);
xor U14980 (N_14980,N_12139,N_10136);
or U14981 (N_14981,N_11916,N_10472);
or U14982 (N_14982,N_11996,N_11600);
or U14983 (N_14983,N_11862,N_11338);
xor U14984 (N_14984,N_10812,N_11979);
xor U14985 (N_14985,N_10285,N_12027);
nor U14986 (N_14986,N_12431,N_10103);
and U14987 (N_14987,N_12160,N_12034);
xnor U14988 (N_14988,N_11465,N_10856);
nor U14989 (N_14989,N_10913,N_11503);
and U14990 (N_14990,N_10992,N_12371);
and U14991 (N_14991,N_11379,N_11267);
or U14992 (N_14992,N_12043,N_12486);
nor U14993 (N_14993,N_10688,N_11670);
and U14994 (N_14994,N_10327,N_10087);
and U14995 (N_14995,N_10626,N_11018);
nand U14996 (N_14996,N_12419,N_10446);
and U14997 (N_14997,N_10997,N_10128);
xor U14998 (N_14998,N_11086,N_12454);
nand U14999 (N_14999,N_12415,N_12098);
nor U15000 (N_15000,N_13227,N_14765);
nor U15001 (N_15001,N_13915,N_12548);
nand U15002 (N_15002,N_14806,N_14907);
nor U15003 (N_15003,N_14874,N_13493);
nand U15004 (N_15004,N_12722,N_13640);
nor U15005 (N_15005,N_13471,N_13279);
nor U15006 (N_15006,N_14039,N_14361);
or U15007 (N_15007,N_14957,N_12628);
nand U15008 (N_15008,N_14367,N_13341);
and U15009 (N_15009,N_14536,N_13872);
xor U15010 (N_15010,N_13753,N_14509);
xor U15011 (N_15011,N_13989,N_13707);
and U15012 (N_15012,N_13808,N_14935);
nor U15013 (N_15013,N_12750,N_14748);
or U15014 (N_15014,N_14326,N_14510);
nand U15015 (N_15015,N_14081,N_14459);
nor U15016 (N_15016,N_12696,N_13647);
nand U15017 (N_15017,N_14940,N_14445);
xor U15018 (N_15018,N_13099,N_13906);
or U15019 (N_15019,N_14391,N_12665);
nor U15020 (N_15020,N_12820,N_13170);
or U15021 (N_15021,N_14207,N_14966);
and U15022 (N_15022,N_12523,N_13096);
nand U15023 (N_15023,N_13444,N_12909);
nand U15024 (N_15024,N_12976,N_12887);
nor U15025 (N_15025,N_14743,N_14041);
nor U15026 (N_15026,N_14673,N_14153);
or U15027 (N_15027,N_12922,N_12651);
xor U15028 (N_15028,N_14527,N_14357);
or U15029 (N_15029,N_14864,N_13933);
or U15030 (N_15030,N_14863,N_13089);
and U15031 (N_15031,N_13787,N_14561);
or U15032 (N_15032,N_13593,N_13675);
or U15033 (N_15033,N_14151,N_12791);
or U15034 (N_15034,N_14782,N_14483);
nor U15035 (N_15035,N_14046,N_13583);
or U15036 (N_15036,N_14195,N_13169);
and U15037 (N_15037,N_12658,N_12657);
or U15038 (N_15038,N_12588,N_13931);
xor U15039 (N_15039,N_14197,N_12731);
and U15040 (N_15040,N_14511,N_13442);
and U15041 (N_15041,N_14001,N_13581);
or U15042 (N_15042,N_14463,N_14789);
nand U15043 (N_15043,N_14978,N_13422);
nor U15044 (N_15044,N_12507,N_13244);
or U15045 (N_15045,N_14160,N_14420);
nor U15046 (N_15046,N_14904,N_14764);
nand U15047 (N_15047,N_13241,N_13695);
and U15048 (N_15048,N_14914,N_12752);
and U15049 (N_15049,N_14921,N_12927);
xnor U15050 (N_15050,N_12527,N_12577);
and U15051 (N_15051,N_12712,N_14530);
xnor U15052 (N_15052,N_14264,N_14328);
or U15053 (N_15053,N_14019,N_13761);
and U15054 (N_15054,N_13226,N_14828);
xor U15055 (N_15055,N_13252,N_12753);
nand U15056 (N_15056,N_13667,N_12785);
nand U15057 (N_15057,N_14034,N_13970);
or U15058 (N_15058,N_13396,N_14289);
nor U15059 (N_15059,N_13268,N_13440);
nor U15060 (N_15060,N_13569,N_14987);
nor U15061 (N_15061,N_14517,N_14755);
xnor U15062 (N_15062,N_12622,N_12938);
xnor U15063 (N_15063,N_13044,N_14523);
xor U15064 (N_15064,N_13446,N_14570);
or U15065 (N_15065,N_13214,N_14559);
xnor U15066 (N_15066,N_14735,N_12743);
xnor U15067 (N_15067,N_13194,N_14659);
nor U15068 (N_15068,N_14913,N_13621);
or U15069 (N_15069,N_14088,N_12794);
and U15070 (N_15070,N_13469,N_14891);
xnor U15071 (N_15071,N_13159,N_12705);
xor U15072 (N_15072,N_13339,N_12584);
nand U15073 (N_15073,N_13610,N_13634);
nor U15074 (N_15074,N_14549,N_14223);
nand U15075 (N_15075,N_13649,N_13353);
nor U15076 (N_15076,N_13239,N_14879);
nand U15077 (N_15077,N_14679,N_12849);
nand U15078 (N_15078,N_13280,N_12798);
and U15079 (N_15079,N_13137,N_12990);
xor U15080 (N_15080,N_14339,N_13415);
nand U15081 (N_15081,N_13532,N_12506);
nand U15082 (N_15082,N_12851,N_13187);
xnor U15083 (N_15083,N_13255,N_12510);
xor U15084 (N_15084,N_13542,N_13413);
and U15085 (N_15085,N_14473,N_12508);
nor U15086 (N_15086,N_12988,N_14777);
or U15087 (N_15087,N_13917,N_14329);
and U15088 (N_15088,N_13988,N_12757);
and U15089 (N_15089,N_13014,N_12636);
xor U15090 (N_15090,N_13288,N_13855);
nor U15091 (N_15091,N_14291,N_14836);
and U15092 (N_15092,N_13777,N_13778);
xor U15093 (N_15093,N_12975,N_12806);
nand U15094 (N_15094,N_12906,N_14991);
nor U15095 (N_15095,N_12830,N_12550);
nor U15096 (N_15096,N_14902,N_13365);
xor U15097 (N_15097,N_13193,N_13368);
nand U15098 (N_15098,N_13077,N_14432);
or U15099 (N_15099,N_14520,N_14422);
nor U15100 (N_15100,N_12686,N_14456);
nand U15101 (N_15101,N_13069,N_13489);
nand U15102 (N_15102,N_12900,N_12702);
or U15103 (N_15103,N_14890,N_13780);
or U15104 (N_15104,N_13627,N_13217);
xnor U15105 (N_15105,N_13402,N_14824);
or U15106 (N_15106,N_14350,N_12866);
or U15107 (N_15107,N_13393,N_13369);
and U15108 (N_15108,N_12983,N_14807);
xor U15109 (N_15109,N_12566,N_12559);
nand U15110 (N_15110,N_14490,N_13507);
or U15111 (N_15111,N_14155,N_12637);
and U15112 (N_15112,N_13470,N_13483);
xnor U15113 (N_15113,N_13876,N_14279);
nor U15114 (N_15114,N_13846,N_13122);
nor U15115 (N_15115,N_13091,N_14932);
or U15116 (N_15116,N_12553,N_14993);
and U15117 (N_15117,N_14388,N_13463);
xor U15118 (N_15118,N_12525,N_13531);
or U15119 (N_15119,N_12649,N_14167);
or U15120 (N_15120,N_14919,N_13038);
or U15121 (N_15121,N_14332,N_13597);
or U15122 (N_15122,N_14644,N_13421);
xor U15123 (N_15123,N_14680,N_12847);
xnor U15124 (N_15124,N_12714,N_13171);
xor U15125 (N_15125,N_14783,N_13395);
xnor U15126 (N_15126,N_13494,N_14047);
or U15127 (N_15127,N_13768,N_14898);
nand U15128 (N_15128,N_14192,N_13847);
and U15129 (N_15129,N_13937,N_13809);
xnor U15130 (N_15130,N_14277,N_14905);
xor U15131 (N_15131,N_14933,N_12500);
nor U15132 (N_15132,N_14851,N_13403);
nor U15133 (N_15133,N_13033,N_14116);
and U15134 (N_15134,N_13690,N_14754);
xor U15135 (N_15135,N_13423,N_13701);
or U15136 (N_15136,N_14150,N_14687);
and U15137 (N_15137,N_13433,N_13886);
nand U15138 (N_15138,N_13559,N_13766);
nor U15139 (N_15139,N_14002,N_13203);
or U15140 (N_15140,N_13998,N_13303);
nand U15141 (N_15141,N_14119,N_13999);
or U15142 (N_15142,N_13405,N_14453);
nand U15143 (N_15143,N_13930,N_13139);
or U15144 (N_15144,N_14964,N_13950);
nand U15145 (N_15145,N_13282,N_13974);
and U15146 (N_15146,N_13063,N_13020);
or U15147 (N_15147,N_14196,N_14613);
nor U15148 (N_15148,N_13565,N_12602);
nor U15149 (N_15149,N_14372,N_13208);
or U15150 (N_15150,N_13875,N_13052);
nand U15151 (N_15151,N_14056,N_12756);
nand U15152 (N_15152,N_13158,N_14936);
xnor U15153 (N_15153,N_12641,N_13448);
nand U15154 (N_15154,N_14564,N_13716);
nor U15155 (N_15155,N_14396,N_13606);
or U15156 (N_15156,N_13455,N_12853);
xnor U15157 (N_15157,N_14747,N_14354);
and U15158 (N_15158,N_14746,N_14437);
and U15159 (N_15159,N_14513,N_13673);
and U15160 (N_15160,N_13696,N_13845);
nand U15161 (N_15161,N_14537,N_14281);
nor U15162 (N_15162,N_13224,N_14717);
nand U15163 (N_15163,N_14796,N_14946);
nand U15164 (N_15164,N_13892,N_14937);
and U15165 (N_15165,N_12595,N_14501);
nor U15166 (N_15166,N_14825,N_12792);
nand U15167 (N_15167,N_13111,N_14431);
or U15168 (N_15168,N_13262,N_14736);
nor U15169 (N_15169,N_13076,N_13347);
or U15170 (N_15170,N_12799,N_13258);
nor U15171 (N_15171,N_13617,N_14258);
or U15172 (N_15172,N_12958,N_13744);
and U15173 (N_15173,N_14610,N_14685);
nor U15174 (N_15174,N_14959,N_14705);
and U15175 (N_15175,N_14591,N_14389);
and U15176 (N_15176,N_14263,N_12583);
and U15177 (N_15177,N_13880,N_13719);
nor U15178 (N_15178,N_12761,N_12700);
xnor U15179 (N_15179,N_13088,N_12765);
nor U15180 (N_15180,N_14148,N_13043);
nand U15181 (N_15181,N_14022,N_13460);
nand U15182 (N_15182,N_12611,N_13580);
xnor U15183 (N_15183,N_13090,N_14867);
nand U15184 (N_15184,N_13791,N_13399);
and U15185 (N_15185,N_12949,N_14468);
nor U15186 (N_15186,N_13049,N_13284);
xnor U15187 (N_15187,N_13773,N_14665);
xor U15188 (N_15188,N_14908,N_13671);
and U15189 (N_15189,N_13685,N_13555);
nor U15190 (N_15190,N_14773,N_13884);
nand U15191 (N_15191,N_14548,N_14236);
and U15192 (N_15192,N_13447,N_14609);
and U15193 (N_15193,N_13418,N_14224);
xnor U15194 (N_15194,N_14878,N_14286);
nor U15195 (N_15195,N_13485,N_12932);
nor U15196 (N_15196,N_12552,N_13688);
xnor U15197 (N_15197,N_13461,N_14401);
nor U15198 (N_15198,N_13290,N_13591);
xnor U15199 (N_15199,N_12740,N_14496);
or U15200 (N_15200,N_13926,N_13296);
xnor U15201 (N_15201,N_12529,N_13115);
and U15202 (N_15202,N_12824,N_13045);
xor U15203 (N_15203,N_14838,N_12687);
xnor U15204 (N_15204,N_14062,N_12864);
xnor U15205 (N_15205,N_14776,N_14666);
xnor U15206 (N_15206,N_13568,N_13358);
nand U15207 (N_15207,N_12675,N_14753);
and U15208 (N_15208,N_14597,N_14278);
or U15209 (N_15209,N_14906,N_14784);
xor U15210 (N_15210,N_13822,N_14615);
or U15211 (N_15211,N_14226,N_14374);
nand U15212 (N_15212,N_14928,N_12617);
and U15213 (N_15213,N_14604,N_13238);
nor U15214 (N_15214,N_12982,N_13518);
xnor U15215 (N_15215,N_13980,N_14174);
xnor U15216 (N_15216,N_14481,N_14020);
and U15217 (N_15217,N_13117,N_13372);
and U15218 (N_15218,N_13804,N_12998);
nor U15219 (N_15219,N_14512,N_14572);
and U15220 (N_15220,N_12633,N_13292);
xnor U15221 (N_15221,N_13703,N_13990);
nand U15222 (N_15222,N_14611,N_13453);
nor U15223 (N_15223,N_13916,N_13031);
or U15224 (N_15224,N_14926,N_14706);
nor U15225 (N_15225,N_12981,N_14364);
nand U15226 (N_15226,N_14573,N_13965);
xor U15227 (N_15227,N_13397,N_13592);
nand U15228 (N_15228,N_12838,N_14653);
and U15229 (N_15229,N_14010,N_12681);
or U15230 (N_15230,N_14800,N_13150);
and U15231 (N_15231,N_14060,N_12653);
nand U15232 (N_15232,N_13912,N_14467);
nor U15233 (N_15233,N_12968,N_13769);
or U15234 (N_15234,N_14267,N_13449);
and U15235 (N_15235,N_13981,N_14288);
or U15236 (N_15236,N_13545,N_14628);
xnor U15237 (N_15237,N_14025,N_13281);
nand U15238 (N_15238,N_13272,N_14311);
nand U15239 (N_15239,N_14647,N_13835);
nor U15240 (N_15240,N_14742,N_14156);
xor U15241 (N_15241,N_12913,N_14065);
nand U15242 (N_15242,N_13196,N_12728);
xnor U15243 (N_15243,N_13220,N_13398);
nor U15244 (N_15244,N_14469,N_12616);
or U15245 (N_15245,N_14027,N_12967);
nand U15246 (N_15246,N_13225,N_13725);
nand U15247 (N_15247,N_12669,N_14111);
xor U15248 (N_15248,N_14474,N_13589);
or U15249 (N_15249,N_13560,N_14127);
nor U15250 (N_15250,N_14818,N_14115);
and U15251 (N_15251,N_12883,N_13888);
or U15252 (N_15252,N_14566,N_13746);
nor U15253 (N_15253,N_14066,N_12762);
nand U15254 (N_15254,N_12797,N_14532);
xnor U15255 (N_15255,N_14285,N_14418);
nand U15256 (N_15256,N_14727,N_13924);
nor U15257 (N_15257,N_13514,N_14147);
nand U15258 (N_15258,N_12995,N_13704);
and U15259 (N_15259,N_14662,N_14560);
nor U15260 (N_15260,N_12671,N_13953);
or U15261 (N_15261,N_14865,N_13012);
nand U15262 (N_15262,N_14341,N_14953);
and U15263 (N_15263,N_12903,N_14883);
xor U15264 (N_15264,N_12661,N_14333);
nand U15265 (N_15265,N_13186,N_12694);
nor U15266 (N_15266,N_14255,N_13904);
or U15267 (N_15267,N_13082,N_13141);
nor U15268 (N_15268,N_13788,N_13711);
nor U15269 (N_15269,N_14620,N_14299);
or U15270 (N_15270,N_14857,N_12736);
and U15271 (N_15271,N_14528,N_13179);
nor U15272 (N_15272,N_13271,N_12754);
xnor U15273 (N_15273,N_13902,N_14663);
or U15274 (N_15274,N_14232,N_13819);
nand U15275 (N_15275,N_13541,N_12629);
xnor U15276 (N_15276,N_14827,N_12989);
or U15277 (N_15277,N_12570,N_13414);
or U15278 (N_15278,N_14442,N_14077);
xnor U15279 (N_15279,N_14786,N_14541);
or U15280 (N_15280,N_13969,N_13278);
nor U15281 (N_15281,N_13182,N_13000);
nand U15282 (N_15282,N_14975,N_14227);
nor U15283 (N_15283,N_14063,N_14045);
xnor U15284 (N_15284,N_14312,N_14208);
or U15285 (N_15285,N_14252,N_14318);
and U15286 (N_15286,N_13384,N_12936);
nor U15287 (N_15287,N_14449,N_13342);
nor U15288 (N_15288,N_14382,N_13144);
or U15289 (N_15289,N_14028,N_12678);
nor U15290 (N_15290,N_12748,N_13248);
nand U15291 (N_15291,N_14538,N_12943);
xnor U15292 (N_15292,N_13730,N_14596);
nor U15293 (N_15293,N_12620,N_14812);
nor U15294 (N_15294,N_13806,N_13452);
nor U15295 (N_15295,N_12572,N_12815);
nor U15296 (N_15296,N_13135,N_14657);
and U15297 (N_15297,N_14406,N_13600);
and U15298 (N_15298,N_14871,N_14454);
nand U15299 (N_15299,N_13897,N_12813);
xor U15300 (N_15300,N_14131,N_14268);
nand U15301 (N_15301,N_14545,N_13001);
xor U15302 (N_15302,N_13246,N_13661);
nand U15303 (N_15303,N_13259,N_14962);
xor U15304 (N_15304,N_13923,N_13645);
nor U15305 (N_15305,N_13301,N_13860);
nand U15306 (N_15306,N_13046,N_14213);
or U15307 (N_15307,N_14648,N_14164);
xor U15308 (N_15308,N_14669,N_13445);
or U15309 (N_15309,N_12638,N_13213);
or U15310 (N_15310,N_13106,N_13834);
and U15311 (N_15311,N_14270,N_13491);
and U15312 (N_15312,N_13658,N_14390);
and U15313 (N_15313,N_14228,N_14133);
or U15314 (N_15314,N_13073,N_13513);
nand U15315 (N_15315,N_14804,N_14497);
and U15316 (N_15316,N_13827,N_13336);
nor U15317 (N_15317,N_12727,N_13266);
or U15318 (N_15318,N_14592,N_14884);
nor U15319 (N_15319,N_13315,N_14096);
xor U15320 (N_15320,N_12827,N_13830);
xnor U15321 (N_15321,N_13665,N_13997);
xnor U15322 (N_15322,N_14494,N_14385);
nand U15323 (N_15323,N_14106,N_14756);
nor U15324 (N_15324,N_14349,N_13047);
nor U15325 (N_15325,N_14029,N_13120);
xor U15326 (N_15326,N_14426,N_14443);
nor U15327 (N_15327,N_14729,N_14927);
and U15328 (N_15328,N_14169,N_13670);
or U15329 (N_15329,N_13588,N_14014);
xor U15330 (N_15330,N_14308,N_13154);
nand U15331 (N_15331,N_13623,N_13401);
nand U15332 (N_15332,N_14626,N_13682);
nand U15333 (N_15333,N_13891,N_13613);
nor U15334 (N_15334,N_13816,N_13134);
nand U15335 (N_15335,N_13375,N_13466);
nor U15336 (N_15336,N_13624,N_14085);
nand U15337 (N_15337,N_12537,N_12786);
nand U15338 (N_15338,N_13011,N_13802);
and U15339 (N_15339,N_13192,N_14275);
and U15340 (N_15340,N_13307,N_12873);
and U15341 (N_15341,N_13853,N_13717);
and U15342 (N_15342,N_13216,N_14108);
xnor U15343 (N_15343,N_12612,N_13210);
nand U15344 (N_15344,N_12571,N_13253);
nor U15345 (N_15345,N_13409,N_14184);
nor U15346 (N_15346,N_12737,N_13938);
or U15347 (N_15347,N_14451,N_13803);
and U15348 (N_15348,N_13550,N_14760);
nor U15349 (N_15349,N_14099,N_12544);
and U15350 (N_15350,N_13464,N_12541);
or U15351 (N_15351,N_13496,N_13863);
nand U15352 (N_15352,N_14144,N_13814);
and U15353 (N_15353,N_14375,N_12946);
nand U15354 (N_15354,N_14641,N_14023);
and U15355 (N_15355,N_12939,N_13364);
nor U15356 (N_15356,N_14204,N_13681);
xnor U15357 (N_15357,N_13492,N_13710);
or U15358 (N_15358,N_13859,N_14245);
and U15359 (N_15359,N_13166,N_12895);
nand U15360 (N_15360,N_14290,N_13877);
nand U15361 (N_15361,N_14949,N_14939);
and U15362 (N_15362,N_14216,N_13810);
or U15363 (N_15363,N_13850,N_14790);
and U15364 (N_15364,N_13242,N_13006);
xor U15365 (N_15365,N_12954,N_12993);
and U15366 (N_15366,N_14918,N_14071);
or U15367 (N_15367,N_12645,N_14846);
or U15368 (N_15368,N_13918,N_14911);
nor U15369 (N_15369,N_12905,N_14452);
nand U15370 (N_15370,N_14059,N_14321);
and U15371 (N_15371,N_13331,N_14187);
xnor U15372 (N_15372,N_13986,N_13407);
nor U15373 (N_15373,N_12941,N_12626);
xor U15374 (N_15374,N_14831,N_14672);
and U15375 (N_15375,N_13826,N_14157);
nor U15376 (N_15376,N_14097,N_13388);
nand U15377 (N_15377,N_12805,N_14745);
or U15378 (N_15378,N_14915,N_12920);
and U15379 (N_15379,N_12590,N_13865);
nand U15380 (N_15380,N_14661,N_14324);
xor U15381 (N_15381,N_14798,N_12625);
and U15382 (N_15382,N_13913,N_14811);
nor U15383 (N_15383,N_13519,N_14708);
and U15384 (N_15384,N_12543,N_14072);
xor U15385 (N_15385,N_14325,N_14580);
or U15386 (N_15386,N_14552,N_13270);
xor U15387 (N_15387,N_12929,N_13456);
and U15388 (N_15388,N_13350,N_13286);
or U15389 (N_15389,N_13838,N_14404);
and U15390 (N_15390,N_13503,N_12979);
nor U15391 (N_15391,N_14415,N_12679);
and U15392 (N_15392,N_14380,N_13003);
or U15393 (N_15393,N_13320,N_12667);
nand U15394 (N_15394,N_14677,N_13479);
and U15395 (N_15395,N_14583,N_13429);
nand U15396 (N_15396,N_14539,N_13871);
or U15397 (N_15397,N_12601,N_14006);
nand U15398 (N_15398,N_13854,N_13306);
nand U15399 (N_15399,N_14860,N_14858);
nand U15400 (N_15400,N_12999,N_14785);
and U15401 (N_15401,N_13297,N_14362);
nor U15402 (N_15402,N_14938,N_12837);
nand U15403 (N_15403,N_12632,N_12648);
or U15404 (N_15404,N_14651,N_12844);
xnor U15405 (N_15405,N_13202,N_14810);
xnor U15406 (N_15406,N_14612,N_13944);
nand U15407 (N_15407,N_12840,N_12944);
nor U15408 (N_15408,N_12885,N_14813);
or U15409 (N_15409,N_14035,N_14688);
nand U15410 (N_15410,N_12646,N_12518);
nand U15411 (N_15411,N_13551,N_14897);
and U15412 (N_15412,N_14994,N_14120);
or U15413 (N_15413,N_13007,N_13772);
or U15414 (N_15414,N_14486,N_12763);
xnor U15415 (N_15415,N_14185,N_14466);
and U15416 (N_15416,N_13636,N_12801);
or U15417 (N_15417,N_13434,N_13939);
xnor U15418 (N_15418,N_13321,N_14220);
and U15419 (N_15419,N_14606,N_13361);
and U15420 (N_15420,N_14681,N_13651);
nand U15421 (N_15421,N_14634,N_12841);
nand U15422 (N_15422,N_13495,N_13656);
or U15423 (N_15423,N_14498,N_13209);
and U15424 (N_15424,N_14242,N_14061);
or U15425 (N_15425,N_14877,N_13967);
or U15426 (N_15426,N_13390,N_14082);
or U15427 (N_15427,N_14394,N_13066);
xor U15428 (N_15428,N_14887,N_13952);
xnor U15429 (N_15429,N_13714,N_14142);
and U15430 (N_15430,N_12817,N_12787);
and U15431 (N_15431,N_13818,N_13343);
and U15432 (N_15432,N_14584,N_13660);
xor U15433 (N_15433,N_13180,N_13737);
nor U15434 (N_15434,N_12603,N_14042);
and U15435 (N_15435,N_13611,N_14000);
or U15436 (N_15436,N_12862,N_13586);
xor U15437 (N_15437,N_14849,N_14575);
nand U15438 (N_15438,N_14912,N_13757);
or U15439 (N_15439,N_13363,N_13946);
nor U15440 (N_15440,N_14392,N_13895);
and U15441 (N_15441,N_14778,N_13692);
and U15442 (N_15442,N_13157,N_14343);
nor U15443 (N_15443,N_13468,N_14670);
xnor U15444 (N_15444,N_13724,N_14433);
or U15445 (N_15445,N_14733,N_14594);
and U15446 (N_15446,N_13153,N_13273);
xnor U15447 (N_15447,N_14054,N_13638);
nand U15448 (N_15448,N_14386,N_12746);
xor U15449 (N_15449,N_13475,N_14462);
or U15450 (N_15450,N_13858,N_14011);
and U15451 (N_15451,N_12621,N_14974);
nor U15452 (N_15452,N_13702,N_13957);
xnor U15453 (N_15453,N_12513,N_13932);
nand U15454 (N_15454,N_13867,N_14519);
or U15455 (N_15455,N_14668,N_12908);
or U15456 (N_15456,N_13700,N_13861);
nand U15457 (N_15457,N_14191,N_12876);
nor U15458 (N_15458,N_14676,N_13506);
or U15459 (N_15459,N_14305,N_14992);
nor U15460 (N_15460,N_14876,N_13484);
nand U15461 (N_15461,N_13779,N_13005);
nor U15462 (N_15462,N_12574,N_14698);
nand U15463 (N_15463,N_13098,N_12962);
or U15464 (N_15464,N_14750,N_13247);
and U15465 (N_15465,N_14221,N_14231);
nand U15466 (N_15466,N_13438,N_14159);
nand U15467 (N_15467,N_13474,N_14287);
or U15468 (N_15468,N_14985,N_13662);
or U15469 (N_15469,N_13057,N_14408);
nor U15470 (N_15470,N_13709,N_12768);
and U15471 (N_15471,N_13961,N_14143);
nand U15472 (N_15472,N_13380,N_12919);
or U15473 (N_15473,N_12779,N_13512);
or U15474 (N_15474,N_13812,N_12959);
nand U15475 (N_15475,N_13498,N_14013);
nor U15476 (N_15476,N_13302,N_14585);
and U15477 (N_15477,N_13143,N_14546);
and U15478 (N_15478,N_13112,N_13813);
and U15479 (N_15479,N_12618,N_14274);
or U15480 (N_15480,N_14043,N_13622);
nand U15481 (N_15481,N_14068,N_13116);
or U15482 (N_15482,N_14900,N_13837);
nor U15483 (N_15483,N_13960,N_13008);
nand U15484 (N_15484,N_13529,N_13298);
and U15485 (N_15485,N_13893,N_13308);
nor U15486 (N_15486,N_14441,N_14005);
or U15487 (N_15487,N_14684,N_13108);
xnor U15488 (N_15488,N_14749,N_12869);
xor U15489 (N_15489,N_12843,N_13207);
nand U15490 (N_15490,N_14979,N_14440);
and U15491 (N_15491,N_14924,N_14734);
nor U15492 (N_15492,N_12901,N_13328);
nand U15493 (N_15493,N_14487,N_13473);
nor U15494 (N_15494,N_14909,N_14700);
and U15495 (N_15495,N_13832,N_14799);
xnor U15496 (N_15496,N_14320,N_12615);
nor U15497 (N_15497,N_12778,N_14319);
and U15498 (N_15498,N_14322,N_12888);
xor U15499 (N_15499,N_14709,N_14856);
nand U15500 (N_15500,N_13079,N_13570);
nand U15501 (N_15501,N_14917,N_13732);
nand U15502 (N_15502,N_13553,N_13508);
xnor U15503 (N_15503,N_12524,N_13729);
or U15504 (N_15504,N_12732,N_13971);
nor U15505 (N_15505,N_14493,N_14737);
nand U15506 (N_15506,N_13333,N_13740);
nor U15507 (N_15507,N_14531,N_13481);
or U15508 (N_15508,N_12812,N_14089);
nor U15509 (N_15509,N_14716,N_14193);
xor U15510 (N_15510,N_14740,N_14635);
or U15511 (N_15511,N_14759,N_13105);
nand U15512 (N_15512,N_14639,N_13502);
nand U15513 (N_15513,N_12915,N_13684);
and U15514 (N_15514,N_14488,N_13392);
or U15515 (N_15515,N_12565,N_14847);
or U15516 (N_15516,N_13686,N_14843);
nand U15517 (N_15517,N_14499,N_12904);
or U15518 (N_15518,N_14981,N_14303);
nand U15519 (N_15519,N_14457,N_13130);
xnor U15520 (N_15520,N_14896,N_14313);
and U15521 (N_15521,N_14916,N_13929);
nand U15522 (N_15522,N_14057,N_14237);
nand U15523 (N_15523,N_14310,N_12751);
xnor U15524 (N_15524,N_14282,N_13594);
xor U15525 (N_15525,N_14105,N_14752);
nand U15526 (N_15526,N_14558,N_13533);
xnor U15527 (N_15527,N_12684,N_13821);
nand U15528 (N_15528,N_13383,N_14861);
xnor U15529 (N_15529,N_14791,N_14446);
xor U15530 (N_15530,N_12854,N_13800);
or U15531 (N_15531,N_13607,N_13412);
nor U15532 (N_15532,N_14038,N_14870);
nand U15533 (N_15533,N_13985,N_14788);
and U15534 (N_15534,N_13878,N_13124);
xor U15535 (N_15535,N_13269,N_14823);
xor U15536 (N_15536,N_12558,N_13945);
xnor U15537 (N_15537,N_13973,N_14003);
or U15538 (N_15538,N_13603,N_14533);
nor U15539 (N_15539,N_14690,N_13679);
and U15540 (N_15540,N_13417,N_14833);
nor U15541 (N_15541,N_12692,N_12512);
nor U15542 (N_15542,N_13018,N_13748);
or U15543 (N_15543,N_13478,N_14229);
xnor U15544 (N_15544,N_13678,N_12781);
or U15545 (N_15545,N_13616,N_14910);
and U15546 (N_15546,N_14098,N_13996);
xor U15547 (N_15547,N_13454,N_14428);
or U15548 (N_15548,N_14276,N_13628);
nor U15549 (N_15549,N_12729,N_14083);
nor U15550 (N_15550,N_12826,N_14567);
xor U15551 (N_15551,N_13815,N_14210);
xor U15552 (N_15552,N_14413,N_14982);
and U15553 (N_15553,N_14976,N_14682);
and U15554 (N_15554,N_14205,N_13092);
nand U15555 (N_15555,N_14781,N_13752);
nor U15556 (N_15556,N_12914,N_12725);
or U15557 (N_15557,N_12970,N_14787);
xnor U15558 (N_15558,N_13776,N_14271);
nor U15559 (N_15559,N_12807,N_14090);
xnor U15560 (N_15560,N_14145,N_13465);
nand U15561 (N_15561,N_13081,N_14129);
nand U15562 (N_15562,N_13760,N_14424);
nand U15563 (N_15563,N_13019,N_13200);
and U15564 (N_15564,N_14901,N_14990);
and U15565 (N_15565,N_13713,N_13335);
nand U15566 (N_15566,N_13516,N_14176);
and U15567 (N_15567,N_14427,N_13840);
and U15568 (N_15568,N_12822,N_12764);
nor U15569 (N_15569,N_14630,N_13326);
and U15570 (N_15570,N_14724,N_14489);
xor U15571 (N_15571,N_12592,N_13026);
and U15572 (N_15572,N_12576,N_13820);
xnor U15573 (N_15573,N_13206,N_14899);
nor U15574 (N_15574,N_13500,N_14803);
nand U15575 (N_15575,N_13316,N_14862);
nor U15576 (N_15576,N_14686,N_12707);
and U15577 (N_15577,N_12502,N_13071);
xor U15578 (N_15578,N_12957,N_14563);
or U15579 (N_15579,N_12788,N_12889);
nor U15580 (N_15580,N_13344,N_14730);
or U15581 (N_15581,N_14829,N_13749);
xnor U15582 (N_15582,N_13528,N_13215);
nor U15583 (N_15583,N_13118,N_14149);
nor U15584 (N_15584,N_12770,N_12672);
nor U15585 (N_15585,N_14347,N_13882);
or U15586 (N_15586,N_14298,N_13404);
nand U15587 (N_15587,N_12880,N_14351);
nand U15588 (N_15588,N_13083,N_12660);
nor U15589 (N_15589,N_14365,N_13385);
and U15590 (N_15590,N_14762,N_14925);
nor U15591 (N_15591,N_14017,N_13608);
or U15592 (N_15592,N_13431,N_12769);
xor U15593 (N_15593,N_12814,N_14363);
and U15594 (N_15594,N_12832,N_14058);
or U15595 (N_15595,N_13146,N_14186);
nand U15596 (N_15596,N_14300,N_14140);
or U15597 (N_15597,N_13056,N_13763);
nor U15598 (N_15598,N_12829,N_14342);
xor U15599 (N_15599,N_12991,N_14977);
and U15600 (N_15600,N_13476,N_13218);
xnor U15601 (N_15601,N_13577,N_12530);
nand U15602 (N_15602,N_14175,N_12878);
and U15603 (N_15603,N_13523,N_13992);
nor U15604 (N_15604,N_13123,N_13705);
or U15605 (N_15605,N_13764,N_14190);
nor U15606 (N_15606,N_14625,N_13305);
nor U15607 (N_15607,N_12789,N_13156);
xnor U15608 (N_15608,N_12758,N_13334);
or U15609 (N_15609,N_12969,N_12540);
nor U15610 (N_15610,N_13657,N_14033);
or U15611 (N_15611,N_14886,N_14366);
nand U15612 (N_15612,N_13524,N_13889);
and U15613 (N_15613,N_14516,N_13068);
and U15614 (N_15614,N_13504,N_14198);
xor U15615 (N_15615,N_12685,N_13697);
nand U15616 (N_15616,N_13067,N_13175);
nor U15617 (N_15617,N_12708,N_12921);
or U15618 (N_15618,N_14348,N_14165);
or U15619 (N_15619,N_14302,N_14067);
xnor U15620 (N_15620,N_13609,N_12997);
nand U15621 (N_15621,N_14809,N_13612);
nand U15622 (N_15622,N_14557,N_13467);
xor U15623 (N_15623,N_13199,N_14036);
nor U15624 (N_15624,N_12662,N_14774);
or U15625 (N_15625,N_13870,N_13313);
and U15626 (N_15626,N_12777,N_13095);
and U15627 (N_15627,N_14075,N_13275);
nor U15628 (N_15628,N_12604,N_14244);
xor U15629 (N_15629,N_12693,N_14885);
nand U15630 (N_15630,N_13230,N_13002);
and U15631 (N_15631,N_14587,N_14859);
nor U15632 (N_15632,N_13741,N_14358);
and U15633 (N_15633,N_13360,N_14576);
and U15634 (N_15634,N_12634,N_14868);
xnor U15635 (N_15635,N_14225,N_13107);
xor U15636 (N_15636,N_14447,N_12974);
or U15637 (N_15637,N_14234,N_14888);
or U15638 (N_15638,N_14699,N_13534);
xor U15639 (N_15639,N_13222,N_13626);
nand U15640 (N_15640,N_14421,N_14114);
nor U15641 (N_15641,N_14021,N_12511);
xor U15642 (N_15642,N_12655,N_12713);
and U15643 (N_15643,N_14243,N_13605);
xor U15644 (N_15644,N_13984,N_14893);
and U15645 (N_15645,N_13291,N_14645);
nor U15646 (N_15646,N_13629,N_13659);
nor U15647 (N_15647,N_13899,N_12845);
nand U15648 (N_15648,N_14168,N_13021);
nor U15649 (N_15649,N_13852,N_12774);
or U15650 (N_15650,N_14438,N_13055);
or U15651 (N_15651,N_13751,N_13499);
xnor U15652 (N_15652,N_14779,N_14118);
nand U15653 (N_15653,N_12551,N_14547);
xnor U15654 (N_15654,N_12613,N_13293);
and U15655 (N_15655,N_13520,N_13894);
xor U15656 (N_15656,N_13024,N_12749);
nor U15657 (N_15657,N_13100,N_14079);
or U15658 (N_15658,N_13097,N_14439);
nand U15659 (N_15659,N_13669,N_14403);
xnor U15660 (N_15660,N_14608,N_13547);
nor U15661 (N_15661,N_14955,N_14125);
nor U15662 (N_15662,N_13437,N_13652);
xnor U15663 (N_15663,N_12690,N_12809);
nor U15664 (N_15664,N_14840,N_13786);
nor U15665 (N_15665,N_13515,N_12894);
or U15666 (N_15666,N_14922,N_13110);
nor U15667 (N_15667,N_14769,N_13976);
nor U15668 (N_15668,N_12780,N_13048);
and U15669 (N_15669,N_13131,N_13549);
xnor U15670 (N_15670,N_13994,N_13311);
and U15671 (N_15671,N_13903,N_14970);
xnor U15672 (N_15672,N_13354,N_12952);
xnor U15673 (N_15673,N_12872,N_14854);
xor U15674 (N_15674,N_14405,N_13190);
nor U15675 (N_15675,N_13979,N_14044);
or U15676 (N_15676,N_14491,N_12600);
nor U15677 (N_15677,N_14757,N_14605);
or U15678 (N_15678,N_13172,N_13625);
and U15679 (N_15679,N_13432,N_14654);
nor U15680 (N_15680,N_14632,N_13260);
nor U15681 (N_15681,N_14795,N_13420);
or U15682 (N_15682,N_13191,N_13371);
xnor U15683 (N_15683,N_13126,N_13511);
xnor U15684 (N_15684,N_14235,N_14306);
nor U15685 (N_15685,N_13543,N_13377);
nand U15686 (N_15686,N_13136,N_12893);
xor U15687 (N_15687,N_12771,N_14095);
nor U15688 (N_15688,N_12673,N_14455);
nor U15689 (N_15689,N_14866,N_14658);
or U15690 (N_15690,N_13229,N_13323);
xnor U15691 (N_15691,N_14507,N_13576);
nand U15692 (N_15692,N_14074,N_12721);
or U15693 (N_15693,N_13908,N_13578);
xnor U15694 (N_15694,N_13964,N_14598);
or U15695 (N_15695,N_13346,N_13948);
and U15696 (N_15696,N_12767,N_14214);
or U15697 (N_15697,N_13666,N_13128);
and U15698 (N_15698,N_13942,N_14980);
nand U15699 (N_15699,N_13650,N_12554);
nand U15700 (N_15700,N_14616,N_14173);
xnor U15701 (N_15701,N_14640,N_13319);
and U15702 (N_15702,N_13155,N_14248);
or U15703 (N_15703,N_13085,N_14397);
or U15704 (N_15704,N_12709,N_13486);
xor U15705 (N_15705,N_14711,N_12773);
xnor U15706 (N_15706,N_13956,N_13632);
xor U15707 (N_15707,N_13329,N_13522);
or U15708 (N_15708,N_14808,N_12627);
xor U15709 (N_15709,N_13868,N_13731);
nor U15710 (N_15710,N_14535,N_13037);
nor U15711 (N_15711,N_14622,N_14177);
and U15712 (N_15712,N_13811,N_14246);
nand U15713 (N_15713,N_13721,N_13771);
and U15714 (N_15714,N_13173,N_12925);
and U15715 (N_15715,N_14881,N_13641);
xnor U15716 (N_15716,N_14222,N_13619);
and U15717 (N_15717,N_13635,N_14758);
or U15718 (N_15718,N_12591,N_14624);
nand U15719 (N_15719,N_14534,N_13029);
nand U15720 (N_15720,N_12596,N_13604);
nor U15721 (N_15721,N_13501,N_14948);
or U15722 (N_15722,N_14674,N_13546);
nand U15723 (N_15723,N_13164,N_13557);
nand U15724 (N_15724,N_14816,N_13739);
and U15725 (N_15725,N_12803,N_12987);
xnor U15726 (N_15726,N_13304,N_12842);
nor U15727 (N_15727,N_14503,N_13587);
or U15728 (N_15728,N_12892,N_13699);
nor U15729 (N_15729,N_13968,N_14104);
and U15730 (N_15730,N_12664,N_13911);
nor U15731 (N_15731,N_13338,N_12861);
nor U15732 (N_15732,N_14732,N_12886);
or U15733 (N_15733,N_14923,N_13955);
or U15734 (N_15734,N_13790,N_13574);
or U15735 (N_15735,N_13907,N_14819);
and U15736 (N_15736,N_14815,N_12945);
nor U15737 (N_15737,N_13537,N_12755);
nand U15738 (N_15738,N_14051,N_14841);
and U15739 (N_15739,N_13035,N_14134);
or U15740 (N_15740,N_14377,N_14331);
nand U15741 (N_15741,N_13795,N_13920);
and U15742 (N_15742,N_14554,N_13458);
and U15743 (N_15743,N_13836,N_14942);
nand U15744 (N_15744,N_14579,N_13276);
nand U15745 (N_15745,N_13527,N_12726);
nand U15746 (N_15746,N_14617,N_12759);
and U15747 (N_15747,N_14425,N_13138);
nand U15748 (N_15748,N_12735,N_14500);
nand U15749 (N_15749,N_12808,N_13742);
nor U15750 (N_15750,N_12747,N_12573);
nor U15751 (N_15751,N_13646,N_14621);
or U15752 (N_15752,N_12966,N_14436);
nand U15753 (N_15753,N_13849,N_14336);
or U15754 (N_15754,N_14470,N_14307);
xnor U15755 (N_15755,N_13833,N_14947);
xor U15756 (N_15756,N_12795,N_14113);
xnor U15757 (N_15757,N_14599,N_14007);
and U15758 (N_15758,N_13767,N_13406);
xnor U15759 (N_15759,N_13219,N_14112);
xnor U15760 (N_15760,N_12609,N_14475);
nand U15761 (N_15761,N_14110,N_13283);
nand U15762 (N_15762,N_14693,N_12828);
nor U15763 (N_15763,N_12972,N_13324);
and U15764 (N_15764,N_12528,N_13927);
nor U15765 (N_15765,N_14410,N_13977);
or U15766 (N_15766,N_14929,N_13424);
or U15767 (N_15767,N_13677,N_14409);
and U15768 (N_15768,N_13036,N_13579);
nor U15769 (N_15769,N_14801,N_14952);
nor U15770 (N_15770,N_13921,N_13851);
and U15771 (N_15771,N_12937,N_12724);
or U15772 (N_15772,N_13723,N_14999);
or U15773 (N_15773,N_13544,N_13023);
nand U15774 (N_15774,N_13410,N_13905);
nand U15775 (N_15775,N_14217,N_12556);
xor U15776 (N_15776,N_14069,N_14219);
nor U15777 (N_15777,N_12926,N_14166);
nand U15778 (N_15778,N_13928,N_12699);
nand U15779 (N_15779,N_14954,N_12956);
and U15780 (N_15780,N_14154,N_14965);
nand U15781 (N_15781,N_13536,N_14960);
nor U15782 (N_15782,N_12631,N_12984);
and U15783 (N_15783,N_13376,N_12859);
nor U15784 (N_15784,N_12668,N_13548);
nor U15785 (N_15785,N_14853,N_14505);
nand U15786 (N_15786,N_13330,N_14722);
nand U15787 (N_15787,N_12689,N_13736);
or U15788 (N_15788,N_14767,N_12663);
xor U15789 (N_15789,N_14338,N_14461);
nor U15790 (N_15790,N_12891,N_12833);
nor U15791 (N_15791,N_13103,N_14542);
nand U15792 (N_15792,N_14696,N_12857);
xnor U15793 (N_15793,N_14162,N_12516);
nor U15794 (N_15794,N_13152,N_13630);
nand U15795 (N_15795,N_13183,N_14544);
nand U15796 (N_15796,N_13104,N_14052);
nor U15797 (N_15797,N_14792,N_13824);
xor U15798 (N_15798,N_12867,N_14763);
nand U15799 (N_15799,N_14464,N_14650);
and U15800 (N_15800,N_14988,N_14262);
xnor U15801 (N_15801,N_14247,N_12585);
and U15802 (N_15802,N_13250,N_13575);
nand U15803 (N_15803,N_12642,N_13345);
xor U15804 (N_15804,N_14543,N_13715);
and U15805 (N_15805,N_12928,N_14053);
nor U15806 (N_15806,N_14969,N_14805);
nand U15807 (N_15807,N_12582,N_14691);
nand U15808 (N_15808,N_14340,N_12619);
xnor U15809 (N_15809,N_14101,N_13966);
xor U15810 (N_15810,N_14109,N_12654);
nand U15811 (N_15811,N_14667,N_13535);
or U15812 (N_15812,N_13526,N_14212);
and U15813 (N_15813,N_13505,N_14233);
nand U15814 (N_15814,N_14578,N_13844);
nand U15815 (N_15815,N_13400,N_14444);
and U15816 (N_15816,N_13914,N_13941);
xor U15817 (N_15817,N_14703,N_12882);
and U15818 (N_15818,N_14093,N_12580);
xor U15819 (N_15819,N_13801,N_14577);
nor U15820 (N_15820,N_13025,N_13234);
and U15821 (N_15821,N_13362,N_12963);
and U15822 (N_15822,N_13086,N_13718);
nor U15823 (N_15823,N_14179,N_14768);
nand U15824 (N_15824,N_13439,N_13053);
nor U15825 (N_15825,N_13691,N_14200);
and U15826 (N_15826,N_13762,N_14373);
nand U15827 (N_15827,N_12688,N_13256);
xor U15828 (N_15828,N_14850,N_13734);
and U15829 (N_15829,N_13954,N_12526);
nor U15830 (N_15830,N_14266,N_12977);
or U15831 (N_15831,N_12561,N_12640);
xor U15832 (N_15832,N_13357,N_13240);
or U15833 (N_15833,N_12519,N_13178);
xor U15834 (N_15834,N_13770,N_14032);
and U15835 (N_15835,N_12695,N_13857);
or U15836 (N_15836,N_14450,N_13140);
nand U15837 (N_15837,N_12624,N_14304);
and U15838 (N_15838,N_14379,N_13925);
or U15839 (N_15839,N_12947,N_13087);
nand U15840 (N_15840,N_12793,N_14903);
and U15841 (N_15841,N_12711,N_14834);
xnor U15842 (N_15842,N_12608,N_13841);
nor U15843 (N_15843,N_13490,N_13829);
or U15844 (N_15844,N_14294,N_12910);
nor U15845 (N_15845,N_14943,N_14842);
xor U15846 (N_15846,N_14309,N_14117);
xnor U15847 (N_15847,N_14832,N_14376);
or U15848 (N_15848,N_14086,N_14423);
or U15849 (N_15849,N_14820,N_12676);
or U15850 (N_15850,N_13197,N_14772);
nand U15851 (N_15851,N_12994,N_13462);
nand U15852 (N_15852,N_13598,N_13792);
nor U15853 (N_15853,N_14181,N_13680);
or U15854 (N_15854,N_14770,N_13901);
and U15855 (N_15855,N_12531,N_13540);
nand U15856 (N_15856,N_14723,N_13951);
xor U15857 (N_15857,N_14138,N_13181);
nor U15858 (N_15858,N_14702,N_12902);
or U15859 (N_15859,N_13267,N_14581);
nor U15860 (N_15860,N_14435,N_14484);
xnor U15861 (N_15861,N_13995,N_14283);
nor U15862 (N_15862,N_13743,N_13883);
nand U15863 (N_15863,N_12831,N_12501);
or U15864 (N_15864,N_12564,N_13349);
nand U15865 (N_15865,N_13864,N_12545);
nand U15866 (N_15866,N_14713,N_14821);
and U15867 (N_15867,N_13382,N_12589);
nor U15868 (N_15868,N_12539,N_13805);
nor U15869 (N_15869,N_14565,N_13784);
nand U15870 (N_15870,N_12534,N_14107);
nor U15871 (N_15871,N_13602,N_14430);
and U15872 (N_15872,N_14084,N_13148);
nand U15873 (N_15873,N_14508,N_14553);
xnor U15874 (N_15874,N_12715,N_14614);
nor U15875 (N_15875,N_12796,N_14967);
and U15876 (N_15876,N_13887,N_14623);
and U15877 (N_15877,N_13698,N_13972);
and U15878 (N_15878,N_14369,N_13185);
or U15879 (N_15879,N_13596,N_14419);
xor U15880 (N_15880,N_14230,N_13590);
xnor U15881 (N_15881,N_14875,N_13869);
or U15882 (N_15882,N_12606,N_12630);
nor U15883 (N_15883,N_13102,N_13530);
or U15884 (N_15884,N_14845,N_13351);
xnor U15885 (N_15885,N_12911,N_14971);
nand U15886 (N_15886,N_13340,N_14472);
and U15887 (N_15887,N_12935,N_12691);
and U15888 (N_15888,N_14720,N_13327);
nor U15889 (N_15889,N_14171,N_13643);
nor U15890 (N_15890,N_14797,N_14360);
and U15891 (N_15891,N_14826,N_14963);
or U15892 (N_15892,N_12623,N_13317);
and U15893 (N_15893,N_14257,N_12639);
nor U15894 (N_15894,N_14458,N_14848);
and U15895 (N_15895,N_12575,N_12930);
nor U15896 (N_15896,N_12874,N_13664);
and U15897 (N_15897,N_13381,N_13631);
or U15898 (N_15898,N_14844,N_14715);
or U15899 (N_15899,N_12848,N_12503);
nor U15900 (N_15900,N_14238,N_14920);
and U15901 (N_15901,N_14889,N_14692);
nand U15902 (N_15902,N_14710,N_14951);
xnor U15903 (N_15903,N_12597,N_14412);
or U15904 (N_15904,N_13663,N_13300);
nand U15905 (N_15905,N_14250,N_14064);
xor U15906 (N_15906,N_13257,N_13416);
nand U15907 (N_15907,N_13084,N_14731);
or U15908 (N_15908,N_13428,N_12775);
nand U15909 (N_15909,N_12931,N_14741);
nand U15910 (N_15910,N_13785,N_14352);
nor U15911 (N_15911,N_12579,N_14619);
nand U15912 (N_15912,N_14675,N_14158);
xor U15913 (N_15913,N_14315,N_12933);
nor U15914 (N_15914,N_13310,N_12647);
nor U15915 (N_15915,N_13051,N_13142);
and U15916 (N_15916,N_13881,N_13188);
nor U15917 (N_15917,N_13221,N_13042);
nand U15918 (N_15918,N_13796,N_12560);
xor U15919 (N_15919,N_14368,N_13765);
nor U15920 (N_15920,N_14371,N_13982);
xnor U15921 (N_15921,N_14590,N_14353);
nor U15922 (N_15922,N_13251,N_14480);
xor U15923 (N_15923,N_13254,N_14049);
and U15924 (N_15924,N_14837,N_14574);
nor U15925 (N_15925,N_13759,N_12877);
nor U15926 (N_15926,N_12980,N_13487);
nor U15927 (N_15927,N_13599,N_13563);
xor U15928 (N_15928,N_13538,N_12701);
xor U15929 (N_15929,N_14751,N_12953);
and U15930 (N_15930,N_12916,N_14240);
or U15931 (N_15931,N_14163,N_13750);
and U15932 (N_15932,N_14346,N_12835);
xor U15933 (N_15933,N_14894,N_14189);
or U15934 (N_15934,N_14337,N_12825);
or U15935 (N_15935,N_13212,N_13573);
or U15936 (N_15936,N_13078,N_14260);
and U15937 (N_15937,N_14514,N_12871);
xor U15938 (N_15938,N_13058,N_13848);
or U15939 (N_15939,N_13425,N_14384);
nor U15940 (N_15940,N_13318,N_12898);
xnor U15941 (N_15941,N_13232,N_13694);
xnor U15942 (N_15942,N_14618,N_14139);
nor U15943 (N_15943,N_12783,N_12536);
or U15944 (N_15944,N_13022,N_14822);
xnor U15945 (N_15945,N_12718,N_13963);
and U15946 (N_15946,N_14643,N_13299);
or U15947 (N_15947,N_14103,N_13265);
nor U15948 (N_15948,N_14636,N_12782);
nor U15949 (N_15949,N_14128,N_12674);
nor U15950 (N_15950,N_13165,N_14671);
or U15951 (N_15951,N_14256,N_12563);
or U15952 (N_15952,N_14471,N_14526);
and U15953 (N_15953,N_14009,N_14293);
or U15954 (N_15954,N_14460,N_14314);
or U15955 (N_15955,N_14301,N_14714);
xnor U15956 (N_15956,N_14972,N_14525);
or U15957 (N_15957,N_12567,N_14393);
and U15958 (N_15958,N_13245,N_14269);
or U15959 (N_15959,N_12776,N_13620);
or U15960 (N_15960,N_13648,N_14211);
nor U15961 (N_15961,N_13582,N_12716);
or U15962 (N_15962,N_13109,N_13910);
xnor U15963 (N_15963,N_14448,N_12868);
and U15964 (N_15964,N_13521,N_12996);
and U15965 (N_15965,N_13391,N_13539);
nor U15966 (N_15966,N_13919,N_14855);
and U15967 (N_15967,N_14070,N_12504);
xor U15968 (N_15968,N_14345,N_14180);
and U15969 (N_15969,N_12598,N_14524);
xnor U15970 (N_15970,N_14869,N_13295);
nand U15971 (N_15971,N_13755,N_12804);
nand U15972 (N_15972,N_13633,N_13119);
and U15973 (N_15973,N_13285,N_14334);
nand U15974 (N_15974,N_13027,N_14414);
or U15975 (N_15975,N_12978,N_13922);
nor U15976 (N_15976,N_13289,N_12802);
xor U15977 (N_15977,N_13825,N_12568);
or U15978 (N_15978,N_12766,N_12652);
nand U15979 (N_15979,N_14330,N_14830);
xor U15980 (N_15980,N_12899,N_13584);
nand U15981 (N_15981,N_13233,N_14506);
or U15982 (N_15982,N_14793,N_14280);
and U15983 (N_15983,N_14695,N_14188);
xnor U15984 (N_15984,N_14400,N_12971);
or U15985 (N_15985,N_13909,N_13862);
xnor U15986 (N_15986,N_12520,N_12907);
or U15987 (N_15987,N_14586,N_14146);
nor U15988 (N_15988,N_14582,N_14637);
xnor U15989 (N_15989,N_14872,N_14121);
and U15990 (N_15990,N_14895,N_13898);
xor U15991 (N_15991,N_12918,N_14984);
or U15992 (N_15992,N_14102,N_14728);
and U15993 (N_15993,N_13184,N_14664);
and U15994 (N_15994,N_12973,N_12790);
nor U15995 (N_15995,N_14944,N_13693);
nand U15996 (N_15996,N_13793,N_13228);
nand U15997 (N_15997,N_14766,N_13287);
xor U15998 (N_15998,N_12992,N_14378);
and U15999 (N_15999,N_13167,N_13644);
and U16000 (N_16000,N_13552,N_14178);
nor U16001 (N_16001,N_13789,N_13149);
nand U16002 (N_16002,N_13064,N_13373);
or U16003 (N_16003,N_14030,N_12569);
nand U16004 (N_16004,N_14555,N_13009);
xnor U16005 (N_16005,N_14297,N_12821);
and U16006 (N_16006,N_14087,N_12733);
nand U16007 (N_16007,N_12677,N_14356);
and U16008 (N_16008,N_12650,N_14251);
xnor U16009 (N_16009,N_14694,N_13831);
nor U16010 (N_16010,N_13348,N_14292);
and U16011 (N_16011,N_12562,N_13080);
nand U16012 (N_16012,N_12719,N_13807);
xnor U16013 (N_16013,N_13249,N_12836);
xnor U16014 (N_16014,N_14744,N_13041);
nand U16015 (N_16015,N_12533,N_13211);
nor U16016 (N_16016,N_13572,N_13797);
nand U16017 (N_16017,N_12917,N_12555);
nor U16018 (N_16018,N_13783,N_13712);
and U16019 (N_16019,N_13756,N_12863);
nor U16020 (N_16020,N_13205,N_14495);
nor U16021 (N_16021,N_13733,N_13004);
xor U16022 (N_16022,N_13615,N_12879);
nor U16023 (N_16023,N_13309,N_13450);
or U16024 (N_16024,N_14521,N_14721);
nand U16025 (N_16025,N_13728,N_13936);
xor U16026 (N_16026,N_14627,N_13722);
nor U16027 (N_16027,N_12897,N_13885);
xor U16028 (N_16028,N_14249,N_13571);
xnor U16029 (N_16029,N_13497,N_13195);
and U16030 (N_16030,N_12960,N_13129);
nor U16031 (N_16031,N_12745,N_13873);
nor U16032 (N_16032,N_12961,N_14050);
nor U16033 (N_16033,N_14031,N_13151);
and U16034 (N_16034,N_14602,N_14550);
xor U16035 (N_16035,N_12614,N_13457);
or U16036 (N_16036,N_13016,N_13387);
xor U16037 (N_16037,N_14476,N_14296);
or U16038 (N_16038,N_12542,N_14218);
nor U16039 (N_16039,N_12800,N_13060);
or U16040 (N_16040,N_13983,N_13030);
or U16041 (N_16041,N_13655,N_13947);
nor U16042 (N_16042,N_13934,N_14206);
nor U16043 (N_16043,N_13775,N_12846);
nand U16044 (N_16044,N_12710,N_12810);
or U16045 (N_16045,N_12547,N_13509);
xor U16046 (N_16046,N_13017,N_14556);
and U16047 (N_16047,N_13828,N_14638);
xnor U16048 (N_16048,N_13145,N_12818);
or U16049 (N_16049,N_13618,N_12538);
xnor U16050 (N_16050,N_13231,N_14652);
or U16051 (N_16051,N_14986,N_14265);
and U16052 (N_16052,N_13817,N_14950);
and U16053 (N_16053,N_14416,N_13263);
xnor U16054 (N_16054,N_13223,N_13394);
and U16055 (N_16055,N_13672,N_14381);
and U16056 (N_16056,N_13039,N_12896);
nor U16057 (N_16057,N_14215,N_14930);
nor U16058 (N_16058,N_14383,N_13426);
nor U16059 (N_16059,N_13013,N_14998);
or U16060 (N_16060,N_13430,N_13676);
or U16061 (N_16061,N_14123,N_14562);
xor U16062 (N_16062,N_13355,N_13378);
or U16063 (N_16063,N_14712,N_14124);
xor U16064 (N_16064,N_13010,N_12772);
or U16065 (N_16065,N_12955,N_12704);
and U16066 (N_16066,N_14656,N_13482);
or U16067 (N_16067,N_14814,N_12964);
nor U16068 (N_16068,N_14254,N_14261);
nand U16069 (N_16069,N_14370,N_13161);
or U16070 (N_16070,N_13879,N_12744);
nor U16071 (N_16071,N_14429,N_13794);
nor U16072 (N_16072,N_14004,N_13558);
and U16073 (N_16073,N_12742,N_13727);
or U16074 (N_16074,N_14316,N_13900);
nand U16075 (N_16075,N_14655,N_12811);
and U16076 (N_16076,N_13176,N_14137);
xor U16077 (N_16077,N_13566,N_14958);
or U16078 (N_16078,N_13061,N_12819);
xnor U16079 (N_16079,N_12659,N_12610);
and U16080 (N_16080,N_12521,N_13720);
or U16081 (N_16081,N_14259,N_13408);
xor U16082 (N_16082,N_13204,N_14719);
nand U16083 (N_16083,N_13040,N_13322);
nand U16084 (N_16084,N_13781,N_12834);
and U16085 (N_16085,N_13639,N_14522);
or U16086 (N_16086,N_14203,N_12586);
or U16087 (N_16087,N_13032,N_14725);
nor U16088 (N_16088,N_13556,N_14996);
and U16089 (N_16089,N_12682,N_14761);
nor U16090 (N_16090,N_13352,N_13162);
nor U16091 (N_16091,N_13754,N_14478);
xor U16092 (N_16092,N_13798,N_13561);
xor U16093 (N_16093,N_13379,N_14780);
xor U16094 (N_16094,N_14956,N_13054);
nand U16095 (N_16095,N_14239,N_12517);
and U16096 (N_16096,N_14983,N_13668);
nor U16097 (N_16097,N_13163,N_14152);
xor U16098 (N_16098,N_12823,N_14026);
and U16099 (N_16099,N_12697,N_12680);
nand U16100 (N_16100,N_13689,N_14593);
or U16101 (N_16101,N_14678,N_13477);
xor U16102 (N_16102,N_13034,N_13274);
or U16103 (N_16103,N_13747,N_13459);
and U16104 (N_16104,N_13738,N_13093);
xnor U16105 (N_16105,N_13133,N_13480);
and U16106 (N_16106,N_12942,N_13101);
or U16107 (N_16107,N_12965,N_14355);
nand U16108 (N_16108,N_12635,N_13189);
xnor U16109 (N_16109,N_14253,N_14504);
nor U16110 (N_16110,N_13890,N_12760);
and U16111 (N_16111,N_13708,N_12923);
nor U16112 (N_16112,N_12581,N_13987);
nor U16113 (N_16113,N_14048,N_13940);
nand U16114 (N_16114,N_13745,N_12950);
and U16115 (N_16115,N_13359,N_13367);
or U16116 (N_16116,N_12870,N_14387);
nand U16117 (N_16117,N_14892,N_14873);
nor U16118 (N_16118,N_14398,N_14989);
nand U16119 (N_16119,N_13962,N_12587);
xor U16120 (N_16120,N_12670,N_14100);
and U16121 (N_16121,N_13427,N_12924);
or U16122 (N_16122,N_14502,N_14395);
nand U16123 (N_16123,N_13866,N_13125);
nor U16124 (N_16124,N_13842,N_14852);
nor U16125 (N_16125,N_13896,N_13654);
or U16126 (N_16126,N_13958,N_13370);
and U16127 (N_16127,N_14092,N_13435);
and U16128 (N_16128,N_13451,N_12852);
xnor U16129 (N_16129,N_14738,N_14327);
nor U16130 (N_16130,N_14775,N_14477);
and U16131 (N_16131,N_12730,N_14571);
xor U16132 (N_16132,N_14707,N_14182);
xor U16133 (N_16133,N_12890,N_13168);
nand U16134 (N_16134,N_13510,N_14931);
xor U16135 (N_16135,N_13637,N_12816);
and U16136 (N_16136,N_14465,N_12599);
and U16137 (N_16137,N_13554,N_13525);
xor U16138 (N_16138,N_13564,N_14601);
xnor U16139 (N_16139,N_13443,N_13674);
xnor U16140 (N_16140,N_12549,N_13419);
and U16141 (N_16141,N_13114,N_12856);
or U16142 (N_16142,N_12717,N_13562);
and U16143 (N_16143,N_13839,N_12643);
or U16144 (N_16144,N_14934,N_14882);
nand U16145 (N_16145,N_14076,N_13687);
and U16146 (N_16146,N_13653,N_12720);
and U16147 (N_16147,N_14479,N_14718);
nand U16148 (N_16148,N_12948,N_13991);
and U16149 (N_16149,N_14660,N_13978);
nor U16150 (N_16150,N_14880,N_13975);
nand U16151 (N_16151,N_14202,N_13856);
nor U16152 (N_16152,N_13237,N_14073);
xnor U16153 (N_16153,N_13567,N_14492);
or U16154 (N_16154,N_13799,N_13015);
and U16155 (N_16155,N_14012,N_14589);
xnor U16156 (N_16156,N_12875,N_12850);
xor U16157 (N_16157,N_14771,N_13198);
xor U16158 (N_16158,N_12546,N_14683);
and U16159 (N_16159,N_14317,N_14132);
nor U16160 (N_16160,N_14130,N_13949);
nor U16161 (N_16161,N_14629,N_13436);
and U16162 (N_16162,N_13201,N_12940);
nor U16163 (N_16163,N_14024,N_12951);
nand U16164 (N_16164,N_13132,N_14595);
nand U16165 (N_16165,N_12557,N_12698);
xnor U16166 (N_16166,N_14016,N_13147);
or U16167 (N_16167,N_12723,N_13074);
nand U16168 (N_16168,N_14997,N_14817);
xor U16169 (N_16169,N_14794,N_12784);
nor U16170 (N_16170,N_13028,N_14015);
nand U16171 (N_16171,N_14323,N_13517);
xnor U16172 (N_16172,N_14417,N_13332);
xor U16173 (N_16173,N_13683,N_12739);
and U16174 (N_16174,N_12532,N_13062);
xor U16175 (N_16175,N_14689,N_14273);
nor U16176 (N_16176,N_14136,N_14402);
xnor U16177 (N_16177,N_13488,N_14540);
nand U16178 (N_16178,N_13277,N_14094);
or U16179 (N_16179,N_13235,N_13325);
xor U16180 (N_16180,N_14272,N_12706);
xor U16181 (N_16181,N_14802,N_14551);
xnor U16182 (N_16182,N_13441,N_14122);
nor U16183 (N_16183,N_13959,N_14588);
and U16184 (N_16184,N_13374,N_13642);
or U16185 (N_16185,N_13411,N_14008);
nand U16186 (N_16186,N_13585,N_12593);
xnor U16187 (N_16187,N_14529,N_14961);
nand U16188 (N_16188,N_14485,N_13312);
or U16189 (N_16189,N_14091,N_14141);
or U16190 (N_16190,N_13993,N_14040);
or U16191 (N_16191,N_13113,N_12734);
and U16192 (N_16192,N_12912,N_14359);
and U16193 (N_16193,N_14642,N_14515);
xnor U16194 (N_16194,N_12860,N_14633);
nand U16195 (N_16195,N_14399,N_13236);
xor U16196 (N_16196,N_14161,N_14607);
and U16197 (N_16197,N_12683,N_13065);
xor U16198 (N_16198,N_14434,N_13177);
xor U16199 (N_16199,N_14407,N_12578);
and U16200 (N_16200,N_14411,N_13366);
or U16201 (N_16201,N_14080,N_13614);
nor U16202 (N_16202,N_12605,N_14839);
nand U16203 (N_16203,N_12865,N_13075);
xnor U16204 (N_16204,N_13072,N_13601);
or U16205 (N_16205,N_14194,N_14201);
and U16206 (N_16206,N_13758,N_14646);
and U16207 (N_16207,N_14739,N_12509);
and U16208 (N_16208,N_14335,N_12666);
nor U16209 (N_16209,N_13595,N_14482);
xnor U16210 (N_16210,N_13389,N_14973);
or U16211 (N_16211,N_14701,N_14170);
or U16212 (N_16212,N_13726,N_14835);
nand U16213 (N_16213,N_13935,N_12855);
nor U16214 (N_16214,N_13774,N_12703);
or U16215 (N_16215,N_14568,N_12644);
or U16216 (N_16216,N_14995,N_13337);
and U16217 (N_16217,N_14055,N_14078);
or U16218 (N_16218,N_12741,N_13094);
or U16219 (N_16219,N_13472,N_14941);
xor U16220 (N_16220,N_12522,N_14241);
nor U16221 (N_16221,N_12934,N_14704);
nor U16222 (N_16222,N_12839,N_12858);
xnor U16223 (N_16223,N_14344,N_13050);
nor U16224 (N_16224,N_13782,N_14697);
nor U16225 (N_16225,N_13261,N_12607);
nor U16226 (N_16226,N_14209,N_14037);
nor U16227 (N_16227,N_12514,N_13294);
or U16228 (N_16228,N_14284,N_13070);
xnor U16229 (N_16229,N_13127,N_13174);
nand U16230 (N_16230,N_12535,N_13735);
or U16231 (N_16231,N_14631,N_13121);
nor U16232 (N_16232,N_12881,N_12594);
xnor U16233 (N_16233,N_14600,N_14295);
and U16234 (N_16234,N_13314,N_12985);
nor U16235 (N_16235,N_14018,N_14126);
nor U16236 (N_16236,N_12515,N_14945);
and U16237 (N_16237,N_14518,N_14183);
or U16238 (N_16238,N_14968,N_13160);
nand U16239 (N_16239,N_12738,N_13243);
and U16240 (N_16240,N_14172,N_12656);
xnor U16241 (N_16241,N_12505,N_13843);
nand U16242 (N_16242,N_13386,N_13823);
and U16243 (N_16243,N_13059,N_13874);
nor U16244 (N_16244,N_13943,N_14726);
nor U16245 (N_16245,N_14135,N_12884);
xnor U16246 (N_16246,N_14649,N_12986);
nor U16247 (N_16247,N_13356,N_14569);
or U16248 (N_16248,N_13264,N_13706);
nand U16249 (N_16249,N_14199,N_14603);
xor U16250 (N_16250,N_14311,N_13731);
or U16251 (N_16251,N_12835,N_13316);
nand U16252 (N_16252,N_13050,N_13875);
or U16253 (N_16253,N_14214,N_13347);
xor U16254 (N_16254,N_14575,N_13904);
xnor U16255 (N_16255,N_12862,N_13631);
and U16256 (N_16256,N_13343,N_13922);
nand U16257 (N_16257,N_14814,N_13601);
nand U16258 (N_16258,N_14536,N_13528);
or U16259 (N_16259,N_12973,N_14861);
nor U16260 (N_16260,N_13187,N_14854);
nand U16261 (N_16261,N_14250,N_14343);
or U16262 (N_16262,N_12884,N_13838);
or U16263 (N_16263,N_12940,N_14298);
nand U16264 (N_16264,N_14271,N_12581);
nor U16265 (N_16265,N_12972,N_13218);
nor U16266 (N_16266,N_13485,N_14117);
or U16267 (N_16267,N_14336,N_13984);
or U16268 (N_16268,N_13963,N_13094);
and U16269 (N_16269,N_12980,N_13502);
nand U16270 (N_16270,N_14397,N_12539);
and U16271 (N_16271,N_13105,N_13524);
or U16272 (N_16272,N_14323,N_12972);
nand U16273 (N_16273,N_13780,N_12852);
xor U16274 (N_16274,N_12619,N_13447);
and U16275 (N_16275,N_14049,N_13457);
and U16276 (N_16276,N_13479,N_12970);
xor U16277 (N_16277,N_13135,N_13646);
xnor U16278 (N_16278,N_13000,N_12579);
or U16279 (N_16279,N_12856,N_13722);
or U16280 (N_16280,N_13921,N_14644);
nand U16281 (N_16281,N_12899,N_12985);
xnor U16282 (N_16282,N_14787,N_13988);
nor U16283 (N_16283,N_13951,N_14409);
xor U16284 (N_16284,N_12794,N_13895);
xor U16285 (N_16285,N_12824,N_13994);
or U16286 (N_16286,N_13813,N_12543);
xor U16287 (N_16287,N_13054,N_14138);
nor U16288 (N_16288,N_13164,N_14690);
xor U16289 (N_16289,N_13458,N_13895);
nand U16290 (N_16290,N_13650,N_14306);
xnor U16291 (N_16291,N_14573,N_13479);
nor U16292 (N_16292,N_14601,N_12825);
and U16293 (N_16293,N_13654,N_14421);
xor U16294 (N_16294,N_14286,N_13567);
and U16295 (N_16295,N_13864,N_13057);
nor U16296 (N_16296,N_13587,N_13833);
or U16297 (N_16297,N_14512,N_13521);
xnor U16298 (N_16298,N_14369,N_13775);
nand U16299 (N_16299,N_13558,N_13306);
nor U16300 (N_16300,N_14084,N_14064);
or U16301 (N_16301,N_13982,N_14378);
and U16302 (N_16302,N_14815,N_12583);
nand U16303 (N_16303,N_13633,N_12627);
nand U16304 (N_16304,N_12772,N_12698);
nand U16305 (N_16305,N_14192,N_14761);
and U16306 (N_16306,N_14082,N_13167);
nor U16307 (N_16307,N_14258,N_13222);
xnor U16308 (N_16308,N_13440,N_13290);
nand U16309 (N_16309,N_14535,N_12869);
xor U16310 (N_16310,N_14176,N_14552);
nand U16311 (N_16311,N_12763,N_12518);
nor U16312 (N_16312,N_13854,N_12577);
xnor U16313 (N_16313,N_13872,N_13570);
or U16314 (N_16314,N_13585,N_12857);
xor U16315 (N_16315,N_12941,N_13148);
xnor U16316 (N_16316,N_14716,N_14132);
xor U16317 (N_16317,N_14485,N_14868);
nor U16318 (N_16318,N_13398,N_14261);
and U16319 (N_16319,N_14934,N_13008);
nand U16320 (N_16320,N_12870,N_13813);
or U16321 (N_16321,N_14775,N_14523);
xor U16322 (N_16322,N_13841,N_13139);
nand U16323 (N_16323,N_13472,N_14907);
or U16324 (N_16324,N_12824,N_14613);
or U16325 (N_16325,N_14598,N_14124);
nand U16326 (N_16326,N_14047,N_13643);
nor U16327 (N_16327,N_14157,N_12736);
xor U16328 (N_16328,N_14552,N_14674);
nand U16329 (N_16329,N_13207,N_13190);
nor U16330 (N_16330,N_13930,N_13112);
or U16331 (N_16331,N_13984,N_13625);
or U16332 (N_16332,N_14369,N_14556);
nand U16333 (N_16333,N_14993,N_13694);
or U16334 (N_16334,N_12519,N_12751);
nand U16335 (N_16335,N_14933,N_13931);
nand U16336 (N_16336,N_13462,N_13639);
and U16337 (N_16337,N_13164,N_13509);
nor U16338 (N_16338,N_13596,N_14753);
and U16339 (N_16339,N_14476,N_14236);
nand U16340 (N_16340,N_13150,N_13570);
or U16341 (N_16341,N_13180,N_12871);
xnor U16342 (N_16342,N_13483,N_14610);
nand U16343 (N_16343,N_12811,N_12557);
nor U16344 (N_16344,N_14329,N_13325);
and U16345 (N_16345,N_13124,N_13221);
nand U16346 (N_16346,N_13957,N_14942);
xor U16347 (N_16347,N_14409,N_14454);
nand U16348 (N_16348,N_14249,N_13370);
or U16349 (N_16349,N_13444,N_12578);
nand U16350 (N_16350,N_14553,N_14595);
xor U16351 (N_16351,N_14704,N_13503);
or U16352 (N_16352,N_12517,N_13173);
or U16353 (N_16353,N_13103,N_12869);
nor U16354 (N_16354,N_13653,N_13534);
or U16355 (N_16355,N_14203,N_13264);
and U16356 (N_16356,N_14059,N_13108);
and U16357 (N_16357,N_13780,N_13395);
and U16358 (N_16358,N_14571,N_13383);
or U16359 (N_16359,N_14466,N_13717);
nor U16360 (N_16360,N_14286,N_13178);
or U16361 (N_16361,N_14497,N_13103);
or U16362 (N_16362,N_14969,N_13429);
and U16363 (N_16363,N_13443,N_14804);
nor U16364 (N_16364,N_13346,N_13408);
or U16365 (N_16365,N_12763,N_13814);
and U16366 (N_16366,N_14399,N_12748);
or U16367 (N_16367,N_14829,N_12706);
xor U16368 (N_16368,N_14056,N_13132);
nor U16369 (N_16369,N_14624,N_14386);
and U16370 (N_16370,N_13274,N_14752);
nand U16371 (N_16371,N_12920,N_12523);
nor U16372 (N_16372,N_12607,N_14440);
nor U16373 (N_16373,N_13688,N_12663);
nor U16374 (N_16374,N_13429,N_13053);
and U16375 (N_16375,N_14044,N_13887);
nand U16376 (N_16376,N_14680,N_13413);
and U16377 (N_16377,N_14478,N_12999);
and U16378 (N_16378,N_14347,N_14304);
nor U16379 (N_16379,N_13209,N_14641);
xor U16380 (N_16380,N_13213,N_13431);
or U16381 (N_16381,N_12508,N_14573);
nor U16382 (N_16382,N_13553,N_13069);
nor U16383 (N_16383,N_13641,N_14954);
nand U16384 (N_16384,N_14150,N_13095);
nor U16385 (N_16385,N_12612,N_14985);
xor U16386 (N_16386,N_13003,N_14549);
nand U16387 (N_16387,N_13666,N_13070);
nand U16388 (N_16388,N_13095,N_13411);
nor U16389 (N_16389,N_13277,N_14873);
xor U16390 (N_16390,N_12523,N_13476);
nand U16391 (N_16391,N_12634,N_13707);
nor U16392 (N_16392,N_12631,N_14954);
or U16393 (N_16393,N_13117,N_13046);
and U16394 (N_16394,N_13689,N_12532);
xor U16395 (N_16395,N_13994,N_14249);
xnor U16396 (N_16396,N_13088,N_14613);
nand U16397 (N_16397,N_12863,N_12637);
nand U16398 (N_16398,N_12579,N_12636);
nand U16399 (N_16399,N_12527,N_12969);
xor U16400 (N_16400,N_14114,N_12536);
and U16401 (N_16401,N_14712,N_14661);
or U16402 (N_16402,N_14090,N_13127);
or U16403 (N_16403,N_13564,N_13916);
xnor U16404 (N_16404,N_13892,N_13176);
and U16405 (N_16405,N_12783,N_13485);
nand U16406 (N_16406,N_13696,N_13227);
nor U16407 (N_16407,N_12903,N_12786);
nand U16408 (N_16408,N_13143,N_13350);
nor U16409 (N_16409,N_12594,N_13176);
nand U16410 (N_16410,N_13067,N_12640);
or U16411 (N_16411,N_12682,N_13879);
xnor U16412 (N_16412,N_14949,N_13147);
xnor U16413 (N_16413,N_14194,N_12888);
and U16414 (N_16414,N_13645,N_13812);
nor U16415 (N_16415,N_14717,N_13371);
or U16416 (N_16416,N_13749,N_13805);
nand U16417 (N_16417,N_13883,N_14560);
nand U16418 (N_16418,N_13539,N_13497);
xnor U16419 (N_16419,N_12718,N_14654);
and U16420 (N_16420,N_12835,N_13847);
and U16421 (N_16421,N_14136,N_14828);
nor U16422 (N_16422,N_14723,N_12518);
nor U16423 (N_16423,N_13396,N_12794);
or U16424 (N_16424,N_13540,N_13159);
xor U16425 (N_16425,N_14952,N_13982);
nand U16426 (N_16426,N_12971,N_13128);
xor U16427 (N_16427,N_14306,N_12921);
xnor U16428 (N_16428,N_13654,N_14459);
or U16429 (N_16429,N_12718,N_13187);
and U16430 (N_16430,N_14320,N_12539);
or U16431 (N_16431,N_12820,N_14568);
or U16432 (N_16432,N_14764,N_14603);
nand U16433 (N_16433,N_13846,N_14465);
nor U16434 (N_16434,N_14938,N_13395);
xnor U16435 (N_16435,N_14912,N_14567);
xor U16436 (N_16436,N_12957,N_13072);
and U16437 (N_16437,N_13964,N_14339);
or U16438 (N_16438,N_13291,N_14998);
xnor U16439 (N_16439,N_14161,N_14705);
xor U16440 (N_16440,N_13116,N_13306);
nand U16441 (N_16441,N_13240,N_13393);
nand U16442 (N_16442,N_13402,N_14693);
and U16443 (N_16443,N_14887,N_12657);
or U16444 (N_16444,N_14243,N_12601);
xnor U16445 (N_16445,N_14173,N_13097);
xor U16446 (N_16446,N_13015,N_12938);
or U16447 (N_16447,N_14759,N_13030);
xnor U16448 (N_16448,N_14070,N_13539);
or U16449 (N_16449,N_13259,N_14537);
nor U16450 (N_16450,N_13352,N_14672);
or U16451 (N_16451,N_13714,N_14080);
or U16452 (N_16452,N_14822,N_13528);
xnor U16453 (N_16453,N_13569,N_12940);
nor U16454 (N_16454,N_12610,N_12666);
xnor U16455 (N_16455,N_14693,N_13897);
nand U16456 (N_16456,N_13189,N_13987);
nand U16457 (N_16457,N_14754,N_13939);
nand U16458 (N_16458,N_12703,N_13621);
and U16459 (N_16459,N_14473,N_14005);
xor U16460 (N_16460,N_14612,N_13893);
nand U16461 (N_16461,N_13907,N_14103);
xor U16462 (N_16462,N_12991,N_14116);
xnor U16463 (N_16463,N_12961,N_12824);
xnor U16464 (N_16464,N_14093,N_14424);
nand U16465 (N_16465,N_13405,N_13076);
nor U16466 (N_16466,N_12955,N_13786);
nand U16467 (N_16467,N_12712,N_14695);
xor U16468 (N_16468,N_14005,N_13304);
nor U16469 (N_16469,N_14630,N_14438);
or U16470 (N_16470,N_14956,N_14197);
nand U16471 (N_16471,N_14794,N_14680);
and U16472 (N_16472,N_13172,N_14643);
nand U16473 (N_16473,N_13414,N_13476);
nor U16474 (N_16474,N_14876,N_12555);
nor U16475 (N_16475,N_14271,N_13198);
and U16476 (N_16476,N_13910,N_12858);
or U16477 (N_16477,N_12953,N_13600);
nand U16478 (N_16478,N_13252,N_14306);
or U16479 (N_16479,N_13533,N_14468);
and U16480 (N_16480,N_12813,N_13552);
and U16481 (N_16481,N_13632,N_14668);
and U16482 (N_16482,N_14209,N_13486);
or U16483 (N_16483,N_14606,N_13927);
nor U16484 (N_16484,N_14392,N_12644);
nor U16485 (N_16485,N_14152,N_14734);
xnor U16486 (N_16486,N_13071,N_13366);
xnor U16487 (N_16487,N_13667,N_14950);
nand U16488 (N_16488,N_13738,N_14355);
and U16489 (N_16489,N_14898,N_13171);
nand U16490 (N_16490,N_12941,N_13360);
xnor U16491 (N_16491,N_14155,N_14491);
and U16492 (N_16492,N_14289,N_13533);
xnor U16493 (N_16493,N_13062,N_14623);
nor U16494 (N_16494,N_12987,N_12732);
xor U16495 (N_16495,N_14886,N_14547);
nand U16496 (N_16496,N_14099,N_13557);
or U16497 (N_16497,N_14399,N_14400);
xor U16498 (N_16498,N_12781,N_14928);
nand U16499 (N_16499,N_13367,N_14245);
and U16500 (N_16500,N_13266,N_12719);
or U16501 (N_16501,N_13225,N_12900);
and U16502 (N_16502,N_12593,N_14706);
xnor U16503 (N_16503,N_13398,N_12697);
or U16504 (N_16504,N_14883,N_13513);
and U16505 (N_16505,N_12547,N_13728);
and U16506 (N_16506,N_12949,N_14696);
or U16507 (N_16507,N_14258,N_14572);
nor U16508 (N_16508,N_13923,N_14746);
and U16509 (N_16509,N_14093,N_12548);
or U16510 (N_16510,N_13740,N_13315);
nand U16511 (N_16511,N_14309,N_13084);
nand U16512 (N_16512,N_13592,N_13142);
nor U16513 (N_16513,N_14430,N_12591);
nor U16514 (N_16514,N_14124,N_12811);
nand U16515 (N_16515,N_12659,N_14911);
nand U16516 (N_16516,N_14810,N_12850);
and U16517 (N_16517,N_12798,N_14381);
or U16518 (N_16518,N_12823,N_12610);
xnor U16519 (N_16519,N_13023,N_14565);
nand U16520 (N_16520,N_14509,N_12706);
xor U16521 (N_16521,N_13131,N_13281);
xor U16522 (N_16522,N_13912,N_14909);
and U16523 (N_16523,N_14931,N_12560);
or U16524 (N_16524,N_14783,N_14347);
nor U16525 (N_16525,N_14205,N_13554);
nor U16526 (N_16526,N_13750,N_13836);
nand U16527 (N_16527,N_13719,N_14588);
xnor U16528 (N_16528,N_14434,N_12649);
or U16529 (N_16529,N_13192,N_13464);
nor U16530 (N_16530,N_14877,N_13333);
or U16531 (N_16531,N_13826,N_12922);
nand U16532 (N_16532,N_14432,N_14621);
xnor U16533 (N_16533,N_13576,N_13120);
nand U16534 (N_16534,N_14341,N_13132);
or U16535 (N_16535,N_14119,N_13431);
nand U16536 (N_16536,N_13249,N_14276);
nand U16537 (N_16537,N_12735,N_12819);
and U16538 (N_16538,N_13331,N_13304);
nor U16539 (N_16539,N_14729,N_14482);
and U16540 (N_16540,N_12565,N_14804);
and U16541 (N_16541,N_12995,N_13204);
xor U16542 (N_16542,N_13525,N_14467);
nand U16543 (N_16543,N_13276,N_14182);
nor U16544 (N_16544,N_13009,N_14560);
and U16545 (N_16545,N_13314,N_14944);
xor U16546 (N_16546,N_14519,N_12707);
xnor U16547 (N_16547,N_13163,N_13958);
nor U16548 (N_16548,N_14313,N_13531);
nand U16549 (N_16549,N_14551,N_13042);
and U16550 (N_16550,N_14366,N_13232);
nand U16551 (N_16551,N_13655,N_14545);
nor U16552 (N_16552,N_14033,N_13074);
nand U16553 (N_16553,N_13736,N_12815);
nand U16554 (N_16554,N_13425,N_13026);
and U16555 (N_16555,N_12727,N_14450);
nand U16556 (N_16556,N_13538,N_12651);
xor U16557 (N_16557,N_14009,N_13225);
or U16558 (N_16558,N_14283,N_13167);
or U16559 (N_16559,N_14332,N_14008);
and U16560 (N_16560,N_13872,N_13443);
and U16561 (N_16561,N_14863,N_14846);
and U16562 (N_16562,N_13074,N_14048);
or U16563 (N_16563,N_14681,N_13265);
and U16564 (N_16564,N_13918,N_13500);
and U16565 (N_16565,N_13888,N_14219);
nand U16566 (N_16566,N_13205,N_14479);
xnor U16567 (N_16567,N_12964,N_14792);
or U16568 (N_16568,N_12905,N_13636);
xor U16569 (N_16569,N_13106,N_13172);
nor U16570 (N_16570,N_14934,N_14677);
and U16571 (N_16571,N_14330,N_13815);
or U16572 (N_16572,N_14984,N_12605);
or U16573 (N_16573,N_12947,N_13352);
xor U16574 (N_16574,N_13356,N_14046);
nor U16575 (N_16575,N_14752,N_13079);
xnor U16576 (N_16576,N_12676,N_14995);
nand U16577 (N_16577,N_14270,N_13539);
or U16578 (N_16578,N_13786,N_13057);
xor U16579 (N_16579,N_13242,N_13263);
nand U16580 (N_16580,N_14338,N_14697);
nand U16581 (N_16581,N_14404,N_14891);
xor U16582 (N_16582,N_14086,N_14631);
xor U16583 (N_16583,N_14320,N_13435);
xor U16584 (N_16584,N_14428,N_12849);
nor U16585 (N_16585,N_14351,N_12973);
nand U16586 (N_16586,N_14756,N_14474);
xor U16587 (N_16587,N_13796,N_14833);
or U16588 (N_16588,N_13367,N_13360);
and U16589 (N_16589,N_14920,N_12666);
or U16590 (N_16590,N_14628,N_14014);
and U16591 (N_16591,N_12715,N_14361);
nor U16592 (N_16592,N_12981,N_14186);
and U16593 (N_16593,N_14096,N_13646);
nand U16594 (N_16594,N_13712,N_12626);
nand U16595 (N_16595,N_14046,N_13827);
nand U16596 (N_16596,N_13872,N_12582);
and U16597 (N_16597,N_12739,N_13737);
nand U16598 (N_16598,N_12779,N_12800);
nor U16599 (N_16599,N_14309,N_12844);
or U16600 (N_16600,N_13868,N_14228);
nor U16601 (N_16601,N_13916,N_13368);
nand U16602 (N_16602,N_14325,N_13533);
and U16603 (N_16603,N_12616,N_14926);
xor U16604 (N_16604,N_14427,N_14429);
xor U16605 (N_16605,N_14215,N_14328);
nor U16606 (N_16606,N_14921,N_13072);
nor U16607 (N_16607,N_13771,N_14499);
and U16608 (N_16608,N_14994,N_12727);
nand U16609 (N_16609,N_14151,N_14284);
or U16610 (N_16610,N_14290,N_13853);
nor U16611 (N_16611,N_14751,N_12875);
and U16612 (N_16612,N_13489,N_14019);
xor U16613 (N_16613,N_13285,N_13465);
nand U16614 (N_16614,N_14996,N_14567);
or U16615 (N_16615,N_14137,N_12542);
nand U16616 (N_16616,N_14811,N_12850);
nor U16617 (N_16617,N_13329,N_14438);
or U16618 (N_16618,N_12916,N_14724);
xnor U16619 (N_16619,N_13328,N_12608);
or U16620 (N_16620,N_14254,N_13922);
and U16621 (N_16621,N_13874,N_14959);
and U16622 (N_16622,N_14204,N_12503);
nand U16623 (N_16623,N_14981,N_14794);
and U16624 (N_16624,N_14695,N_13256);
xnor U16625 (N_16625,N_14416,N_12902);
xor U16626 (N_16626,N_12934,N_14708);
and U16627 (N_16627,N_14027,N_13437);
nor U16628 (N_16628,N_13399,N_14723);
xor U16629 (N_16629,N_13364,N_14469);
and U16630 (N_16630,N_14151,N_14513);
or U16631 (N_16631,N_13623,N_13359);
or U16632 (N_16632,N_14772,N_13568);
nand U16633 (N_16633,N_13202,N_14352);
xor U16634 (N_16634,N_14184,N_12749);
and U16635 (N_16635,N_13613,N_13412);
nand U16636 (N_16636,N_12709,N_14340);
nor U16637 (N_16637,N_13706,N_12940);
or U16638 (N_16638,N_14803,N_14104);
nor U16639 (N_16639,N_14828,N_14289);
and U16640 (N_16640,N_13872,N_14507);
nand U16641 (N_16641,N_12934,N_13140);
and U16642 (N_16642,N_13015,N_12681);
xnor U16643 (N_16643,N_13438,N_13141);
or U16644 (N_16644,N_13391,N_14440);
nand U16645 (N_16645,N_13127,N_13589);
xor U16646 (N_16646,N_13433,N_13184);
nand U16647 (N_16647,N_12555,N_13535);
nor U16648 (N_16648,N_13508,N_14925);
xor U16649 (N_16649,N_14710,N_13246);
xor U16650 (N_16650,N_13057,N_12575);
nor U16651 (N_16651,N_14692,N_14305);
nor U16652 (N_16652,N_13175,N_14155);
xnor U16653 (N_16653,N_14794,N_13829);
xnor U16654 (N_16654,N_14471,N_14358);
nor U16655 (N_16655,N_14427,N_14970);
or U16656 (N_16656,N_13993,N_14683);
and U16657 (N_16657,N_13800,N_12769);
xor U16658 (N_16658,N_14684,N_14510);
nand U16659 (N_16659,N_14912,N_14615);
xnor U16660 (N_16660,N_13408,N_12870);
or U16661 (N_16661,N_14844,N_14461);
or U16662 (N_16662,N_13917,N_14602);
and U16663 (N_16663,N_13997,N_13681);
nor U16664 (N_16664,N_14462,N_14218);
nand U16665 (N_16665,N_14255,N_12916);
or U16666 (N_16666,N_12933,N_13257);
or U16667 (N_16667,N_14285,N_13484);
or U16668 (N_16668,N_14711,N_13853);
xnor U16669 (N_16669,N_13979,N_12830);
nor U16670 (N_16670,N_13287,N_13010);
nand U16671 (N_16671,N_14249,N_13308);
nor U16672 (N_16672,N_14347,N_13716);
or U16673 (N_16673,N_14814,N_12725);
nand U16674 (N_16674,N_13420,N_13827);
nor U16675 (N_16675,N_14459,N_14312);
nor U16676 (N_16676,N_13264,N_14360);
and U16677 (N_16677,N_14192,N_12812);
or U16678 (N_16678,N_12612,N_14753);
nand U16679 (N_16679,N_14041,N_13230);
nor U16680 (N_16680,N_12595,N_13533);
and U16681 (N_16681,N_14743,N_14845);
and U16682 (N_16682,N_13469,N_14026);
xnor U16683 (N_16683,N_13118,N_12825);
nor U16684 (N_16684,N_14362,N_13233);
or U16685 (N_16685,N_13178,N_13711);
nor U16686 (N_16686,N_14989,N_14484);
nor U16687 (N_16687,N_13030,N_13503);
nand U16688 (N_16688,N_14801,N_12739);
nand U16689 (N_16689,N_13508,N_13818);
nand U16690 (N_16690,N_13526,N_14796);
or U16691 (N_16691,N_13759,N_13781);
xnor U16692 (N_16692,N_13863,N_13515);
nand U16693 (N_16693,N_14420,N_12806);
nor U16694 (N_16694,N_14763,N_14675);
or U16695 (N_16695,N_13916,N_14601);
nand U16696 (N_16696,N_14561,N_14572);
nor U16697 (N_16697,N_14330,N_12990);
xnor U16698 (N_16698,N_13865,N_13214);
nand U16699 (N_16699,N_13333,N_14223);
or U16700 (N_16700,N_14506,N_13290);
or U16701 (N_16701,N_14436,N_13177);
nand U16702 (N_16702,N_13999,N_13271);
or U16703 (N_16703,N_14478,N_14997);
or U16704 (N_16704,N_13386,N_13441);
nand U16705 (N_16705,N_13743,N_13607);
xnor U16706 (N_16706,N_14698,N_14598);
xor U16707 (N_16707,N_13779,N_14275);
or U16708 (N_16708,N_14493,N_13409);
or U16709 (N_16709,N_14420,N_14613);
xnor U16710 (N_16710,N_13324,N_12558);
xor U16711 (N_16711,N_12825,N_14639);
xnor U16712 (N_16712,N_12519,N_14011);
nor U16713 (N_16713,N_13342,N_13839);
nand U16714 (N_16714,N_13865,N_13054);
or U16715 (N_16715,N_13891,N_12784);
xor U16716 (N_16716,N_14489,N_12561);
xor U16717 (N_16717,N_13762,N_13265);
nor U16718 (N_16718,N_12663,N_13714);
nor U16719 (N_16719,N_13400,N_13016);
xnor U16720 (N_16720,N_14415,N_14642);
nor U16721 (N_16721,N_14197,N_12771);
xnor U16722 (N_16722,N_13942,N_13845);
xnor U16723 (N_16723,N_14795,N_14385);
nand U16724 (N_16724,N_13778,N_13845);
and U16725 (N_16725,N_14470,N_12709);
xnor U16726 (N_16726,N_13547,N_13304);
xor U16727 (N_16727,N_13664,N_12578);
and U16728 (N_16728,N_13510,N_13103);
and U16729 (N_16729,N_14477,N_12984);
and U16730 (N_16730,N_12801,N_13590);
or U16731 (N_16731,N_13520,N_13603);
and U16732 (N_16732,N_13028,N_13301);
nand U16733 (N_16733,N_14938,N_13987);
xnor U16734 (N_16734,N_13362,N_13019);
nand U16735 (N_16735,N_13441,N_12873);
nand U16736 (N_16736,N_13964,N_13071);
nand U16737 (N_16737,N_14354,N_14415);
nor U16738 (N_16738,N_14904,N_14342);
xnor U16739 (N_16739,N_12778,N_14432);
or U16740 (N_16740,N_14793,N_14934);
or U16741 (N_16741,N_13903,N_14465);
nand U16742 (N_16742,N_13526,N_14567);
nand U16743 (N_16743,N_13590,N_14161);
xnor U16744 (N_16744,N_14426,N_13085);
and U16745 (N_16745,N_14440,N_14776);
and U16746 (N_16746,N_14931,N_14418);
and U16747 (N_16747,N_14640,N_13279);
and U16748 (N_16748,N_14918,N_14235);
nand U16749 (N_16749,N_14639,N_14075);
nand U16750 (N_16750,N_13131,N_14257);
xor U16751 (N_16751,N_14308,N_14340);
xnor U16752 (N_16752,N_12675,N_14607);
or U16753 (N_16753,N_14326,N_12793);
nand U16754 (N_16754,N_12711,N_14669);
nand U16755 (N_16755,N_12755,N_12655);
nand U16756 (N_16756,N_12543,N_14121);
and U16757 (N_16757,N_13032,N_14726);
nor U16758 (N_16758,N_14725,N_14670);
and U16759 (N_16759,N_13180,N_13178);
xnor U16760 (N_16760,N_14824,N_12823);
xor U16761 (N_16761,N_14286,N_12722);
xnor U16762 (N_16762,N_14451,N_13191);
xnor U16763 (N_16763,N_14682,N_14617);
and U16764 (N_16764,N_13344,N_14900);
xor U16765 (N_16765,N_13876,N_14390);
and U16766 (N_16766,N_13165,N_12677);
or U16767 (N_16767,N_12858,N_12547);
or U16768 (N_16768,N_14750,N_14156);
nand U16769 (N_16769,N_14392,N_13959);
nand U16770 (N_16770,N_13890,N_12613);
or U16771 (N_16771,N_13688,N_13888);
nand U16772 (N_16772,N_14249,N_14994);
nor U16773 (N_16773,N_14252,N_12552);
and U16774 (N_16774,N_14165,N_13535);
and U16775 (N_16775,N_14968,N_13210);
and U16776 (N_16776,N_13320,N_14835);
nor U16777 (N_16777,N_13356,N_12864);
and U16778 (N_16778,N_13333,N_12929);
xor U16779 (N_16779,N_12510,N_13973);
or U16780 (N_16780,N_13426,N_14451);
nand U16781 (N_16781,N_14906,N_14643);
nor U16782 (N_16782,N_13189,N_13470);
xor U16783 (N_16783,N_12759,N_13899);
and U16784 (N_16784,N_14727,N_14623);
and U16785 (N_16785,N_13821,N_13305);
xnor U16786 (N_16786,N_14362,N_14577);
xnor U16787 (N_16787,N_14267,N_14251);
xnor U16788 (N_16788,N_12682,N_12728);
nor U16789 (N_16789,N_13393,N_12898);
or U16790 (N_16790,N_14870,N_13104);
and U16791 (N_16791,N_12524,N_14324);
and U16792 (N_16792,N_14671,N_12770);
and U16793 (N_16793,N_13813,N_13422);
or U16794 (N_16794,N_14452,N_13556);
xor U16795 (N_16795,N_14362,N_13744);
and U16796 (N_16796,N_14745,N_14719);
and U16797 (N_16797,N_13027,N_13286);
or U16798 (N_16798,N_14001,N_13084);
and U16799 (N_16799,N_12741,N_14919);
or U16800 (N_16800,N_14965,N_14570);
and U16801 (N_16801,N_12946,N_14521);
nor U16802 (N_16802,N_13888,N_14595);
nor U16803 (N_16803,N_13046,N_14022);
nor U16804 (N_16804,N_14856,N_14344);
and U16805 (N_16805,N_14920,N_14349);
and U16806 (N_16806,N_14566,N_13131);
and U16807 (N_16807,N_12581,N_13280);
nor U16808 (N_16808,N_14770,N_14761);
nor U16809 (N_16809,N_14216,N_14064);
and U16810 (N_16810,N_14001,N_14148);
and U16811 (N_16811,N_12579,N_14907);
or U16812 (N_16812,N_14778,N_13622);
or U16813 (N_16813,N_13248,N_13165);
or U16814 (N_16814,N_13121,N_14087);
or U16815 (N_16815,N_12822,N_13641);
and U16816 (N_16816,N_12604,N_12963);
and U16817 (N_16817,N_13532,N_13167);
nor U16818 (N_16818,N_14107,N_14543);
nand U16819 (N_16819,N_12609,N_14221);
xnor U16820 (N_16820,N_13159,N_14205);
or U16821 (N_16821,N_14745,N_13664);
and U16822 (N_16822,N_14968,N_14550);
xnor U16823 (N_16823,N_13439,N_14490);
or U16824 (N_16824,N_14921,N_13793);
and U16825 (N_16825,N_14940,N_14583);
and U16826 (N_16826,N_13628,N_12634);
nand U16827 (N_16827,N_12596,N_13469);
or U16828 (N_16828,N_14318,N_13355);
nand U16829 (N_16829,N_13386,N_13844);
and U16830 (N_16830,N_13194,N_14676);
nand U16831 (N_16831,N_13155,N_12975);
nand U16832 (N_16832,N_13375,N_14821);
or U16833 (N_16833,N_13687,N_13311);
nor U16834 (N_16834,N_12986,N_14128);
nand U16835 (N_16835,N_13668,N_13706);
or U16836 (N_16836,N_14815,N_12658);
and U16837 (N_16837,N_12760,N_13881);
nor U16838 (N_16838,N_12824,N_13252);
xor U16839 (N_16839,N_13475,N_13166);
nand U16840 (N_16840,N_13436,N_14641);
or U16841 (N_16841,N_12996,N_14317);
xor U16842 (N_16842,N_12995,N_13707);
nand U16843 (N_16843,N_14345,N_14150);
and U16844 (N_16844,N_14087,N_14425);
nand U16845 (N_16845,N_13761,N_13080);
xor U16846 (N_16846,N_13425,N_14347);
nor U16847 (N_16847,N_13609,N_13518);
or U16848 (N_16848,N_14803,N_14901);
xor U16849 (N_16849,N_12624,N_14581);
and U16850 (N_16850,N_13132,N_12791);
nor U16851 (N_16851,N_14847,N_14365);
nor U16852 (N_16852,N_14829,N_12830);
nand U16853 (N_16853,N_14613,N_14780);
and U16854 (N_16854,N_13537,N_12668);
nand U16855 (N_16855,N_12807,N_13240);
nand U16856 (N_16856,N_13092,N_13664);
nand U16857 (N_16857,N_12673,N_14661);
or U16858 (N_16858,N_12633,N_12878);
xnor U16859 (N_16859,N_13034,N_13270);
xnor U16860 (N_16860,N_12769,N_13243);
nand U16861 (N_16861,N_14479,N_13602);
or U16862 (N_16862,N_12614,N_12920);
and U16863 (N_16863,N_13846,N_14498);
or U16864 (N_16864,N_12537,N_12650);
nand U16865 (N_16865,N_14048,N_13880);
or U16866 (N_16866,N_14665,N_14242);
nand U16867 (N_16867,N_12592,N_13704);
xor U16868 (N_16868,N_14267,N_13867);
and U16869 (N_16869,N_13232,N_13807);
and U16870 (N_16870,N_12542,N_12521);
xnor U16871 (N_16871,N_12793,N_14591);
or U16872 (N_16872,N_13124,N_13322);
and U16873 (N_16873,N_12644,N_13119);
xor U16874 (N_16874,N_12945,N_14566);
xnor U16875 (N_16875,N_12977,N_12660);
xor U16876 (N_16876,N_13588,N_12951);
nand U16877 (N_16877,N_14554,N_13896);
nor U16878 (N_16878,N_13207,N_14875);
nor U16879 (N_16879,N_13728,N_14259);
nor U16880 (N_16880,N_13095,N_13126);
nor U16881 (N_16881,N_14305,N_14587);
nand U16882 (N_16882,N_14034,N_13769);
nand U16883 (N_16883,N_14956,N_13565);
and U16884 (N_16884,N_13908,N_13758);
or U16885 (N_16885,N_13287,N_14165);
xor U16886 (N_16886,N_13584,N_14388);
xnor U16887 (N_16887,N_14609,N_14546);
xnor U16888 (N_16888,N_13285,N_14755);
and U16889 (N_16889,N_13808,N_14263);
and U16890 (N_16890,N_12610,N_12679);
and U16891 (N_16891,N_13891,N_13310);
and U16892 (N_16892,N_13869,N_13259);
nand U16893 (N_16893,N_14638,N_13663);
xor U16894 (N_16894,N_13310,N_14366);
nor U16895 (N_16895,N_13785,N_14574);
nor U16896 (N_16896,N_13621,N_13697);
xnor U16897 (N_16897,N_13398,N_12777);
or U16898 (N_16898,N_14388,N_14266);
nor U16899 (N_16899,N_13892,N_14273);
nand U16900 (N_16900,N_13043,N_13100);
or U16901 (N_16901,N_14042,N_12785);
xnor U16902 (N_16902,N_13933,N_12995);
and U16903 (N_16903,N_13286,N_14788);
xor U16904 (N_16904,N_14526,N_13965);
and U16905 (N_16905,N_12986,N_13924);
xnor U16906 (N_16906,N_13791,N_14153);
xnor U16907 (N_16907,N_13069,N_14595);
xor U16908 (N_16908,N_12822,N_13278);
and U16909 (N_16909,N_13878,N_12610);
or U16910 (N_16910,N_13593,N_14149);
nand U16911 (N_16911,N_13420,N_14029);
nor U16912 (N_16912,N_13303,N_13095);
and U16913 (N_16913,N_12622,N_14201);
xor U16914 (N_16914,N_14281,N_14679);
nor U16915 (N_16915,N_12760,N_14932);
or U16916 (N_16916,N_13403,N_14459);
nand U16917 (N_16917,N_13804,N_14246);
or U16918 (N_16918,N_14462,N_12577);
xor U16919 (N_16919,N_14270,N_14184);
and U16920 (N_16920,N_14587,N_14665);
and U16921 (N_16921,N_14309,N_14505);
and U16922 (N_16922,N_12664,N_13610);
nand U16923 (N_16923,N_12983,N_14661);
xor U16924 (N_16924,N_14845,N_14953);
or U16925 (N_16925,N_12935,N_13530);
or U16926 (N_16926,N_13044,N_14737);
or U16927 (N_16927,N_13110,N_14947);
nand U16928 (N_16928,N_14869,N_13396);
or U16929 (N_16929,N_13835,N_13319);
xor U16930 (N_16930,N_14522,N_14687);
and U16931 (N_16931,N_12880,N_14609);
nand U16932 (N_16932,N_13758,N_14040);
nand U16933 (N_16933,N_13402,N_13860);
or U16934 (N_16934,N_13826,N_12586);
or U16935 (N_16935,N_13454,N_13278);
xnor U16936 (N_16936,N_13580,N_14307);
or U16937 (N_16937,N_14078,N_14985);
nand U16938 (N_16938,N_13503,N_14548);
xnor U16939 (N_16939,N_13324,N_14765);
or U16940 (N_16940,N_12945,N_12606);
nand U16941 (N_16941,N_14408,N_13758);
nand U16942 (N_16942,N_14147,N_13474);
xnor U16943 (N_16943,N_14772,N_14024);
xor U16944 (N_16944,N_13364,N_14076);
nand U16945 (N_16945,N_13850,N_13987);
and U16946 (N_16946,N_12822,N_13333);
nand U16947 (N_16947,N_14180,N_14663);
xor U16948 (N_16948,N_13725,N_14147);
and U16949 (N_16949,N_14953,N_13871);
nor U16950 (N_16950,N_13946,N_14037);
nor U16951 (N_16951,N_12637,N_13432);
and U16952 (N_16952,N_14377,N_12601);
xor U16953 (N_16953,N_12689,N_14798);
and U16954 (N_16954,N_14000,N_14933);
nand U16955 (N_16955,N_12684,N_14094);
nand U16956 (N_16956,N_12589,N_14884);
and U16957 (N_16957,N_13703,N_14708);
nor U16958 (N_16958,N_13615,N_12897);
nor U16959 (N_16959,N_13124,N_13264);
nand U16960 (N_16960,N_14656,N_14756);
or U16961 (N_16961,N_13320,N_14870);
or U16962 (N_16962,N_14366,N_14744);
and U16963 (N_16963,N_13568,N_14347);
xor U16964 (N_16964,N_13455,N_12693);
and U16965 (N_16965,N_13216,N_12915);
or U16966 (N_16966,N_12785,N_13041);
nand U16967 (N_16967,N_14509,N_13556);
nor U16968 (N_16968,N_13518,N_12883);
nor U16969 (N_16969,N_13831,N_13422);
or U16970 (N_16970,N_13258,N_13678);
and U16971 (N_16971,N_13935,N_14409);
nor U16972 (N_16972,N_13015,N_13290);
nor U16973 (N_16973,N_14554,N_12774);
nor U16974 (N_16974,N_14047,N_13759);
and U16975 (N_16975,N_13624,N_14652);
or U16976 (N_16976,N_13429,N_13516);
or U16977 (N_16977,N_12673,N_14869);
and U16978 (N_16978,N_13026,N_14074);
nand U16979 (N_16979,N_14331,N_13817);
nand U16980 (N_16980,N_14640,N_13165);
xor U16981 (N_16981,N_13496,N_13089);
nand U16982 (N_16982,N_12677,N_12502);
xor U16983 (N_16983,N_13239,N_12561);
xor U16984 (N_16984,N_13935,N_13163);
nand U16985 (N_16985,N_13403,N_13349);
xor U16986 (N_16986,N_12519,N_13037);
nor U16987 (N_16987,N_14671,N_13550);
or U16988 (N_16988,N_14972,N_12864);
xnor U16989 (N_16989,N_13479,N_13398);
nand U16990 (N_16990,N_13026,N_14186);
xnor U16991 (N_16991,N_12788,N_14512);
and U16992 (N_16992,N_13385,N_12732);
nor U16993 (N_16993,N_13802,N_14838);
and U16994 (N_16994,N_14970,N_14506);
nand U16995 (N_16995,N_13814,N_13074);
nand U16996 (N_16996,N_14934,N_13372);
nand U16997 (N_16997,N_13043,N_14131);
and U16998 (N_16998,N_12519,N_12655);
nand U16999 (N_16999,N_12567,N_14722);
nand U17000 (N_17000,N_12877,N_14936);
and U17001 (N_17001,N_12808,N_12895);
and U17002 (N_17002,N_13023,N_13252);
or U17003 (N_17003,N_14164,N_12988);
or U17004 (N_17004,N_13095,N_14765);
and U17005 (N_17005,N_12682,N_13537);
nor U17006 (N_17006,N_13222,N_13827);
or U17007 (N_17007,N_14678,N_14890);
or U17008 (N_17008,N_13668,N_13997);
nor U17009 (N_17009,N_12907,N_14050);
xnor U17010 (N_17010,N_12641,N_14416);
or U17011 (N_17011,N_14630,N_13344);
or U17012 (N_17012,N_13725,N_13854);
nor U17013 (N_17013,N_13320,N_14758);
and U17014 (N_17014,N_14711,N_14149);
xnor U17015 (N_17015,N_13391,N_13599);
nor U17016 (N_17016,N_13644,N_13506);
nand U17017 (N_17017,N_13623,N_12718);
and U17018 (N_17018,N_12833,N_13132);
nor U17019 (N_17019,N_13174,N_14541);
or U17020 (N_17020,N_14490,N_13031);
and U17021 (N_17021,N_13825,N_14337);
nor U17022 (N_17022,N_13032,N_12557);
nor U17023 (N_17023,N_14749,N_13602);
nor U17024 (N_17024,N_12818,N_12611);
or U17025 (N_17025,N_13690,N_13407);
or U17026 (N_17026,N_14523,N_14356);
nor U17027 (N_17027,N_12940,N_13925);
or U17028 (N_17028,N_13459,N_12568);
nand U17029 (N_17029,N_14399,N_14314);
xor U17030 (N_17030,N_13976,N_14294);
or U17031 (N_17031,N_12641,N_12580);
xor U17032 (N_17032,N_12787,N_13529);
xnor U17033 (N_17033,N_12981,N_14096);
nand U17034 (N_17034,N_14412,N_13827);
xnor U17035 (N_17035,N_13240,N_14661);
xnor U17036 (N_17036,N_14096,N_12661);
xor U17037 (N_17037,N_13691,N_13179);
xnor U17038 (N_17038,N_12705,N_12986);
nand U17039 (N_17039,N_13038,N_13416);
and U17040 (N_17040,N_14830,N_12541);
nand U17041 (N_17041,N_14137,N_13470);
nor U17042 (N_17042,N_14382,N_14994);
nor U17043 (N_17043,N_13580,N_14629);
and U17044 (N_17044,N_13919,N_14260);
xor U17045 (N_17045,N_14244,N_14896);
nand U17046 (N_17046,N_12943,N_13906);
nor U17047 (N_17047,N_12959,N_13352);
and U17048 (N_17048,N_14147,N_13488);
and U17049 (N_17049,N_12604,N_13773);
nand U17050 (N_17050,N_13499,N_13176);
nor U17051 (N_17051,N_13939,N_14308);
nor U17052 (N_17052,N_12881,N_12621);
nor U17053 (N_17053,N_13953,N_14850);
xnor U17054 (N_17054,N_13987,N_12630);
nor U17055 (N_17055,N_14938,N_14434);
or U17056 (N_17056,N_14168,N_13698);
xnor U17057 (N_17057,N_12555,N_12872);
and U17058 (N_17058,N_13582,N_14648);
xnor U17059 (N_17059,N_14077,N_13138);
xnor U17060 (N_17060,N_14870,N_14672);
and U17061 (N_17061,N_14224,N_13904);
xor U17062 (N_17062,N_14854,N_13247);
nor U17063 (N_17063,N_13916,N_13659);
or U17064 (N_17064,N_14687,N_14048);
nor U17065 (N_17065,N_12966,N_12993);
xnor U17066 (N_17066,N_14794,N_13580);
nand U17067 (N_17067,N_14091,N_14012);
and U17068 (N_17068,N_13958,N_14278);
xor U17069 (N_17069,N_13156,N_12699);
nor U17070 (N_17070,N_14458,N_14174);
and U17071 (N_17071,N_13333,N_13011);
xor U17072 (N_17072,N_14187,N_12785);
nor U17073 (N_17073,N_14020,N_13560);
nand U17074 (N_17074,N_14205,N_12792);
nor U17075 (N_17075,N_12602,N_13655);
or U17076 (N_17076,N_12861,N_14644);
nor U17077 (N_17077,N_12821,N_14035);
nor U17078 (N_17078,N_14250,N_14998);
xor U17079 (N_17079,N_12854,N_13164);
nor U17080 (N_17080,N_14545,N_14364);
nand U17081 (N_17081,N_14759,N_14205);
and U17082 (N_17082,N_13970,N_13812);
xnor U17083 (N_17083,N_12966,N_12767);
or U17084 (N_17084,N_14812,N_12822);
xor U17085 (N_17085,N_14875,N_14690);
nor U17086 (N_17086,N_13667,N_13801);
xor U17087 (N_17087,N_14022,N_12865);
and U17088 (N_17088,N_12785,N_14146);
nand U17089 (N_17089,N_14391,N_13425);
and U17090 (N_17090,N_14865,N_14495);
xor U17091 (N_17091,N_12943,N_14248);
or U17092 (N_17092,N_13041,N_14482);
or U17093 (N_17093,N_12840,N_13252);
nor U17094 (N_17094,N_13712,N_14631);
and U17095 (N_17095,N_14752,N_14836);
xnor U17096 (N_17096,N_13039,N_13579);
and U17097 (N_17097,N_14699,N_12579);
and U17098 (N_17098,N_13122,N_13884);
xor U17099 (N_17099,N_12778,N_14785);
nand U17100 (N_17100,N_14203,N_13512);
or U17101 (N_17101,N_12541,N_13718);
and U17102 (N_17102,N_14326,N_13582);
xor U17103 (N_17103,N_14517,N_13783);
nand U17104 (N_17104,N_12975,N_12671);
xor U17105 (N_17105,N_14320,N_13123);
and U17106 (N_17106,N_14732,N_13071);
nand U17107 (N_17107,N_14311,N_14053);
nor U17108 (N_17108,N_13471,N_12954);
and U17109 (N_17109,N_12540,N_14589);
or U17110 (N_17110,N_12712,N_14296);
and U17111 (N_17111,N_14542,N_13206);
nor U17112 (N_17112,N_14301,N_13887);
nor U17113 (N_17113,N_13198,N_13217);
nand U17114 (N_17114,N_13974,N_12730);
nor U17115 (N_17115,N_13240,N_14986);
nand U17116 (N_17116,N_13826,N_12961);
nand U17117 (N_17117,N_13357,N_13422);
nand U17118 (N_17118,N_14019,N_13474);
or U17119 (N_17119,N_13359,N_14747);
nor U17120 (N_17120,N_14402,N_14178);
or U17121 (N_17121,N_13746,N_13790);
xnor U17122 (N_17122,N_14007,N_12909);
and U17123 (N_17123,N_12918,N_13456);
and U17124 (N_17124,N_13969,N_13918);
or U17125 (N_17125,N_12661,N_13101);
or U17126 (N_17126,N_12536,N_14400);
nor U17127 (N_17127,N_12922,N_14780);
nand U17128 (N_17128,N_14113,N_14000);
xnor U17129 (N_17129,N_13680,N_13381);
nand U17130 (N_17130,N_14970,N_14444);
or U17131 (N_17131,N_14524,N_13333);
and U17132 (N_17132,N_14466,N_14898);
nand U17133 (N_17133,N_13194,N_14587);
xor U17134 (N_17134,N_12797,N_13721);
xor U17135 (N_17135,N_12898,N_14440);
and U17136 (N_17136,N_12890,N_14090);
or U17137 (N_17137,N_14141,N_13423);
nand U17138 (N_17138,N_12984,N_14516);
nand U17139 (N_17139,N_14425,N_12597);
nor U17140 (N_17140,N_14118,N_14461);
and U17141 (N_17141,N_12941,N_12999);
and U17142 (N_17142,N_13937,N_13903);
nor U17143 (N_17143,N_12990,N_12892);
or U17144 (N_17144,N_12673,N_13102);
nand U17145 (N_17145,N_13089,N_14295);
nand U17146 (N_17146,N_13645,N_14585);
nand U17147 (N_17147,N_13087,N_13262);
xnor U17148 (N_17148,N_14029,N_13040);
or U17149 (N_17149,N_14266,N_13624);
or U17150 (N_17150,N_14297,N_13073);
nand U17151 (N_17151,N_13920,N_14374);
xnor U17152 (N_17152,N_14517,N_13031);
and U17153 (N_17153,N_13323,N_14718);
and U17154 (N_17154,N_13388,N_14112);
and U17155 (N_17155,N_14949,N_14733);
and U17156 (N_17156,N_13228,N_13684);
xnor U17157 (N_17157,N_13854,N_13562);
and U17158 (N_17158,N_13525,N_14165);
or U17159 (N_17159,N_14595,N_14575);
or U17160 (N_17160,N_12581,N_13006);
and U17161 (N_17161,N_13268,N_13776);
nor U17162 (N_17162,N_14272,N_13933);
or U17163 (N_17163,N_12675,N_13904);
or U17164 (N_17164,N_13181,N_14028);
nand U17165 (N_17165,N_12552,N_13008);
nand U17166 (N_17166,N_14142,N_13128);
or U17167 (N_17167,N_14466,N_12595);
xnor U17168 (N_17168,N_13444,N_14731);
or U17169 (N_17169,N_14404,N_13003);
nor U17170 (N_17170,N_14794,N_13362);
xor U17171 (N_17171,N_12985,N_13446);
or U17172 (N_17172,N_13629,N_12567);
nand U17173 (N_17173,N_14871,N_14412);
nor U17174 (N_17174,N_12529,N_13107);
nand U17175 (N_17175,N_14845,N_14291);
xnor U17176 (N_17176,N_12587,N_13997);
xor U17177 (N_17177,N_12695,N_13670);
xnor U17178 (N_17178,N_13524,N_12821);
nand U17179 (N_17179,N_14976,N_13159);
nor U17180 (N_17180,N_13527,N_13803);
xnor U17181 (N_17181,N_13477,N_14281);
nand U17182 (N_17182,N_13701,N_12968);
nand U17183 (N_17183,N_14693,N_14716);
and U17184 (N_17184,N_12661,N_12687);
nor U17185 (N_17185,N_13438,N_14229);
and U17186 (N_17186,N_14316,N_12514);
and U17187 (N_17187,N_13796,N_13008);
and U17188 (N_17188,N_14387,N_14075);
nand U17189 (N_17189,N_12905,N_13658);
or U17190 (N_17190,N_14662,N_13613);
xnor U17191 (N_17191,N_12695,N_12788);
and U17192 (N_17192,N_13041,N_12968);
nor U17193 (N_17193,N_13313,N_12844);
or U17194 (N_17194,N_13690,N_13676);
nor U17195 (N_17195,N_13507,N_14545);
nor U17196 (N_17196,N_14554,N_13048);
nor U17197 (N_17197,N_13861,N_12825);
nand U17198 (N_17198,N_14848,N_14466);
or U17199 (N_17199,N_12788,N_12982);
nor U17200 (N_17200,N_13121,N_14037);
and U17201 (N_17201,N_14749,N_12641);
or U17202 (N_17202,N_13994,N_13151);
and U17203 (N_17203,N_13602,N_12522);
xnor U17204 (N_17204,N_13520,N_14993);
nand U17205 (N_17205,N_13785,N_14659);
or U17206 (N_17206,N_14548,N_14888);
xor U17207 (N_17207,N_13700,N_13014);
nor U17208 (N_17208,N_13259,N_14474);
nand U17209 (N_17209,N_14248,N_14009);
nand U17210 (N_17210,N_12924,N_14227);
or U17211 (N_17211,N_12623,N_13705);
nand U17212 (N_17212,N_14986,N_12850);
or U17213 (N_17213,N_14912,N_14132);
and U17214 (N_17214,N_13363,N_14201);
nor U17215 (N_17215,N_14136,N_14547);
nand U17216 (N_17216,N_13839,N_14787);
and U17217 (N_17217,N_13483,N_14561);
nand U17218 (N_17218,N_14102,N_14476);
nand U17219 (N_17219,N_13576,N_12517);
and U17220 (N_17220,N_13845,N_13017);
or U17221 (N_17221,N_13384,N_12852);
nand U17222 (N_17222,N_13874,N_13247);
or U17223 (N_17223,N_12844,N_13717);
nor U17224 (N_17224,N_12755,N_13353);
nand U17225 (N_17225,N_14838,N_13341);
nand U17226 (N_17226,N_13377,N_12783);
nand U17227 (N_17227,N_13496,N_13601);
and U17228 (N_17228,N_13502,N_12551);
nand U17229 (N_17229,N_14304,N_12813);
xnor U17230 (N_17230,N_14346,N_14734);
nor U17231 (N_17231,N_14783,N_14852);
nand U17232 (N_17232,N_13592,N_14776);
nand U17233 (N_17233,N_14924,N_13150);
nand U17234 (N_17234,N_14658,N_12634);
nor U17235 (N_17235,N_14198,N_14860);
nor U17236 (N_17236,N_13740,N_13449);
nand U17237 (N_17237,N_12695,N_14996);
nor U17238 (N_17238,N_13560,N_14715);
nor U17239 (N_17239,N_14681,N_13889);
xnor U17240 (N_17240,N_13881,N_12610);
nand U17241 (N_17241,N_13456,N_12888);
or U17242 (N_17242,N_13567,N_13886);
nand U17243 (N_17243,N_12711,N_13463);
nand U17244 (N_17244,N_14995,N_13999);
xor U17245 (N_17245,N_13088,N_14432);
and U17246 (N_17246,N_14296,N_12640);
nor U17247 (N_17247,N_13450,N_13473);
nand U17248 (N_17248,N_14139,N_12904);
or U17249 (N_17249,N_13834,N_14659);
and U17250 (N_17250,N_12730,N_13063);
and U17251 (N_17251,N_13261,N_12662);
nor U17252 (N_17252,N_13255,N_13857);
nand U17253 (N_17253,N_14909,N_13945);
and U17254 (N_17254,N_13606,N_14566);
nand U17255 (N_17255,N_14137,N_14657);
xnor U17256 (N_17256,N_14750,N_13767);
nor U17257 (N_17257,N_12556,N_13275);
nor U17258 (N_17258,N_14228,N_14594);
xnor U17259 (N_17259,N_14983,N_14513);
nand U17260 (N_17260,N_13566,N_13634);
or U17261 (N_17261,N_13888,N_13714);
and U17262 (N_17262,N_12721,N_12906);
xor U17263 (N_17263,N_13848,N_12882);
xor U17264 (N_17264,N_14442,N_14665);
and U17265 (N_17265,N_13810,N_12846);
xnor U17266 (N_17266,N_12516,N_14332);
nand U17267 (N_17267,N_14046,N_14281);
nand U17268 (N_17268,N_13048,N_12721);
nor U17269 (N_17269,N_12992,N_12830);
xnor U17270 (N_17270,N_14742,N_13771);
nor U17271 (N_17271,N_13916,N_13828);
or U17272 (N_17272,N_12581,N_13631);
nor U17273 (N_17273,N_13224,N_13516);
nor U17274 (N_17274,N_13293,N_13960);
and U17275 (N_17275,N_13991,N_13719);
nor U17276 (N_17276,N_13686,N_14190);
and U17277 (N_17277,N_13267,N_13854);
and U17278 (N_17278,N_14395,N_12814);
nor U17279 (N_17279,N_14098,N_13413);
and U17280 (N_17280,N_13043,N_13540);
or U17281 (N_17281,N_14000,N_14042);
or U17282 (N_17282,N_13448,N_14578);
xnor U17283 (N_17283,N_14227,N_13097);
and U17284 (N_17284,N_13278,N_12966);
nor U17285 (N_17285,N_14271,N_14739);
and U17286 (N_17286,N_13406,N_12853);
and U17287 (N_17287,N_14492,N_12961);
nor U17288 (N_17288,N_13967,N_12843);
or U17289 (N_17289,N_13624,N_14702);
and U17290 (N_17290,N_14318,N_13958);
nand U17291 (N_17291,N_13130,N_12882);
or U17292 (N_17292,N_13784,N_13497);
nor U17293 (N_17293,N_14913,N_12672);
and U17294 (N_17294,N_13081,N_14891);
nor U17295 (N_17295,N_14376,N_12674);
xnor U17296 (N_17296,N_14330,N_13747);
and U17297 (N_17297,N_13699,N_12610);
or U17298 (N_17298,N_13033,N_13824);
or U17299 (N_17299,N_14595,N_14263);
or U17300 (N_17300,N_14685,N_14039);
xor U17301 (N_17301,N_14880,N_14911);
xor U17302 (N_17302,N_14495,N_14818);
nand U17303 (N_17303,N_12788,N_14937);
or U17304 (N_17304,N_14885,N_13258);
xor U17305 (N_17305,N_14134,N_13242);
or U17306 (N_17306,N_13433,N_14763);
xnor U17307 (N_17307,N_13070,N_12742);
or U17308 (N_17308,N_14423,N_14100);
nor U17309 (N_17309,N_14047,N_12696);
and U17310 (N_17310,N_13931,N_14872);
nor U17311 (N_17311,N_13173,N_13697);
nor U17312 (N_17312,N_13181,N_13083);
xnor U17313 (N_17313,N_12713,N_14366);
or U17314 (N_17314,N_12890,N_14437);
or U17315 (N_17315,N_14312,N_13156);
and U17316 (N_17316,N_14800,N_14319);
nand U17317 (N_17317,N_14311,N_13424);
xor U17318 (N_17318,N_12882,N_12689);
nor U17319 (N_17319,N_13022,N_13327);
nand U17320 (N_17320,N_14904,N_12933);
and U17321 (N_17321,N_12649,N_14550);
nor U17322 (N_17322,N_13279,N_13680);
and U17323 (N_17323,N_14145,N_13809);
or U17324 (N_17324,N_12999,N_13701);
nand U17325 (N_17325,N_13729,N_14224);
and U17326 (N_17326,N_13030,N_14757);
and U17327 (N_17327,N_14868,N_13188);
and U17328 (N_17328,N_14769,N_13062);
nor U17329 (N_17329,N_14072,N_14786);
or U17330 (N_17330,N_14891,N_13303);
and U17331 (N_17331,N_12710,N_14986);
and U17332 (N_17332,N_13213,N_14547);
nor U17333 (N_17333,N_12903,N_14191);
and U17334 (N_17334,N_13516,N_14175);
nor U17335 (N_17335,N_12726,N_12963);
and U17336 (N_17336,N_13154,N_14819);
nor U17337 (N_17337,N_14901,N_13483);
or U17338 (N_17338,N_13746,N_12732);
xor U17339 (N_17339,N_13086,N_13012);
xor U17340 (N_17340,N_14326,N_13653);
nor U17341 (N_17341,N_14348,N_14793);
or U17342 (N_17342,N_14122,N_14414);
nor U17343 (N_17343,N_13839,N_14776);
nand U17344 (N_17344,N_13508,N_13185);
and U17345 (N_17345,N_12746,N_12563);
or U17346 (N_17346,N_13940,N_14900);
nor U17347 (N_17347,N_13151,N_13188);
xor U17348 (N_17348,N_14887,N_13486);
xor U17349 (N_17349,N_14768,N_12559);
xor U17350 (N_17350,N_13575,N_14248);
or U17351 (N_17351,N_13471,N_13796);
nor U17352 (N_17352,N_12569,N_13972);
nor U17353 (N_17353,N_14983,N_14025);
and U17354 (N_17354,N_14762,N_12554);
xnor U17355 (N_17355,N_13255,N_13125);
nor U17356 (N_17356,N_12886,N_13601);
nor U17357 (N_17357,N_14650,N_14951);
xor U17358 (N_17358,N_14356,N_13569);
or U17359 (N_17359,N_14458,N_14836);
and U17360 (N_17360,N_13108,N_13974);
nor U17361 (N_17361,N_14167,N_13900);
nor U17362 (N_17362,N_14750,N_14392);
nor U17363 (N_17363,N_14650,N_14873);
or U17364 (N_17364,N_13138,N_13716);
nor U17365 (N_17365,N_14301,N_13136);
or U17366 (N_17366,N_13247,N_13092);
or U17367 (N_17367,N_13630,N_14676);
or U17368 (N_17368,N_13591,N_14964);
nand U17369 (N_17369,N_13971,N_13752);
nand U17370 (N_17370,N_13845,N_13060);
nand U17371 (N_17371,N_14203,N_13794);
nand U17372 (N_17372,N_12901,N_14853);
xnor U17373 (N_17373,N_14723,N_13623);
nor U17374 (N_17374,N_14248,N_13619);
or U17375 (N_17375,N_13572,N_14243);
xnor U17376 (N_17376,N_12909,N_13123);
and U17377 (N_17377,N_14392,N_14089);
nor U17378 (N_17378,N_14803,N_12757);
nor U17379 (N_17379,N_12570,N_13618);
or U17380 (N_17380,N_14396,N_13039);
or U17381 (N_17381,N_14924,N_13115);
and U17382 (N_17382,N_13393,N_12684);
and U17383 (N_17383,N_14834,N_12822);
xnor U17384 (N_17384,N_13636,N_13126);
nor U17385 (N_17385,N_13517,N_14178);
nand U17386 (N_17386,N_12979,N_12960);
and U17387 (N_17387,N_13137,N_12525);
nand U17388 (N_17388,N_12983,N_13278);
xor U17389 (N_17389,N_12752,N_12945);
nand U17390 (N_17390,N_14590,N_13457);
nand U17391 (N_17391,N_14097,N_14324);
xnor U17392 (N_17392,N_12610,N_14075);
or U17393 (N_17393,N_14436,N_13065);
nor U17394 (N_17394,N_13673,N_14814);
nand U17395 (N_17395,N_14724,N_14093);
xnor U17396 (N_17396,N_13865,N_14230);
nor U17397 (N_17397,N_14737,N_13154);
nand U17398 (N_17398,N_13199,N_12707);
or U17399 (N_17399,N_12745,N_13548);
nand U17400 (N_17400,N_14555,N_12731);
nand U17401 (N_17401,N_14315,N_14093);
nor U17402 (N_17402,N_12789,N_14581);
nand U17403 (N_17403,N_14570,N_14039);
xnor U17404 (N_17404,N_14686,N_14691);
or U17405 (N_17405,N_12658,N_14668);
nor U17406 (N_17406,N_14820,N_14413);
nand U17407 (N_17407,N_12889,N_12768);
or U17408 (N_17408,N_12591,N_12595);
or U17409 (N_17409,N_14661,N_14587);
nand U17410 (N_17410,N_14268,N_13880);
or U17411 (N_17411,N_13147,N_12510);
and U17412 (N_17412,N_14694,N_14159);
nand U17413 (N_17413,N_14411,N_12987);
xnor U17414 (N_17414,N_13111,N_14561);
nand U17415 (N_17415,N_13363,N_14114);
and U17416 (N_17416,N_13300,N_14934);
nor U17417 (N_17417,N_12629,N_13750);
nor U17418 (N_17418,N_12586,N_14359);
or U17419 (N_17419,N_13137,N_12512);
xor U17420 (N_17420,N_13057,N_13111);
or U17421 (N_17421,N_12597,N_12756);
or U17422 (N_17422,N_14286,N_13815);
nand U17423 (N_17423,N_13380,N_14560);
nor U17424 (N_17424,N_13454,N_13099);
nand U17425 (N_17425,N_13084,N_14079);
xnor U17426 (N_17426,N_14186,N_13336);
nand U17427 (N_17427,N_13068,N_13554);
nand U17428 (N_17428,N_12575,N_14415);
or U17429 (N_17429,N_12513,N_14899);
and U17430 (N_17430,N_13437,N_13235);
nand U17431 (N_17431,N_14838,N_14303);
or U17432 (N_17432,N_13360,N_14435);
nor U17433 (N_17433,N_14089,N_13868);
nor U17434 (N_17434,N_14019,N_14279);
or U17435 (N_17435,N_14278,N_13771);
or U17436 (N_17436,N_13999,N_14359);
nor U17437 (N_17437,N_13559,N_13145);
xnor U17438 (N_17438,N_13821,N_14373);
and U17439 (N_17439,N_13834,N_14533);
nand U17440 (N_17440,N_13757,N_12948);
or U17441 (N_17441,N_14269,N_12511);
nor U17442 (N_17442,N_13708,N_14956);
or U17443 (N_17443,N_14602,N_12796);
or U17444 (N_17444,N_14020,N_13300);
nor U17445 (N_17445,N_13604,N_14186);
and U17446 (N_17446,N_13366,N_13643);
xnor U17447 (N_17447,N_14001,N_14271);
or U17448 (N_17448,N_14943,N_13141);
nand U17449 (N_17449,N_13994,N_14803);
and U17450 (N_17450,N_12931,N_12727);
nand U17451 (N_17451,N_14607,N_13321);
or U17452 (N_17452,N_14810,N_13192);
or U17453 (N_17453,N_14261,N_12824);
nand U17454 (N_17454,N_13630,N_12577);
and U17455 (N_17455,N_12878,N_12520);
nand U17456 (N_17456,N_14660,N_13168);
and U17457 (N_17457,N_14145,N_14873);
nand U17458 (N_17458,N_14516,N_14317);
nor U17459 (N_17459,N_12515,N_13948);
nand U17460 (N_17460,N_13261,N_14644);
nand U17461 (N_17461,N_12724,N_13073);
and U17462 (N_17462,N_14891,N_13234);
or U17463 (N_17463,N_14694,N_12611);
xnor U17464 (N_17464,N_13762,N_14213);
nand U17465 (N_17465,N_14931,N_14967);
nand U17466 (N_17466,N_12500,N_13384);
nor U17467 (N_17467,N_13768,N_13517);
nor U17468 (N_17468,N_12690,N_13211);
xor U17469 (N_17469,N_13155,N_13439);
or U17470 (N_17470,N_14435,N_13999);
or U17471 (N_17471,N_14111,N_13743);
xnor U17472 (N_17472,N_12957,N_14069);
or U17473 (N_17473,N_13553,N_14708);
xnor U17474 (N_17474,N_12607,N_13010);
or U17475 (N_17475,N_12562,N_13786);
xnor U17476 (N_17476,N_14537,N_12521);
xnor U17477 (N_17477,N_13959,N_13135);
nand U17478 (N_17478,N_14620,N_13200);
xor U17479 (N_17479,N_14626,N_13872);
or U17480 (N_17480,N_13041,N_14480);
xnor U17481 (N_17481,N_13056,N_14122);
and U17482 (N_17482,N_13175,N_14751);
nor U17483 (N_17483,N_13770,N_14638);
nor U17484 (N_17484,N_12696,N_14439);
xnor U17485 (N_17485,N_13472,N_14822);
or U17486 (N_17486,N_13879,N_14251);
and U17487 (N_17487,N_13401,N_12798);
nand U17488 (N_17488,N_13925,N_14281);
and U17489 (N_17489,N_14841,N_14637);
and U17490 (N_17490,N_13804,N_14714);
or U17491 (N_17491,N_13129,N_13412);
nand U17492 (N_17492,N_14241,N_12808);
and U17493 (N_17493,N_13250,N_14993);
and U17494 (N_17494,N_14905,N_12936);
nand U17495 (N_17495,N_12569,N_12717);
or U17496 (N_17496,N_14972,N_13080);
or U17497 (N_17497,N_13453,N_13281);
or U17498 (N_17498,N_13865,N_12786);
nand U17499 (N_17499,N_12806,N_13072);
and U17500 (N_17500,N_15455,N_16699);
or U17501 (N_17501,N_15305,N_16513);
xnor U17502 (N_17502,N_16966,N_16934);
nand U17503 (N_17503,N_15125,N_15683);
nor U17504 (N_17504,N_15597,N_17243);
and U17505 (N_17505,N_16256,N_15576);
or U17506 (N_17506,N_15556,N_16127);
or U17507 (N_17507,N_16314,N_16840);
nand U17508 (N_17508,N_16382,N_16079);
nand U17509 (N_17509,N_15417,N_15191);
xnor U17510 (N_17510,N_16827,N_16643);
and U17511 (N_17511,N_16979,N_15278);
nand U17512 (N_17512,N_15520,N_17419);
and U17513 (N_17513,N_16989,N_16284);
nor U17514 (N_17514,N_17148,N_15533);
nor U17515 (N_17515,N_15512,N_15812);
and U17516 (N_17516,N_17150,N_16512);
xnor U17517 (N_17517,N_15905,N_16747);
nor U17518 (N_17518,N_15044,N_16907);
or U17519 (N_17519,N_16549,N_17047);
nand U17520 (N_17520,N_15988,N_15953);
and U17521 (N_17521,N_15565,N_16520);
and U17522 (N_17522,N_15386,N_16004);
or U17523 (N_17523,N_17038,N_16442);
and U17524 (N_17524,N_17286,N_15684);
xor U17525 (N_17525,N_16764,N_16250);
nand U17526 (N_17526,N_16420,N_16164);
xnor U17527 (N_17527,N_16338,N_17266);
and U17528 (N_17528,N_15303,N_16854);
nor U17529 (N_17529,N_15767,N_17016);
or U17530 (N_17530,N_15972,N_15977);
or U17531 (N_17531,N_15122,N_15699);
xor U17532 (N_17532,N_17379,N_16807);
nor U17533 (N_17533,N_16388,N_15243);
and U17534 (N_17534,N_16012,N_15105);
and U17535 (N_17535,N_15523,N_15898);
and U17536 (N_17536,N_15548,N_15844);
nor U17537 (N_17537,N_15215,N_17043);
or U17538 (N_17538,N_17453,N_15101);
or U17539 (N_17539,N_17474,N_16637);
and U17540 (N_17540,N_16589,N_16060);
xor U17541 (N_17541,N_15840,N_16550);
or U17542 (N_17542,N_15820,N_16812);
or U17543 (N_17543,N_15677,N_17054);
xnor U17544 (N_17544,N_16066,N_15255);
and U17545 (N_17545,N_16571,N_17022);
xor U17546 (N_17546,N_17028,N_15049);
or U17547 (N_17547,N_15161,N_16475);
xor U17548 (N_17548,N_15100,N_15273);
and U17549 (N_17549,N_15950,N_15685);
and U17550 (N_17550,N_16150,N_15630);
or U17551 (N_17551,N_15747,N_17133);
nand U17552 (N_17552,N_15909,N_15661);
and U17553 (N_17553,N_16304,N_15458);
nand U17554 (N_17554,N_15194,N_15642);
nor U17555 (N_17555,N_15516,N_16581);
xnor U17556 (N_17556,N_17198,N_16514);
and U17557 (N_17557,N_16358,N_15230);
and U17558 (N_17558,N_15078,N_17300);
and U17559 (N_17559,N_17007,N_17230);
xor U17560 (N_17560,N_15061,N_15599);
nor U17561 (N_17561,N_17153,N_16819);
and U17562 (N_17562,N_17174,N_15018);
and U17563 (N_17563,N_16678,N_15221);
nor U17564 (N_17564,N_16748,N_15394);
nand U17565 (N_17565,N_16786,N_16599);
and U17566 (N_17566,N_15934,N_15427);
and U17567 (N_17567,N_16009,N_16644);
nand U17568 (N_17568,N_15709,N_17437);
nand U17569 (N_17569,N_16887,N_16462);
or U17570 (N_17570,N_15181,N_17181);
nand U17571 (N_17571,N_16290,N_15140);
and U17572 (N_17572,N_15223,N_15942);
and U17573 (N_17573,N_16558,N_17440);
or U17574 (N_17574,N_15325,N_15829);
xor U17575 (N_17575,N_16553,N_17147);
and U17576 (N_17576,N_16479,N_16305);
nor U17577 (N_17577,N_16945,N_16321);
nor U17578 (N_17578,N_16226,N_16929);
and U17579 (N_17579,N_16158,N_15131);
or U17580 (N_17580,N_15262,N_16183);
or U17581 (N_17581,N_16441,N_16114);
or U17582 (N_17582,N_15979,N_16774);
and U17583 (N_17583,N_15527,N_17163);
and U17584 (N_17584,N_15744,N_16869);
nor U17585 (N_17585,N_16604,N_16974);
and U17586 (N_17586,N_17081,N_16387);
nand U17587 (N_17587,N_16610,N_15153);
or U17588 (N_17588,N_15041,N_17210);
xor U17589 (N_17589,N_16364,N_16179);
or U17590 (N_17590,N_17141,N_17255);
nand U17591 (N_17591,N_17018,N_15593);
xor U17592 (N_17592,N_17308,N_15773);
xnor U17593 (N_17593,N_17143,N_16204);
nor U17594 (N_17594,N_17185,N_16700);
and U17595 (N_17595,N_15819,N_17132);
nor U17596 (N_17596,N_17349,N_15207);
xor U17597 (N_17597,N_17472,N_15600);
xor U17598 (N_17598,N_15231,N_15169);
and U17599 (N_17599,N_16115,N_16283);
nor U17600 (N_17600,N_17068,N_16718);
xor U17601 (N_17601,N_16524,N_15948);
nand U17602 (N_17602,N_16689,N_16405);
and U17603 (N_17603,N_15722,N_16279);
nor U17604 (N_17604,N_15434,N_17162);
and U17605 (N_17605,N_16768,N_16815);
xnor U17606 (N_17606,N_15004,N_15232);
nand U17607 (N_17607,N_16094,N_16389);
nor U17608 (N_17608,N_16316,N_15851);
or U17609 (N_17609,N_15856,N_16662);
xnor U17610 (N_17610,N_16241,N_17443);
nand U17611 (N_17611,N_16577,N_17469);
or U17612 (N_17612,N_16765,N_15269);
nor U17613 (N_17613,N_15496,N_17160);
and U17614 (N_17614,N_15931,N_16449);
nor U17615 (N_17615,N_17244,N_17091);
or U17616 (N_17616,N_15992,N_15333);
nor U17617 (N_17617,N_16126,N_15206);
nand U17618 (N_17618,N_15892,N_15121);
xnor U17619 (N_17619,N_17214,N_15841);
or U17620 (N_17620,N_15476,N_16735);
xor U17621 (N_17621,N_15497,N_17173);
or U17622 (N_17622,N_17053,N_15023);
nand U17623 (N_17623,N_15713,N_16519);
xor U17624 (N_17624,N_15911,N_16476);
and U17625 (N_17625,N_16752,N_15257);
nor U17626 (N_17626,N_15658,N_15254);
nor U17627 (N_17627,N_16121,N_16848);
xnor U17628 (N_17628,N_16510,N_17129);
and U17629 (N_17629,N_16984,N_15771);
xor U17630 (N_17630,N_17357,N_16814);
or U17631 (N_17631,N_16049,N_16697);
or U17632 (N_17632,N_17267,N_16457);
xor U17633 (N_17633,N_17090,N_15885);
nor U17634 (N_17634,N_16077,N_15359);
nor U17635 (N_17635,N_15341,N_16086);
or U17636 (N_17636,N_17227,N_15678);
or U17637 (N_17637,N_16922,N_16638);
and U17638 (N_17638,N_15768,N_16269);
nor U17639 (N_17639,N_15432,N_15987);
nor U17640 (N_17640,N_15757,N_16953);
or U17641 (N_17641,N_15784,N_16704);
or U17642 (N_17642,N_17478,N_15149);
xor U17643 (N_17643,N_15390,N_16556);
nor U17644 (N_17644,N_15688,N_16156);
or U17645 (N_17645,N_17427,N_15200);
and U17646 (N_17646,N_15077,N_17454);
xor U17647 (N_17647,N_15261,N_17380);
or U17648 (N_17648,N_16210,N_15788);
nor U17649 (N_17649,N_17191,N_15016);
and U17650 (N_17650,N_15936,N_15906);
and U17651 (N_17651,N_16563,N_15939);
nor U17652 (N_17652,N_15726,N_16386);
xor U17653 (N_17653,N_15368,N_15995);
or U17654 (N_17654,N_15634,N_15800);
nand U17655 (N_17655,N_17445,N_16046);
nand U17656 (N_17656,N_17456,N_15542);
xor U17657 (N_17657,N_15088,N_16603);
xor U17658 (N_17658,N_15251,N_17428);
or U17659 (N_17659,N_15838,N_15863);
nor U17660 (N_17660,N_16265,N_15227);
or U17661 (N_17661,N_16749,N_15886);
nand U17662 (N_17662,N_17183,N_17390);
or U17663 (N_17663,N_17476,N_16598);
or U17664 (N_17664,N_15845,N_15259);
nor U17665 (N_17665,N_16824,N_17331);
or U17666 (N_17666,N_16890,N_16022);
xnor U17667 (N_17667,N_16285,N_15351);
nor U17668 (N_17668,N_15021,N_17395);
xor U17669 (N_17669,N_15705,N_15967);
nor U17670 (N_17670,N_17358,N_17079);
nand U17671 (N_17671,N_16935,N_17259);
and U17672 (N_17672,N_16010,N_15239);
nand U17673 (N_17673,N_15772,N_15090);
xnor U17674 (N_17674,N_16227,N_16404);
and U17675 (N_17675,N_15855,N_16138);
nand U17676 (N_17676,N_15756,N_15406);
xor U17677 (N_17677,N_16467,N_15324);
and U17678 (N_17678,N_16236,N_16507);
xnor U17679 (N_17679,N_15681,N_15913);
xor U17680 (N_17680,N_16874,N_16946);
and U17681 (N_17681,N_16048,N_16790);
nor U17682 (N_17682,N_17446,N_15138);
and U17683 (N_17683,N_17320,N_15361);
and U17684 (N_17684,N_15505,N_15103);
and U17685 (N_17685,N_16855,N_16918);
xor U17686 (N_17686,N_17050,N_16354);
nand U17687 (N_17687,N_16137,N_15952);
and U17688 (N_17688,N_17480,N_17055);
nand U17689 (N_17689,N_15258,N_15792);
xnor U17690 (N_17690,N_16853,N_17123);
nand U17691 (N_17691,N_15037,N_16008);
or U17692 (N_17692,N_17275,N_17186);
or U17693 (N_17693,N_16772,N_17101);
xor U17694 (N_17694,N_15479,N_15724);
nand U17695 (N_17695,N_15062,N_16642);
xnor U17696 (N_17696,N_15618,N_16287);
xor U17697 (N_17697,N_16175,N_16542);
nor U17698 (N_17698,N_16160,N_16731);
nor U17699 (N_17699,N_16111,N_16097);
or U17700 (N_17700,N_16818,N_17017);
or U17701 (N_17701,N_16185,N_16797);
xor U17702 (N_17702,N_15859,N_15787);
and U17703 (N_17703,N_17494,N_16417);
nand U17704 (N_17704,N_17295,N_15842);
and U17705 (N_17705,N_15382,N_15495);
or U17706 (N_17706,N_15112,N_15204);
nor U17707 (N_17707,N_16348,N_17346);
or U17708 (N_17708,N_17444,N_15235);
and U17709 (N_17709,N_17231,N_15999);
or U17710 (N_17710,N_15422,N_16882);
nor U17711 (N_17711,N_15641,N_15731);
and U17712 (N_17712,N_16844,N_16654);
nand U17713 (N_17713,N_15353,N_16851);
nand U17714 (N_17714,N_15344,N_16091);
nor U17715 (N_17715,N_15435,N_15299);
xor U17716 (N_17716,N_17188,N_16342);
or U17717 (N_17717,N_15968,N_16756);
xor U17718 (N_17718,N_16493,N_17491);
and U17719 (N_17719,N_16745,N_17058);
and U17720 (N_17720,N_16540,N_16761);
and U17721 (N_17721,N_17325,N_15289);
nor U17722 (N_17722,N_16845,N_15890);
and U17723 (N_17723,N_15954,N_16280);
or U17724 (N_17724,N_17364,N_16013);
xor U17725 (N_17725,N_17296,N_16026);
or U17726 (N_17726,N_17251,N_16968);
nand U17727 (N_17727,N_17288,N_15040);
and U17728 (N_17728,N_15826,N_15068);
or U17729 (N_17729,N_17106,N_17299);
nand U17730 (N_17730,N_17199,N_16042);
xor U17731 (N_17731,N_17413,N_16736);
nor U17732 (N_17732,N_16167,N_16368);
and U17733 (N_17733,N_16623,N_15917);
and U17734 (N_17734,N_16532,N_15810);
xnor U17735 (N_17735,N_15914,N_15391);
xor U17736 (N_17736,N_16973,N_17430);
nand U17737 (N_17737,N_15084,N_15392);
nor U17738 (N_17738,N_16205,N_15183);
nor U17739 (N_17739,N_15236,N_16289);
nor U17740 (N_17740,N_16633,N_16596);
nand U17741 (N_17741,N_15091,N_15291);
nor U17742 (N_17742,N_15164,N_15625);
xnor U17743 (N_17743,N_16559,N_17070);
and U17744 (N_17744,N_17415,N_17481);
and U17745 (N_17745,N_16548,N_16072);
nor U17746 (N_17746,N_16809,N_15431);
and U17747 (N_17747,N_16903,N_16412);
xor U17748 (N_17748,N_15009,N_16237);
xnor U17749 (N_17749,N_17011,N_16278);
and U17750 (N_17750,N_16792,N_15594);
nand U17751 (N_17751,N_15943,N_15793);
or U17752 (N_17752,N_15580,N_17350);
and U17753 (N_17753,N_17212,N_16607);
nor U17754 (N_17754,N_16419,N_16120);
and U17755 (N_17755,N_15835,N_16703);
or U17756 (N_17756,N_17277,N_16207);
xor U17757 (N_17757,N_16313,N_15837);
and U17758 (N_17758,N_15424,N_17120);
and U17759 (N_17759,N_17146,N_16339);
and U17760 (N_17760,N_17180,N_16193);
xnor U17761 (N_17761,N_17082,N_15963);
nor U17762 (N_17762,N_15312,N_16406);
nor U17763 (N_17763,N_16927,N_16397);
xnor U17764 (N_17764,N_16355,N_16605);
nor U17765 (N_17765,N_15912,N_15371);
and U17766 (N_17766,N_15447,N_16336);
and U17767 (N_17767,N_15607,N_17239);
xor U17768 (N_17768,N_16239,N_15654);
nor U17769 (N_17769,N_16334,N_15660);
xor U17770 (N_17770,N_16763,N_16229);
nand U17771 (N_17771,N_17057,N_15033);
nor U17772 (N_17772,N_16232,N_16029);
nand U17773 (N_17773,N_17176,N_17093);
nand U17774 (N_17774,N_17086,N_15623);
nand U17775 (N_17775,N_16011,N_16143);
nand U17776 (N_17776,N_16569,N_17126);
and U17777 (N_17777,N_15657,N_16883);
or U17778 (N_17778,N_15277,N_17392);
nand U17779 (N_17779,N_16410,N_16400);
xnor U17780 (N_17780,N_17327,N_16378);
nand U17781 (N_17781,N_16561,N_16690);
and U17782 (N_17782,N_16987,N_16119);
xor U17783 (N_17783,N_16852,N_15094);
or U17784 (N_17784,N_16568,N_17152);
nor U17785 (N_17785,N_17363,N_16465);
or U17786 (N_17786,N_16393,N_16455);
xor U17787 (N_17787,N_15581,N_15983);
xnor U17788 (N_17788,N_16857,N_16490);
nand U17789 (N_17789,N_15160,N_15464);
nor U17790 (N_17790,N_17439,N_16600);
xor U17791 (N_17791,N_16862,N_16168);
nor U17792 (N_17792,N_17045,N_16053);
xnor U17793 (N_17793,N_15689,N_16714);
xor U17794 (N_17794,N_15861,N_15192);
and U17795 (N_17795,N_17064,N_16025);
nor U17796 (N_17796,N_16459,N_16116);
and U17797 (N_17797,N_15414,N_17382);
and U17798 (N_17798,N_16362,N_15998);
nand U17799 (N_17799,N_16155,N_15986);
and U17800 (N_17800,N_15143,N_16954);
nor U17801 (N_17801,N_16351,N_15484);
nor U17802 (N_17802,N_16988,N_15349);
and U17803 (N_17803,N_16440,N_16257);
nor U17804 (N_17804,N_16629,N_17013);
nand U17805 (N_17805,N_15604,N_16875);
nor U17806 (N_17806,N_17383,N_15266);
xnor U17807 (N_17807,N_15478,N_17423);
nand U17808 (N_17808,N_15416,N_15467);
or U17809 (N_17809,N_15375,N_16067);
nand U17810 (N_17810,N_15737,N_17073);
and U17811 (N_17811,N_16893,N_15765);
nand U17812 (N_17812,N_16881,N_17071);
xor U17813 (N_17813,N_16565,N_15358);
nor U17814 (N_17814,N_16609,N_16031);
and U17815 (N_17815,N_15442,N_17482);
xor U17816 (N_17816,N_15538,N_16880);
xnor U17817 (N_17817,N_17448,N_16525);
nand U17818 (N_17818,N_15165,N_15794);
nor U17819 (N_17819,N_15853,N_16213);
nor U17820 (N_17820,N_17305,N_16648);
or U17821 (N_17821,N_16751,N_17246);
and U17822 (N_17822,N_15339,N_15471);
nor U17823 (N_17823,N_16335,N_15240);
nand U17824 (N_17824,N_15201,N_15318);
xnor U17825 (N_17825,N_16647,N_16482);
and U17826 (N_17826,N_16833,N_16502);
nor U17827 (N_17827,N_16312,N_15896);
or U17828 (N_17828,N_16724,N_16595);
nand U17829 (N_17829,N_16760,N_15430);
nor U17830 (N_17830,N_17004,N_16742);
xor U17831 (N_17831,N_15663,N_16640);
nor U17832 (N_17832,N_15867,N_17435);
xor U17833 (N_17833,N_16795,N_17077);
nand U17834 (N_17834,N_15309,N_16407);
xnor U17835 (N_17835,N_15904,N_16377);
nand U17836 (N_17836,N_15734,N_16602);
nor U17837 (N_17837,N_17115,N_16744);
nor U17838 (N_17838,N_17434,N_17222);
nor U17839 (N_17839,N_16949,N_16757);
or U17840 (N_17840,N_16032,N_16970);
nor U17841 (N_17841,N_16076,N_15397);
and U17842 (N_17842,N_15753,N_16508);
nor U17843 (N_17843,N_16800,N_16353);
xnor U17844 (N_17844,N_16650,N_17409);
or U17845 (N_17845,N_15976,N_16839);
xor U17846 (N_17846,N_16021,N_17194);
or U17847 (N_17847,N_15067,N_15609);
and U17848 (N_17848,N_16383,N_15880);
xnor U17849 (N_17849,N_17475,N_15111);
xor U17850 (N_17850,N_15321,N_16789);
or U17851 (N_17851,N_16661,N_15676);
xnor U17852 (N_17852,N_17204,N_16715);
nor U17853 (N_17853,N_16162,N_16017);
and U17854 (N_17854,N_16247,N_15510);
nand U17855 (N_17855,N_16211,N_16930);
xor U17856 (N_17856,N_15690,N_15462);
nand U17857 (N_17857,N_15546,N_15456);
nor U17858 (N_17858,N_15453,N_17220);
and U17859 (N_17859,N_17278,N_15878);
nor U17860 (N_17860,N_15485,N_16593);
nor U17861 (N_17861,N_17121,N_16904);
and U17862 (N_17862,N_15927,N_15005);
and U17863 (N_17863,N_15568,N_15865);
or U17864 (N_17864,N_15488,N_16359);
nand U17865 (N_17865,N_16246,N_15739);
or U17866 (N_17866,N_17362,N_15446);
or U17867 (N_17867,N_15099,N_16919);
xnor U17868 (N_17868,N_17003,N_16014);
nor U17869 (N_17869,N_16165,N_15758);
nor U17870 (N_17870,N_17381,N_16435);
nand U17871 (N_17871,N_17483,N_16430);
and U17872 (N_17872,N_16743,N_17303);
nor U17873 (N_17873,N_17361,N_16983);
xor U17874 (N_17874,N_15978,N_17464);
nor U17875 (N_17875,N_15136,N_15283);
or U17876 (N_17876,N_17490,N_17458);
and U17877 (N_17877,N_15355,N_16416);
or U17878 (N_17878,N_16537,N_15352);
and U17879 (N_17879,N_17012,N_17159);
nand U17880 (N_17880,N_15852,N_15933);
and U17881 (N_17881,N_15096,N_15082);
nor U17882 (N_17882,N_15334,N_17021);
nand U17883 (N_17883,N_15144,N_17328);
and U17884 (N_17884,N_15650,N_15736);
nor U17885 (N_17885,N_16309,N_15069);
nor U17886 (N_17886,N_15058,N_17042);
xor U17887 (N_17887,N_17084,N_16990);
nand U17888 (N_17888,N_17027,N_15779);
and U17889 (N_17889,N_16361,N_15602);
nor U17890 (N_17890,N_15601,N_16144);
nand U17891 (N_17891,N_15668,N_16635);
or U17892 (N_17892,N_16492,N_16776);
xor U17893 (N_17893,N_17046,N_17279);
nor U17894 (N_17894,N_16912,N_16617);
nor U17895 (N_17895,N_16737,N_16594);
nor U17896 (N_17896,N_15970,N_16102);
nor U17897 (N_17897,N_15760,N_15123);
or U17898 (N_17898,N_16972,N_15379);
or U17899 (N_17899,N_16228,N_15071);
or U17900 (N_17900,N_15635,N_17030);
or U17901 (N_17901,N_15899,N_15376);
or U17902 (N_17902,N_17006,N_16473);
or U17903 (N_17903,N_15854,N_17138);
or U17904 (N_17904,N_16346,N_16978);
xor U17905 (N_17905,N_17417,N_16641);
and U17906 (N_17906,N_17374,N_17497);
xnor U17907 (N_17907,N_17355,N_15189);
and U17908 (N_17908,N_15876,N_15585);
nand U17909 (N_17909,N_16999,N_16319);
or U17910 (N_17910,N_16834,N_17466);
xor U17911 (N_17911,N_16371,N_17149);
xor U17912 (N_17912,N_16310,N_17433);
and U17913 (N_17913,N_15778,N_15525);
nor U17914 (N_17914,N_16277,N_16045);
and U17915 (N_17915,N_16775,N_15174);
nand U17916 (N_17916,N_16130,N_16055);
and U17917 (N_17917,N_16439,N_15649);
and U17918 (N_17918,N_16679,N_16263);
and U17919 (N_17919,N_15811,N_16341);
nor U17920 (N_17920,N_15666,N_16695);
xnor U17921 (N_17921,N_15212,N_15322);
or U17922 (N_17922,N_15238,N_16992);
xnor U17923 (N_17923,N_15213,N_15893);
nor U17924 (N_17924,N_16961,N_15443);
xor U17925 (N_17925,N_16135,N_16431);
nor U17926 (N_17926,N_17353,N_17309);
and U17927 (N_17927,N_15648,N_16317);
and U17928 (N_17928,N_16885,N_16959);
xor U17929 (N_17929,N_15966,N_16666);
xnor U17930 (N_17930,N_16154,N_17324);
xor U17931 (N_17931,N_15958,N_15108);
nor U17932 (N_17932,N_16657,N_16147);
nor U17933 (N_17933,N_17301,N_16948);
or U17934 (N_17934,N_15761,N_16981);
nor U17935 (N_17935,N_17312,N_16157);
nand U17936 (N_17936,N_15437,N_16868);
and U17937 (N_17937,N_16709,N_17098);
nor U17938 (N_17938,N_16218,N_17157);
nand U17939 (N_17939,N_16522,N_16813);
and U17940 (N_17940,N_15219,N_15452);
nor U17941 (N_17941,N_16347,N_16499);
and U17942 (N_17942,N_15847,N_16732);
xor U17943 (N_17943,N_15571,N_15588);
nand U17944 (N_17944,N_15749,N_15117);
and U17945 (N_17945,N_15610,N_16141);
nor U17946 (N_17946,N_15065,N_15515);
or U17947 (N_17947,N_16932,N_15962);
or U17948 (N_17948,N_17001,N_17302);
and U17949 (N_17949,N_16253,N_15036);
nor U17950 (N_17950,N_15552,N_15002);
or U17951 (N_17951,N_16301,N_16293);
and U17952 (N_17952,N_15524,N_15193);
nor U17953 (N_17953,N_15407,N_16913);
nand U17954 (N_17954,N_17099,N_16971);
nand U17955 (N_17955,N_17424,N_15719);
nor U17956 (N_17956,N_15307,N_15957);
nor U17957 (N_17957,N_16823,N_15451);
and U17958 (N_17958,N_16688,N_15244);
and U17959 (N_17959,N_15367,N_15319);
xnor U17960 (N_17960,N_17175,N_17321);
or U17961 (N_17961,N_16923,N_16423);
and U17962 (N_17962,N_16740,N_16159);
nand U17963 (N_17963,N_15545,N_15613);
and U17964 (N_17964,N_16245,N_16184);
nand U17965 (N_17965,N_16496,N_16261);
nor U17966 (N_17966,N_15225,N_16621);
or U17967 (N_17967,N_16235,N_15292);
xnor U17968 (N_17968,N_17356,N_15955);
xnor U17969 (N_17969,N_16924,N_16655);
xor U17970 (N_17970,N_17359,N_17124);
nand U17971 (N_17971,N_17271,N_17369);
or U17972 (N_17972,N_15474,N_16333);
or U17973 (N_17973,N_15048,N_17112);
or U17974 (N_17974,N_16952,N_15203);
xor U17975 (N_17975,N_15864,N_15190);
xor U17976 (N_17976,N_17488,N_17241);
nand U17977 (N_17977,N_16489,N_16521);
xnor U17978 (N_17978,N_16259,N_16065);
nor U17979 (N_17979,N_15714,N_15045);
xnor U17980 (N_17980,N_15871,N_15014);
xnor U17981 (N_17981,N_15460,N_15572);
nand U17982 (N_17982,N_15679,N_17370);
nor U17983 (N_17983,N_15064,N_15282);
nand U17984 (N_17984,N_16876,N_17113);
nor U17985 (N_17985,N_15872,N_15107);
xnor U17986 (N_17986,N_16171,N_16035);
and U17987 (N_17987,N_15499,N_15031);
xor U17988 (N_17988,N_16681,N_15866);
and U17989 (N_17989,N_16541,N_15664);
xnor U17990 (N_17990,N_16613,N_15109);
and U17991 (N_17991,N_16230,N_15172);
nor U17992 (N_17992,N_15486,N_16258);
nand U17993 (N_17993,N_16276,N_16075);
or U17994 (N_17994,N_17118,N_15583);
nor U17995 (N_17995,N_17144,N_16487);
xnor U17996 (N_17996,N_17169,N_17062);
or U17997 (N_17997,N_15157,N_15074);
xnor U17998 (N_17998,N_15740,N_16081);
and U17999 (N_17999,N_15393,N_17347);
or U18000 (N_18000,N_15175,N_15764);
and U18001 (N_18001,N_15420,N_15302);
or U18002 (N_18002,N_16574,N_16888);
xnor U18003 (N_18003,N_16849,N_16296);
and U18004 (N_18004,N_17063,N_16197);
and U18005 (N_18005,N_17499,N_15260);
or U18006 (N_18006,N_16418,N_16707);
and U18007 (N_18007,N_15547,N_15554);
nor U18008 (N_18008,N_15463,N_17293);
xnor U18009 (N_18009,N_16163,N_16686);
nand U18010 (N_18010,N_15081,N_15821);
nor U18011 (N_18011,N_16495,N_16056);
or U18012 (N_18012,N_16717,N_15517);
nor U18013 (N_18013,N_16132,N_16373);
nor U18014 (N_18014,N_16039,N_15901);
xor U18015 (N_18015,N_17203,N_17345);
or U18016 (N_18016,N_15294,N_15636);
or U18017 (N_18017,N_17224,N_16625);
or U18018 (N_18018,N_16480,N_15669);
or U18019 (N_18019,N_15869,N_16329);
xor U18020 (N_18020,N_17228,N_17348);
xor U18021 (N_18021,N_15900,N_15996);
xnor U18022 (N_18022,N_16370,N_16762);
or U18023 (N_18023,N_16799,N_17292);
xnor U18024 (N_18024,N_16891,N_15754);
or U18025 (N_18025,N_15528,N_16659);
xor U18026 (N_18026,N_16402,N_17280);
xor U18027 (N_18027,N_15830,N_17052);
xnor U18028 (N_18028,N_16831,N_15015);
nand U18029 (N_18029,N_17388,N_15895);
nor U18030 (N_18030,N_16209,N_15628);
xnor U18031 (N_18031,N_16415,N_16863);
xnor U18032 (N_18032,N_15626,N_16318);
or U18033 (N_18033,N_15092,N_15466);
nand U18034 (N_18034,N_15195,N_15621);
nand U18035 (N_18035,N_17461,N_16000);
or U18036 (N_18036,N_16052,N_16033);
and U18037 (N_18037,N_15530,N_15306);
nand U18038 (N_18038,N_17283,N_15922);
xnor U18039 (N_18039,N_17338,N_17116);
xor U18040 (N_18040,N_16585,N_15897);
nor U18041 (N_18041,N_16723,N_15295);
nand U18042 (N_18042,N_15271,N_16687);
xnor U18043 (N_18043,N_16136,N_17449);
nor U18044 (N_18044,N_15708,N_15032);
nor U18045 (N_18045,N_15335,N_16837);
nand U18046 (N_18046,N_16526,N_16306);
nand U18047 (N_18047,N_16248,N_15057);
nand U18048 (N_18048,N_17365,N_15670);
xor U18049 (N_18049,N_17489,N_15448);
and U18050 (N_18050,N_15275,N_17452);
or U18051 (N_18051,N_17467,N_16054);
xnor U18052 (N_18052,N_15924,N_16592);
nor U18053 (N_18053,N_15205,N_16078);
nand U18054 (N_18054,N_15323,N_15245);
and U18055 (N_18055,N_15587,N_16829);
xnor U18056 (N_18056,N_16722,N_16991);
nand U18057 (N_18057,N_15624,N_16536);
nand U18058 (N_18058,N_15971,N_17104);
and U18059 (N_18059,N_16805,N_15710);
xnor U18060 (N_18060,N_15211,N_15148);
and U18061 (N_18061,N_16427,N_16716);
and U18062 (N_18062,N_15742,N_16766);
and U18063 (N_18063,N_16803,N_17307);
nor U18064 (N_18064,N_16281,N_17039);
nor U18065 (N_18065,N_16591,N_15469);
and U18066 (N_18066,N_15700,N_15655);
nand U18067 (N_18067,N_15725,N_16244);
xnor U18068 (N_18068,N_17479,N_15646);
or U18069 (N_18069,N_17202,N_15168);
or U18070 (N_18070,N_15582,N_15550);
or U18071 (N_18071,N_15951,N_15481);
xor U18072 (N_18072,N_15789,N_16082);
nor U18073 (N_18073,N_15513,N_16360);
and U18074 (N_18074,N_17397,N_15862);
and U18075 (N_18075,N_16702,N_15696);
or U18076 (N_18076,N_15330,N_16651);
and U18077 (N_18077,N_15285,N_15146);
nor U18078 (N_18078,N_15526,N_16425);
xor U18079 (N_18079,N_16582,N_17114);
nand U18080 (N_18080,N_15730,N_15475);
xor U18081 (N_18081,N_16785,N_16024);
nand U18082 (N_18082,N_16836,N_17051);
and U18083 (N_18083,N_17268,N_16315);
or U18084 (N_18084,N_15365,N_15293);
or U18085 (N_18085,N_16590,N_17207);
nand U18086 (N_18086,N_17368,N_15214);
xor U18087 (N_18087,N_15770,N_15766);
nand U18088 (N_18088,N_16960,N_16345);
xnor U18089 (N_18089,N_16859,N_15347);
and U18090 (N_18090,N_15997,N_15620);
and U18091 (N_18091,N_15457,N_17219);
nor U18092 (N_18092,N_16251,N_15461);
or U18093 (N_18093,N_16399,N_16331);
nor U18094 (N_18094,N_16200,N_16461);
xnor U18095 (N_18095,N_17425,N_15555);
nor U18096 (N_18096,N_16584,N_16421);
xnor U18097 (N_18097,N_16727,N_17196);
or U18098 (N_18098,N_16178,N_15385);
nor U18099 (N_18099,N_15929,N_15637);
xnor U18100 (N_18100,N_16693,N_17360);
nor U18101 (N_18101,N_16062,N_16109);
nand U18102 (N_18102,N_17407,N_15220);
nand U18103 (N_18103,N_15176,N_15741);
and U18104 (N_18104,N_15301,N_17056);
nand U18105 (N_18105,N_16685,N_16433);
and U18106 (N_18106,N_16028,N_15631);
or U18107 (N_18107,N_16129,N_17264);
nor U18108 (N_18108,N_17217,N_16445);
nor U18109 (N_18109,N_16083,N_15472);
xor U18110 (N_18110,N_16963,N_15027);
nor U18111 (N_18111,N_15489,N_16649);
nor U18112 (N_18112,N_15373,N_15357);
or U18113 (N_18113,N_17083,N_15281);
or U18114 (N_18114,N_16931,N_15540);
nor U18115 (N_18115,N_15252,N_15815);
nand U18116 (N_18116,N_16089,N_17201);
or U18117 (N_18117,N_17412,N_16453);
or U18118 (N_18118,N_16392,N_15774);
nand U18119 (N_18119,N_15799,N_17285);
and U18120 (N_18120,N_15732,N_15218);
xor U18121 (N_18121,N_16509,N_15606);
and U18122 (N_18122,N_17037,N_16460);
xor U18123 (N_18123,N_16908,N_15154);
nor U18124 (N_18124,N_16734,N_15209);
xnor U18125 (N_18125,N_16486,N_16720);
or U18126 (N_18126,N_17245,N_15314);
xor U18127 (N_18127,N_15017,N_15401);
xor U18128 (N_18128,N_17002,N_15762);
xnor U18129 (N_18129,N_15127,N_16057);
or U18130 (N_18130,N_16534,N_16307);
nand U18131 (N_18131,N_15234,N_15264);
xnor U18132 (N_18132,N_16886,N_16104);
and U18133 (N_18133,N_15825,N_16286);
or U18134 (N_18134,N_16993,N_15504);
nor U18135 (N_18135,N_15384,N_16394);
or U18136 (N_18136,N_15562,N_15128);
or U18137 (N_18137,N_17177,N_16212);
xor U18138 (N_18138,N_16456,N_17105);
and U18139 (N_18139,N_16630,N_16125);
nor U18140 (N_18140,N_15804,N_16472);
nand U18141 (N_18141,N_16498,N_15561);
nand U18142 (N_18142,N_17462,N_15534);
and U18143 (N_18143,N_16866,N_15079);
and U18144 (N_18144,N_15824,N_16216);
nand U18145 (N_18145,N_16544,N_15250);
nand U18146 (N_18146,N_17375,N_15544);
or U18147 (N_18147,N_15818,N_15807);
and U18148 (N_18148,N_16432,N_17495);
or U18149 (N_18149,N_15296,N_15142);
nand U18150 (N_18150,N_16064,N_16494);
xnor U18151 (N_18151,N_16937,N_15147);
nand U18152 (N_18152,N_16587,N_15519);
or U18153 (N_18153,N_15902,N_16614);
nor U18154 (N_18154,N_15877,N_15256);
xnor U18155 (N_18155,N_16941,N_15487);
nand U18156 (N_18156,N_16413,N_16517);
and U18157 (N_18157,N_15263,N_15106);
xor U18158 (N_18158,N_16275,N_15398);
or U18159 (N_18159,N_15060,N_17208);
nor U18160 (N_18160,N_17384,N_17438);
and U18161 (N_18161,N_15622,N_16369);
nand U18162 (N_18162,N_15944,N_15055);
xnor U18163 (N_18163,N_17313,N_15560);
and U18164 (N_18164,N_15216,N_16426);
nor U18165 (N_18165,N_17298,N_16220);
and U18166 (N_18166,N_16428,N_15493);
and U18167 (N_18167,N_17284,N_16260);
xnor U18168 (N_18168,N_16835,N_15870);
nor U18169 (N_18169,N_15000,N_17117);
nor U18170 (N_18170,N_15196,N_15763);
or U18171 (N_18171,N_16463,N_16298);
xor U18172 (N_18172,N_16955,N_16505);
nand U18173 (N_18173,N_16485,N_16282);
and U18174 (N_18174,N_16741,N_16942);
xor U18175 (N_18175,N_17033,N_16926);
nor U18176 (N_18176,N_15806,N_15617);
nand U18177 (N_18177,N_16767,N_15786);
xor U18178 (N_18178,N_17317,N_17460);
nor U18179 (N_18179,N_17140,N_16551);
or U18180 (N_18180,N_15008,N_15536);
or U18181 (N_18181,N_17270,N_16573);
and U18182 (N_18182,N_16817,N_17418);
nor U18183 (N_18183,N_16671,N_15752);
nand U18184 (N_18184,N_16073,N_17273);
and U18185 (N_18185,N_17229,N_15454);
nand U18186 (N_18186,N_15177,N_16580);
or U18187 (N_18187,N_15383,N_15956);
nor U18188 (N_18188,N_16958,N_16153);
nand U18189 (N_18189,N_15605,N_15381);
nand U18190 (N_18190,N_15611,N_16787);
xnor U18191 (N_18191,N_15716,N_15881);
nand U18192 (N_18192,N_17310,N_15797);
nor U18193 (N_18193,N_15403,N_15627);
nor U18194 (N_18194,N_16570,N_17168);
nor U18195 (N_18195,N_16325,N_15249);
and U18196 (N_18196,N_15173,N_16701);
and U18197 (N_18197,N_16096,N_15468);
xnor U18198 (N_18198,N_15846,N_16071);
xor U18199 (N_18199,N_16676,N_17421);
and U18200 (N_18200,N_16186,N_15695);
nand U18201 (N_18201,N_16806,N_16779);
nand U18202 (N_18202,N_16957,N_15574);
or U18203 (N_18203,N_16195,N_15210);
and U18204 (N_18204,N_16915,N_15419);
nor U18205 (N_18205,N_15985,N_16936);
nand U18206 (N_18206,N_15570,N_16523);
and U18207 (N_18207,N_16170,N_16552);
nor U18208 (N_18208,N_15051,N_16443);
nand U18209 (N_18209,N_17457,N_16344);
and U18210 (N_18210,N_16636,N_16243);
and U18211 (N_18211,N_16798,N_15369);
nor U18212 (N_18212,N_15640,N_16458);
or U18213 (N_18213,N_15087,N_15551);
xnor U18214 (N_18214,N_15492,N_16148);
and U18215 (N_18215,N_16889,N_16543);
nor U18216 (N_18216,N_17074,N_17289);
or U18217 (N_18217,N_15908,N_17322);
nand U18218 (N_18218,N_16719,N_15233);
nor U18219 (N_18219,N_17094,N_16106);
nor U18220 (N_18220,N_16739,N_15120);
nor U18221 (N_18221,N_17125,N_16698);
and U18222 (N_18222,N_16268,N_16327);
nand U18223 (N_18223,N_16546,N_17274);
or U18224 (N_18224,N_16531,N_15030);
or U18225 (N_18225,N_16098,N_17253);
nor U18226 (N_18226,N_15947,N_16295);
nand U18227 (N_18227,N_15313,N_15498);
or U18228 (N_18228,N_15399,N_16192);
nor U18229 (N_18229,N_15662,N_17109);
nand U18230 (N_18230,N_16374,N_16446);
nor U18231 (N_18231,N_15364,N_17405);
nand U18232 (N_18232,N_15199,N_15268);
nor U18233 (N_18233,N_15659,N_15054);
nor U18234 (N_18234,N_16322,N_15409);
or U18235 (N_18235,N_17252,N_16092);
or U18236 (N_18236,N_17178,N_16645);
nand U18237 (N_18237,N_16198,N_16665);
nor U18238 (N_18238,N_15687,N_16464);
or U18239 (N_18239,N_17393,N_16673);
nand U18240 (N_18240,N_17455,N_15832);
nand U18241 (N_18241,N_16323,N_16469);
nor U18242 (N_18242,N_15080,N_15848);
or U18243 (N_18243,N_16471,N_17484);
and U18244 (N_18244,N_16846,N_15857);
xnor U18245 (N_18245,N_15152,N_16780);
nand U18246 (N_18246,N_15891,N_15803);
nor U18247 (N_18247,N_16255,N_16043);
xor U18248 (N_18248,N_16084,N_16980);
or U18249 (N_18249,N_17432,N_16450);
or U18250 (N_18250,N_16262,N_16597);
nand U18251 (N_18251,N_16139,N_15354);
and U18252 (N_18252,N_15059,N_15186);
nor U18253 (N_18253,N_16811,N_16710);
or U18254 (N_18254,N_17334,N_15110);
or U18255 (N_18255,N_15980,N_17378);
xnor U18256 (N_18256,N_17248,N_15632);
nand U18257 (N_18257,N_17076,N_17394);
nor U18258 (N_18258,N_16555,N_17403);
xor U18259 (N_18259,N_15946,N_15916);
nand U18260 (N_18260,N_15001,N_15836);
or U18261 (N_18261,N_16670,N_17377);
nand U18262 (N_18262,N_15284,N_15817);
or U18263 (N_18263,N_15290,N_16895);
nand U18264 (N_18264,N_16291,N_16504);
nor U18265 (N_18265,N_15509,N_16996);
and U18266 (N_18266,N_16518,N_15095);
and U18267 (N_18267,N_16511,N_15348);
or U18268 (N_18268,N_15822,N_15072);
xnor U18269 (N_18269,N_15097,N_16628);
nor U18270 (N_18270,N_17025,N_16843);
or U18271 (N_18271,N_15188,N_17250);
nand U18272 (N_18272,N_15180,N_16340);
xor U18273 (N_18273,N_16667,N_16755);
xnor U18274 (N_18274,N_17410,N_15038);
and U18275 (N_18275,N_15873,N_16203);
xnor U18276 (N_18276,N_17089,N_15874);
nand U18277 (N_18277,N_16822,N_17486);
or U18278 (N_18278,N_15717,N_16311);
xor U18279 (N_18279,N_16769,N_17107);
nand U18280 (N_18280,N_15643,N_16409);
nand U18281 (N_18281,N_16632,N_15715);
or U18282 (N_18282,N_17297,N_15444);
xnor U18283 (N_18283,N_17318,N_15178);
or U18284 (N_18284,N_16746,N_16847);
or U18285 (N_18285,N_15056,N_17130);
nand U18286 (N_18286,N_17154,N_15198);
or U18287 (N_18287,N_16879,N_15343);
and U18288 (N_18288,N_15445,N_15411);
and U18289 (N_18289,N_15039,N_17391);
nand U18290 (N_18290,N_15521,N_16214);
nand U18291 (N_18291,N_16023,N_17386);
and U18292 (N_18292,N_16206,N_17487);
nor U18293 (N_18293,N_17195,N_15795);
xor U18294 (N_18294,N_16808,N_16123);
nand U18295 (N_18295,N_16773,N_17179);
or U18296 (N_18296,N_16982,N_15421);
xnor U18297 (N_18297,N_15674,N_15723);
nor U18298 (N_18298,N_15482,N_15267);
and U18299 (N_18299,N_15494,N_15653);
and U18300 (N_18300,N_16576,N_16965);
or U18301 (N_18301,N_16007,N_15346);
xnor U18302 (N_18302,N_16016,N_17087);
nor U18303 (N_18303,N_15940,N_15400);
xnor U18304 (N_18304,N_16330,N_17352);
xor U18305 (N_18305,N_15918,N_15656);
and U18306 (N_18306,N_16770,N_15288);
nor U18307 (N_18307,N_17213,N_15025);
xor U18308 (N_18308,N_16867,N_17182);
nand U18309 (N_18309,N_16986,N_17209);
and U18310 (N_18310,N_15984,N_15532);
nor U18311 (N_18311,N_17385,N_15336);
xor U18312 (N_18312,N_15828,N_16664);
or U18313 (N_18313,N_15704,N_16611);
and U18314 (N_18314,N_17128,N_16481);
or U18315 (N_18315,N_15511,N_16669);
nor U18316 (N_18316,N_16821,N_15702);
nor U18317 (N_18317,N_15814,N_17240);
and U18318 (N_18318,N_15919,N_15915);
and U18319 (N_18319,N_17000,N_16500);
nor U18320 (N_18320,N_17078,N_17026);
or U18321 (N_18321,N_17100,N_17333);
nor U18322 (N_18322,N_16328,N_17451);
xor U18323 (N_18323,N_15459,N_15868);
or U18324 (N_18324,N_15720,N_15801);
or U18325 (N_18325,N_15569,N_16515);
xor U18326 (N_18326,N_17339,N_16349);
nor U18327 (N_18327,N_15553,N_15426);
nor U18328 (N_18328,N_16692,N_15834);
xor U18329 (N_18329,N_16050,N_15706);
and U18330 (N_18330,N_17032,N_15166);
and U18331 (N_18331,N_16068,N_15781);
xnor U18332 (N_18332,N_16199,N_17335);
nand U18333 (N_18333,N_15328,N_16588);
nand U18334 (N_18334,N_15035,N_17493);
and U18335 (N_18335,N_17072,N_15721);
nand U18336 (N_18336,N_15104,N_15418);
nor U18337 (N_18337,N_16539,N_17184);
xnor U18338 (N_18338,N_17238,N_16242);
and U18339 (N_18339,N_16917,N_15053);
nand U18340 (N_18340,N_16215,N_17319);
nand U18341 (N_18341,N_15387,N_16838);
xor U18342 (N_18342,N_16434,N_16272);
nand U18343 (N_18343,N_16466,N_17258);
nand U18344 (N_18344,N_15738,N_16976);
xnor U18345 (N_18345,N_16771,N_15139);
and U18346 (N_18346,N_15647,N_16801);
nand U18347 (N_18347,N_16564,N_17366);
nand U18348 (N_18348,N_17408,N_16483);
nor U18349 (N_18349,N_16985,N_17097);
or U18350 (N_18350,N_15701,N_16221);
xnor U18351 (N_18351,N_15675,N_15543);
and U18352 (N_18352,N_16782,N_16090);
xnor U18353 (N_18353,N_15694,N_16950);
nor U18354 (N_18354,N_16639,N_15395);
or U18355 (N_18355,N_16122,N_16173);
or U18356 (N_18356,N_17036,N_15733);
nor U18357 (N_18357,N_15644,N_15404);
nor U18358 (N_18358,N_17354,N_17372);
xor U18359 (N_18359,N_15712,N_16047);
nor U18360 (N_18360,N_16529,N_16474);
nor U18361 (N_18361,N_17015,N_16612);
nand U18362 (N_18362,N_17167,N_17463);
xor U18363 (N_18363,N_15473,N_17276);
nor U18364 (N_18364,N_15860,N_15428);
xnor U18365 (N_18365,N_16390,N_16380);
nand U18366 (N_18366,N_15119,N_16391);
or U18367 (N_18367,N_16217,N_15162);
nor U18368 (N_18368,N_15135,N_17400);
and U18369 (N_18369,N_15402,N_16759);
nand U18370 (N_18370,N_16385,N_17092);
nor U18371 (N_18371,N_17340,N_15748);
and U18372 (N_18372,N_15595,N_15529);
and U18373 (N_18373,N_16451,N_16516);
xnor U18374 (N_18374,N_16303,N_16006);
and U18375 (N_18375,N_16906,N_16015);
nand U18376 (N_18376,N_16873,N_17447);
and U18377 (N_18377,N_17436,N_15046);
and U18378 (N_18378,N_15615,N_16300);
nor U18379 (N_18379,N_16951,N_15522);
nor U18380 (N_18380,N_16027,N_15729);
nor U18381 (N_18381,N_16858,N_16995);
nand U18382 (N_18382,N_15300,N_16118);
and U18383 (N_18383,N_16606,N_16326);
xnor U18384 (N_18384,N_15308,N_15735);
or U18385 (N_18385,N_16964,N_16219);
nand U18386 (N_18386,N_15298,N_16832);
nor U18387 (N_18387,N_16019,N_16545);
xor U18388 (N_18388,N_15134,N_16302);
and U18389 (N_18389,N_16566,N_15350);
xor U18390 (N_18390,N_15707,N_15989);
and U18391 (N_18391,N_16788,N_15063);
nand U18392 (N_18392,N_16962,N_16367);
and U18393 (N_18393,N_16728,N_15113);
and U18394 (N_18394,N_16100,N_15026);
nand U18395 (N_18395,N_17401,N_16497);
and U18396 (N_18396,N_17134,N_16020);
or U18397 (N_18397,N_17166,N_15673);
xnor U18398 (N_18398,N_15247,N_15539);
and U18399 (N_18399,N_15651,N_15412);
and U18400 (N_18400,N_17019,N_17470);
xor U18401 (N_18401,N_15578,N_16051);
nor U18402 (N_18402,N_15246,N_16151);
nand U18403 (N_18403,N_16448,N_15020);
nor U18404 (N_18404,N_15423,N_16675);
nand U18405 (N_18405,N_15366,N_15884);
xor U18406 (N_18406,N_15589,N_15286);
or U18407 (N_18407,N_17215,N_17189);
or U18408 (N_18408,N_15809,N_15782);
and U18409 (N_18409,N_15926,N_16530);
nor U18410 (N_18410,N_16134,N_16208);
nor U18411 (N_18411,N_16411,N_17373);
and U18412 (N_18412,N_16861,N_15531);
and U18413 (N_18413,N_15429,N_15629);
nand U18414 (N_18414,N_16712,N_17216);
xnor U18415 (N_18415,N_16429,N_16061);
and U18416 (N_18416,N_17048,N_17014);
and U18417 (N_18417,N_15310,N_16058);
xnor U18418 (N_18418,N_15237,N_16124);
or U18419 (N_18419,N_15185,N_17197);
nor U18420 (N_18420,N_16706,N_15316);
and U18421 (N_18421,N_16299,N_15270);
xor U18422 (N_18422,N_16730,N_15331);
nand U18423 (N_18423,N_15133,N_15242);
nor U18424 (N_18424,N_16905,N_16352);
nand U18425 (N_18425,N_15502,N_15279);
nand U18426 (N_18426,N_17414,N_17341);
nand U18427 (N_18427,N_15894,N_15377);
or U18428 (N_18428,N_15248,N_16826);
nand U18429 (N_18429,N_16101,N_16080);
and U18430 (N_18430,N_16646,N_16187);
xnor U18431 (N_18431,N_16928,N_16194);
xor U18432 (N_18432,N_15759,N_16249);
xor U18433 (N_18433,N_16560,N_16624);
or U18434 (N_18434,N_16099,N_16395);
nor U18435 (N_18435,N_16133,N_15440);
xor U18436 (N_18436,N_16977,N_15746);
and U18437 (N_18437,N_15086,N_16224);
nand U18438 (N_18438,N_15925,N_16274);
xor U18439 (N_18439,N_15396,N_15274);
nand U18440 (N_18440,N_16668,N_16816);
and U18441 (N_18441,N_16088,N_16713);
nand U18442 (N_18442,N_15483,N_17102);
and U18443 (N_18443,N_15450,N_15652);
nand U18444 (N_18444,N_16372,N_17272);
and U18445 (N_18445,N_17110,N_16297);
nand U18446 (N_18446,N_16484,N_16997);
xnor U18447 (N_18447,N_16188,N_15614);
nand U18448 (N_18448,N_16356,N_15579);
nor U18449 (N_18449,N_15363,N_16506);
and U18450 (N_18450,N_16579,N_17145);
xnor U18451 (N_18451,N_17416,N_15541);
or U18452 (N_18452,N_15066,N_15360);
xor U18453 (N_18453,N_15370,N_15598);
nand U18454 (N_18454,N_15374,N_15993);
or U18455 (N_18455,N_16146,N_17406);
or U18456 (N_18456,N_16363,N_16401);
nor U18457 (N_18457,N_15969,N_16894);
or U18458 (N_18458,N_15557,N_15728);
nand U18459 (N_18459,N_16436,N_15612);
or U18460 (N_18460,N_15964,N_17294);
nand U18461 (N_18461,N_15777,N_16074);
nand U18462 (N_18462,N_16572,N_15141);
and U18463 (N_18463,N_16161,N_17249);
and U18464 (N_18464,N_17108,N_16444);
and U18465 (N_18465,N_16149,N_15151);
and U18466 (N_18466,N_15170,N_15839);
nand U18467 (N_18467,N_16169,N_17291);
or U18468 (N_18468,N_15253,N_17009);
nor U18469 (N_18469,N_16131,N_17477);
xor U18470 (N_18470,N_16914,N_16454);
xnor U18471 (N_18471,N_17330,N_16040);
or U18472 (N_18472,N_15137,N_17468);
nand U18473 (N_18473,N_16796,N_16266);
nand U18474 (N_18474,N_16884,N_16586);
nor U18475 (N_18475,N_15564,N_16503);
and U18476 (N_18476,N_15276,N_16841);
nor U18477 (N_18477,N_15973,N_15197);
nor U18478 (N_18478,N_17450,N_15050);
nor U18479 (N_18479,N_16308,N_15575);
nand U18480 (N_18480,N_15070,N_15116);
nand U18481 (N_18481,N_16112,N_17257);
and U18482 (N_18482,N_16758,N_17190);
or U18483 (N_18483,N_15785,N_16933);
or U18484 (N_18484,N_15465,N_16608);
or U18485 (N_18485,N_15888,N_15043);
nand U18486 (N_18486,N_16182,N_15342);
nand U18487 (N_18487,N_16113,N_15849);
nand U18488 (N_18488,N_15130,N_15228);
nand U18489 (N_18489,N_15408,N_16292);
or U18490 (N_18490,N_16820,N_16231);
nor U18491 (N_18491,N_16860,N_15790);
or U18492 (N_18492,N_17165,N_15920);
xnor U18493 (N_18493,N_16107,N_15577);
and U18494 (N_18494,N_16729,N_17234);
nor U18495 (N_18495,N_16802,N_16191);
nor U18496 (N_18496,N_15727,N_15665);
or U18497 (N_18497,N_16943,N_16180);
or U18498 (N_18498,N_15960,N_15798);
or U18499 (N_18499,N_16622,N_17311);
xnor U18500 (N_18500,N_17066,N_16142);
and U18501 (N_18501,N_17265,N_16095);
or U18502 (N_18502,N_16332,N_17088);
nand U18503 (N_18503,N_15047,N_16181);
xnor U18504 (N_18504,N_17398,N_15686);
or U18505 (N_18505,N_17024,N_16896);
and U18506 (N_18506,N_16396,N_16947);
and U18507 (N_18507,N_16562,N_16398);
and U18508 (N_18508,N_16781,N_17135);
nand U18509 (N_18509,N_17236,N_16850);
xnor U18510 (N_18510,N_16865,N_15930);
nor U18511 (N_18511,N_16778,N_16898);
or U18512 (N_18512,N_15808,N_15490);
xnor U18513 (N_18513,N_16616,N_17065);
nor U18514 (N_18514,N_15990,N_15155);
nor U18515 (N_18515,N_15439,N_15645);
nor U18516 (N_18516,N_16252,N_17256);
or U18517 (N_18517,N_15697,N_15372);
xor U18518 (N_18518,N_15012,N_17211);
nor U18519 (N_18519,N_15003,N_17187);
nand U18520 (N_18520,N_15937,N_16005);
nand U18521 (N_18521,N_15907,N_15802);
xor U18522 (N_18522,N_17306,N_15320);
and U18523 (N_18523,N_15769,N_16864);
nor U18524 (N_18524,N_15356,N_16108);
nor U18525 (N_18525,N_16956,N_17387);
nand U18526 (N_18526,N_17059,N_15241);
xor U18527 (N_18527,N_15796,N_16384);
nand U18528 (N_18528,N_16233,N_17262);
and U18529 (N_18529,N_15265,N_17399);
or U18530 (N_18530,N_17142,N_16087);
nand U18531 (N_18531,N_16528,N_16527);
nor U18532 (N_18532,N_17471,N_16825);
and U18533 (N_18533,N_15743,N_15150);
xnor U18534 (N_18534,N_15935,N_17221);
and U18535 (N_18535,N_17315,N_16680);
or U18536 (N_18536,N_15680,N_17290);
nand U18537 (N_18537,N_15167,N_16810);
nor U18538 (N_18538,N_15506,N_17459);
nor U18539 (N_18539,N_15433,N_16842);
or U18540 (N_18540,N_17156,N_15159);
nand U18541 (N_18541,N_15503,N_17075);
nor U18542 (N_18542,N_17281,N_15875);
nor U18543 (N_18543,N_16110,N_15994);
nor U18544 (N_18544,N_16631,N_16916);
or U18545 (N_18545,N_15226,N_15501);
and U18546 (N_18546,N_16938,N_15672);
xnor U18547 (N_18547,N_16620,N_17218);
xor U18548 (N_18548,N_16270,N_15858);
nor U18549 (N_18549,N_16998,N_17155);
or U18550 (N_18550,N_15590,N_16177);
nor U18551 (N_18551,N_16618,N_16222);
nand U18552 (N_18552,N_15833,N_15558);
and U18553 (N_18553,N_17005,N_15338);
xnor U18554 (N_18554,N_16117,N_16478);
or U18555 (N_18555,N_17069,N_16288);
or U18556 (N_18556,N_15596,N_15217);
nor U18557 (N_18557,N_16791,N_16828);
nor U18558 (N_18558,N_16626,N_16128);
or U18559 (N_18559,N_15362,N_15780);
nor U18560 (N_18560,N_15132,N_16470);
xor U18561 (N_18561,N_15991,N_16003);
and U18562 (N_18562,N_15083,N_17008);
and U18563 (N_18563,N_17085,N_16754);
and U18564 (N_18564,N_16038,N_15883);
and U18565 (N_18565,N_15229,N_17232);
nand U18566 (N_18566,N_16575,N_17422);
or U18567 (N_18567,N_17465,N_17420);
nor U18568 (N_18568,N_16656,N_15187);
nand U18569 (N_18569,N_17035,N_16683);
nor U18570 (N_18570,N_15102,N_15791);
and U18571 (N_18571,N_15981,N_15075);
or U18572 (N_18572,N_16660,N_16658);
xor U18573 (N_18573,N_17067,N_17485);
xor U18574 (N_18574,N_16902,N_16909);
nor U18575 (N_18575,N_15158,N_16897);
or U18576 (N_18576,N_16911,N_16376);
and U18577 (N_18577,N_17161,N_15449);
xor U18578 (N_18578,N_17139,N_16105);
nand U18579 (N_18579,N_16910,N_17496);
nand U18580 (N_18580,N_17287,N_16018);
nor U18581 (N_18581,N_15823,N_16001);
nand U18582 (N_18582,N_17172,N_16176);
nor U18583 (N_18583,N_16653,N_17103);
nand U18584 (N_18584,N_15805,N_17304);
or U18585 (N_18585,N_17260,N_16152);
or U18586 (N_18586,N_17034,N_15843);
nand U18587 (N_18587,N_15011,N_17404);
and U18588 (N_18588,N_16892,N_15941);
or U18589 (N_18589,N_16350,N_17171);
or U18590 (N_18590,N_15184,N_15345);
or U18591 (N_18591,N_17205,N_16174);
xor U18592 (N_18592,N_15441,N_17351);
and U18593 (N_18593,N_15813,N_16725);
xor U18594 (N_18594,N_16994,N_17023);
and U18595 (N_18595,N_16145,N_15124);
and U18596 (N_18596,N_15563,N_17396);
or U18597 (N_18597,N_15006,N_15480);
nor U18598 (N_18598,N_16601,N_16708);
xnor U18599 (N_18599,N_16103,N_15639);
and U18600 (N_18600,N_15436,N_15887);
nor U18601 (N_18601,N_15783,N_16294);
or U18602 (N_18602,N_17342,N_15380);
xor U18603 (N_18603,N_16343,N_17119);
and U18604 (N_18604,N_16856,N_16940);
and U18605 (N_18605,N_16452,N_17111);
nand U18606 (N_18606,N_15633,N_15129);
or U18607 (N_18607,N_17020,N_16677);
nor U18608 (N_18608,N_17402,N_16267);
nor U18609 (N_18609,N_15156,N_15638);
xnor U18610 (N_18610,N_16872,N_17080);
or U18611 (N_18611,N_15691,N_17237);
and U18612 (N_18612,N_15491,N_15608);
nand U18613 (N_18613,N_15566,N_16324);
nor U18614 (N_18614,N_15567,N_16901);
nor U18615 (N_18615,N_17158,N_16804);
or U18616 (N_18616,N_17282,N_15287);
and U18617 (N_18617,N_16920,N_15208);
and U18618 (N_18618,N_16696,N_15961);
nor U18619 (N_18619,N_16059,N_16403);
or U18620 (N_18620,N_16794,N_15425);
nor U18621 (N_18621,N_16784,N_16684);
and U18622 (N_18622,N_15317,N_15202);
and U18623 (N_18623,N_16422,N_15537);
nand U18624 (N_18624,N_15470,N_15573);
nor U18625 (N_18625,N_15076,N_17031);
or U18626 (N_18626,N_17151,N_15179);
nand U18627 (N_18627,N_17441,N_16557);
or U18628 (N_18628,N_16357,N_15028);
or U18629 (N_18629,N_16753,N_16870);
nor U18630 (N_18630,N_15182,N_15477);
and U18631 (N_18631,N_16533,N_16172);
nand U18632 (N_18632,N_15438,N_17170);
and U18633 (N_18633,N_15332,N_15923);
xnor U18634 (N_18634,N_15938,N_16925);
nand U18635 (N_18635,N_17492,N_16273);
nand U18636 (N_18636,N_15118,N_17473);
nor U18637 (N_18637,N_15280,N_15698);
and U18638 (N_18638,N_16627,N_15098);
and U18639 (N_18639,N_16069,N_15692);
nor U18640 (N_18640,N_16567,N_16975);
or U18641 (N_18641,N_16202,N_16437);
or U18642 (N_18642,N_17332,N_17367);
nand U18643 (N_18643,N_16240,N_16002);
and U18644 (N_18644,N_16037,N_17426);
and U18645 (N_18645,N_16578,N_17096);
and U18646 (N_18646,N_15304,N_17316);
nand U18647 (N_18647,N_16721,N_16477);
nor U18648 (N_18648,N_16878,N_16830);
xor U18649 (N_18649,N_16264,N_15340);
or U18650 (N_18650,N_15297,N_16468);
xor U18651 (N_18651,N_15315,N_16877);
xnor U18652 (N_18652,N_15827,N_16320);
xnor U18653 (N_18653,N_15052,N_15222);
nand U18654 (N_18654,N_15042,N_16234);
xor U18655 (N_18655,N_17164,N_16871);
and U18656 (N_18656,N_15745,N_16070);
xnor U18657 (N_18657,N_15126,N_17010);
xnor U18658 (N_18658,N_15010,N_17254);
and U18659 (N_18659,N_15089,N_15224);
nor U18660 (N_18660,N_15013,N_15272);
or U18661 (N_18661,N_17044,N_16921);
xnor U18662 (N_18662,N_15879,N_17127);
or U18663 (N_18663,N_16414,N_17131);
nand U18664 (N_18664,N_17442,N_15850);
xor U18665 (N_18665,N_15535,N_17326);
nand U18666 (N_18666,N_15410,N_17235);
nor U18667 (N_18667,N_16408,N_15775);
xor U18668 (N_18668,N_15022,N_16036);
nor U18669 (N_18669,N_17136,N_16063);
or U18670 (N_18670,N_16619,N_16201);
xnor U18671 (N_18671,N_17137,N_16694);
or U18672 (N_18672,N_16366,N_16381);
or U18673 (N_18673,N_16447,N_16583);
or U18674 (N_18674,N_16672,N_17263);
nand U18675 (N_18675,N_15508,N_15337);
xor U18676 (N_18676,N_15750,N_16379);
and U18677 (N_18677,N_16034,N_15755);
nand U18678 (N_18678,N_15145,N_17337);
xor U18679 (N_18679,N_16375,N_15928);
nor U18680 (N_18680,N_17343,N_15093);
nand U18681 (N_18681,N_16944,N_15518);
nand U18682 (N_18682,N_16501,N_17269);
nor U18683 (N_18683,N_16674,N_15415);
xnor U18684 (N_18684,N_15592,N_15114);
nand U18685 (N_18685,N_17314,N_15945);
nor U18686 (N_18686,N_15603,N_15329);
nor U18687 (N_18687,N_17095,N_17376);
nor U18688 (N_18688,N_15882,N_15965);
and U18689 (N_18689,N_15327,N_16254);
and U18690 (N_18690,N_15982,N_15591);
nand U18691 (N_18691,N_17122,N_17192);
nand U18692 (N_18692,N_16271,N_17371);
and U18693 (N_18693,N_16967,N_17498);
nor U18694 (N_18694,N_15559,N_15949);
xor U18695 (N_18695,N_16939,N_15007);
nand U18696 (N_18696,N_15932,N_15326);
and U18697 (N_18697,N_15903,N_15034);
nand U18698 (N_18698,N_16491,N_15718);
xor U18699 (N_18699,N_17329,N_16705);
xnor U18700 (N_18700,N_15024,N_17225);
or U18701 (N_18701,N_15619,N_15975);
and U18702 (N_18702,N_16900,N_16634);
nor U18703 (N_18703,N_15115,N_17040);
nor U18704 (N_18704,N_16535,N_17247);
nand U18705 (N_18705,N_17200,N_16238);
and U18706 (N_18706,N_15703,N_16777);
nor U18707 (N_18707,N_16189,N_15073);
nor U18708 (N_18708,N_15389,N_15671);
xnor U18709 (N_18709,N_17060,N_17041);
xnor U18710 (N_18710,N_17206,N_15171);
xnor U18711 (N_18711,N_15776,N_16793);
xor U18712 (N_18712,N_16691,N_16682);
nor U18713 (N_18713,N_16750,N_15711);
nor U18714 (N_18714,N_15667,N_16726);
xnor U18715 (N_18715,N_17242,N_15085);
or U18716 (N_18716,N_16652,N_17261);
and U18717 (N_18717,N_15751,N_15616);
xor U18718 (N_18718,N_16969,N_17193);
nor U18719 (N_18719,N_16140,N_15921);
and U18720 (N_18720,N_17029,N_16030);
or U18721 (N_18721,N_15831,N_17233);
xnor U18722 (N_18722,N_15974,N_16783);
xnor U18723 (N_18723,N_16711,N_15549);
or U18724 (N_18724,N_16899,N_15019);
xnor U18725 (N_18725,N_16738,N_16615);
nor U18726 (N_18726,N_17429,N_16044);
nor U18727 (N_18727,N_16337,N_17049);
and U18728 (N_18728,N_15413,N_16041);
and U18729 (N_18729,N_15586,N_16424);
xnor U18730 (N_18730,N_17061,N_17323);
nor U18731 (N_18731,N_15405,N_16190);
and U18732 (N_18732,N_15388,N_16223);
or U18733 (N_18733,N_15693,N_17226);
or U18734 (N_18734,N_16554,N_15500);
or U18735 (N_18735,N_15311,N_17344);
xnor U18736 (N_18736,N_17223,N_17431);
nor U18737 (N_18737,N_15889,N_15682);
nand U18738 (N_18738,N_16733,N_15816);
xor U18739 (N_18739,N_16663,N_17389);
or U18740 (N_18740,N_15910,N_16538);
or U18741 (N_18741,N_15378,N_15507);
or U18742 (N_18742,N_15029,N_17411);
and U18743 (N_18743,N_16488,N_16438);
nand U18744 (N_18744,N_15959,N_16547);
and U18745 (N_18745,N_16196,N_15163);
or U18746 (N_18746,N_16166,N_16225);
nand U18747 (N_18747,N_16085,N_16093);
or U18748 (N_18748,N_15514,N_17336);
xnor U18749 (N_18749,N_15584,N_16365);
or U18750 (N_18750,N_15983,N_16857);
nor U18751 (N_18751,N_17325,N_17458);
or U18752 (N_18752,N_17384,N_16591);
xnor U18753 (N_18753,N_15960,N_17158);
xor U18754 (N_18754,N_15267,N_15094);
or U18755 (N_18755,N_15614,N_15205);
and U18756 (N_18756,N_17496,N_16426);
xor U18757 (N_18757,N_15055,N_17048);
xnor U18758 (N_18758,N_16886,N_16652);
xor U18759 (N_18759,N_16526,N_16440);
and U18760 (N_18760,N_17310,N_17291);
and U18761 (N_18761,N_16027,N_16813);
nand U18762 (N_18762,N_16893,N_16639);
nand U18763 (N_18763,N_16006,N_17271);
xnor U18764 (N_18764,N_17411,N_15448);
and U18765 (N_18765,N_16083,N_16630);
and U18766 (N_18766,N_17441,N_17230);
nand U18767 (N_18767,N_17073,N_16784);
nand U18768 (N_18768,N_15356,N_15088);
nor U18769 (N_18769,N_15232,N_15178);
xor U18770 (N_18770,N_15142,N_15131);
xor U18771 (N_18771,N_15908,N_15663);
nand U18772 (N_18772,N_17215,N_15004);
and U18773 (N_18773,N_16453,N_16296);
nand U18774 (N_18774,N_16824,N_16891);
nand U18775 (N_18775,N_15103,N_16362);
xnor U18776 (N_18776,N_16840,N_17196);
or U18777 (N_18777,N_15604,N_15583);
xor U18778 (N_18778,N_15327,N_15269);
nor U18779 (N_18779,N_15516,N_15526);
nand U18780 (N_18780,N_15970,N_16730);
xnor U18781 (N_18781,N_15568,N_17316);
xnor U18782 (N_18782,N_17389,N_17475);
xnor U18783 (N_18783,N_16828,N_16180);
or U18784 (N_18784,N_15173,N_16273);
xnor U18785 (N_18785,N_16861,N_16505);
nand U18786 (N_18786,N_17423,N_16904);
and U18787 (N_18787,N_15149,N_16343);
xor U18788 (N_18788,N_15946,N_15422);
or U18789 (N_18789,N_15766,N_15063);
nor U18790 (N_18790,N_16507,N_15313);
nand U18791 (N_18791,N_16160,N_16858);
nor U18792 (N_18792,N_16096,N_17235);
and U18793 (N_18793,N_16029,N_16957);
and U18794 (N_18794,N_15122,N_15250);
or U18795 (N_18795,N_16724,N_15042);
or U18796 (N_18796,N_16190,N_15815);
nand U18797 (N_18797,N_16175,N_15570);
and U18798 (N_18798,N_15147,N_15967);
nand U18799 (N_18799,N_16447,N_15301);
nand U18800 (N_18800,N_17134,N_15689);
or U18801 (N_18801,N_15399,N_16677);
nor U18802 (N_18802,N_15178,N_15978);
and U18803 (N_18803,N_16099,N_15895);
or U18804 (N_18804,N_16506,N_16246);
and U18805 (N_18805,N_16982,N_16037);
and U18806 (N_18806,N_15690,N_15034);
nand U18807 (N_18807,N_16785,N_16469);
or U18808 (N_18808,N_16670,N_15173);
nand U18809 (N_18809,N_15052,N_17101);
nand U18810 (N_18810,N_17080,N_15462);
or U18811 (N_18811,N_17389,N_16863);
xnor U18812 (N_18812,N_15957,N_16942);
and U18813 (N_18813,N_16139,N_17145);
and U18814 (N_18814,N_16941,N_15475);
nor U18815 (N_18815,N_15321,N_15421);
nand U18816 (N_18816,N_15594,N_16729);
nor U18817 (N_18817,N_15132,N_15057);
xnor U18818 (N_18818,N_17194,N_16500);
and U18819 (N_18819,N_15148,N_16858);
nor U18820 (N_18820,N_16999,N_17162);
nor U18821 (N_18821,N_17385,N_16999);
nand U18822 (N_18822,N_15489,N_17366);
nand U18823 (N_18823,N_17499,N_15848);
nand U18824 (N_18824,N_16028,N_16541);
xnor U18825 (N_18825,N_15927,N_15164);
and U18826 (N_18826,N_16966,N_15962);
and U18827 (N_18827,N_15425,N_16133);
xor U18828 (N_18828,N_17387,N_17175);
or U18829 (N_18829,N_16783,N_16310);
nand U18830 (N_18830,N_16602,N_17451);
and U18831 (N_18831,N_15145,N_16710);
nand U18832 (N_18832,N_16727,N_15264);
and U18833 (N_18833,N_17007,N_15192);
nand U18834 (N_18834,N_17231,N_17433);
nor U18835 (N_18835,N_16677,N_15772);
and U18836 (N_18836,N_16177,N_17384);
and U18837 (N_18837,N_15509,N_15613);
and U18838 (N_18838,N_15150,N_15052);
nand U18839 (N_18839,N_16810,N_15058);
nand U18840 (N_18840,N_15359,N_16989);
and U18841 (N_18841,N_17361,N_16076);
xnor U18842 (N_18842,N_16137,N_16579);
or U18843 (N_18843,N_16398,N_17391);
or U18844 (N_18844,N_15903,N_16108);
or U18845 (N_18845,N_16963,N_17324);
nor U18846 (N_18846,N_17152,N_15374);
and U18847 (N_18847,N_17341,N_15364);
xnor U18848 (N_18848,N_15795,N_16190);
or U18849 (N_18849,N_15908,N_16975);
nor U18850 (N_18850,N_16471,N_16344);
nand U18851 (N_18851,N_17320,N_15661);
xor U18852 (N_18852,N_16925,N_15544);
nand U18853 (N_18853,N_15937,N_16269);
or U18854 (N_18854,N_16808,N_16893);
nand U18855 (N_18855,N_16121,N_15757);
and U18856 (N_18856,N_16009,N_15673);
and U18857 (N_18857,N_15254,N_15278);
xor U18858 (N_18858,N_16990,N_16921);
or U18859 (N_18859,N_16628,N_15971);
or U18860 (N_18860,N_15940,N_15964);
xor U18861 (N_18861,N_15982,N_16478);
xor U18862 (N_18862,N_16165,N_15106);
and U18863 (N_18863,N_17259,N_17021);
or U18864 (N_18864,N_16556,N_17186);
nor U18865 (N_18865,N_16114,N_16329);
nor U18866 (N_18866,N_16863,N_15340);
or U18867 (N_18867,N_16953,N_15871);
nand U18868 (N_18868,N_17063,N_15139);
xor U18869 (N_18869,N_15490,N_15684);
and U18870 (N_18870,N_15006,N_15670);
nor U18871 (N_18871,N_17333,N_16855);
xor U18872 (N_18872,N_16900,N_17238);
or U18873 (N_18873,N_16220,N_16185);
nor U18874 (N_18874,N_15405,N_16623);
nand U18875 (N_18875,N_15267,N_15027);
nand U18876 (N_18876,N_17260,N_15692);
nand U18877 (N_18877,N_17368,N_17355);
nand U18878 (N_18878,N_15987,N_16561);
nand U18879 (N_18879,N_16930,N_15318);
nor U18880 (N_18880,N_15686,N_16670);
and U18881 (N_18881,N_16383,N_15753);
nor U18882 (N_18882,N_16843,N_16193);
or U18883 (N_18883,N_17294,N_16979);
xor U18884 (N_18884,N_17162,N_16780);
nor U18885 (N_18885,N_17269,N_17436);
and U18886 (N_18886,N_17405,N_16478);
and U18887 (N_18887,N_17178,N_16563);
xnor U18888 (N_18888,N_17437,N_15344);
xor U18889 (N_18889,N_17226,N_16573);
or U18890 (N_18890,N_16403,N_16717);
and U18891 (N_18891,N_15918,N_15143);
nand U18892 (N_18892,N_16216,N_16031);
or U18893 (N_18893,N_16808,N_15983);
or U18894 (N_18894,N_17464,N_16774);
nor U18895 (N_18895,N_15588,N_16139);
nor U18896 (N_18896,N_17071,N_16073);
nand U18897 (N_18897,N_15991,N_15908);
nor U18898 (N_18898,N_15180,N_15190);
and U18899 (N_18899,N_15540,N_15241);
or U18900 (N_18900,N_16733,N_16988);
or U18901 (N_18901,N_16814,N_15152);
nor U18902 (N_18902,N_16341,N_16364);
nor U18903 (N_18903,N_15022,N_15004);
xor U18904 (N_18904,N_15636,N_16110);
nand U18905 (N_18905,N_15172,N_16047);
nor U18906 (N_18906,N_16938,N_16037);
or U18907 (N_18907,N_15750,N_16570);
xnor U18908 (N_18908,N_15022,N_16125);
nor U18909 (N_18909,N_17056,N_17314);
nor U18910 (N_18910,N_15963,N_15029);
or U18911 (N_18911,N_17375,N_17019);
or U18912 (N_18912,N_15439,N_15089);
nor U18913 (N_18913,N_15077,N_17053);
and U18914 (N_18914,N_15572,N_16111);
and U18915 (N_18915,N_15582,N_16989);
or U18916 (N_18916,N_17427,N_15901);
or U18917 (N_18917,N_15413,N_17047);
and U18918 (N_18918,N_16116,N_16044);
xor U18919 (N_18919,N_16410,N_15569);
or U18920 (N_18920,N_15501,N_15758);
nand U18921 (N_18921,N_15355,N_15071);
nand U18922 (N_18922,N_17434,N_17140);
nor U18923 (N_18923,N_15853,N_15788);
nand U18924 (N_18924,N_16338,N_17326);
or U18925 (N_18925,N_16042,N_15822);
nand U18926 (N_18926,N_15035,N_15754);
or U18927 (N_18927,N_15269,N_17236);
or U18928 (N_18928,N_17402,N_15944);
xor U18929 (N_18929,N_16038,N_16448);
or U18930 (N_18930,N_16797,N_15101);
and U18931 (N_18931,N_17267,N_16189);
nor U18932 (N_18932,N_16465,N_17060);
nor U18933 (N_18933,N_15809,N_16524);
or U18934 (N_18934,N_15468,N_17239);
nand U18935 (N_18935,N_16288,N_17236);
nand U18936 (N_18936,N_16978,N_16457);
or U18937 (N_18937,N_17335,N_15704);
xor U18938 (N_18938,N_16416,N_16787);
nand U18939 (N_18939,N_15065,N_15664);
nand U18940 (N_18940,N_15237,N_17310);
nor U18941 (N_18941,N_17160,N_15342);
nand U18942 (N_18942,N_17014,N_15840);
nor U18943 (N_18943,N_16801,N_15100);
nor U18944 (N_18944,N_15908,N_16663);
xnor U18945 (N_18945,N_17019,N_16158);
nor U18946 (N_18946,N_16973,N_17318);
or U18947 (N_18947,N_16240,N_16522);
and U18948 (N_18948,N_15761,N_16773);
and U18949 (N_18949,N_17348,N_16593);
or U18950 (N_18950,N_15685,N_16647);
nand U18951 (N_18951,N_16477,N_16409);
nor U18952 (N_18952,N_16331,N_15304);
nand U18953 (N_18953,N_16649,N_15255);
xor U18954 (N_18954,N_16698,N_17222);
nand U18955 (N_18955,N_15936,N_15816);
nor U18956 (N_18956,N_16692,N_16570);
xor U18957 (N_18957,N_17419,N_15454);
xor U18958 (N_18958,N_15957,N_15887);
xor U18959 (N_18959,N_16703,N_15958);
or U18960 (N_18960,N_16720,N_15924);
or U18961 (N_18961,N_17322,N_16287);
nand U18962 (N_18962,N_15372,N_16375);
nand U18963 (N_18963,N_15822,N_15915);
nand U18964 (N_18964,N_15880,N_15067);
and U18965 (N_18965,N_15237,N_15169);
nand U18966 (N_18966,N_16688,N_16829);
xnor U18967 (N_18967,N_16471,N_15231);
nor U18968 (N_18968,N_17297,N_15010);
nand U18969 (N_18969,N_16352,N_15795);
xnor U18970 (N_18970,N_17333,N_17348);
nor U18971 (N_18971,N_16340,N_15939);
and U18972 (N_18972,N_15313,N_17063);
and U18973 (N_18973,N_15548,N_15839);
nand U18974 (N_18974,N_15611,N_15872);
or U18975 (N_18975,N_15061,N_16351);
xnor U18976 (N_18976,N_16091,N_17230);
or U18977 (N_18977,N_15701,N_17040);
and U18978 (N_18978,N_17482,N_15210);
or U18979 (N_18979,N_15405,N_16074);
or U18980 (N_18980,N_16091,N_16499);
nand U18981 (N_18981,N_16926,N_15851);
nand U18982 (N_18982,N_17036,N_16780);
or U18983 (N_18983,N_15321,N_17447);
nor U18984 (N_18984,N_15056,N_16007);
and U18985 (N_18985,N_16530,N_15628);
and U18986 (N_18986,N_17085,N_16190);
and U18987 (N_18987,N_17337,N_15324);
xor U18988 (N_18988,N_15542,N_15879);
or U18989 (N_18989,N_17471,N_15411);
nand U18990 (N_18990,N_15422,N_15192);
or U18991 (N_18991,N_15242,N_16542);
xnor U18992 (N_18992,N_15891,N_15544);
nor U18993 (N_18993,N_15126,N_16064);
or U18994 (N_18994,N_15316,N_15705);
or U18995 (N_18995,N_16637,N_17074);
nand U18996 (N_18996,N_16602,N_16985);
nor U18997 (N_18997,N_16761,N_16859);
and U18998 (N_18998,N_16908,N_16837);
xor U18999 (N_18999,N_17210,N_15569);
xor U19000 (N_19000,N_16231,N_15110);
xnor U19001 (N_19001,N_16833,N_17281);
or U19002 (N_19002,N_16797,N_16585);
nand U19003 (N_19003,N_15941,N_16755);
or U19004 (N_19004,N_16829,N_15253);
nand U19005 (N_19005,N_15164,N_17312);
xor U19006 (N_19006,N_15465,N_16402);
nand U19007 (N_19007,N_15255,N_15458);
and U19008 (N_19008,N_17013,N_16360);
xor U19009 (N_19009,N_17376,N_15575);
xor U19010 (N_19010,N_16027,N_16715);
xor U19011 (N_19011,N_17497,N_16168);
nand U19012 (N_19012,N_16975,N_15184);
and U19013 (N_19013,N_15528,N_16231);
or U19014 (N_19014,N_16648,N_16543);
xnor U19015 (N_19015,N_16172,N_15727);
xnor U19016 (N_19016,N_17178,N_15387);
nor U19017 (N_19017,N_17092,N_15648);
nor U19018 (N_19018,N_16100,N_16842);
nor U19019 (N_19019,N_16503,N_16163);
xor U19020 (N_19020,N_15167,N_15693);
and U19021 (N_19021,N_15387,N_15547);
nor U19022 (N_19022,N_17171,N_17031);
nor U19023 (N_19023,N_16745,N_16480);
and U19024 (N_19024,N_15972,N_16643);
xor U19025 (N_19025,N_16393,N_16584);
xnor U19026 (N_19026,N_16169,N_16994);
and U19027 (N_19027,N_16300,N_15586);
and U19028 (N_19028,N_15197,N_16196);
xnor U19029 (N_19029,N_17105,N_15709);
nand U19030 (N_19030,N_15976,N_15957);
xnor U19031 (N_19031,N_15645,N_15363);
nor U19032 (N_19032,N_16745,N_16652);
or U19033 (N_19033,N_15684,N_16543);
or U19034 (N_19034,N_17270,N_15604);
and U19035 (N_19035,N_15426,N_16035);
nand U19036 (N_19036,N_15160,N_17239);
nor U19037 (N_19037,N_17208,N_17372);
nand U19038 (N_19038,N_16190,N_16434);
nand U19039 (N_19039,N_15451,N_16045);
xnor U19040 (N_19040,N_17030,N_17099);
or U19041 (N_19041,N_17433,N_16201);
xor U19042 (N_19042,N_17360,N_17301);
or U19043 (N_19043,N_16843,N_16103);
nand U19044 (N_19044,N_16461,N_15615);
nor U19045 (N_19045,N_16047,N_16969);
and U19046 (N_19046,N_15436,N_17449);
nand U19047 (N_19047,N_15997,N_17041);
or U19048 (N_19048,N_16809,N_15367);
and U19049 (N_19049,N_16939,N_16497);
nand U19050 (N_19050,N_15635,N_15818);
xnor U19051 (N_19051,N_16826,N_17473);
xor U19052 (N_19052,N_15538,N_16303);
xnor U19053 (N_19053,N_15157,N_15591);
nand U19054 (N_19054,N_16941,N_17371);
nand U19055 (N_19055,N_15666,N_17061);
and U19056 (N_19056,N_17345,N_15704);
nand U19057 (N_19057,N_17223,N_15993);
or U19058 (N_19058,N_16609,N_15057);
xor U19059 (N_19059,N_16585,N_15478);
nand U19060 (N_19060,N_16103,N_16128);
and U19061 (N_19061,N_17373,N_15894);
or U19062 (N_19062,N_17182,N_15456);
xnor U19063 (N_19063,N_16538,N_16734);
xor U19064 (N_19064,N_16934,N_15135);
nand U19065 (N_19065,N_16715,N_15465);
xnor U19066 (N_19066,N_16090,N_16783);
and U19067 (N_19067,N_17294,N_15032);
nor U19068 (N_19068,N_17173,N_16356);
and U19069 (N_19069,N_16002,N_17218);
xnor U19070 (N_19070,N_15196,N_16489);
or U19071 (N_19071,N_15577,N_16369);
xnor U19072 (N_19072,N_15905,N_15715);
nand U19073 (N_19073,N_17301,N_16504);
and U19074 (N_19074,N_16028,N_16369);
nor U19075 (N_19075,N_15221,N_17464);
nand U19076 (N_19076,N_17445,N_15977);
nor U19077 (N_19077,N_16969,N_17190);
xor U19078 (N_19078,N_15680,N_17236);
xnor U19079 (N_19079,N_16812,N_15822);
xor U19080 (N_19080,N_15673,N_16748);
xnor U19081 (N_19081,N_15301,N_15164);
nor U19082 (N_19082,N_15291,N_15347);
and U19083 (N_19083,N_16673,N_17059);
nor U19084 (N_19084,N_15786,N_15606);
xor U19085 (N_19085,N_16386,N_15234);
and U19086 (N_19086,N_15998,N_15461);
and U19087 (N_19087,N_15028,N_16557);
xnor U19088 (N_19088,N_15977,N_15547);
nand U19089 (N_19089,N_16410,N_16154);
xnor U19090 (N_19090,N_15601,N_17186);
nor U19091 (N_19091,N_15056,N_15592);
and U19092 (N_19092,N_16738,N_16158);
xnor U19093 (N_19093,N_15742,N_17044);
or U19094 (N_19094,N_17295,N_16774);
or U19095 (N_19095,N_15839,N_17023);
or U19096 (N_19096,N_15444,N_17039);
or U19097 (N_19097,N_16780,N_15571);
and U19098 (N_19098,N_15353,N_15572);
xor U19099 (N_19099,N_16795,N_17308);
nand U19100 (N_19100,N_15246,N_16355);
or U19101 (N_19101,N_16596,N_16651);
xor U19102 (N_19102,N_15539,N_17363);
xor U19103 (N_19103,N_16472,N_16889);
and U19104 (N_19104,N_15576,N_15813);
or U19105 (N_19105,N_16747,N_15774);
or U19106 (N_19106,N_16689,N_15641);
xor U19107 (N_19107,N_15122,N_17221);
nor U19108 (N_19108,N_16913,N_16597);
xnor U19109 (N_19109,N_17453,N_17321);
nand U19110 (N_19110,N_15334,N_17222);
and U19111 (N_19111,N_16686,N_16473);
or U19112 (N_19112,N_16494,N_17251);
and U19113 (N_19113,N_15407,N_15837);
xor U19114 (N_19114,N_15548,N_16693);
nor U19115 (N_19115,N_17261,N_15186);
or U19116 (N_19116,N_17410,N_16572);
xor U19117 (N_19117,N_17082,N_17427);
or U19118 (N_19118,N_16805,N_16267);
nand U19119 (N_19119,N_15854,N_15269);
nand U19120 (N_19120,N_16497,N_16733);
nor U19121 (N_19121,N_17082,N_16331);
or U19122 (N_19122,N_16095,N_16899);
nor U19123 (N_19123,N_16530,N_15559);
nor U19124 (N_19124,N_15720,N_15690);
nand U19125 (N_19125,N_15608,N_15474);
nor U19126 (N_19126,N_16782,N_16939);
and U19127 (N_19127,N_17321,N_16970);
or U19128 (N_19128,N_16699,N_16461);
nand U19129 (N_19129,N_16903,N_15989);
and U19130 (N_19130,N_17166,N_16057);
and U19131 (N_19131,N_15225,N_17126);
nand U19132 (N_19132,N_16344,N_15135);
or U19133 (N_19133,N_15636,N_15781);
and U19134 (N_19134,N_15048,N_16474);
and U19135 (N_19135,N_15055,N_16821);
or U19136 (N_19136,N_17438,N_16922);
and U19137 (N_19137,N_16886,N_15717);
or U19138 (N_19138,N_16425,N_15653);
or U19139 (N_19139,N_15421,N_15400);
nor U19140 (N_19140,N_16456,N_16059);
nor U19141 (N_19141,N_17222,N_17047);
nand U19142 (N_19142,N_17345,N_16849);
and U19143 (N_19143,N_16137,N_16136);
and U19144 (N_19144,N_16749,N_17397);
or U19145 (N_19145,N_15600,N_15099);
and U19146 (N_19146,N_15370,N_16174);
or U19147 (N_19147,N_16677,N_15158);
nand U19148 (N_19148,N_15980,N_17258);
nand U19149 (N_19149,N_16001,N_15561);
or U19150 (N_19150,N_15378,N_15143);
or U19151 (N_19151,N_15938,N_15730);
or U19152 (N_19152,N_17305,N_17354);
and U19153 (N_19153,N_17441,N_15308);
nor U19154 (N_19154,N_16899,N_15705);
nand U19155 (N_19155,N_16301,N_16059);
xnor U19156 (N_19156,N_16719,N_17409);
nand U19157 (N_19157,N_15016,N_17283);
or U19158 (N_19158,N_15721,N_15062);
and U19159 (N_19159,N_16599,N_15562);
nor U19160 (N_19160,N_16525,N_17110);
xor U19161 (N_19161,N_15717,N_15557);
and U19162 (N_19162,N_17255,N_15355);
xor U19163 (N_19163,N_16602,N_15592);
xnor U19164 (N_19164,N_16352,N_16911);
or U19165 (N_19165,N_17020,N_17200);
nand U19166 (N_19166,N_16781,N_15196);
xor U19167 (N_19167,N_16765,N_15119);
and U19168 (N_19168,N_15151,N_15930);
and U19169 (N_19169,N_15916,N_16978);
nor U19170 (N_19170,N_16282,N_16831);
nand U19171 (N_19171,N_15479,N_16799);
nand U19172 (N_19172,N_16552,N_16314);
and U19173 (N_19173,N_17400,N_15345);
nand U19174 (N_19174,N_17282,N_16295);
nor U19175 (N_19175,N_17218,N_15371);
or U19176 (N_19176,N_17459,N_16020);
nand U19177 (N_19177,N_16438,N_15229);
xor U19178 (N_19178,N_15461,N_16790);
xor U19179 (N_19179,N_15585,N_16728);
or U19180 (N_19180,N_16611,N_15481);
nand U19181 (N_19181,N_15894,N_15036);
nand U19182 (N_19182,N_15173,N_16216);
nor U19183 (N_19183,N_15935,N_15914);
or U19184 (N_19184,N_15199,N_16324);
xor U19185 (N_19185,N_16709,N_16855);
nor U19186 (N_19186,N_15482,N_17451);
nand U19187 (N_19187,N_17403,N_16185);
and U19188 (N_19188,N_16395,N_15263);
nand U19189 (N_19189,N_17044,N_17279);
or U19190 (N_19190,N_16663,N_15306);
xor U19191 (N_19191,N_16120,N_15415);
nor U19192 (N_19192,N_15475,N_15782);
xnor U19193 (N_19193,N_16553,N_15783);
xor U19194 (N_19194,N_15304,N_15966);
nor U19195 (N_19195,N_16584,N_16305);
nand U19196 (N_19196,N_16008,N_15680);
nor U19197 (N_19197,N_15476,N_17030);
nand U19198 (N_19198,N_16251,N_16903);
or U19199 (N_19199,N_16756,N_17054);
nor U19200 (N_19200,N_15171,N_15032);
nor U19201 (N_19201,N_17456,N_16417);
xnor U19202 (N_19202,N_15440,N_15289);
nor U19203 (N_19203,N_15788,N_16879);
xor U19204 (N_19204,N_16956,N_16605);
and U19205 (N_19205,N_16980,N_16343);
and U19206 (N_19206,N_15646,N_16488);
xor U19207 (N_19207,N_15360,N_15426);
nor U19208 (N_19208,N_16147,N_17285);
nand U19209 (N_19209,N_17030,N_16858);
nor U19210 (N_19210,N_17287,N_16505);
and U19211 (N_19211,N_15739,N_16381);
and U19212 (N_19212,N_15023,N_15502);
or U19213 (N_19213,N_17206,N_15947);
or U19214 (N_19214,N_17123,N_17008);
nand U19215 (N_19215,N_16540,N_16547);
or U19216 (N_19216,N_16267,N_15659);
xor U19217 (N_19217,N_15536,N_16518);
nand U19218 (N_19218,N_16150,N_17116);
nand U19219 (N_19219,N_17322,N_15884);
nand U19220 (N_19220,N_16540,N_17222);
nor U19221 (N_19221,N_15940,N_17470);
nor U19222 (N_19222,N_15991,N_16953);
xnor U19223 (N_19223,N_15463,N_16641);
and U19224 (N_19224,N_17138,N_15752);
nor U19225 (N_19225,N_15599,N_15050);
xnor U19226 (N_19226,N_15790,N_16685);
and U19227 (N_19227,N_15732,N_16958);
and U19228 (N_19228,N_17422,N_15036);
and U19229 (N_19229,N_16062,N_15625);
or U19230 (N_19230,N_17441,N_16370);
and U19231 (N_19231,N_17462,N_17232);
xnor U19232 (N_19232,N_15138,N_15659);
or U19233 (N_19233,N_16850,N_16020);
nor U19234 (N_19234,N_16737,N_17319);
nand U19235 (N_19235,N_17360,N_17022);
xor U19236 (N_19236,N_15429,N_16836);
nor U19237 (N_19237,N_16885,N_15251);
nor U19238 (N_19238,N_15380,N_15207);
or U19239 (N_19239,N_16093,N_16730);
nand U19240 (N_19240,N_15728,N_15998);
xor U19241 (N_19241,N_15293,N_17063);
and U19242 (N_19242,N_16683,N_16940);
and U19243 (N_19243,N_15925,N_16348);
and U19244 (N_19244,N_16495,N_15430);
and U19245 (N_19245,N_16135,N_17365);
nand U19246 (N_19246,N_15336,N_16787);
and U19247 (N_19247,N_16647,N_16102);
xnor U19248 (N_19248,N_16432,N_16277);
or U19249 (N_19249,N_16456,N_15143);
and U19250 (N_19250,N_15565,N_17488);
and U19251 (N_19251,N_15398,N_16740);
nand U19252 (N_19252,N_16874,N_16284);
nor U19253 (N_19253,N_16067,N_16146);
or U19254 (N_19254,N_15459,N_17367);
xor U19255 (N_19255,N_15351,N_15323);
or U19256 (N_19256,N_15863,N_17072);
or U19257 (N_19257,N_16038,N_17211);
or U19258 (N_19258,N_16739,N_15588);
nor U19259 (N_19259,N_17415,N_15871);
and U19260 (N_19260,N_15169,N_16384);
nand U19261 (N_19261,N_15135,N_15886);
and U19262 (N_19262,N_17094,N_16851);
or U19263 (N_19263,N_16571,N_16295);
nand U19264 (N_19264,N_15183,N_17432);
and U19265 (N_19265,N_17018,N_15938);
or U19266 (N_19266,N_16263,N_15569);
nand U19267 (N_19267,N_16487,N_15043);
nor U19268 (N_19268,N_15419,N_16553);
nand U19269 (N_19269,N_15181,N_17420);
nand U19270 (N_19270,N_15050,N_16988);
xor U19271 (N_19271,N_15200,N_16110);
or U19272 (N_19272,N_17158,N_15142);
or U19273 (N_19273,N_17434,N_15115);
xor U19274 (N_19274,N_16790,N_15371);
or U19275 (N_19275,N_15923,N_16095);
or U19276 (N_19276,N_17392,N_16879);
and U19277 (N_19277,N_17420,N_17250);
and U19278 (N_19278,N_15578,N_16222);
xnor U19279 (N_19279,N_15213,N_16449);
nand U19280 (N_19280,N_17080,N_15424);
and U19281 (N_19281,N_16610,N_15671);
nand U19282 (N_19282,N_16259,N_16369);
xnor U19283 (N_19283,N_15380,N_15773);
xor U19284 (N_19284,N_15354,N_17430);
nor U19285 (N_19285,N_17172,N_16372);
or U19286 (N_19286,N_16239,N_16506);
xnor U19287 (N_19287,N_16918,N_16392);
xor U19288 (N_19288,N_16171,N_15661);
or U19289 (N_19289,N_17185,N_16779);
and U19290 (N_19290,N_15262,N_15580);
and U19291 (N_19291,N_15173,N_16987);
xor U19292 (N_19292,N_15738,N_16901);
and U19293 (N_19293,N_15614,N_15206);
nor U19294 (N_19294,N_16384,N_16112);
xor U19295 (N_19295,N_17054,N_16356);
and U19296 (N_19296,N_15137,N_16157);
nand U19297 (N_19297,N_15547,N_15695);
and U19298 (N_19298,N_15360,N_16420);
nor U19299 (N_19299,N_16208,N_16409);
and U19300 (N_19300,N_16982,N_16051);
nor U19301 (N_19301,N_16606,N_15814);
nor U19302 (N_19302,N_15752,N_15388);
and U19303 (N_19303,N_15615,N_15860);
xor U19304 (N_19304,N_15529,N_15792);
nand U19305 (N_19305,N_15115,N_15947);
nor U19306 (N_19306,N_16339,N_17047);
nand U19307 (N_19307,N_17112,N_17160);
nor U19308 (N_19308,N_15345,N_15972);
nor U19309 (N_19309,N_17020,N_16559);
nor U19310 (N_19310,N_16790,N_17013);
nor U19311 (N_19311,N_16891,N_17438);
or U19312 (N_19312,N_16594,N_15797);
or U19313 (N_19313,N_16293,N_16933);
nor U19314 (N_19314,N_16973,N_17009);
nand U19315 (N_19315,N_15482,N_15455);
nand U19316 (N_19316,N_15529,N_15785);
or U19317 (N_19317,N_16329,N_16963);
or U19318 (N_19318,N_16041,N_15514);
xnor U19319 (N_19319,N_16745,N_15254);
nand U19320 (N_19320,N_15599,N_15383);
nor U19321 (N_19321,N_15294,N_16660);
nand U19322 (N_19322,N_17435,N_16171);
or U19323 (N_19323,N_16754,N_17384);
nor U19324 (N_19324,N_16659,N_17181);
nor U19325 (N_19325,N_16470,N_15987);
and U19326 (N_19326,N_15905,N_15133);
or U19327 (N_19327,N_15886,N_15241);
nand U19328 (N_19328,N_17386,N_16811);
xor U19329 (N_19329,N_15792,N_15794);
or U19330 (N_19330,N_15026,N_17421);
and U19331 (N_19331,N_15560,N_16919);
or U19332 (N_19332,N_15569,N_17477);
xnor U19333 (N_19333,N_16061,N_16198);
or U19334 (N_19334,N_16420,N_16777);
and U19335 (N_19335,N_15654,N_17464);
nor U19336 (N_19336,N_15474,N_16256);
nor U19337 (N_19337,N_16742,N_17060);
nor U19338 (N_19338,N_15115,N_17499);
nor U19339 (N_19339,N_17423,N_15891);
or U19340 (N_19340,N_16413,N_17071);
or U19341 (N_19341,N_15940,N_16041);
xnor U19342 (N_19342,N_15285,N_16436);
and U19343 (N_19343,N_17130,N_15259);
and U19344 (N_19344,N_15600,N_16385);
nor U19345 (N_19345,N_15076,N_15829);
nor U19346 (N_19346,N_16457,N_17152);
and U19347 (N_19347,N_17442,N_16313);
nand U19348 (N_19348,N_16960,N_17204);
nor U19349 (N_19349,N_16935,N_15380);
xnor U19350 (N_19350,N_16268,N_16023);
nor U19351 (N_19351,N_16433,N_15396);
and U19352 (N_19352,N_16834,N_16865);
nor U19353 (N_19353,N_15655,N_16371);
and U19354 (N_19354,N_16515,N_17031);
or U19355 (N_19355,N_16946,N_16259);
xor U19356 (N_19356,N_17263,N_16114);
nor U19357 (N_19357,N_17409,N_17404);
xor U19358 (N_19358,N_15850,N_16438);
or U19359 (N_19359,N_15293,N_15808);
and U19360 (N_19360,N_16938,N_16906);
nand U19361 (N_19361,N_15553,N_17442);
nand U19362 (N_19362,N_16621,N_17368);
or U19363 (N_19363,N_15542,N_16870);
nor U19364 (N_19364,N_16022,N_16251);
and U19365 (N_19365,N_16569,N_15127);
nor U19366 (N_19366,N_17295,N_15321);
nand U19367 (N_19367,N_15588,N_15951);
nand U19368 (N_19368,N_15797,N_16746);
nand U19369 (N_19369,N_15215,N_15243);
or U19370 (N_19370,N_17443,N_17197);
xnor U19371 (N_19371,N_15639,N_15051);
or U19372 (N_19372,N_15552,N_16317);
or U19373 (N_19373,N_15277,N_16651);
nor U19374 (N_19374,N_15474,N_17141);
and U19375 (N_19375,N_16820,N_16210);
or U19376 (N_19376,N_15906,N_17135);
or U19377 (N_19377,N_16201,N_16935);
and U19378 (N_19378,N_15706,N_15898);
nor U19379 (N_19379,N_17147,N_16081);
nand U19380 (N_19380,N_16802,N_16830);
nor U19381 (N_19381,N_17339,N_16249);
or U19382 (N_19382,N_16345,N_15254);
nand U19383 (N_19383,N_15094,N_15525);
nor U19384 (N_19384,N_15746,N_16690);
or U19385 (N_19385,N_17092,N_17019);
nor U19386 (N_19386,N_16473,N_17356);
and U19387 (N_19387,N_16656,N_16827);
nand U19388 (N_19388,N_16320,N_15389);
and U19389 (N_19389,N_15076,N_17177);
nand U19390 (N_19390,N_16295,N_16499);
nor U19391 (N_19391,N_15558,N_15842);
or U19392 (N_19392,N_15293,N_15473);
or U19393 (N_19393,N_15483,N_16768);
and U19394 (N_19394,N_15123,N_16770);
nor U19395 (N_19395,N_15758,N_16264);
or U19396 (N_19396,N_16414,N_17481);
xnor U19397 (N_19397,N_15624,N_17077);
nand U19398 (N_19398,N_15371,N_15692);
nor U19399 (N_19399,N_17273,N_17264);
nor U19400 (N_19400,N_16285,N_16765);
nor U19401 (N_19401,N_16349,N_17162);
or U19402 (N_19402,N_17192,N_16695);
or U19403 (N_19403,N_16513,N_15975);
nor U19404 (N_19404,N_17207,N_16584);
nor U19405 (N_19405,N_15285,N_15672);
nor U19406 (N_19406,N_16070,N_16475);
and U19407 (N_19407,N_16287,N_16205);
nand U19408 (N_19408,N_17310,N_15647);
xor U19409 (N_19409,N_15007,N_16189);
nor U19410 (N_19410,N_16802,N_16088);
xnor U19411 (N_19411,N_16248,N_16082);
and U19412 (N_19412,N_15402,N_15792);
nor U19413 (N_19413,N_16135,N_16021);
nand U19414 (N_19414,N_15713,N_15549);
and U19415 (N_19415,N_16745,N_15835);
xor U19416 (N_19416,N_15972,N_15125);
xor U19417 (N_19417,N_16846,N_17360);
or U19418 (N_19418,N_15397,N_16955);
nor U19419 (N_19419,N_16825,N_16787);
nand U19420 (N_19420,N_15308,N_15299);
nand U19421 (N_19421,N_15017,N_15925);
and U19422 (N_19422,N_16440,N_17202);
or U19423 (N_19423,N_15428,N_15433);
nand U19424 (N_19424,N_15682,N_17348);
and U19425 (N_19425,N_16369,N_15051);
nand U19426 (N_19426,N_16976,N_16464);
xor U19427 (N_19427,N_15902,N_17112);
or U19428 (N_19428,N_15941,N_15705);
and U19429 (N_19429,N_15698,N_16800);
nor U19430 (N_19430,N_15166,N_15428);
and U19431 (N_19431,N_15788,N_15213);
nor U19432 (N_19432,N_17305,N_15875);
nand U19433 (N_19433,N_15309,N_15921);
xnor U19434 (N_19434,N_15982,N_15796);
and U19435 (N_19435,N_15324,N_16973);
or U19436 (N_19436,N_15180,N_16747);
nor U19437 (N_19437,N_16950,N_17210);
or U19438 (N_19438,N_15659,N_17305);
xor U19439 (N_19439,N_15026,N_15088);
nor U19440 (N_19440,N_16960,N_15495);
nand U19441 (N_19441,N_17209,N_17010);
or U19442 (N_19442,N_16870,N_15079);
nor U19443 (N_19443,N_15623,N_16412);
nor U19444 (N_19444,N_15341,N_15789);
or U19445 (N_19445,N_16831,N_15834);
nor U19446 (N_19446,N_16901,N_17464);
nor U19447 (N_19447,N_17405,N_16102);
nor U19448 (N_19448,N_16653,N_15610);
or U19449 (N_19449,N_16198,N_17044);
nand U19450 (N_19450,N_15606,N_16119);
nand U19451 (N_19451,N_15819,N_16287);
nand U19452 (N_19452,N_15043,N_16726);
nand U19453 (N_19453,N_16192,N_17271);
xnor U19454 (N_19454,N_17266,N_16413);
xor U19455 (N_19455,N_16079,N_17341);
nand U19456 (N_19456,N_15289,N_16643);
or U19457 (N_19457,N_15858,N_17320);
nor U19458 (N_19458,N_17102,N_15850);
and U19459 (N_19459,N_17339,N_15934);
and U19460 (N_19460,N_15411,N_15636);
nand U19461 (N_19461,N_15352,N_17170);
nor U19462 (N_19462,N_15293,N_15949);
xor U19463 (N_19463,N_15741,N_16108);
nand U19464 (N_19464,N_17490,N_15720);
and U19465 (N_19465,N_15119,N_15542);
nor U19466 (N_19466,N_16118,N_16576);
nor U19467 (N_19467,N_15145,N_15677);
nand U19468 (N_19468,N_15085,N_16474);
nand U19469 (N_19469,N_16525,N_15196);
nor U19470 (N_19470,N_16198,N_17029);
or U19471 (N_19471,N_16068,N_15762);
xor U19472 (N_19472,N_15658,N_15061);
and U19473 (N_19473,N_16506,N_15347);
xnor U19474 (N_19474,N_16172,N_16980);
nor U19475 (N_19475,N_15601,N_16171);
and U19476 (N_19476,N_16947,N_16999);
xnor U19477 (N_19477,N_15867,N_15605);
and U19478 (N_19478,N_17262,N_16622);
nor U19479 (N_19479,N_15260,N_17107);
nand U19480 (N_19480,N_15201,N_15021);
xor U19481 (N_19481,N_15164,N_15023);
nor U19482 (N_19482,N_15602,N_15349);
or U19483 (N_19483,N_16266,N_15672);
xor U19484 (N_19484,N_16101,N_16203);
and U19485 (N_19485,N_16991,N_16440);
and U19486 (N_19486,N_16189,N_16786);
or U19487 (N_19487,N_15398,N_16351);
nor U19488 (N_19488,N_16528,N_17005);
nor U19489 (N_19489,N_17111,N_17012);
xor U19490 (N_19490,N_15425,N_16902);
and U19491 (N_19491,N_15725,N_16193);
and U19492 (N_19492,N_16087,N_16593);
or U19493 (N_19493,N_15281,N_16586);
and U19494 (N_19494,N_16629,N_16411);
nand U19495 (N_19495,N_16757,N_16504);
and U19496 (N_19496,N_15636,N_16993);
xor U19497 (N_19497,N_16675,N_15831);
or U19498 (N_19498,N_17306,N_16143);
and U19499 (N_19499,N_16275,N_15052);
nor U19500 (N_19500,N_16246,N_16486);
or U19501 (N_19501,N_15741,N_16198);
nor U19502 (N_19502,N_17499,N_15618);
xor U19503 (N_19503,N_15391,N_15160);
and U19504 (N_19504,N_16707,N_16781);
nand U19505 (N_19505,N_15398,N_15041);
nand U19506 (N_19506,N_15228,N_17152);
and U19507 (N_19507,N_16589,N_16412);
or U19508 (N_19508,N_15420,N_16977);
and U19509 (N_19509,N_16997,N_16648);
nand U19510 (N_19510,N_16281,N_15560);
nor U19511 (N_19511,N_17443,N_15450);
nor U19512 (N_19512,N_15942,N_17228);
nand U19513 (N_19513,N_15494,N_17071);
and U19514 (N_19514,N_17296,N_15714);
or U19515 (N_19515,N_16950,N_17333);
nor U19516 (N_19516,N_16842,N_15899);
nand U19517 (N_19517,N_16004,N_17306);
nor U19518 (N_19518,N_15143,N_16556);
nand U19519 (N_19519,N_16673,N_16559);
or U19520 (N_19520,N_16707,N_15735);
nand U19521 (N_19521,N_17454,N_15306);
xor U19522 (N_19522,N_16537,N_17461);
nand U19523 (N_19523,N_17034,N_16392);
and U19524 (N_19524,N_15481,N_17390);
or U19525 (N_19525,N_16185,N_16616);
xor U19526 (N_19526,N_16991,N_17075);
or U19527 (N_19527,N_15922,N_16981);
xnor U19528 (N_19528,N_15020,N_15832);
or U19529 (N_19529,N_15767,N_16211);
xnor U19530 (N_19530,N_15823,N_15737);
or U19531 (N_19531,N_17457,N_15581);
nor U19532 (N_19532,N_16580,N_16852);
xor U19533 (N_19533,N_15230,N_17294);
and U19534 (N_19534,N_16352,N_15660);
and U19535 (N_19535,N_16369,N_15849);
nand U19536 (N_19536,N_17452,N_16773);
or U19537 (N_19537,N_17129,N_16512);
xnor U19538 (N_19538,N_17264,N_15369);
nor U19539 (N_19539,N_15244,N_16820);
nand U19540 (N_19540,N_15383,N_15206);
xor U19541 (N_19541,N_15121,N_16281);
xor U19542 (N_19542,N_17023,N_15112);
and U19543 (N_19543,N_15679,N_15373);
nor U19544 (N_19544,N_15700,N_16892);
and U19545 (N_19545,N_17384,N_16535);
xnor U19546 (N_19546,N_16262,N_15159);
nand U19547 (N_19547,N_15897,N_15443);
xor U19548 (N_19548,N_16828,N_15553);
xor U19549 (N_19549,N_16231,N_15668);
and U19550 (N_19550,N_16724,N_16203);
nand U19551 (N_19551,N_17021,N_15317);
nand U19552 (N_19552,N_16215,N_16859);
nor U19553 (N_19553,N_15705,N_17026);
xnor U19554 (N_19554,N_15786,N_16552);
nor U19555 (N_19555,N_16190,N_16762);
and U19556 (N_19556,N_15445,N_16596);
nand U19557 (N_19557,N_16564,N_16256);
nor U19558 (N_19558,N_15654,N_17235);
nor U19559 (N_19559,N_16477,N_17032);
nand U19560 (N_19560,N_15045,N_16005);
nand U19561 (N_19561,N_15745,N_16951);
or U19562 (N_19562,N_16288,N_16901);
nor U19563 (N_19563,N_15032,N_15099);
xor U19564 (N_19564,N_16038,N_16624);
xor U19565 (N_19565,N_16171,N_17443);
and U19566 (N_19566,N_17109,N_15919);
xnor U19567 (N_19567,N_16511,N_15993);
and U19568 (N_19568,N_16656,N_16289);
and U19569 (N_19569,N_15405,N_16795);
nor U19570 (N_19570,N_16676,N_16079);
nand U19571 (N_19571,N_15781,N_16911);
nand U19572 (N_19572,N_15442,N_15036);
or U19573 (N_19573,N_17399,N_16006);
nand U19574 (N_19574,N_16821,N_15198);
nand U19575 (N_19575,N_15432,N_15303);
nand U19576 (N_19576,N_17197,N_16822);
nand U19577 (N_19577,N_17040,N_17252);
or U19578 (N_19578,N_15984,N_16115);
nand U19579 (N_19579,N_15291,N_16037);
or U19580 (N_19580,N_16520,N_15232);
nand U19581 (N_19581,N_15371,N_16773);
xnor U19582 (N_19582,N_15122,N_15510);
nor U19583 (N_19583,N_16882,N_16511);
nor U19584 (N_19584,N_15441,N_16192);
nor U19585 (N_19585,N_16264,N_16682);
nor U19586 (N_19586,N_15327,N_16557);
and U19587 (N_19587,N_15499,N_16585);
and U19588 (N_19588,N_15694,N_15524);
nand U19589 (N_19589,N_15619,N_15463);
nand U19590 (N_19590,N_16976,N_15752);
and U19591 (N_19591,N_16374,N_15434);
or U19592 (N_19592,N_15346,N_16288);
or U19593 (N_19593,N_15431,N_16389);
or U19594 (N_19594,N_16608,N_17340);
nand U19595 (N_19595,N_17201,N_16382);
nand U19596 (N_19596,N_15764,N_16013);
or U19597 (N_19597,N_16264,N_15047);
nand U19598 (N_19598,N_16605,N_15706);
xnor U19599 (N_19599,N_17367,N_16825);
xnor U19600 (N_19600,N_17145,N_15991);
nor U19601 (N_19601,N_15789,N_15578);
nor U19602 (N_19602,N_16716,N_17011);
or U19603 (N_19603,N_17104,N_17090);
nor U19604 (N_19604,N_16825,N_17122);
nand U19605 (N_19605,N_17365,N_17071);
nor U19606 (N_19606,N_15539,N_16841);
xor U19607 (N_19607,N_16391,N_17201);
and U19608 (N_19608,N_15237,N_15879);
nor U19609 (N_19609,N_15261,N_15944);
nor U19610 (N_19610,N_15233,N_16562);
nor U19611 (N_19611,N_17312,N_15899);
and U19612 (N_19612,N_16808,N_15051);
or U19613 (N_19613,N_15634,N_17400);
and U19614 (N_19614,N_17197,N_16190);
or U19615 (N_19615,N_15952,N_16585);
or U19616 (N_19616,N_16537,N_15979);
and U19617 (N_19617,N_16668,N_15928);
nor U19618 (N_19618,N_16666,N_15752);
or U19619 (N_19619,N_17400,N_16301);
and U19620 (N_19620,N_15082,N_15638);
and U19621 (N_19621,N_15370,N_15164);
nor U19622 (N_19622,N_16815,N_15142);
nor U19623 (N_19623,N_16600,N_16276);
nor U19624 (N_19624,N_16439,N_16325);
nor U19625 (N_19625,N_16995,N_17048);
nor U19626 (N_19626,N_15936,N_15996);
nand U19627 (N_19627,N_15664,N_17268);
nand U19628 (N_19628,N_17496,N_16411);
or U19629 (N_19629,N_15675,N_16143);
nor U19630 (N_19630,N_17310,N_17035);
xnor U19631 (N_19631,N_15997,N_17032);
and U19632 (N_19632,N_17208,N_15945);
and U19633 (N_19633,N_16157,N_16177);
or U19634 (N_19634,N_16403,N_15683);
nor U19635 (N_19635,N_16867,N_15249);
and U19636 (N_19636,N_16148,N_16223);
and U19637 (N_19637,N_16200,N_15847);
nand U19638 (N_19638,N_15902,N_15091);
and U19639 (N_19639,N_15619,N_16252);
nor U19640 (N_19640,N_15774,N_16369);
nor U19641 (N_19641,N_16886,N_15689);
xnor U19642 (N_19642,N_16051,N_15161);
and U19643 (N_19643,N_15788,N_17308);
nor U19644 (N_19644,N_16128,N_16759);
xnor U19645 (N_19645,N_16312,N_15738);
xnor U19646 (N_19646,N_15264,N_16868);
or U19647 (N_19647,N_15478,N_17081);
xnor U19648 (N_19648,N_17094,N_16862);
or U19649 (N_19649,N_15557,N_15941);
or U19650 (N_19650,N_15332,N_15425);
nor U19651 (N_19651,N_16695,N_15502);
and U19652 (N_19652,N_17253,N_16613);
nand U19653 (N_19653,N_15504,N_17249);
and U19654 (N_19654,N_16029,N_16534);
or U19655 (N_19655,N_16398,N_16717);
xor U19656 (N_19656,N_16437,N_16719);
nand U19657 (N_19657,N_17308,N_15476);
xor U19658 (N_19658,N_15799,N_15881);
nor U19659 (N_19659,N_15922,N_16860);
xnor U19660 (N_19660,N_15928,N_15035);
nand U19661 (N_19661,N_17464,N_15632);
nor U19662 (N_19662,N_15155,N_15735);
or U19663 (N_19663,N_15306,N_15578);
nor U19664 (N_19664,N_16015,N_16891);
or U19665 (N_19665,N_15728,N_15680);
xnor U19666 (N_19666,N_15721,N_16938);
xor U19667 (N_19667,N_15684,N_15638);
xnor U19668 (N_19668,N_15708,N_16379);
nand U19669 (N_19669,N_17405,N_16544);
nand U19670 (N_19670,N_16347,N_16134);
nor U19671 (N_19671,N_15944,N_16254);
nand U19672 (N_19672,N_15410,N_16325);
xor U19673 (N_19673,N_15806,N_17252);
nor U19674 (N_19674,N_16860,N_15743);
or U19675 (N_19675,N_16156,N_15198);
xnor U19676 (N_19676,N_15453,N_16293);
xor U19677 (N_19677,N_15984,N_17315);
and U19678 (N_19678,N_17096,N_16554);
xor U19679 (N_19679,N_15147,N_15042);
xnor U19680 (N_19680,N_16590,N_15378);
or U19681 (N_19681,N_16216,N_17251);
and U19682 (N_19682,N_15196,N_17480);
xor U19683 (N_19683,N_17434,N_17406);
nand U19684 (N_19684,N_17275,N_15007);
nor U19685 (N_19685,N_15048,N_15211);
and U19686 (N_19686,N_15730,N_15402);
nor U19687 (N_19687,N_16799,N_15782);
nand U19688 (N_19688,N_16438,N_17203);
nand U19689 (N_19689,N_17348,N_16971);
or U19690 (N_19690,N_17499,N_17470);
nand U19691 (N_19691,N_15964,N_15506);
nand U19692 (N_19692,N_15124,N_16476);
xor U19693 (N_19693,N_16910,N_16690);
or U19694 (N_19694,N_17351,N_16305);
or U19695 (N_19695,N_15511,N_15722);
nor U19696 (N_19696,N_17429,N_15739);
or U19697 (N_19697,N_17430,N_17432);
nand U19698 (N_19698,N_16497,N_15359);
nand U19699 (N_19699,N_16922,N_17013);
nand U19700 (N_19700,N_15498,N_17440);
or U19701 (N_19701,N_16856,N_17183);
nand U19702 (N_19702,N_15139,N_16642);
nand U19703 (N_19703,N_16867,N_16063);
xor U19704 (N_19704,N_15681,N_15601);
nand U19705 (N_19705,N_16206,N_15897);
xnor U19706 (N_19706,N_17351,N_15118);
nor U19707 (N_19707,N_16698,N_16878);
and U19708 (N_19708,N_17071,N_16361);
and U19709 (N_19709,N_15987,N_15228);
xor U19710 (N_19710,N_15690,N_17293);
nand U19711 (N_19711,N_17381,N_16715);
xnor U19712 (N_19712,N_17439,N_15742);
or U19713 (N_19713,N_17428,N_15098);
and U19714 (N_19714,N_15532,N_16002);
nand U19715 (N_19715,N_17315,N_16059);
and U19716 (N_19716,N_17257,N_16289);
xnor U19717 (N_19717,N_17262,N_15828);
and U19718 (N_19718,N_15811,N_16605);
xor U19719 (N_19719,N_15336,N_15206);
nand U19720 (N_19720,N_17220,N_16486);
nand U19721 (N_19721,N_16647,N_16914);
nor U19722 (N_19722,N_16401,N_15582);
or U19723 (N_19723,N_15783,N_17458);
and U19724 (N_19724,N_17044,N_16178);
and U19725 (N_19725,N_16810,N_17246);
nand U19726 (N_19726,N_17472,N_17277);
nand U19727 (N_19727,N_15392,N_16964);
and U19728 (N_19728,N_15031,N_15265);
nand U19729 (N_19729,N_15235,N_15814);
and U19730 (N_19730,N_17039,N_15387);
nor U19731 (N_19731,N_16772,N_17282);
nor U19732 (N_19732,N_15932,N_16571);
nor U19733 (N_19733,N_15930,N_16500);
nand U19734 (N_19734,N_15071,N_15313);
nand U19735 (N_19735,N_16754,N_16618);
nand U19736 (N_19736,N_16088,N_16773);
nor U19737 (N_19737,N_15729,N_15560);
or U19738 (N_19738,N_16311,N_16373);
or U19739 (N_19739,N_15791,N_15018);
nand U19740 (N_19740,N_16491,N_17123);
or U19741 (N_19741,N_16738,N_16943);
or U19742 (N_19742,N_17039,N_15755);
or U19743 (N_19743,N_17403,N_17126);
nand U19744 (N_19744,N_15539,N_16771);
nor U19745 (N_19745,N_15703,N_16392);
nor U19746 (N_19746,N_15410,N_15470);
xor U19747 (N_19747,N_15564,N_16305);
nor U19748 (N_19748,N_17178,N_15853);
nand U19749 (N_19749,N_16747,N_16269);
nand U19750 (N_19750,N_16489,N_17480);
and U19751 (N_19751,N_17328,N_15868);
nand U19752 (N_19752,N_15434,N_15940);
xnor U19753 (N_19753,N_16621,N_16845);
or U19754 (N_19754,N_17052,N_15005);
nand U19755 (N_19755,N_17318,N_15021);
and U19756 (N_19756,N_15100,N_17225);
nand U19757 (N_19757,N_15440,N_17224);
xnor U19758 (N_19758,N_17338,N_15145);
xor U19759 (N_19759,N_17392,N_16066);
or U19760 (N_19760,N_17048,N_15479);
nor U19761 (N_19761,N_16196,N_17259);
or U19762 (N_19762,N_15143,N_16575);
and U19763 (N_19763,N_17364,N_16341);
and U19764 (N_19764,N_15826,N_15609);
nand U19765 (N_19765,N_17364,N_16003);
nand U19766 (N_19766,N_16309,N_16352);
and U19767 (N_19767,N_16842,N_15177);
or U19768 (N_19768,N_16565,N_16922);
nor U19769 (N_19769,N_16206,N_17462);
and U19770 (N_19770,N_15124,N_15326);
xor U19771 (N_19771,N_15258,N_17346);
nand U19772 (N_19772,N_15490,N_15838);
and U19773 (N_19773,N_17268,N_16248);
nand U19774 (N_19774,N_17401,N_15104);
or U19775 (N_19775,N_17086,N_15092);
xor U19776 (N_19776,N_16604,N_15303);
and U19777 (N_19777,N_16514,N_15761);
xnor U19778 (N_19778,N_15337,N_17361);
nand U19779 (N_19779,N_17096,N_16664);
nor U19780 (N_19780,N_15883,N_16526);
or U19781 (N_19781,N_16058,N_16980);
or U19782 (N_19782,N_16416,N_17175);
nor U19783 (N_19783,N_15756,N_15574);
and U19784 (N_19784,N_15503,N_15976);
or U19785 (N_19785,N_16357,N_16173);
and U19786 (N_19786,N_16523,N_17120);
nand U19787 (N_19787,N_17406,N_17167);
or U19788 (N_19788,N_16858,N_17433);
or U19789 (N_19789,N_16375,N_16184);
xnor U19790 (N_19790,N_16511,N_17441);
nand U19791 (N_19791,N_15291,N_15974);
nand U19792 (N_19792,N_15078,N_16000);
or U19793 (N_19793,N_15031,N_16940);
or U19794 (N_19794,N_17375,N_16034);
or U19795 (N_19795,N_16206,N_15504);
and U19796 (N_19796,N_16257,N_17378);
nand U19797 (N_19797,N_16711,N_16300);
nand U19798 (N_19798,N_15024,N_16480);
nand U19799 (N_19799,N_17014,N_17132);
nor U19800 (N_19800,N_15706,N_17179);
and U19801 (N_19801,N_15534,N_16045);
nand U19802 (N_19802,N_15855,N_16276);
or U19803 (N_19803,N_15927,N_16053);
nor U19804 (N_19804,N_15865,N_15974);
nand U19805 (N_19805,N_16237,N_15233);
nor U19806 (N_19806,N_15542,N_16558);
xor U19807 (N_19807,N_17192,N_17229);
nand U19808 (N_19808,N_17144,N_15391);
or U19809 (N_19809,N_17245,N_15795);
nor U19810 (N_19810,N_15659,N_17224);
or U19811 (N_19811,N_16678,N_16055);
nand U19812 (N_19812,N_16581,N_15052);
nand U19813 (N_19813,N_16963,N_16670);
and U19814 (N_19814,N_16325,N_17207);
nor U19815 (N_19815,N_15944,N_15063);
nor U19816 (N_19816,N_17204,N_16688);
nor U19817 (N_19817,N_17125,N_16561);
and U19818 (N_19818,N_15771,N_17155);
xor U19819 (N_19819,N_15415,N_16852);
and U19820 (N_19820,N_16525,N_17475);
nor U19821 (N_19821,N_17213,N_16320);
nand U19822 (N_19822,N_15254,N_15453);
nand U19823 (N_19823,N_16563,N_17101);
xnor U19824 (N_19824,N_16501,N_17060);
xnor U19825 (N_19825,N_16141,N_15193);
or U19826 (N_19826,N_16824,N_16046);
or U19827 (N_19827,N_15896,N_16541);
and U19828 (N_19828,N_16260,N_15103);
and U19829 (N_19829,N_16020,N_17328);
nor U19830 (N_19830,N_16351,N_15128);
nand U19831 (N_19831,N_16353,N_16830);
or U19832 (N_19832,N_16815,N_16209);
or U19833 (N_19833,N_15511,N_15780);
or U19834 (N_19834,N_15224,N_16227);
and U19835 (N_19835,N_17368,N_15232);
xnor U19836 (N_19836,N_17270,N_15480);
and U19837 (N_19837,N_16234,N_16013);
xnor U19838 (N_19838,N_17022,N_17116);
nor U19839 (N_19839,N_15231,N_15546);
or U19840 (N_19840,N_16646,N_16046);
nand U19841 (N_19841,N_16921,N_16082);
or U19842 (N_19842,N_17373,N_15488);
or U19843 (N_19843,N_17321,N_16783);
nand U19844 (N_19844,N_15211,N_15711);
and U19845 (N_19845,N_15186,N_16481);
nor U19846 (N_19846,N_16335,N_16902);
or U19847 (N_19847,N_17157,N_16256);
nand U19848 (N_19848,N_15809,N_16896);
nand U19849 (N_19849,N_15868,N_15711);
nor U19850 (N_19850,N_15190,N_16043);
xor U19851 (N_19851,N_16002,N_17139);
nor U19852 (N_19852,N_15860,N_16849);
and U19853 (N_19853,N_15875,N_15512);
nand U19854 (N_19854,N_15899,N_15235);
and U19855 (N_19855,N_17121,N_17352);
and U19856 (N_19856,N_15049,N_16889);
nor U19857 (N_19857,N_16330,N_16904);
or U19858 (N_19858,N_17121,N_15807);
or U19859 (N_19859,N_15757,N_17338);
nand U19860 (N_19860,N_16869,N_15334);
and U19861 (N_19861,N_15018,N_15937);
or U19862 (N_19862,N_15337,N_16266);
nor U19863 (N_19863,N_15537,N_16208);
xor U19864 (N_19864,N_16285,N_16414);
or U19865 (N_19865,N_16002,N_15007);
nor U19866 (N_19866,N_17349,N_16224);
and U19867 (N_19867,N_17191,N_16405);
nor U19868 (N_19868,N_15617,N_15396);
nand U19869 (N_19869,N_17102,N_17221);
nor U19870 (N_19870,N_16734,N_15734);
nor U19871 (N_19871,N_16776,N_16280);
xor U19872 (N_19872,N_15029,N_15413);
and U19873 (N_19873,N_16573,N_16221);
nand U19874 (N_19874,N_17310,N_16516);
or U19875 (N_19875,N_15245,N_16160);
or U19876 (N_19876,N_15358,N_15908);
or U19877 (N_19877,N_16746,N_15385);
nor U19878 (N_19878,N_16058,N_16725);
nor U19879 (N_19879,N_15115,N_16340);
nand U19880 (N_19880,N_15789,N_16794);
and U19881 (N_19881,N_17121,N_16646);
nand U19882 (N_19882,N_16820,N_16897);
or U19883 (N_19883,N_15845,N_15515);
nor U19884 (N_19884,N_15779,N_15140);
or U19885 (N_19885,N_16980,N_16212);
or U19886 (N_19886,N_16602,N_16526);
nand U19887 (N_19887,N_15804,N_15286);
nand U19888 (N_19888,N_15290,N_15914);
nand U19889 (N_19889,N_17330,N_16197);
or U19890 (N_19890,N_16113,N_16443);
nand U19891 (N_19891,N_16637,N_16110);
xor U19892 (N_19892,N_15826,N_16187);
nor U19893 (N_19893,N_16428,N_16437);
nor U19894 (N_19894,N_17443,N_17001);
nand U19895 (N_19895,N_15487,N_15274);
nor U19896 (N_19896,N_17050,N_16703);
nor U19897 (N_19897,N_15474,N_16746);
nor U19898 (N_19898,N_16790,N_17037);
xnor U19899 (N_19899,N_16656,N_15858);
nand U19900 (N_19900,N_16345,N_17462);
nand U19901 (N_19901,N_17440,N_16951);
xor U19902 (N_19902,N_16308,N_17066);
and U19903 (N_19903,N_15292,N_15552);
and U19904 (N_19904,N_16138,N_16352);
or U19905 (N_19905,N_17078,N_16051);
xor U19906 (N_19906,N_15035,N_16467);
nor U19907 (N_19907,N_17175,N_15255);
xnor U19908 (N_19908,N_16316,N_16759);
xnor U19909 (N_19909,N_15257,N_15384);
nand U19910 (N_19910,N_16884,N_16315);
or U19911 (N_19911,N_15528,N_15078);
or U19912 (N_19912,N_16046,N_15152);
nand U19913 (N_19913,N_16409,N_15760);
nor U19914 (N_19914,N_16075,N_15971);
nor U19915 (N_19915,N_16334,N_15105);
nand U19916 (N_19916,N_16972,N_16789);
nand U19917 (N_19917,N_16749,N_16438);
nor U19918 (N_19918,N_17380,N_15764);
nand U19919 (N_19919,N_15351,N_15283);
nor U19920 (N_19920,N_16007,N_15673);
nand U19921 (N_19921,N_16549,N_15307);
xor U19922 (N_19922,N_16510,N_16099);
nor U19923 (N_19923,N_16809,N_17474);
nand U19924 (N_19924,N_15889,N_15713);
xor U19925 (N_19925,N_16090,N_16355);
xor U19926 (N_19926,N_15931,N_15666);
xor U19927 (N_19927,N_16476,N_16328);
and U19928 (N_19928,N_16482,N_16916);
nand U19929 (N_19929,N_15360,N_15641);
xor U19930 (N_19930,N_16390,N_16610);
nor U19931 (N_19931,N_15507,N_16313);
and U19932 (N_19932,N_15360,N_16059);
nand U19933 (N_19933,N_17373,N_15971);
xnor U19934 (N_19934,N_15071,N_16414);
and U19935 (N_19935,N_17419,N_15624);
and U19936 (N_19936,N_16282,N_16664);
and U19937 (N_19937,N_15718,N_15664);
nand U19938 (N_19938,N_16383,N_16470);
xnor U19939 (N_19939,N_16172,N_15419);
or U19940 (N_19940,N_15682,N_16022);
xnor U19941 (N_19941,N_15532,N_15551);
xnor U19942 (N_19942,N_16911,N_15257);
nor U19943 (N_19943,N_16987,N_15097);
or U19944 (N_19944,N_16303,N_17023);
nand U19945 (N_19945,N_15399,N_16669);
nand U19946 (N_19946,N_16025,N_17374);
or U19947 (N_19947,N_15233,N_15782);
and U19948 (N_19948,N_16235,N_15122);
nand U19949 (N_19949,N_17480,N_16787);
xor U19950 (N_19950,N_15893,N_15080);
nand U19951 (N_19951,N_15572,N_16611);
and U19952 (N_19952,N_15412,N_16488);
or U19953 (N_19953,N_15532,N_15545);
nand U19954 (N_19954,N_16889,N_16139);
nand U19955 (N_19955,N_17263,N_16781);
nor U19956 (N_19956,N_16758,N_15163);
or U19957 (N_19957,N_17074,N_17430);
or U19958 (N_19958,N_16368,N_15510);
or U19959 (N_19959,N_15730,N_16254);
nor U19960 (N_19960,N_15718,N_16367);
and U19961 (N_19961,N_16569,N_16882);
or U19962 (N_19962,N_17483,N_16763);
nand U19963 (N_19963,N_16638,N_15820);
or U19964 (N_19964,N_15409,N_15377);
xnor U19965 (N_19965,N_15322,N_15213);
nor U19966 (N_19966,N_16566,N_17290);
nand U19967 (N_19967,N_16642,N_15373);
xor U19968 (N_19968,N_15413,N_16650);
and U19969 (N_19969,N_17113,N_15048);
nor U19970 (N_19970,N_16114,N_15733);
nand U19971 (N_19971,N_17394,N_16375);
nor U19972 (N_19972,N_17417,N_16612);
nand U19973 (N_19973,N_16818,N_17026);
xor U19974 (N_19974,N_16562,N_16801);
or U19975 (N_19975,N_17123,N_15708);
or U19976 (N_19976,N_16045,N_17352);
and U19977 (N_19977,N_17350,N_15276);
xor U19978 (N_19978,N_16219,N_16524);
nand U19979 (N_19979,N_16108,N_16704);
nand U19980 (N_19980,N_15337,N_15679);
xnor U19981 (N_19981,N_16828,N_15762);
xor U19982 (N_19982,N_16519,N_16117);
nor U19983 (N_19983,N_16282,N_16128);
nor U19984 (N_19984,N_16339,N_16669);
nand U19985 (N_19985,N_17399,N_16814);
and U19986 (N_19986,N_15616,N_15353);
nand U19987 (N_19987,N_17257,N_15289);
nand U19988 (N_19988,N_15513,N_15097);
and U19989 (N_19989,N_16263,N_16480);
or U19990 (N_19990,N_17445,N_16104);
nor U19991 (N_19991,N_15892,N_16644);
nand U19992 (N_19992,N_15844,N_15207);
or U19993 (N_19993,N_16903,N_16051);
or U19994 (N_19994,N_16692,N_17290);
or U19995 (N_19995,N_15231,N_15310);
and U19996 (N_19996,N_15598,N_17002);
xor U19997 (N_19997,N_16428,N_15728);
nor U19998 (N_19998,N_17233,N_16441);
or U19999 (N_19999,N_16025,N_17056);
and U20000 (N_20000,N_19822,N_17942);
or U20001 (N_20001,N_19922,N_19683);
nand U20002 (N_20002,N_18276,N_19705);
xor U20003 (N_20003,N_17612,N_19275);
nor U20004 (N_20004,N_19145,N_19377);
and U20005 (N_20005,N_19345,N_19589);
nor U20006 (N_20006,N_19941,N_19294);
nand U20007 (N_20007,N_19694,N_18028);
and U20008 (N_20008,N_18754,N_18376);
nor U20009 (N_20009,N_19086,N_18725);
nand U20010 (N_20010,N_18964,N_19506);
nor U20011 (N_20011,N_17684,N_17875);
nand U20012 (N_20012,N_17518,N_17729);
and U20013 (N_20013,N_19936,N_17688);
nor U20014 (N_20014,N_19007,N_19419);
and U20015 (N_20015,N_19513,N_17540);
nor U20016 (N_20016,N_18357,N_19659);
nand U20017 (N_20017,N_17772,N_19119);
or U20018 (N_20018,N_17714,N_19350);
or U20019 (N_20019,N_18269,N_19792);
xnor U20020 (N_20020,N_18402,N_19503);
nand U20021 (N_20021,N_19805,N_19697);
nor U20022 (N_20022,N_18597,N_18022);
xor U20023 (N_20023,N_18427,N_18046);
xor U20024 (N_20024,N_19985,N_18946);
or U20025 (N_20025,N_17666,N_17639);
nand U20026 (N_20026,N_18462,N_19576);
and U20027 (N_20027,N_18898,N_18832);
nor U20028 (N_20028,N_18998,N_17662);
nor U20029 (N_20029,N_19718,N_19994);
or U20030 (N_20030,N_19573,N_18076);
nand U20031 (N_20031,N_18840,N_17584);
xnor U20032 (N_20032,N_18524,N_19742);
or U20033 (N_20033,N_18612,N_17732);
and U20034 (N_20034,N_19632,N_19093);
nand U20035 (N_20035,N_17669,N_19990);
xnor U20036 (N_20036,N_17730,N_18280);
and U20037 (N_20037,N_19300,N_19339);
nand U20038 (N_20038,N_19611,N_19072);
or U20039 (N_20039,N_19876,N_17727);
nor U20040 (N_20040,N_17889,N_18686);
xor U20041 (N_20041,N_18650,N_18669);
nand U20042 (N_20042,N_17756,N_17615);
nand U20043 (N_20043,N_17759,N_19411);
nor U20044 (N_20044,N_19098,N_17689);
xnor U20045 (N_20045,N_17902,N_19527);
nand U20046 (N_20046,N_19290,N_18654);
xor U20047 (N_20047,N_19753,N_17509);
or U20048 (N_20048,N_19963,N_19899);
xor U20049 (N_20049,N_19172,N_19715);
xnor U20050 (N_20050,N_17678,N_18024);
nor U20051 (N_20051,N_17629,N_19486);
nand U20052 (N_20052,N_18884,N_18311);
xnor U20053 (N_20053,N_19128,N_17698);
and U20054 (N_20054,N_17646,N_18041);
and U20055 (N_20055,N_19826,N_18331);
nor U20056 (N_20056,N_18468,N_19819);
or U20057 (N_20057,N_18708,N_18823);
nor U20058 (N_20058,N_19130,N_18585);
or U20059 (N_20059,N_19518,N_17716);
nor U20060 (N_20060,N_19144,N_17681);
nor U20061 (N_20061,N_19712,N_19592);
or U20062 (N_20062,N_19771,N_19153);
nor U20063 (N_20063,N_19192,N_19522);
or U20064 (N_20064,N_19523,N_18348);
nor U20065 (N_20065,N_17950,N_18851);
nor U20066 (N_20066,N_17601,N_18474);
or U20067 (N_20067,N_18140,N_17631);
or U20068 (N_20068,N_19030,N_18662);
nand U20069 (N_20069,N_19544,N_17828);
or U20070 (N_20070,N_18342,N_19642);
xnor U20071 (N_20071,N_19921,N_19295);
nand U20072 (N_20072,N_17816,N_19695);
xnor U20073 (N_20073,N_19997,N_17933);
or U20074 (N_20074,N_18991,N_19443);
or U20075 (N_20075,N_19241,N_19399);
or U20076 (N_20076,N_19686,N_19422);
nor U20077 (N_20077,N_18992,N_18798);
or U20078 (N_20078,N_18497,N_18383);
nand U20079 (N_20079,N_17944,N_18382);
and U20080 (N_20080,N_18476,N_19635);
nor U20081 (N_20081,N_18846,N_19949);
or U20082 (N_20082,N_18002,N_19099);
or U20083 (N_20083,N_18627,N_18525);
and U20084 (N_20084,N_18172,N_19863);
xor U20085 (N_20085,N_18567,N_18271);
nand U20086 (N_20086,N_19674,N_17578);
nor U20087 (N_20087,N_19862,N_18407);
nand U20088 (N_20088,N_19005,N_17938);
nor U20089 (N_20089,N_17948,N_18515);
nand U20090 (N_20090,N_18417,N_18976);
or U20091 (N_20091,N_19626,N_18859);
nand U20092 (N_20092,N_18935,N_19171);
xnor U20093 (N_20093,N_18575,N_18475);
nor U20094 (N_20094,N_18503,N_19424);
nor U20095 (N_20095,N_17943,N_19239);
and U20096 (N_20096,N_17625,N_18444);
or U20097 (N_20097,N_19152,N_19918);
and U20098 (N_20098,N_19854,N_17620);
or U20099 (N_20099,N_17892,N_17535);
nand U20100 (N_20100,N_19579,N_19406);
and U20101 (N_20101,N_19616,N_17651);
or U20102 (N_20102,N_18029,N_19500);
xor U20103 (N_20103,N_17847,N_17715);
and U20104 (N_20104,N_18435,N_19268);
nand U20105 (N_20105,N_19673,N_19227);
and U20106 (N_20106,N_19105,N_19956);
or U20107 (N_20107,N_18709,N_19559);
nor U20108 (N_20108,N_17537,N_18732);
nor U20109 (N_20109,N_18239,N_17758);
xor U20110 (N_20110,N_17774,N_17965);
xor U20111 (N_20111,N_19050,N_18431);
nand U20112 (N_20112,N_19006,N_18337);
nand U20113 (N_20113,N_19911,N_18107);
and U20114 (N_20114,N_17663,N_18541);
or U20115 (N_20115,N_19657,N_19379);
xor U20116 (N_20116,N_17825,N_18792);
xor U20117 (N_20117,N_19542,N_19925);
nand U20118 (N_20118,N_18275,N_19230);
or U20119 (N_20119,N_18071,N_19586);
xor U20120 (N_20120,N_18428,N_17574);
nand U20121 (N_20121,N_18031,N_17528);
nor U20122 (N_20122,N_17827,N_18129);
or U20123 (N_20123,N_19610,N_17692);
or U20124 (N_20124,N_17947,N_18096);
nand U20125 (N_20125,N_18550,N_19881);
and U20126 (N_20126,N_19408,N_18498);
nand U20127 (N_20127,N_18943,N_18278);
xor U20128 (N_20128,N_18023,N_18176);
nand U20129 (N_20129,N_17534,N_19371);
nor U20130 (N_20130,N_19211,N_19008);
nand U20131 (N_20131,N_19165,N_19568);
or U20132 (N_20132,N_19692,N_17973);
nand U20133 (N_20133,N_18090,N_18443);
nand U20134 (N_20134,N_17582,N_17740);
or U20135 (N_20135,N_18739,N_18756);
xnor U20136 (N_20136,N_18381,N_17876);
nand U20137 (N_20137,N_19034,N_18349);
or U20138 (N_20138,N_18600,N_19120);
or U20139 (N_20139,N_17953,N_19627);
and U20140 (N_20140,N_18098,N_19136);
nand U20141 (N_20141,N_19235,N_18328);
xnor U20142 (N_20142,N_18319,N_18522);
xnor U20143 (N_20143,N_18863,N_19681);
nor U20144 (N_20144,N_17926,N_17568);
or U20145 (N_20145,N_18640,N_18582);
nand U20146 (N_20146,N_18747,N_18584);
nand U20147 (N_20147,N_18235,N_18472);
or U20148 (N_20148,N_18665,N_18405);
or U20149 (N_20149,N_18562,N_19018);
xor U20150 (N_20150,N_19721,N_18897);
nor U20151 (N_20151,N_19209,N_18393);
or U20152 (N_20152,N_19440,N_17585);
or U20153 (N_20153,N_18369,N_19009);
or U20154 (N_20154,N_17810,N_17526);
nor U20155 (N_20155,N_17762,N_19534);
nor U20156 (N_20156,N_19717,N_18481);
and U20157 (N_20157,N_19930,N_19395);
nor U20158 (N_20158,N_17867,N_19597);
nor U20159 (N_20159,N_19217,N_18656);
and U20160 (N_20160,N_19601,N_17626);
nand U20161 (N_20161,N_18950,N_19474);
nand U20162 (N_20162,N_18658,N_18642);
and U20163 (N_20163,N_18529,N_19426);
xnor U20164 (N_20164,N_19582,N_17768);
and U20165 (N_20165,N_19510,N_19979);
nor U20166 (N_20166,N_19388,N_18788);
nor U20167 (N_20167,N_17807,N_18543);
nor U20168 (N_20168,N_18735,N_19807);
nand U20169 (N_20169,N_19306,N_17508);
nand U20170 (N_20170,N_19070,N_18359);
or U20171 (N_20171,N_18360,N_19279);
nand U20172 (N_20172,N_18063,N_17635);
nor U20173 (N_20173,N_17981,N_19106);
or U20174 (N_20174,N_19427,N_18557);
or U20175 (N_20175,N_17549,N_17776);
and U20176 (N_20176,N_19647,N_18212);
xor U20177 (N_20177,N_18100,N_18253);
nor U20178 (N_20178,N_19001,N_18972);
xor U20179 (N_20179,N_19855,N_18317);
or U20180 (N_20180,N_19434,N_19969);
and U20181 (N_20181,N_19351,N_19374);
nand U20182 (N_20182,N_17909,N_17991);
xnor U20183 (N_20183,N_17580,N_18890);
nand U20184 (N_20184,N_19556,N_19679);
xor U20185 (N_20185,N_17751,N_19829);
nor U20186 (N_20186,N_17562,N_18777);
and U20187 (N_20187,N_19947,N_18323);
xor U20188 (N_20188,N_19957,N_19287);
xnor U20189 (N_20189,N_19740,N_18601);
or U20190 (N_20190,N_17804,N_19107);
xor U20191 (N_20191,N_19469,N_18691);
or U20192 (N_20192,N_17788,N_18088);
and U20193 (N_20193,N_19360,N_18716);
nor U20194 (N_20194,N_18839,N_18354);
or U20195 (N_20195,N_19902,N_17990);
nand U20196 (N_20196,N_19430,N_19314);
nor U20197 (N_20197,N_19977,N_18891);
and U20198 (N_20198,N_19968,N_17918);
nor U20199 (N_20199,N_18746,N_17643);
and U20200 (N_20200,N_19233,N_17739);
or U20201 (N_20201,N_17900,N_17815);
xnor U20202 (N_20202,N_19044,N_18807);
and U20203 (N_20203,N_18980,N_18711);
or U20204 (N_20204,N_18085,N_17809);
nor U20205 (N_20205,N_18762,N_17849);
or U20206 (N_20206,N_19507,N_17752);
nor U20207 (N_20207,N_18936,N_18161);
xor U20208 (N_20208,N_18429,N_17718);
and U20209 (N_20209,N_18255,N_19067);
xnor U20210 (N_20210,N_17887,N_19250);
nor U20211 (N_20211,N_19877,N_17690);
and U20212 (N_20212,N_17648,N_18881);
or U20213 (N_20213,N_17608,N_18406);
or U20214 (N_20214,N_18900,N_17932);
xnor U20215 (N_20215,N_19464,N_18307);
nor U20216 (N_20216,N_17848,N_19931);
nor U20217 (N_20217,N_17711,N_17667);
nor U20218 (N_20218,N_18868,N_19160);
and U20219 (N_20219,N_19061,N_18463);
or U20220 (N_20220,N_17823,N_19085);
nand U20221 (N_20221,N_19210,N_18268);
and U20222 (N_20222,N_17930,N_18379);
and U20223 (N_20223,N_18175,N_19967);
or U20224 (N_20224,N_18855,N_18358);
xnor U20225 (N_20225,N_19833,N_19852);
nor U20226 (N_20226,N_17783,N_18048);
xor U20227 (N_20227,N_18516,N_18791);
xor U20228 (N_20228,N_18467,N_18835);
nor U20229 (N_20229,N_19555,N_19569);
nand U20230 (N_20230,N_17954,N_19139);
nor U20231 (N_20231,N_18929,N_18568);
nand U20232 (N_20232,N_19475,N_17747);
and U20233 (N_20233,N_19776,N_19613);
or U20234 (N_20234,N_19380,N_17682);
and U20235 (N_20235,N_18153,N_19384);
xor U20236 (N_20236,N_18482,N_17888);
nor U20237 (N_20237,N_19958,N_18785);
xnor U20238 (N_20238,N_18534,N_19668);
and U20239 (N_20239,N_19177,N_18888);
nor U20240 (N_20240,N_19780,N_18385);
nand U20241 (N_20241,N_18492,N_17616);
nand U20242 (N_20242,N_19441,N_17680);
or U20243 (N_20243,N_18953,N_19342);
and U20244 (N_20244,N_19751,N_18802);
nand U20245 (N_20245,N_19788,N_18147);
or U20246 (N_20246,N_19784,N_19935);
or U20247 (N_20247,N_18194,N_19281);
xor U20248 (N_20248,N_19069,N_17845);
and U20249 (N_20249,N_18892,N_19491);
or U20250 (N_20250,N_19914,N_18014);
nor U20251 (N_20251,N_18346,N_19373);
and U20252 (N_20252,N_19646,N_19472);
or U20253 (N_20253,N_19915,N_17674);
or U20254 (N_20254,N_19433,N_19129);
and U20255 (N_20255,N_17861,N_19983);
and U20256 (N_20256,N_19907,N_19452);
nand U20257 (N_20257,N_17993,N_19298);
nand U20258 (N_20258,N_17637,N_19270);
xor U20259 (N_20259,N_17858,N_19671);
nand U20260 (N_20260,N_18952,N_18027);
xnor U20261 (N_20261,N_18659,N_18056);
nand U20262 (N_20262,N_19293,N_19398);
nor U20263 (N_20263,N_18774,N_18740);
nor U20264 (N_20264,N_17693,N_19872);
xor U20265 (N_20265,N_19511,N_19261);
nor U20266 (N_20266,N_18668,N_19328);
xor U20267 (N_20267,N_18415,N_17710);
or U20268 (N_20268,N_19769,N_17664);
nand U20269 (N_20269,N_19154,N_18648);
or U20270 (N_20270,N_18160,N_19179);
and U20271 (N_20271,N_19035,N_18822);
or U20272 (N_20272,N_19460,N_19574);
nor U20273 (N_20273,N_19421,N_17874);
xor U20274 (N_20274,N_17723,N_18157);
nor U20275 (N_20275,N_18909,N_17552);
and U20276 (N_20276,N_18591,N_19397);
nand U20277 (N_20277,N_19396,N_18920);
nor U20278 (N_20278,N_19502,N_18963);
xor U20279 (N_20279,N_18574,N_19473);
or U20280 (N_20280,N_18563,N_17589);
xnor U20281 (N_20281,N_19887,N_18386);
and U20282 (N_20282,N_19162,N_19104);
or U20283 (N_20283,N_18272,N_19766);
nand U20284 (N_20284,N_18343,N_18208);
nand U20285 (N_20285,N_19546,N_19847);
and U20286 (N_20286,N_18453,N_18246);
nor U20287 (N_20287,N_19909,N_17782);
nor U20288 (N_20288,N_18166,N_17988);
or U20289 (N_20289,N_19309,N_19484);
or U20290 (N_20290,N_19884,N_19791);
nor U20291 (N_20291,N_18850,N_19663);
and U20292 (N_20292,N_18592,N_17779);
nand U20293 (N_20293,N_19340,N_18264);
or U20294 (N_20294,N_19820,N_17724);
or U20295 (N_20295,N_18389,N_19614);
and U20296 (N_20296,N_18095,N_19512);
nor U20297 (N_20297,N_19536,N_19823);
nor U20298 (N_20298,N_18291,N_17818);
nor U20299 (N_20299,N_18940,N_18351);
or U20300 (N_20300,N_18238,N_19191);
nor U20301 (N_20301,N_18185,N_18501);
xnor U20302 (N_20302,N_19370,N_19330);
and U20303 (N_20303,N_17922,N_18199);
and U20304 (N_20304,N_19514,N_18566);
xnor U20305 (N_20305,N_18731,N_19828);
or U20306 (N_20306,N_19133,N_18603);
and U20307 (N_20307,N_19738,N_18103);
and U20308 (N_20308,N_19416,N_19140);
nand U20309 (N_20309,N_17691,N_17530);
xor U20310 (N_20310,N_18126,N_19974);
nand U20311 (N_20311,N_17513,N_17520);
and U20312 (N_20312,N_19763,N_18795);
nand U20313 (N_20313,N_19643,N_18596);
nand U20314 (N_20314,N_17638,N_18934);
xnor U20315 (N_20315,N_17879,N_18871);
and U20316 (N_20316,N_19942,N_18580);
nand U20317 (N_20317,N_18532,N_19337);
xor U20318 (N_20318,N_18226,N_18139);
xnor U20319 (N_20319,N_19048,N_17654);
xor U20320 (N_20320,N_17541,N_19188);
and U20321 (N_20321,N_17559,N_19773);
and U20322 (N_20322,N_17904,N_18152);
nand U20323 (N_20323,N_18032,N_17855);
nor U20324 (N_20324,N_18365,N_19381);
nand U20325 (N_20325,N_18770,N_17743);
and U20326 (N_20326,N_18388,N_17696);
nor U20327 (N_20327,N_17560,N_19840);
and U20328 (N_20328,N_19449,N_18545);
and U20329 (N_20329,N_19720,N_18174);
xor U20330 (N_20330,N_18364,N_18979);
nand U20331 (N_20331,N_18971,N_18367);
or U20332 (N_20332,N_18615,N_18292);
and U20333 (N_20333,N_19801,N_19937);
nor U20334 (N_20334,N_18030,N_18676);
or U20335 (N_20335,N_19885,N_18589);
nor U20336 (N_20336,N_18217,N_19658);
and U20337 (N_20337,N_18813,N_19781);
nand U20338 (N_20338,N_17713,N_18769);
xor U20339 (N_20339,N_18408,N_18675);
or U20340 (N_20340,N_17566,N_19848);
nand U20341 (N_20341,N_18672,N_19950);
xor U20342 (N_20342,N_19183,N_19739);
or U20343 (N_20343,N_19036,N_17986);
xnor U20344 (N_20344,N_17806,N_19567);
nand U20345 (N_20345,N_19831,N_18702);
or U20346 (N_20346,N_19258,N_17567);
or U20347 (N_20347,N_18981,N_19238);
nand U20348 (N_20348,N_19410,N_18794);
xor U20349 (N_20349,N_18706,N_18906);
and U20350 (N_20350,N_19584,N_19201);
xor U20351 (N_20351,N_19091,N_19505);
xor U20352 (N_20352,N_18968,N_18052);
and U20353 (N_20353,N_18397,N_18723);
nor U20354 (N_20354,N_17974,N_18690);
nand U20355 (N_20355,N_19897,N_17781);
or U20356 (N_20356,N_19839,N_17555);
and U20357 (N_20357,N_17767,N_19053);
or U20358 (N_20358,N_19866,N_17945);
or U20359 (N_20359,N_19796,N_19553);
or U20360 (N_20360,N_18914,N_18999);
nor U20361 (N_20361,N_19895,N_18222);
nand U20362 (N_20362,N_18939,N_19732);
or U20363 (N_20363,N_18223,N_19101);
nor U20364 (N_20364,N_18699,N_19110);
xor U20365 (N_20365,N_17824,N_19237);
and U20366 (N_20366,N_18078,N_19735);
nand U20367 (N_20367,N_18436,N_17908);
nand U20368 (N_20368,N_18645,N_19622);
or U20369 (N_20369,N_19869,N_17576);
nor U20370 (N_20370,N_17898,N_17676);
or U20371 (N_20371,N_19680,N_19456);
or U20372 (N_20372,N_18183,N_18125);
nor U20373 (N_20373,N_19603,N_18738);
nor U20374 (N_20374,N_19468,N_18209);
xor U20375 (N_20375,N_19499,N_17927);
nand U20376 (N_20376,N_18105,N_19992);
nand U20377 (N_20377,N_18277,N_17500);
nand U20378 (N_20378,N_19303,N_17746);
nor U20379 (N_20379,N_19311,N_17734);
nor U20380 (N_20380,N_18069,N_17961);
nor U20381 (N_20381,N_17706,N_18380);
and U20382 (N_20382,N_19509,N_19334);
nand U20383 (N_20383,N_17775,N_18197);
or U20384 (N_20384,N_19630,N_17645);
or U20385 (N_20385,N_18637,N_18712);
and U20386 (N_20386,N_17545,N_19962);
or U20387 (N_20387,N_17812,N_19109);
or U20388 (N_20388,N_19770,N_18975);
nand U20389 (N_20389,N_18778,N_19100);
and U20390 (N_20390,N_19096,N_18141);
xnor U20391 (N_20391,N_18893,N_18520);
or U20392 (N_20392,N_18755,N_18886);
or U20393 (N_20393,N_19538,N_19605);
nor U20394 (N_20394,N_19322,N_18985);
nand U20395 (N_20395,N_18293,N_18314);
nor U20396 (N_20396,N_18483,N_18633);
nand U20397 (N_20397,N_19021,N_17622);
or U20398 (N_20398,N_19481,N_18454);
nor U20399 (N_20399,N_17554,N_19856);
or U20400 (N_20400,N_18412,N_19244);
nand U20401 (N_20401,N_18047,N_19489);
or U20402 (N_20402,N_18652,N_19187);
or U20403 (N_20403,N_18190,N_18335);
or U20404 (N_20404,N_18378,N_18512);
xor U20405 (N_20405,N_19012,N_19708);
or U20406 (N_20406,N_18375,N_19461);
or U20407 (N_20407,N_19369,N_19917);
xor U20408 (N_20408,N_17935,N_17836);
xor U20409 (N_20409,N_18609,N_18248);
nor U20410 (N_20410,N_17737,N_18911);
nor U20411 (N_20411,N_19178,N_18213);
xnor U20412 (N_20412,N_18679,N_18345);
and U20413 (N_20413,N_19117,N_19515);
nor U20414 (N_20414,N_19134,N_19637);
xor U20415 (N_20415,N_18101,N_19762);
and U20416 (N_20416,N_17628,N_18338);
xnor U20417 (N_20417,N_19193,N_19182);
xnor U20418 (N_20418,N_18198,N_18179);
xor U20419 (N_20419,N_17708,N_19944);
xor U20420 (N_20420,N_19492,N_19767);
and U20421 (N_20421,N_19633,N_18649);
xnor U20422 (N_20422,N_19901,N_17984);
nand U20423 (N_20423,N_18167,N_19383);
xor U20424 (N_20424,N_18553,N_18352);
and U20425 (N_20425,N_19273,N_18355);
nand U20426 (N_20426,N_19321,N_19903);
nor U20427 (N_20427,N_17780,N_19073);
xor U20428 (N_20428,N_19625,N_18678);
nor U20429 (N_20429,N_19689,N_17998);
and U20430 (N_20430,N_18689,N_19777);
or U20431 (N_20431,N_18719,N_18083);
nor U20432 (N_20432,N_19205,N_19746);
xor U20433 (N_20433,N_19636,N_17665);
nor U20434 (N_20434,N_19485,N_18558);
nand U20435 (N_20435,N_19861,N_19927);
and U20436 (N_20436,N_18634,N_18510);
and U20437 (N_20437,N_19793,N_19447);
and U20438 (N_20438,N_19127,N_19757);
nand U20439 (N_20439,N_19463,N_18480);
or U20440 (N_20440,N_18681,N_19696);
nor U20441 (N_20441,N_18961,N_19810);
xor U20442 (N_20442,N_19253,N_18599);
and U20443 (N_20443,N_18043,N_19458);
nand U20444 (N_20444,N_18720,N_18200);
nand U20445 (N_20445,N_19690,N_18853);
nor U20446 (N_20446,N_18544,N_18049);
and U20447 (N_20447,N_18165,N_19756);
nor U20448 (N_20448,N_19808,N_17523);
xor U20449 (N_20449,N_18455,N_18995);
xor U20450 (N_20450,N_19644,N_19835);
nor U20451 (N_20451,N_17700,N_19719);
xor U20452 (N_20452,N_19482,N_19064);
nor U20453 (N_20453,N_18279,N_19789);
nand U20454 (N_20454,N_18202,N_19455);
xnor U20455 (N_20455,N_18604,N_19890);
xnor U20456 (N_20456,N_17593,N_18613);
nor U20457 (N_20457,N_19470,N_19400);
or U20458 (N_20458,N_19271,N_17603);
xor U20459 (N_20459,N_18821,N_17915);
nor U20460 (N_20460,N_17839,N_19704);
and U20461 (N_20461,N_19471,N_19954);
nor U20462 (N_20462,N_18146,N_19973);
and U20463 (N_20463,N_17685,N_18489);
xor U20464 (N_20464,N_19961,N_19598);
xor U20465 (N_20465,N_19158,N_18787);
nand U20466 (N_20466,N_18372,N_19873);
xnor U20467 (N_20467,N_19612,N_19478);
and U20468 (N_20468,N_18586,N_18045);
nor U20469 (N_20469,N_17817,N_19361);
nand U20470 (N_20470,N_19640,N_19483);
and U20471 (N_20471,N_19078,N_18684);
and U20472 (N_20472,N_19394,N_19764);
or U20473 (N_20473,N_19075,N_19344);
xnor U20474 (N_20474,N_19058,N_18825);
and U20475 (N_20475,N_18326,N_18546);
nor U20476 (N_20476,N_19056,N_19772);
xnor U20477 (N_20477,N_17979,N_17569);
xor U20478 (N_20478,N_18521,N_17983);
nor U20479 (N_20479,N_18874,N_19565);
nand U20480 (N_20480,N_18977,N_17744);
nor U20481 (N_20481,N_19317,N_18211);
nor U20482 (N_20482,N_19024,N_17840);
nand U20483 (N_20483,N_18526,N_17968);
and U20484 (N_20484,N_18815,N_17633);
or U20485 (N_20485,N_17725,N_19661);
nand U20486 (N_20486,N_17595,N_17618);
nand U20487 (N_20487,N_18858,N_17583);
nor U20488 (N_20488,N_19585,N_17542);
nand U20489 (N_20489,N_18925,N_18163);
xnor U20490 (N_20490,N_18461,N_18322);
xor U20491 (N_20491,N_19439,N_19112);
and U20492 (N_20492,N_17641,N_17581);
nand U20493 (N_20493,N_17844,N_19867);
and U20494 (N_20494,N_18058,N_19254);
or U20495 (N_20495,N_19818,N_19849);
and U20496 (N_20496,N_18000,N_19137);
and U20497 (N_20497,N_19020,N_18715);
xor U20498 (N_20498,N_19375,N_17760);
nand U20499 (N_20499,N_19286,N_19786);
nand U20500 (N_20500,N_17709,N_19540);
nand U20501 (N_20501,N_19016,N_17778);
xor U20502 (N_20502,N_18320,N_18955);
nor U20503 (N_20503,N_19147,N_18162);
nand U20504 (N_20504,N_18879,N_17683);
nor U20505 (N_20505,N_18646,N_18053);
xor U20506 (N_20506,N_19545,N_19864);
nand U20507 (N_20507,N_18445,N_18717);
nor U20508 (N_20508,N_18518,N_19282);
nor U20509 (N_20509,N_19418,N_17573);
nor U20510 (N_20510,N_19623,N_18620);
and U20511 (N_20511,N_19049,N_18965);
or U20512 (N_20512,N_17558,N_19602);
xor U20513 (N_20513,N_19865,N_18647);
xor U20514 (N_20514,N_18254,N_17850);
or U20515 (N_20515,N_19889,N_18290);
xnor U20516 (N_20516,N_19945,N_18064);
nand U20517 (N_20517,N_18536,N_19621);
and U20518 (N_20518,N_18873,N_17661);
xnor U20519 (N_20519,N_19263,N_17784);
xor U20520 (N_20520,N_19348,N_18164);
and U20521 (N_20521,N_19617,N_19138);
xor U20522 (N_20522,N_17524,N_17797);
xnor U20523 (N_20523,N_17911,N_18019);
or U20524 (N_20524,N_17987,N_19905);
nor U20525 (N_20525,N_18232,N_19413);
nand U20526 (N_20526,N_19066,N_17786);
nor U20527 (N_20527,N_18924,N_19754);
or U20528 (N_20528,N_19459,N_17717);
xor U20529 (N_20529,N_18302,N_18782);
nand U20530 (N_20530,N_18598,N_18695);
nand U20531 (N_20531,N_17941,N_18333);
nor U20532 (N_20532,N_19929,N_17539);
xor U20533 (N_20533,N_19023,N_18234);
or U20534 (N_20534,N_19315,N_17557);
or U20535 (N_20535,N_18169,N_19026);
nor U20536 (N_20536,N_18607,N_17869);
or U20537 (N_20537,N_18131,N_18274);
or U20538 (N_20538,N_19022,N_18974);
or U20539 (N_20539,N_18733,N_19844);
xnor U20540 (N_20540,N_19530,N_18551);
xor U20541 (N_20541,N_17966,N_18270);
and U20542 (N_20542,N_17653,N_19924);
and U20543 (N_20543,N_18554,N_19331);
nand U20544 (N_20544,N_19996,N_19528);
or U20545 (N_20545,N_19089,N_19457);
nand U20546 (N_20546,N_19428,N_18632);
xnor U20547 (N_20547,N_18915,N_19186);
xnor U20548 (N_20548,N_17596,N_18789);
nand U20549 (N_20549,N_18781,N_17697);
and U20550 (N_20550,N_19678,N_18506);
and U20551 (N_20551,N_18707,N_18856);
nor U20552 (N_20552,N_18587,N_19723);
or U20553 (N_20553,N_17634,N_17916);
or U20554 (N_20554,N_19462,N_19255);
xnor U20555 (N_20555,N_17738,N_18870);
or U20556 (N_20556,N_19759,N_17590);
and U20557 (N_20557,N_17591,N_17859);
or U20558 (N_20558,N_19677,N_18362);
nand U20559 (N_20559,N_19548,N_18340);
or U20560 (N_20560,N_17771,N_19355);
or U20561 (N_20561,N_18962,N_19562);
nor U20562 (N_20562,N_19734,N_18299);
xnor U20563 (N_20563,N_19296,N_18764);
and U20564 (N_20564,N_19043,N_17512);
or U20565 (N_20565,N_17885,N_19707);
and U20566 (N_20566,N_18724,N_19564);
nand U20567 (N_20567,N_19670,N_19660);
and U20568 (N_20568,N_17884,N_19288);
or U20569 (N_20569,N_18757,N_19948);
or U20570 (N_20570,N_17923,N_19900);
nand U20571 (N_20571,N_18772,N_18865);
and U20572 (N_20572,N_19412,N_19600);
nand U20573 (N_20573,N_19076,N_19225);
xnor U20574 (N_20574,N_19040,N_19516);
nand U20575 (N_20575,N_18932,N_19932);
xnor U20576 (N_20576,N_17870,N_19593);
or U20577 (N_20577,N_19338,N_17668);
xor U20578 (N_20578,N_19445,N_18460);
or U20579 (N_20579,N_17597,N_19656);
xnor U20580 (N_20580,N_18228,N_18666);
nand U20581 (N_20581,N_19648,N_18593);
nor U20582 (N_20582,N_18555,N_18084);
nor U20583 (N_20583,N_19804,N_19693);
and U20584 (N_20584,N_17600,N_18989);
nand U20585 (N_20585,N_19417,N_18542);
nand U20586 (N_20586,N_18579,N_19940);
or U20587 (N_20587,N_19223,N_17514);
and U20588 (N_20588,N_19980,N_18168);
nand U20589 (N_20589,N_19799,N_18826);
nor U20590 (N_20590,N_17865,N_18828);
nor U20591 (N_20591,N_19779,N_18082);
nor U20592 (N_20592,N_17733,N_19713);
and U20593 (N_20593,N_18673,N_17936);
nor U20594 (N_20594,N_18171,N_18796);
xnor U20595 (N_20595,N_18857,N_17613);
nor U20596 (N_20596,N_19236,N_18094);
nor U20597 (N_20597,N_18219,N_19624);
xnor U20598 (N_20598,N_18494,N_19387);
xnor U20599 (N_20599,N_17532,N_18931);
or U20600 (N_20600,N_17547,N_17677);
nand U20601 (N_20601,N_17572,N_19214);
xor U20602 (N_20602,N_18771,N_19208);
nand U20603 (N_20603,N_18148,N_19652);
nor U20604 (N_20604,N_18187,N_19557);
nand U20605 (N_20605,N_18334,N_18124);
nor U20606 (N_20606,N_19359,N_17919);
nand U20607 (N_20607,N_19057,N_17720);
nor U20608 (N_20608,N_19815,N_17602);
or U20609 (N_20609,N_19743,N_18119);
or U20610 (N_20610,N_19993,N_18450);
xnor U20611 (N_20611,N_19376,N_19906);
nand U20612 (N_20612,N_17877,N_17536);
nor U20613 (N_20613,N_19800,N_18286);
xnor U20614 (N_20614,N_18350,N_18973);
and U20615 (N_20615,N_17962,N_19667);
nand U20616 (N_20616,N_18509,N_17834);
and U20617 (N_20617,N_19207,N_18751);
and U20618 (N_20618,N_18294,N_19292);
and U20619 (N_20619,N_17891,N_19700);
nand U20620 (N_20620,N_18128,N_17754);
xor U20621 (N_20621,N_17890,N_18075);
and U20622 (N_20622,N_18416,N_18422);
nor U20623 (N_20623,N_19971,N_18864);
and U20624 (N_20624,N_18411,N_18465);
xor U20625 (N_20625,N_19390,N_19846);
and U20626 (N_20626,N_18245,N_18204);
nor U20627 (N_20627,N_17846,N_18849);
nand U20628 (N_20628,N_17505,N_17975);
and U20629 (N_20629,N_18296,N_18588);
and U20630 (N_20630,N_18097,N_18252);
xor U20631 (N_20631,N_19688,N_18507);
or U20632 (N_20632,N_18800,N_19817);
or U20633 (N_20633,N_19495,N_17763);
or U20634 (N_20634,N_17872,N_18305);
nor U20635 (N_20635,N_19879,N_17630);
or U20636 (N_20636,N_19000,N_19017);
or U20637 (N_20637,N_19893,N_19665);
or U20638 (N_20638,N_17862,N_19180);
and U20639 (N_20639,N_18298,N_19146);
or U20640 (N_20640,N_18425,N_18576);
and U20641 (N_20641,N_18811,N_18638);
xnor U20642 (N_20642,N_18479,N_18282);
xnor U20643 (N_20643,N_19741,N_17982);
nand U20644 (N_20644,N_18437,N_19368);
or U20645 (N_20645,N_19552,N_17929);
and U20646 (N_20646,N_17656,N_19265);
nand U20647 (N_20647,N_18370,N_19389);
xor U20648 (N_20648,N_19323,N_18390);
and U20649 (N_20649,N_18745,N_18556);
or U20650 (N_20650,N_18631,N_17906);
xor U20651 (N_20651,N_18395,N_18984);
and U20652 (N_20652,N_18816,N_18667);
nor U20653 (N_20653,N_17719,N_19547);
and U20654 (N_20654,N_18805,N_17832);
and U20655 (N_20655,N_18227,N_18663);
nand U20656 (N_20656,N_17531,N_17790);
or U20657 (N_20657,N_18773,N_18606);
nor U20658 (N_20658,N_18937,N_19382);
nand U20659 (N_20659,N_18396,N_18683);
xnor U20660 (N_20660,N_18758,N_18523);
xor U20661 (N_20661,N_19122,N_19289);
nand U20662 (N_20662,N_18267,N_18957);
or U20663 (N_20663,N_18414,N_19853);
or U20664 (N_20664,N_19014,N_19782);
nand U20665 (N_20665,N_19203,N_19539);
or U20666 (N_20666,N_17701,N_18639);
or U20667 (N_20667,N_19526,N_17992);
or U20668 (N_20668,N_17561,N_19071);
nor U20669 (N_20669,N_18374,N_18448);
nand U20670 (N_20670,N_18004,N_19834);
or U20671 (N_20671,N_19631,N_18215);
xnor U20672 (N_20672,N_18449,N_19662);
or U20673 (N_20673,N_18363,N_18261);
nor U20674 (N_20674,N_19749,N_17910);
nand U20675 (N_20675,N_17548,N_19259);
nor U20676 (N_20676,N_18173,N_18866);
or U20677 (N_20677,N_19045,N_18619);
nor U20678 (N_20678,N_17735,N_19332);
or U20679 (N_20679,N_19157,N_19278);
nand U20680 (N_20680,N_19729,N_18026);
or U20681 (N_20681,N_18419,N_19190);
and U20682 (N_20682,N_17617,N_19039);
xor U20683 (N_20683,N_17880,N_18493);
xnor U20684 (N_20684,N_18181,N_18201);
nand U20685 (N_20685,N_19033,N_18852);
and U20686 (N_20686,N_19634,N_17853);
xnor U20687 (N_20687,N_19761,N_18700);
or U20688 (N_20688,N_18116,N_17694);
nand U20689 (N_20689,N_17516,N_18025);
or U20690 (N_20690,N_18013,N_18113);
xnor U20691 (N_20691,N_17946,N_18983);
xnor U20692 (N_20692,N_18533,N_17605);
and U20693 (N_20693,N_18471,N_17736);
or U20694 (N_20694,N_19095,N_19803);
nand U20695 (N_20695,N_19806,N_18970);
or U20696 (N_20696,N_18714,N_18867);
nor U20697 (N_20697,N_19838,N_18643);
or U20698 (N_20698,N_19249,N_18761);
nand U20699 (N_20699,N_18966,N_19149);
xnor U20700 (N_20700,N_19896,N_19081);
nor U20701 (N_20701,N_17978,N_19982);
or U20702 (N_20702,N_18423,N_19578);
nand U20703 (N_20703,N_17907,N_19194);
or U20704 (N_20704,N_17795,N_19830);
nor U20705 (N_20705,N_18701,N_19378);
and U20706 (N_20706,N_18921,N_19619);
or U20707 (N_20707,N_17527,N_18927);
or U20708 (N_20708,N_19159,N_17873);
or U20709 (N_20709,N_19451,N_17995);
and U20710 (N_20710,N_17777,N_19431);
and U20711 (N_20711,N_18426,N_19532);
nand U20712 (N_20712,N_19701,N_18134);
nand U20713 (N_20713,N_19031,N_18595);
or U20714 (N_20714,N_18549,N_19976);
and U20715 (N_20715,N_18812,N_19813);
and U20716 (N_20716,N_18062,N_18913);
nand U20717 (N_20717,N_17604,N_19346);
and U20718 (N_20718,N_18067,N_19403);
and U20719 (N_20719,N_18692,N_18003);
nor U20720 (N_20720,N_18624,N_18766);
nor U20721 (N_20721,N_18535,N_19310);
and U20722 (N_20722,N_17999,N_19090);
nor U20723 (N_20723,N_18616,N_19200);
or U20724 (N_20724,N_18111,N_19591);
xor U20725 (N_20725,N_17611,N_18469);
xnor U20726 (N_20726,N_18021,N_19466);
nor U20727 (N_20727,N_18225,N_19995);
xor U20728 (N_20728,N_19283,N_19563);
xor U20729 (N_20729,N_18949,N_19032);
xor U20730 (N_20730,N_17955,N_17921);
and U20731 (N_20731,N_18783,N_19596);
xnor U20732 (N_20732,N_18262,N_19079);
nor U20733 (N_20733,N_17640,N_18741);
nor U20734 (N_20734,N_19156,N_18926);
xnor U20735 (N_20735,N_17675,N_19174);
or U20736 (N_20736,N_18203,N_19519);
nand U20737 (N_20737,N_18137,N_19698);
and U20738 (N_20738,N_17652,N_18573);
and U20739 (N_20739,N_19736,N_18432);
nand U20740 (N_20740,N_19711,N_17814);
or U20741 (N_20741,N_19731,N_19143);
nand U20742 (N_20742,N_19920,N_19164);
or U20743 (N_20743,N_18108,N_18674);
nor U20744 (N_20744,N_19758,N_18086);
or U20745 (N_20745,N_18329,N_18178);
nand U20746 (N_20746,N_17980,N_17791);
nor U20747 (N_20747,N_19047,N_19984);
or U20748 (N_20748,N_19357,N_17658);
and U20749 (N_20749,N_18410,N_17920);
xor U20750 (N_20750,N_17939,N_17985);
or U20751 (N_20751,N_19521,N_19161);
nor U20752 (N_20752,N_18572,N_19124);
nand U20753 (N_20753,N_18318,N_19725);
and U20754 (N_20754,N_19004,N_18836);
xor U20755 (N_20755,N_17949,N_18464);
nand U20756 (N_20756,N_18117,N_18916);
and U20757 (N_20757,N_19946,N_19185);
nand U20758 (N_20758,N_18055,N_19103);
xnor U20759 (N_20759,N_19912,N_18861);
nor U20760 (N_20760,N_18803,N_17882);
and U20761 (N_20761,N_18860,N_17749);
xor U20762 (N_20762,N_19010,N_18847);
or U20763 (N_20763,N_18316,N_19077);
xor U20764 (N_20764,N_19204,N_17588);
and U20765 (N_20765,N_19604,N_18006);
or U20766 (N_20766,N_17994,N_18622);
nor U20767 (N_20767,N_17820,N_19685);
nor U20768 (N_20768,N_17996,N_19755);
nand U20769 (N_20769,N_17905,N_19797);
nor U20770 (N_20770,N_19349,N_17579);
nand U20771 (N_20771,N_19892,N_18749);
xnor U20772 (N_20772,N_19606,N_17897);
nor U20773 (N_20773,N_17679,N_19226);
nor U20774 (N_20774,N_18258,N_18438);
and U20775 (N_20775,N_19088,N_17819);
and U20776 (N_20776,N_17934,N_19438);
nor U20777 (N_20777,N_18682,N_18705);
or U20778 (N_20778,N_19572,N_18186);
nand U20779 (N_20779,N_17960,N_19083);
or U20780 (N_20780,N_18304,N_18361);
and U20781 (N_20781,N_19131,N_18281);
nor U20782 (N_20782,N_18325,N_18051);
nor U20783 (N_20783,N_18005,N_18283);
or U20784 (N_20784,N_19951,N_19898);
xor U20785 (N_20785,N_17551,N_19615);
and U20786 (N_20786,N_18779,N_19218);
and U20787 (N_20787,N_18833,N_18257);
xor U20788 (N_20788,N_18843,N_17606);
xor U20789 (N_20789,N_18490,N_18150);
or U20790 (N_20790,N_17731,N_17704);
xnor U20791 (N_20791,N_18458,N_18196);
nand U20792 (N_20792,N_18231,N_18680);
or U20793 (N_20793,N_18511,N_19529);
nand U20794 (N_20794,N_19837,N_19220);
nand U20795 (N_20795,N_17883,N_19714);
and U20796 (N_20796,N_18502,N_19111);
or U20797 (N_20797,N_19243,N_19274);
xor U20798 (N_20798,N_19299,N_18605);
or U20799 (N_20799,N_17636,N_19385);
and U20800 (N_20800,N_18180,N_18009);
nand U20801 (N_20801,N_17543,N_17506);
xor U20802 (N_20802,N_17594,N_18499);
nor U20803 (N_20803,N_19319,N_18602);
or U20804 (N_20804,N_18967,N_17957);
nor U20805 (N_20805,N_19307,N_19812);
or U20806 (N_20806,N_19037,N_17519);
nand U20807 (N_20807,N_19125,N_18830);
and U20808 (N_20808,N_19437,N_18285);
nand U20809 (N_20809,N_19027,N_19609);
or U20810 (N_20810,N_18312,N_19312);
nor U20811 (N_20811,N_18990,N_18776);
or U20812 (N_20812,N_19716,N_18373);
xor U20813 (N_20813,N_19537,N_17501);
nor U20814 (N_20814,N_19775,N_18066);
xnor U20815 (N_20815,N_18477,N_18947);
or U20816 (N_20816,N_17755,N_18908);
xor U20817 (N_20817,N_19341,N_17695);
nand U20818 (N_20818,N_19054,N_18528);
and U20819 (N_20819,N_19335,N_19809);
xnor U20820 (N_20820,N_19868,N_17913);
xor U20821 (N_20821,N_18077,N_19392);
and U20822 (N_20822,N_17503,N_17525);
or U20823 (N_20823,N_17925,N_19405);
or U20824 (N_20824,N_19454,N_18121);
nand U20825 (N_20825,N_18273,N_19490);
and U20826 (N_20826,N_18880,N_19222);
nor U20827 (N_20827,N_18184,N_18514);
and U20828 (N_20828,N_18527,N_17852);
or U20829 (N_20829,N_18243,N_18485);
or U20830 (N_20830,N_17644,N_18629);
or U20831 (N_20831,N_17822,N_19498);
or U20832 (N_20832,N_19118,N_18945);
nor U20833 (N_20833,N_18300,N_18842);
nand U20834 (N_20834,N_18882,N_18265);
and U20835 (N_20835,N_19429,N_18994);
nor U20836 (N_20836,N_19029,N_17972);
nand U20837 (N_20837,N_19964,N_18583);
nand U20838 (N_20838,N_18737,N_19065);
and U20839 (N_20839,N_17951,N_19908);
and U20840 (N_20840,N_19860,N_18951);
and U20841 (N_20841,N_18767,N_19508);
nor U20842 (N_20842,N_19975,N_17854);
and U20843 (N_20843,N_19232,N_19966);
and U20844 (N_20844,N_19256,N_19329);
and U20845 (N_20845,N_19324,N_17952);
nor U20846 (N_20846,N_18114,N_18565);
nor U20847 (N_20847,N_18948,N_19504);
xor U20848 (N_20848,N_18907,N_18513);
nand U20849 (N_20849,N_19952,N_18159);
nand U20850 (N_20850,N_18155,N_19987);
or U20851 (N_20851,N_18810,N_18042);
and U20852 (N_20852,N_19561,N_19675);
and U20853 (N_20853,N_19841,N_19116);
nand U20854 (N_20854,N_18608,N_19629);
or U20855 (N_20855,N_17721,N_19229);
nand U20856 (N_20856,N_18987,N_18540);
nor U20857 (N_20857,N_18760,N_18327);
xor U20858 (N_20858,N_19571,N_17741);
and U20859 (N_20859,N_18877,N_19175);
nor U20860 (N_20860,N_19301,N_19257);
nor U20861 (N_20861,N_19765,N_18577);
xor U20862 (N_20862,N_18221,N_18734);
xnor U20863 (N_20863,N_18696,N_17546);
xor U20864 (N_20864,N_19184,N_18093);
nand U20865 (N_20865,N_18387,N_19531);
nor U20866 (N_20866,N_19787,N_19195);
nor U20867 (N_20867,N_18635,N_18614);
nand U20868 (N_20868,N_18775,N_19798);
or U20869 (N_20869,N_17860,N_19988);
nor U20870 (N_20870,N_19938,N_17969);
xor U20871 (N_20871,N_19166,N_19664);
xnor U20872 (N_20872,N_18942,N_17757);
or U20873 (N_20873,N_18430,N_19575);
nor U20874 (N_20874,N_19836,N_18177);
xnor U20875 (N_20875,N_19444,N_18959);
nor U20876 (N_20876,N_19888,N_18743);
or U20877 (N_20877,N_17550,N_18418);
nor U20878 (N_20878,N_18564,N_19645);
and U20879 (N_20879,N_17511,N_17893);
nand U20880 (N_20880,N_19916,N_18250);
nor U20881 (N_20881,N_19087,N_19365);
or U20882 (N_20882,N_18997,N_19883);
nand U20883 (N_20883,N_18233,N_18538);
nor U20884 (N_20884,N_18765,N_19851);
nand U20885 (N_20885,N_19302,N_19494);
or U20886 (N_20886,N_18001,N_19121);
and U20887 (N_20887,N_18784,N_19336);
and U20888 (N_20888,N_19497,N_19939);
nor U20889 (N_20889,N_19737,N_17753);
xor U20890 (N_20890,N_19167,N_19989);
xor U20891 (N_20891,N_17959,N_18401);
nor U20892 (N_20892,N_17794,N_18636);
and U20893 (N_20893,N_17742,N_18889);
nand U20894 (N_20894,N_19404,N_19423);
nor U20895 (N_20895,N_17647,N_18728);
and U20896 (N_20896,N_18306,N_18297);
xnor U20897 (N_20897,N_17728,N_18630);
nor U20898 (N_20898,N_18768,N_18391);
nand U20899 (N_20899,N_19358,N_18848);
or U20900 (N_20900,N_18883,N_18321);
and U20901 (N_20901,N_19224,N_17650);
or U20902 (N_20902,N_18722,N_18205);
and U20903 (N_20903,N_18844,N_18404);
nand U20904 (N_20904,N_18035,N_19886);
and U20905 (N_20905,N_17967,N_17971);
xnor U20906 (N_20906,N_18919,N_18590);
nor U20907 (N_20907,N_18073,N_17837);
and U20908 (N_20908,N_19858,N_17599);
nand U20909 (N_20909,N_17687,N_19965);
or U20910 (N_20910,N_19774,N_18730);
nand U20911 (N_20911,N_17587,N_19202);
nand U20912 (N_20912,N_18136,N_17521);
and U20913 (N_20913,N_17686,N_17510);
xnor U20914 (N_20914,N_18347,N_19262);
nor U20915 (N_20915,N_17997,N_19042);
and U20916 (N_20916,N_18875,N_19981);
or U20917 (N_20917,N_18288,N_19176);
nand U20918 (N_20918,N_19051,N_18664);
nor U20919 (N_20919,N_19215,N_18621);
or U20920 (N_20920,N_17642,N_18301);
or U20921 (N_20921,N_18218,N_17964);
xnor U20922 (N_20922,N_19038,N_19541);
nand U20923 (N_20923,N_19618,N_19277);
and U20924 (N_20924,N_19933,N_18154);
or U20925 (N_20925,N_18251,N_18102);
nor U20926 (N_20926,N_19272,N_19607);
nor U20927 (N_20927,N_19953,N_18303);
nor U20928 (N_20928,N_18531,N_19055);
xnor U20929 (N_20929,N_18470,N_19904);
and U20930 (N_20930,N_18191,N_19978);
nor U20931 (N_20931,N_17796,N_18242);
nor U20932 (N_20932,N_19267,N_18249);
nor U20933 (N_20933,N_18552,N_19181);
or U20934 (N_20934,N_17533,N_19870);
or U20935 (N_20935,N_19219,N_19084);
or U20936 (N_20936,N_18677,N_18158);
nand U20937 (N_20937,N_19448,N_19352);
nor U20938 (N_20938,N_17864,N_18687);
nor U20939 (N_20939,N_19414,N_18537);
nand U20940 (N_20940,N_19435,N_17976);
xor U20941 (N_20941,N_18420,N_19304);
and U20942 (N_20942,N_17878,N_18037);
or U20943 (N_20943,N_19778,N_19533);
nand U20944 (N_20944,N_19354,N_19550);
or U20945 (N_20945,N_18504,N_19760);
and U20946 (N_20946,N_19703,N_19816);
and U20947 (N_20947,N_18895,N_19114);
nor U20948 (N_20948,N_19168,N_19706);
xnor U20949 (N_20949,N_19013,N_17707);
nand U20950 (N_20950,N_19480,N_17671);
xor U20951 (N_20951,N_19850,N_18548);
and U20952 (N_20952,N_19999,N_18452);
nand U20953 (N_20953,N_17831,N_18061);
or U20954 (N_20954,N_19501,N_18827);
xor U20955 (N_20955,N_19913,N_18539);
or U20956 (N_20956,N_18610,N_18726);
xnor U20957 (N_20957,N_18617,N_19062);
or U20958 (N_20958,N_19150,N_18446);
nand U20959 (N_20959,N_19407,N_19080);
nor U20960 (N_20960,N_18081,N_19748);
or U20961 (N_20961,N_17843,N_17799);
xor U20962 (N_20962,N_18341,N_18371);
and U20963 (N_20963,N_18366,N_18015);
or U20964 (N_20964,N_18508,N_19825);
xor U20965 (N_20965,N_18206,N_17726);
xor U20966 (N_20966,N_18074,N_18123);
xor U20967 (N_20967,N_17917,N_17621);
xnor U20968 (N_20968,N_19198,N_18309);
nand U20969 (N_20969,N_19871,N_17702);
and U20970 (N_20970,N_19356,N_18207);
or U20971 (N_20971,N_18007,N_18050);
nor U20972 (N_20972,N_19465,N_18941);
xnor U20973 (N_20973,N_17564,N_19517);
xnor U20974 (N_20974,N_19595,N_17764);
and U20975 (N_20975,N_19752,N_17871);
nor U20976 (N_20976,N_18240,N_17522);
nand U20977 (N_20977,N_17802,N_17504);
nor U20978 (N_20978,N_18887,N_17787);
or U20979 (N_20979,N_18287,N_19126);
and U20980 (N_20980,N_18308,N_18938);
xnor U20981 (N_20981,N_19467,N_18112);
and U20982 (N_20982,N_19811,N_19488);
or U20983 (N_20983,N_19986,N_19269);
nor U20984 (N_20984,N_17866,N_19169);
xnor U20985 (N_20985,N_18896,N_18804);
and U20986 (N_20986,N_18409,N_17750);
nor U20987 (N_20987,N_19432,N_18752);
nand U20988 (N_20988,N_18466,N_19638);
or U20989 (N_20989,N_17765,N_19875);
and U20990 (N_20990,N_18763,N_19814);
nor U20991 (N_20991,N_18660,N_17970);
nand U20992 (N_20992,N_18818,N_18838);
xnor U20993 (N_20993,N_19790,N_18933);
nor U20994 (N_20994,N_19558,N_18653);
xnor U20995 (N_20995,N_17801,N_17610);
or U20996 (N_20996,N_18011,N_17857);
and U20997 (N_20997,N_18954,N_18457);
nor U20998 (N_20998,N_17841,N_17792);
nand U20999 (N_20999,N_17798,N_19366);
xnor U21000 (N_21000,N_17856,N_19570);
and U21001 (N_21001,N_18040,N_17619);
or U21002 (N_21002,N_17529,N_19446);
nand U21003 (N_21003,N_17655,N_17672);
xor U21004 (N_21004,N_18192,N_18993);
nor U21005 (N_21005,N_18626,N_17924);
and U21006 (N_21006,N_17785,N_17703);
nand U21007 (N_21007,N_18671,N_18837);
and U21008 (N_21008,N_18087,N_19199);
xnor U21009 (N_21009,N_18079,N_18189);
nand U21010 (N_21010,N_18115,N_18697);
nor U21011 (N_21011,N_18641,N_18336);
or U21012 (N_21012,N_19442,N_18039);
and U21013 (N_21013,N_19934,N_19728);
nand U21014 (N_21014,N_17575,N_19308);
nor U21015 (N_21015,N_19641,N_19587);
or U21016 (N_21016,N_17515,N_19420);
nand U21017 (N_21017,N_18829,N_18442);
nor U21018 (N_21018,N_18736,N_19583);
or U21019 (N_21019,N_19702,N_18091);
or U21020 (N_21020,N_18487,N_19928);
xor U21021 (N_21021,N_18260,N_17835);
nor U21022 (N_21022,N_19313,N_19425);
and U21023 (N_21023,N_18703,N_18392);
and U21024 (N_21024,N_19135,N_19669);
or U21025 (N_21025,N_17989,N_18247);
nor U21026 (N_21026,N_19651,N_18996);
nor U21027 (N_21027,N_19554,N_17842);
nor U21028 (N_21028,N_17607,N_19991);
or U21029 (N_21029,N_17773,N_18459);
or U21030 (N_21030,N_18033,N_18809);
and U21031 (N_21031,N_19409,N_17903);
and U21032 (N_21032,N_17614,N_18065);
nand U21033 (N_21033,N_19479,N_19525);
nor U21034 (N_21034,N_19266,N_18266);
or U21035 (N_21035,N_18721,N_17826);
nand U21036 (N_21036,N_19401,N_17940);
nand U21037 (N_21037,N_19367,N_18688);
and U21038 (N_21038,N_19196,N_18070);
nand U21039 (N_21039,N_17624,N_18704);
xnor U21040 (N_21040,N_19744,N_17623);
nand U21041 (N_21041,N_18559,N_19691);
nand U21042 (N_21042,N_18801,N_17517);
nor U21043 (N_21043,N_17800,N_19212);
or U21044 (N_21044,N_18956,N_18080);
or U21045 (N_21045,N_18530,N_19318);
or U21046 (N_21046,N_17659,N_18710);
xor U21047 (N_21047,N_18628,N_17507);
or U21048 (N_21048,N_19170,N_18344);
nand U21049 (N_21049,N_18698,N_18295);
and U21050 (N_21050,N_19672,N_19363);
nor U21051 (N_21051,N_19453,N_19821);
nor U21052 (N_21052,N_19845,N_18806);
nand U21053 (N_21053,N_18144,N_18092);
nand U21054 (N_21054,N_19247,N_17712);
or U21055 (N_21055,N_17670,N_18036);
or U21056 (N_21056,N_18905,N_18089);
or U21057 (N_21057,N_19248,N_17571);
nand U21058 (N_21058,N_18413,N_19327);
xor U21059 (N_21059,N_18670,N_17793);
and U21060 (N_21060,N_18878,N_18685);
nand U21061 (N_21061,N_19415,N_17632);
nor U21062 (N_21062,N_17586,N_17803);
and U21063 (N_21063,N_18928,N_17829);
and U21064 (N_21064,N_18122,N_17808);
nor U21065 (N_21065,N_18394,N_18008);
nor U21066 (N_21066,N_19843,N_19894);
or U21067 (N_21067,N_17577,N_18960);
nor U21068 (N_21068,N_18912,N_19393);
nor U21069 (N_21069,N_17556,N_19477);
nor U21070 (N_21070,N_17811,N_18038);
nand U21071 (N_21071,N_19305,N_19794);
nand U21072 (N_21072,N_19291,N_17544);
nor U21073 (N_21073,N_17833,N_18127);
nor U21074 (N_21074,N_19094,N_18368);
nor U21075 (N_21075,N_19768,N_19141);
or U21076 (N_21076,N_19543,N_18903);
xnor U21077 (N_21077,N_19666,N_17627);
and U21078 (N_21078,N_18130,N_18495);
or U21079 (N_21079,N_18744,N_19998);
nand U21080 (N_21080,N_19260,N_19750);
and U21081 (N_21081,N_17894,N_19015);
xor U21082 (N_21082,N_18353,N_17851);
xor U21083 (N_21083,N_19581,N_19724);
xnor U21084 (N_21084,N_19795,N_19362);
nand U21085 (N_21085,N_19649,N_19882);
nor U21086 (N_21086,N_19891,N_19115);
nand U21087 (N_21087,N_18729,N_18356);
nand U21088 (N_21088,N_18986,N_19123);
or U21089 (N_21089,N_17598,N_18237);
or U21090 (N_21090,N_18902,N_19943);
nor U21091 (N_21091,N_17914,N_19028);
and U21092 (N_21092,N_18694,N_19653);
xnor U21093 (N_21093,N_19580,N_19063);
xor U21094 (N_21094,N_19234,N_18899);
or U21095 (N_21095,N_19213,N_18060);
or U21096 (N_21096,N_19082,N_18618);
xor U21097 (N_21097,N_18917,N_17977);
nand U21098 (N_21098,N_19590,N_19386);
and U21099 (N_21099,N_19857,N_19599);
and U21100 (N_21100,N_19650,N_18488);
xor U21101 (N_21101,N_17538,N_18982);
nand U21102 (N_21102,N_19628,N_19343);
or U21103 (N_21103,N_19710,N_18651);
or U21104 (N_21104,N_19155,N_19910);
nand U21105 (N_21105,N_19364,N_18793);
and U21106 (N_21106,N_18017,N_19059);
nor U21107 (N_21107,N_18693,N_18236);
xnor U21108 (N_21108,N_18151,N_18020);
xnor U21109 (N_21109,N_18193,N_18834);
nand U21110 (N_21110,N_19730,N_18310);
and U21111 (N_21111,N_18824,N_18145);
nand U21112 (N_21112,N_19827,N_17592);
or U21113 (N_21113,N_18904,N_19727);
and U21114 (N_21114,N_19052,N_18324);
nand U21115 (N_21115,N_19436,N_19251);
nand U21116 (N_21116,N_19206,N_17881);
and U21117 (N_21117,N_18869,N_18930);
and U21118 (N_21118,N_19970,N_18421);
xnor U21119 (N_21119,N_19108,N_19560);
and U21120 (N_21120,N_18433,N_19608);
and U21121 (N_21121,N_17901,N_19476);
xnor U21122 (N_21122,N_18854,N_18885);
nand U21123 (N_21123,N_19148,N_18727);
xnor U21124 (N_21124,N_18110,N_17766);
nand U21125 (N_21125,N_18569,N_18496);
and U21126 (N_21126,N_19802,N_18068);
xor U21127 (N_21127,N_18759,N_18054);
or U21128 (N_21128,N_19824,N_19594);
and U21129 (N_21129,N_18491,N_18841);
nand U21130 (N_21130,N_17821,N_18120);
nand U21131 (N_21131,N_18753,N_19132);
xor U21132 (N_21132,N_17886,N_18958);
and U21133 (N_21133,N_18808,N_19197);
or U21134 (N_21134,N_19919,N_19551);
or U21135 (N_21135,N_19726,N_17958);
and U21136 (N_21136,N_19880,N_19320);
nor U21137 (N_21137,N_18188,N_19655);
xnor U21138 (N_21138,N_19333,N_18819);
and U21139 (N_21139,N_18988,N_19520);
and U21140 (N_21140,N_18790,N_17805);
or U21141 (N_21141,N_19060,N_18517);
nor U21142 (N_21142,N_19019,N_19216);
nand U21143 (N_21143,N_17956,N_18814);
or U21144 (N_21144,N_19566,N_19783);
nor U21145 (N_21145,N_18313,N_19842);
xor U21146 (N_21146,N_18012,N_18486);
nand U21147 (N_21147,N_18456,N_18845);
nand U21148 (N_21148,N_19347,N_17928);
or U21149 (N_21149,N_19496,N_17649);
nand U21150 (N_21150,N_18138,N_19025);
nand U21151 (N_21151,N_18862,N_18149);
nor U21152 (N_21152,N_18519,N_19878);
nand U21153 (N_21153,N_18944,N_18484);
or U21154 (N_21154,N_19620,N_18505);
nand U21155 (N_21155,N_18750,N_18894);
and U21156 (N_21156,N_18820,N_19832);
and U21157 (N_21157,N_17565,N_18560);
and U21158 (N_21158,N_18384,N_18876);
and U21159 (N_21159,N_18500,N_19487);
and U21160 (N_21160,N_18104,N_18156);
and U21161 (N_21161,N_18780,N_19733);
xnor U21162 (N_21162,N_18923,N_18424);
xnor U21163 (N_21163,N_18216,N_18214);
xor U21164 (N_21164,N_18623,N_19676);
and U21165 (N_21165,N_18229,N_18330);
xor U21166 (N_21166,N_18118,N_19684);
and U21167 (N_21167,N_18434,N_18403);
nand U21168 (N_21168,N_18901,N_17868);
or U21169 (N_21169,N_17705,N_18817);
and U21170 (N_21170,N_17570,N_19242);
nand U21171 (N_21171,N_18256,N_18831);
nand U21172 (N_21172,N_17745,N_18220);
xor U21173 (N_21173,N_18611,N_18263);
nand U21174 (N_21174,N_19549,N_18057);
nor U21175 (N_21175,N_19959,N_17789);
nand U21176 (N_21176,N_19785,N_18918);
and U21177 (N_21177,N_19535,N_18400);
and U21178 (N_21178,N_18099,N_19252);
nor U21179 (N_21179,N_19228,N_19011);
or U21180 (N_21180,N_19353,N_18439);
xnor U21181 (N_21181,N_17895,N_19246);
and U21182 (N_21182,N_17673,N_18547);
nand U21183 (N_21183,N_18718,N_17699);
and U21184 (N_21184,N_18034,N_19745);
or U21185 (N_21185,N_19221,N_17563);
xnor U21186 (N_21186,N_19173,N_18581);
nand U21187 (N_21187,N_17657,N_17896);
nor U21188 (N_21188,N_19639,N_17863);
and U21189 (N_21189,N_18799,N_19002);
xor U21190 (N_21190,N_19041,N_17502);
nand U21191 (N_21191,N_19284,N_19163);
nand U21192 (N_21192,N_18398,N_19074);
nand U21193 (N_21193,N_18315,N_18910);
xor U21194 (N_21194,N_19264,N_17609);
nor U21195 (N_21195,N_17838,N_17912);
xnor U21196 (N_21196,N_19524,N_19097);
or U21197 (N_21197,N_17722,N_19151);
and U21198 (N_21198,N_18059,N_18044);
nand U21199 (N_21199,N_18786,N_18339);
or U21200 (N_21200,N_19297,N_18224);
xnor U21201 (N_21201,N_18578,N_19874);
or U21202 (N_21202,N_17660,N_17937);
xnor U21203 (N_21203,N_17830,N_18655);
nand U21204 (N_21204,N_18284,N_19280);
and U21205 (N_21205,N_17813,N_18259);
xnor U21206 (N_21206,N_18561,N_19450);
nor U21207 (N_21207,N_19722,N_19316);
or U21208 (N_21208,N_18644,N_19747);
and U21209 (N_21209,N_18010,N_19493);
and U21210 (N_21210,N_18447,N_18473);
xor U21211 (N_21211,N_17770,N_18797);
xnor U21212 (N_21212,N_19654,N_19955);
xor U21213 (N_21213,N_19092,N_19245);
xor U21214 (N_21214,N_19926,N_18570);
nor U21215 (N_21215,N_18440,N_19972);
nand U21216 (N_21216,N_18872,N_18142);
and U21217 (N_21217,N_18106,N_18922);
nand U21218 (N_21218,N_19240,N_18289);
and U21219 (N_21219,N_18742,N_17761);
nor U21220 (N_21220,N_18210,N_18132);
nand U21221 (N_21221,N_17748,N_18478);
xor U21222 (N_21222,N_19142,N_19699);
nor U21223 (N_21223,N_18451,N_18969);
nand U21224 (N_21224,N_18133,N_18018);
xnor U21225 (N_21225,N_18143,N_18594);
or U21226 (N_21226,N_18109,N_19687);
or U21227 (N_21227,N_19859,N_18016);
nand U21228 (N_21228,N_19113,N_18377);
nor U21229 (N_21229,N_19276,N_19709);
nand U21230 (N_21230,N_18072,N_18195);
xor U21231 (N_21231,N_18978,N_18182);
or U21232 (N_21232,N_18661,N_18230);
or U21233 (N_21233,N_17553,N_18399);
or U21234 (N_21234,N_19372,N_18657);
or U21235 (N_21235,N_19588,N_19391);
xor U21236 (N_21236,N_18441,N_18571);
nor U21237 (N_21237,N_19102,N_19189);
nand U21238 (N_21238,N_18135,N_17769);
or U21239 (N_21239,N_19923,N_19285);
xnor U21240 (N_21240,N_18625,N_18713);
or U21241 (N_21241,N_17899,N_17963);
nand U21242 (N_21242,N_19682,N_18332);
nor U21243 (N_21243,N_18244,N_19326);
and U21244 (N_21244,N_19003,N_19402);
and U21245 (N_21245,N_18241,N_19960);
nand U21246 (N_21246,N_18170,N_19068);
and U21247 (N_21247,N_19325,N_18748);
or U21248 (N_21248,N_19046,N_19577);
xor U21249 (N_21249,N_17931,N_19231);
nor U21250 (N_21250,N_18604,N_19987);
or U21251 (N_21251,N_17852,N_18710);
xor U21252 (N_21252,N_18006,N_18567);
xnor U21253 (N_21253,N_19580,N_19102);
xnor U21254 (N_21254,N_18021,N_18334);
nor U21255 (N_21255,N_19050,N_18033);
nand U21256 (N_21256,N_17587,N_18909);
nor U21257 (N_21257,N_19417,N_18003);
nor U21258 (N_21258,N_18837,N_19726);
nor U21259 (N_21259,N_18201,N_19187);
and U21260 (N_21260,N_17776,N_18116);
and U21261 (N_21261,N_19916,N_19948);
nand U21262 (N_21262,N_18109,N_19510);
xnor U21263 (N_21263,N_17503,N_18588);
or U21264 (N_21264,N_19930,N_18208);
xnor U21265 (N_21265,N_18095,N_19995);
or U21266 (N_21266,N_19350,N_18730);
xor U21267 (N_21267,N_19512,N_19916);
or U21268 (N_21268,N_19320,N_17756);
and U21269 (N_21269,N_18886,N_18762);
nand U21270 (N_21270,N_18088,N_19519);
xor U21271 (N_21271,N_19979,N_18994);
nand U21272 (N_21272,N_18491,N_17886);
xnor U21273 (N_21273,N_17596,N_19448);
or U21274 (N_21274,N_19551,N_19669);
or U21275 (N_21275,N_19652,N_18502);
nand U21276 (N_21276,N_18682,N_17517);
xor U21277 (N_21277,N_17814,N_19273);
or U21278 (N_21278,N_17575,N_18028);
xor U21279 (N_21279,N_18465,N_18860);
and U21280 (N_21280,N_18956,N_17502);
xor U21281 (N_21281,N_18787,N_19399);
nand U21282 (N_21282,N_19232,N_17698);
or U21283 (N_21283,N_18292,N_18039);
xnor U21284 (N_21284,N_18354,N_18596);
or U21285 (N_21285,N_17663,N_18392);
or U21286 (N_21286,N_19991,N_18441);
and U21287 (N_21287,N_18020,N_18759);
or U21288 (N_21288,N_17638,N_18199);
nand U21289 (N_21289,N_17777,N_19684);
xor U21290 (N_21290,N_19226,N_19584);
and U21291 (N_21291,N_18081,N_18012);
or U21292 (N_21292,N_19598,N_19403);
nand U21293 (N_21293,N_19646,N_19315);
nor U21294 (N_21294,N_18711,N_17713);
and U21295 (N_21295,N_18661,N_17819);
or U21296 (N_21296,N_18004,N_18092);
xor U21297 (N_21297,N_18369,N_18124);
nor U21298 (N_21298,N_17951,N_18591);
or U21299 (N_21299,N_18318,N_18749);
and U21300 (N_21300,N_19586,N_19745);
or U21301 (N_21301,N_19896,N_19948);
xnor U21302 (N_21302,N_19246,N_18613);
or U21303 (N_21303,N_17855,N_18671);
or U21304 (N_21304,N_18938,N_18265);
nor U21305 (N_21305,N_18419,N_19518);
and U21306 (N_21306,N_18317,N_18265);
or U21307 (N_21307,N_18705,N_18499);
or U21308 (N_21308,N_18964,N_19225);
nand U21309 (N_21309,N_17669,N_19068);
xnor U21310 (N_21310,N_19662,N_18940);
and U21311 (N_21311,N_17749,N_18598);
and U21312 (N_21312,N_18394,N_19058);
nor U21313 (N_21313,N_18570,N_19084);
xor U21314 (N_21314,N_17895,N_18815);
xnor U21315 (N_21315,N_19256,N_18053);
nand U21316 (N_21316,N_18310,N_19031);
nand U21317 (N_21317,N_18015,N_17851);
and U21318 (N_21318,N_19864,N_18839);
xor U21319 (N_21319,N_18574,N_18483);
nor U21320 (N_21320,N_19805,N_19699);
nand U21321 (N_21321,N_17757,N_19087);
and U21322 (N_21322,N_19804,N_18662);
nand U21323 (N_21323,N_17557,N_19332);
and U21324 (N_21324,N_19217,N_18369);
xor U21325 (N_21325,N_19870,N_18700);
nor U21326 (N_21326,N_17535,N_18467);
or U21327 (N_21327,N_18453,N_18515);
xor U21328 (N_21328,N_17534,N_17872);
nand U21329 (N_21329,N_17905,N_18568);
and U21330 (N_21330,N_19015,N_18475);
nand U21331 (N_21331,N_18725,N_17832);
and U21332 (N_21332,N_17831,N_18401);
or U21333 (N_21333,N_19756,N_19198);
and U21334 (N_21334,N_18800,N_17754);
and U21335 (N_21335,N_19944,N_17880);
or U21336 (N_21336,N_19553,N_19590);
nand U21337 (N_21337,N_19520,N_18195);
nor U21338 (N_21338,N_18852,N_17554);
or U21339 (N_21339,N_17990,N_19140);
nor U21340 (N_21340,N_18858,N_18102);
or U21341 (N_21341,N_18788,N_18795);
nor U21342 (N_21342,N_18413,N_19179);
nand U21343 (N_21343,N_19434,N_18958);
nor U21344 (N_21344,N_17645,N_17779);
and U21345 (N_21345,N_18587,N_17727);
or U21346 (N_21346,N_18605,N_17665);
and U21347 (N_21347,N_18028,N_17930);
or U21348 (N_21348,N_18429,N_18884);
and U21349 (N_21349,N_18823,N_19307);
nor U21350 (N_21350,N_19017,N_17703);
and U21351 (N_21351,N_19500,N_19635);
xnor U21352 (N_21352,N_19426,N_17705);
nor U21353 (N_21353,N_19145,N_19974);
or U21354 (N_21354,N_19206,N_17635);
xnor U21355 (N_21355,N_18779,N_18383);
or U21356 (N_21356,N_19257,N_18185);
nor U21357 (N_21357,N_17623,N_18608);
xnor U21358 (N_21358,N_17507,N_18696);
or U21359 (N_21359,N_17626,N_18219);
or U21360 (N_21360,N_17969,N_18736);
nor U21361 (N_21361,N_18325,N_18302);
nor U21362 (N_21362,N_18611,N_19532);
or U21363 (N_21363,N_18750,N_18224);
or U21364 (N_21364,N_17806,N_18297);
nand U21365 (N_21365,N_18411,N_19831);
nand U21366 (N_21366,N_17680,N_18141);
nand U21367 (N_21367,N_17540,N_19753);
nand U21368 (N_21368,N_18065,N_19346);
and U21369 (N_21369,N_19764,N_19816);
and U21370 (N_21370,N_17584,N_18831);
and U21371 (N_21371,N_19129,N_19531);
and U21372 (N_21372,N_18549,N_18158);
and U21373 (N_21373,N_19983,N_18979);
xnor U21374 (N_21374,N_19406,N_17929);
and U21375 (N_21375,N_17628,N_18354);
xnor U21376 (N_21376,N_18621,N_18613);
nor U21377 (N_21377,N_19148,N_18330);
xor U21378 (N_21378,N_18128,N_19522);
nor U21379 (N_21379,N_19546,N_17932);
xnor U21380 (N_21380,N_17939,N_18453);
xnor U21381 (N_21381,N_19456,N_17582);
nand U21382 (N_21382,N_17821,N_17913);
nand U21383 (N_21383,N_19609,N_17657);
nand U21384 (N_21384,N_18233,N_18916);
nand U21385 (N_21385,N_19923,N_18341);
or U21386 (N_21386,N_17911,N_19512);
nor U21387 (N_21387,N_19287,N_18200);
and U21388 (N_21388,N_19387,N_19583);
nor U21389 (N_21389,N_18269,N_18898);
nor U21390 (N_21390,N_19619,N_17847);
and U21391 (N_21391,N_19889,N_18750);
xor U21392 (N_21392,N_19776,N_18061);
nor U21393 (N_21393,N_17923,N_18222);
and U21394 (N_21394,N_17544,N_19400);
or U21395 (N_21395,N_17524,N_18276);
nor U21396 (N_21396,N_19419,N_19090);
xnor U21397 (N_21397,N_18948,N_19453);
xnor U21398 (N_21398,N_17885,N_18483);
xor U21399 (N_21399,N_17796,N_19728);
xor U21400 (N_21400,N_18890,N_17631);
or U21401 (N_21401,N_17664,N_18523);
and U21402 (N_21402,N_17929,N_19033);
and U21403 (N_21403,N_19279,N_18129);
xnor U21404 (N_21404,N_19887,N_18544);
nor U21405 (N_21405,N_17953,N_18732);
nand U21406 (N_21406,N_18469,N_18553);
xor U21407 (N_21407,N_18399,N_19902);
or U21408 (N_21408,N_18380,N_19055);
nor U21409 (N_21409,N_18131,N_19753);
and U21410 (N_21410,N_17919,N_17850);
nor U21411 (N_21411,N_18271,N_19175);
or U21412 (N_21412,N_17837,N_19772);
or U21413 (N_21413,N_19203,N_17733);
xor U21414 (N_21414,N_18128,N_19391);
nor U21415 (N_21415,N_18070,N_18627);
nor U21416 (N_21416,N_17562,N_18462);
xnor U21417 (N_21417,N_18313,N_18758);
nand U21418 (N_21418,N_18393,N_18606);
and U21419 (N_21419,N_19687,N_18538);
and U21420 (N_21420,N_17905,N_19964);
or U21421 (N_21421,N_18152,N_17544);
nor U21422 (N_21422,N_19302,N_18397);
xor U21423 (N_21423,N_18957,N_18052);
and U21424 (N_21424,N_19951,N_19106);
and U21425 (N_21425,N_19776,N_17820);
xnor U21426 (N_21426,N_18785,N_17593);
or U21427 (N_21427,N_17999,N_19939);
or U21428 (N_21428,N_18064,N_19616);
nor U21429 (N_21429,N_18533,N_19929);
xor U21430 (N_21430,N_19391,N_19279);
xor U21431 (N_21431,N_18692,N_19740);
nor U21432 (N_21432,N_17535,N_17952);
and U21433 (N_21433,N_17700,N_17716);
and U21434 (N_21434,N_17942,N_18614);
or U21435 (N_21435,N_19302,N_18128);
xor U21436 (N_21436,N_18261,N_17897);
xor U21437 (N_21437,N_19365,N_18814);
nand U21438 (N_21438,N_18308,N_19596);
xnor U21439 (N_21439,N_18821,N_17853);
nand U21440 (N_21440,N_18496,N_17977);
and U21441 (N_21441,N_19083,N_19080);
or U21442 (N_21442,N_18016,N_17552);
and U21443 (N_21443,N_19823,N_18094);
and U21444 (N_21444,N_18404,N_19573);
nand U21445 (N_21445,N_18245,N_18122);
or U21446 (N_21446,N_18153,N_19300);
nand U21447 (N_21447,N_18910,N_17663);
xnor U21448 (N_21448,N_17686,N_19258);
nand U21449 (N_21449,N_18713,N_18685);
and U21450 (N_21450,N_19599,N_17638);
nor U21451 (N_21451,N_17527,N_18519);
nand U21452 (N_21452,N_17846,N_19836);
nor U21453 (N_21453,N_18843,N_18705);
and U21454 (N_21454,N_18859,N_18284);
nand U21455 (N_21455,N_19252,N_18162);
and U21456 (N_21456,N_18561,N_19197);
nand U21457 (N_21457,N_19921,N_19136);
nand U21458 (N_21458,N_18123,N_18472);
nand U21459 (N_21459,N_19821,N_17679);
nand U21460 (N_21460,N_18715,N_18905);
or U21461 (N_21461,N_18616,N_18730);
nor U21462 (N_21462,N_19062,N_17929);
nor U21463 (N_21463,N_18796,N_18251);
xor U21464 (N_21464,N_19805,N_17999);
or U21465 (N_21465,N_18984,N_17593);
nand U21466 (N_21466,N_18523,N_19628);
and U21467 (N_21467,N_18774,N_19115);
or U21468 (N_21468,N_19317,N_19778);
nand U21469 (N_21469,N_19607,N_19992);
nand U21470 (N_21470,N_19003,N_17950);
nor U21471 (N_21471,N_19695,N_18684);
nand U21472 (N_21472,N_18556,N_19587);
nand U21473 (N_21473,N_18916,N_17609);
nor U21474 (N_21474,N_19884,N_19471);
and U21475 (N_21475,N_17932,N_18930);
nand U21476 (N_21476,N_19907,N_18914);
nand U21477 (N_21477,N_18885,N_19279);
nand U21478 (N_21478,N_17612,N_18836);
nor U21479 (N_21479,N_19069,N_18215);
or U21480 (N_21480,N_19014,N_19216);
and U21481 (N_21481,N_17659,N_18048);
xor U21482 (N_21482,N_18070,N_19819);
and U21483 (N_21483,N_19919,N_17636);
and U21484 (N_21484,N_19242,N_18514);
nor U21485 (N_21485,N_17707,N_18264);
nand U21486 (N_21486,N_19925,N_17508);
xnor U21487 (N_21487,N_17591,N_18910);
and U21488 (N_21488,N_19925,N_18628);
nor U21489 (N_21489,N_18010,N_18107);
nand U21490 (N_21490,N_17877,N_19755);
xor U21491 (N_21491,N_19336,N_18493);
nand U21492 (N_21492,N_19381,N_17772);
nor U21493 (N_21493,N_19491,N_19083);
nand U21494 (N_21494,N_19744,N_19370);
nor U21495 (N_21495,N_18325,N_17903);
and U21496 (N_21496,N_18789,N_19173);
nand U21497 (N_21497,N_17739,N_17610);
or U21498 (N_21498,N_18885,N_19753);
nor U21499 (N_21499,N_19123,N_18283);
nor U21500 (N_21500,N_17711,N_18707);
nor U21501 (N_21501,N_19066,N_19909);
nor U21502 (N_21502,N_18212,N_18181);
or U21503 (N_21503,N_19911,N_19145);
or U21504 (N_21504,N_19740,N_18026);
or U21505 (N_21505,N_17761,N_19161);
nor U21506 (N_21506,N_17576,N_18705);
nor U21507 (N_21507,N_19726,N_19091);
or U21508 (N_21508,N_19973,N_17500);
xnor U21509 (N_21509,N_19797,N_19414);
and U21510 (N_21510,N_18934,N_19624);
and U21511 (N_21511,N_19723,N_17935);
or U21512 (N_21512,N_18128,N_19451);
and U21513 (N_21513,N_18460,N_18486);
and U21514 (N_21514,N_19392,N_18330);
xor U21515 (N_21515,N_18739,N_19394);
and U21516 (N_21516,N_18170,N_17781);
nor U21517 (N_21517,N_17976,N_18220);
or U21518 (N_21518,N_19273,N_19098);
nand U21519 (N_21519,N_17796,N_19359);
and U21520 (N_21520,N_18589,N_19942);
or U21521 (N_21521,N_18396,N_18183);
and U21522 (N_21522,N_17903,N_19148);
and U21523 (N_21523,N_18651,N_19426);
or U21524 (N_21524,N_18224,N_18831);
xnor U21525 (N_21525,N_19424,N_19498);
nand U21526 (N_21526,N_19689,N_18761);
or U21527 (N_21527,N_18311,N_19214);
and U21528 (N_21528,N_17889,N_19550);
xor U21529 (N_21529,N_19045,N_19477);
or U21530 (N_21530,N_19527,N_18370);
nor U21531 (N_21531,N_19636,N_19566);
nand U21532 (N_21532,N_17551,N_18455);
nand U21533 (N_21533,N_17720,N_19359);
nand U21534 (N_21534,N_19730,N_19407);
and U21535 (N_21535,N_19474,N_17569);
nor U21536 (N_21536,N_17788,N_19597);
and U21537 (N_21537,N_19649,N_19825);
nor U21538 (N_21538,N_19124,N_18017);
nor U21539 (N_21539,N_18258,N_17795);
nand U21540 (N_21540,N_19867,N_18409);
nor U21541 (N_21541,N_18963,N_19810);
and U21542 (N_21542,N_18857,N_19728);
or U21543 (N_21543,N_18460,N_19488);
nand U21544 (N_21544,N_19150,N_17982);
nand U21545 (N_21545,N_17903,N_19454);
nor U21546 (N_21546,N_19818,N_18427);
or U21547 (N_21547,N_19309,N_18600);
nor U21548 (N_21548,N_19583,N_17702);
and U21549 (N_21549,N_18460,N_18160);
or U21550 (N_21550,N_17785,N_18420);
and U21551 (N_21551,N_17984,N_18180);
nor U21552 (N_21552,N_19530,N_19270);
or U21553 (N_21553,N_18378,N_18271);
nand U21554 (N_21554,N_18638,N_19752);
nand U21555 (N_21555,N_18660,N_18717);
and U21556 (N_21556,N_18484,N_18340);
nand U21557 (N_21557,N_18625,N_18917);
nand U21558 (N_21558,N_18946,N_18828);
nand U21559 (N_21559,N_18504,N_18736);
nand U21560 (N_21560,N_18639,N_19200);
nand U21561 (N_21561,N_18438,N_19637);
nor U21562 (N_21562,N_19895,N_19446);
xor U21563 (N_21563,N_18618,N_17530);
nor U21564 (N_21564,N_17520,N_18408);
nand U21565 (N_21565,N_18090,N_18123);
and U21566 (N_21566,N_18542,N_19732);
or U21567 (N_21567,N_17588,N_19733);
nand U21568 (N_21568,N_18657,N_19960);
and U21569 (N_21569,N_19785,N_17823);
or U21570 (N_21570,N_17589,N_17629);
xnor U21571 (N_21571,N_17881,N_19635);
or U21572 (N_21572,N_19377,N_18524);
xor U21573 (N_21573,N_18607,N_17631);
nor U21574 (N_21574,N_19551,N_18672);
xnor U21575 (N_21575,N_18310,N_18479);
nand U21576 (N_21576,N_19620,N_17900);
nand U21577 (N_21577,N_18490,N_19398);
nand U21578 (N_21578,N_19174,N_18697);
and U21579 (N_21579,N_19552,N_17943);
or U21580 (N_21580,N_18914,N_17663);
xnor U21581 (N_21581,N_17671,N_18722);
or U21582 (N_21582,N_19018,N_19610);
and U21583 (N_21583,N_18352,N_19663);
xor U21584 (N_21584,N_19085,N_17748);
or U21585 (N_21585,N_18475,N_19618);
xnor U21586 (N_21586,N_17521,N_18358);
xor U21587 (N_21587,N_19111,N_19810);
or U21588 (N_21588,N_18235,N_17737);
and U21589 (N_21589,N_19891,N_17910);
or U21590 (N_21590,N_18373,N_19340);
nand U21591 (N_21591,N_18115,N_18719);
and U21592 (N_21592,N_19499,N_18501);
xnor U21593 (N_21593,N_19006,N_17950);
xor U21594 (N_21594,N_19150,N_17588);
nand U21595 (N_21595,N_18287,N_18846);
and U21596 (N_21596,N_17834,N_17556);
nand U21597 (N_21597,N_18623,N_18245);
or U21598 (N_21598,N_19035,N_18065);
xor U21599 (N_21599,N_19065,N_17749);
and U21600 (N_21600,N_19876,N_18959);
nand U21601 (N_21601,N_19396,N_19958);
nor U21602 (N_21602,N_18773,N_18198);
xnor U21603 (N_21603,N_19512,N_17537);
xor U21604 (N_21604,N_18510,N_19194);
and U21605 (N_21605,N_17999,N_17535);
or U21606 (N_21606,N_18021,N_18509);
nand U21607 (N_21607,N_19311,N_19641);
or U21608 (N_21608,N_19889,N_18946);
or U21609 (N_21609,N_18985,N_19131);
nand U21610 (N_21610,N_19019,N_17594);
nor U21611 (N_21611,N_17541,N_17932);
nand U21612 (N_21612,N_18649,N_18884);
nor U21613 (N_21613,N_18421,N_18391);
nor U21614 (N_21614,N_18019,N_18539);
or U21615 (N_21615,N_19384,N_17595);
xnor U21616 (N_21616,N_19152,N_18934);
nand U21617 (N_21617,N_18558,N_18351);
and U21618 (N_21618,N_19801,N_18812);
nand U21619 (N_21619,N_19728,N_18705);
or U21620 (N_21620,N_17891,N_19858);
or U21621 (N_21621,N_17518,N_17781);
nor U21622 (N_21622,N_18179,N_18804);
or U21623 (N_21623,N_18274,N_19927);
nand U21624 (N_21624,N_18762,N_18055);
and U21625 (N_21625,N_19839,N_19185);
xor U21626 (N_21626,N_18711,N_18251);
nand U21627 (N_21627,N_18512,N_19956);
and U21628 (N_21628,N_18265,N_18134);
or U21629 (N_21629,N_19106,N_19930);
nor U21630 (N_21630,N_17668,N_19913);
and U21631 (N_21631,N_19602,N_18151);
xor U21632 (N_21632,N_19844,N_18797);
or U21633 (N_21633,N_18426,N_17580);
or U21634 (N_21634,N_18716,N_18520);
and U21635 (N_21635,N_18025,N_19939);
nand U21636 (N_21636,N_19484,N_19397);
nor U21637 (N_21637,N_18074,N_19459);
xnor U21638 (N_21638,N_19329,N_18293);
and U21639 (N_21639,N_18153,N_19026);
nand U21640 (N_21640,N_19846,N_19081);
nor U21641 (N_21641,N_17573,N_18146);
or U21642 (N_21642,N_17842,N_19664);
nor U21643 (N_21643,N_19342,N_18589);
xor U21644 (N_21644,N_19252,N_17854);
nand U21645 (N_21645,N_19898,N_17564);
nand U21646 (N_21646,N_17820,N_19632);
nor U21647 (N_21647,N_19137,N_19522);
nor U21648 (N_21648,N_18283,N_18168);
and U21649 (N_21649,N_19188,N_19645);
or U21650 (N_21650,N_18145,N_18091);
nand U21651 (N_21651,N_19003,N_17990);
or U21652 (N_21652,N_18845,N_19912);
xnor U21653 (N_21653,N_19786,N_19233);
nand U21654 (N_21654,N_19037,N_18855);
xnor U21655 (N_21655,N_19809,N_19371);
nand U21656 (N_21656,N_18881,N_18494);
xnor U21657 (N_21657,N_18646,N_19041);
and U21658 (N_21658,N_18784,N_18189);
xnor U21659 (N_21659,N_19570,N_19935);
nor U21660 (N_21660,N_19227,N_18513);
xnor U21661 (N_21661,N_18914,N_18785);
or U21662 (N_21662,N_19393,N_18775);
xor U21663 (N_21663,N_19224,N_19364);
or U21664 (N_21664,N_19055,N_18156);
xor U21665 (N_21665,N_18835,N_19437);
xnor U21666 (N_21666,N_19159,N_19305);
nor U21667 (N_21667,N_17615,N_17836);
xnor U21668 (N_21668,N_17939,N_17513);
nand U21669 (N_21669,N_19898,N_19347);
or U21670 (N_21670,N_18703,N_18701);
nand U21671 (N_21671,N_19184,N_18630);
and U21672 (N_21672,N_17874,N_18310);
nor U21673 (N_21673,N_18500,N_17626);
xnor U21674 (N_21674,N_18901,N_19626);
or U21675 (N_21675,N_19150,N_18956);
or U21676 (N_21676,N_19038,N_18045);
and U21677 (N_21677,N_17570,N_17752);
nand U21678 (N_21678,N_19381,N_19127);
nand U21679 (N_21679,N_19286,N_17794);
or U21680 (N_21680,N_19999,N_18806);
and U21681 (N_21681,N_19630,N_19564);
or U21682 (N_21682,N_18208,N_19131);
nand U21683 (N_21683,N_18706,N_19874);
and U21684 (N_21684,N_19904,N_17503);
xor U21685 (N_21685,N_18417,N_19284);
or U21686 (N_21686,N_18799,N_18583);
xor U21687 (N_21687,N_17515,N_19642);
nor U21688 (N_21688,N_18120,N_18370);
nand U21689 (N_21689,N_18010,N_18844);
xnor U21690 (N_21690,N_19946,N_18502);
nand U21691 (N_21691,N_17515,N_19195);
and U21692 (N_21692,N_18136,N_19002);
xnor U21693 (N_21693,N_17781,N_18379);
or U21694 (N_21694,N_19668,N_17748);
nand U21695 (N_21695,N_19893,N_17694);
and U21696 (N_21696,N_19668,N_18744);
or U21697 (N_21697,N_18959,N_18153);
and U21698 (N_21698,N_19125,N_19540);
or U21699 (N_21699,N_17993,N_18763);
nand U21700 (N_21700,N_17697,N_18789);
and U21701 (N_21701,N_19203,N_18025);
xnor U21702 (N_21702,N_18998,N_18739);
nor U21703 (N_21703,N_19220,N_18875);
xor U21704 (N_21704,N_19441,N_19848);
and U21705 (N_21705,N_19136,N_18370);
nand U21706 (N_21706,N_17989,N_17580);
nor U21707 (N_21707,N_17896,N_18811);
xnor U21708 (N_21708,N_17729,N_18439);
nor U21709 (N_21709,N_19704,N_18179);
nand U21710 (N_21710,N_19142,N_17820);
or U21711 (N_21711,N_19497,N_19489);
and U21712 (N_21712,N_17926,N_19668);
xor U21713 (N_21713,N_18199,N_18459);
or U21714 (N_21714,N_19539,N_18442);
nand U21715 (N_21715,N_18559,N_18860);
nand U21716 (N_21716,N_19084,N_18074);
nand U21717 (N_21717,N_18615,N_18540);
or U21718 (N_21718,N_19619,N_19816);
and U21719 (N_21719,N_18748,N_18194);
and U21720 (N_21720,N_17690,N_18789);
and U21721 (N_21721,N_18582,N_17905);
or U21722 (N_21722,N_18095,N_19703);
or U21723 (N_21723,N_18955,N_18746);
nand U21724 (N_21724,N_19247,N_17754);
and U21725 (N_21725,N_18075,N_18111);
nand U21726 (N_21726,N_19316,N_19502);
or U21727 (N_21727,N_18830,N_18440);
nand U21728 (N_21728,N_18670,N_19173);
or U21729 (N_21729,N_17826,N_18916);
or U21730 (N_21730,N_18566,N_19385);
xnor U21731 (N_21731,N_17950,N_19103);
and U21732 (N_21732,N_19127,N_19112);
or U21733 (N_21733,N_18380,N_17505);
nand U21734 (N_21734,N_18761,N_19390);
and U21735 (N_21735,N_19212,N_17810);
or U21736 (N_21736,N_17830,N_19607);
nand U21737 (N_21737,N_18631,N_19090);
nor U21738 (N_21738,N_18890,N_19131);
nand U21739 (N_21739,N_17544,N_19802);
nand U21740 (N_21740,N_19979,N_17704);
xnor U21741 (N_21741,N_18358,N_19731);
xnor U21742 (N_21742,N_17881,N_18160);
and U21743 (N_21743,N_19707,N_17982);
nor U21744 (N_21744,N_18334,N_19665);
and U21745 (N_21745,N_19230,N_18529);
or U21746 (N_21746,N_17898,N_18526);
nor U21747 (N_21747,N_18196,N_18820);
xnor U21748 (N_21748,N_18296,N_17641);
nand U21749 (N_21749,N_17685,N_18897);
or U21750 (N_21750,N_18209,N_17556);
or U21751 (N_21751,N_18100,N_19626);
nand U21752 (N_21752,N_17806,N_17805);
or U21753 (N_21753,N_17810,N_18232);
nor U21754 (N_21754,N_19564,N_17693);
and U21755 (N_21755,N_19310,N_19894);
xor U21756 (N_21756,N_18931,N_17903);
and U21757 (N_21757,N_19796,N_18619);
or U21758 (N_21758,N_19731,N_19625);
nor U21759 (N_21759,N_18657,N_18891);
nand U21760 (N_21760,N_19272,N_18429);
and U21761 (N_21761,N_18288,N_18478);
and U21762 (N_21762,N_19794,N_18725);
or U21763 (N_21763,N_18238,N_18206);
nor U21764 (N_21764,N_19734,N_19016);
xor U21765 (N_21765,N_18543,N_18563);
and U21766 (N_21766,N_19478,N_18795);
nand U21767 (N_21767,N_19139,N_17759);
nand U21768 (N_21768,N_19533,N_19172);
and U21769 (N_21769,N_18201,N_17546);
or U21770 (N_21770,N_19021,N_18918);
nand U21771 (N_21771,N_18592,N_19365);
xnor U21772 (N_21772,N_19399,N_18347);
and U21773 (N_21773,N_19486,N_19243);
or U21774 (N_21774,N_18480,N_19830);
nor U21775 (N_21775,N_18734,N_19114);
or U21776 (N_21776,N_19486,N_19772);
or U21777 (N_21777,N_17904,N_19406);
and U21778 (N_21778,N_18579,N_19857);
nand U21779 (N_21779,N_19850,N_18641);
xnor U21780 (N_21780,N_19654,N_19203);
xnor U21781 (N_21781,N_19452,N_18629);
and U21782 (N_21782,N_17643,N_17571);
xnor U21783 (N_21783,N_18293,N_17825);
or U21784 (N_21784,N_19585,N_18757);
and U21785 (N_21785,N_19381,N_17577);
nand U21786 (N_21786,N_19648,N_19984);
xnor U21787 (N_21787,N_17748,N_18084);
nor U21788 (N_21788,N_18390,N_19032);
nand U21789 (N_21789,N_18984,N_18256);
and U21790 (N_21790,N_18497,N_17753);
xnor U21791 (N_21791,N_19674,N_18732);
and U21792 (N_21792,N_17778,N_19813);
nand U21793 (N_21793,N_19982,N_18232);
xnor U21794 (N_21794,N_19582,N_17703);
nand U21795 (N_21795,N_18865,N_18066);
xor U21796 (N_21796,N_18914,N_18263);
or U21797 (N_21797,N_17701,N_19444);
nand U21798 (N_21798,N_19690,N_17661);
nor U21799 (N_21799,N_18664,N_19946);
nor U21800 (N_21800,N_18732,N_19628);
nor U21801 (N_21801,N_18380,N_19234);
nand U21802 (N_21802,N_17533,N_18589);
or U21803 (N_21803,N_19421,N_18856);
nor U21804 (N_21804,N_18470,N_17509);
nor U21805 (N_21805,N_19702,N_19630);
nor U21806 (N_21806,N_19929,N_19657);
or U21807 (N_21807,N_18270,N_19615);
or U21808 (N_21808,N_18251,N_19204);
or U21809 (N_21809,N_19366,N_19702);
nor U21810 (N_21810,N_19548,N_19667);
nand U21811 (N_21811,N_18287,N_19820);
xnor U21812 (N_21812,N_18436,N_18638);
and U21813 (N_21813,N_18146,N_17721);
and U21814 (N_21814,N_18539,N_19640);
or U21815 (N_21815,N_17962,N_17535);
nor U21816 (N_21816,N_19551,N_19372);
nand U21817 (N_21817,N_18039,N_18099);
xnor U21818 (N_21818,N_17617,N_18638);
nor U21819 (N_21819,N_19763,N_19725);
or U21820 (N_21820,N_18891,N_18843);
nor U21821 (N_21821,N_19916,N_18715);
or U21822 (N_21822,N_17589,N_19384);
nor U21823 (N_21823,N_19812,N_17702);
and U21824 (N_21824,N_18128,N_18549);
nand U21825 (N_21825,N_18081,N_17845);
or U21826 (N_21826,N_19847,N_19421);
xor U21827 (N_21827,N_18388,N_19144);
or U21828 (N_21828,N_19040,N_18543);
and U21829 (N_21829,N_19051,N_19081);
or U21830 (N_21830,N_17875,N_18563);
xnor U21831 (N_21831,N_18763,N_19799);
nor U21832 (N_21832,N_19976,N_18944);
nor U21833 (N_21833,N_17987,N_17761);
nor U21834 (N_21834,N_18507,N_17644);
nor U21835 (N_21835,N_18486,N_18563);
or U21836 (N_21836,N_19184,N_19681);
xor U21837 (N_21837,N_18027,N_18365);
nand U21838 (N_21838,N_17620,N_19220);
or U21839 (N_21839,N_17844,N_18816);
nor U21840 (N_21840,N_18080,N_17565);
nand U21841 (N_21841,N_19464,N_19186);
xnor U21842 (N_21842,N_19174,N_17877);
nand U21843 (N_21843,N_19100,N_19722);
xor U21844 (N_21844,N_18734,N_19101);
xnor U21845 (N_21845,N_17858,N_18369);
xor U21846 (N_21846,N_18717,N_17776);
nor U21847 (N_21847,N_19017,N_17580);
or U21848 (N_21848,N_19299,N_18951);
xor U21849 (N_21849,N_18589,N_17668);
nand U21850 (N_21850,N_17940,N_18972);
nor U21851 (N_21851,N_17686,N_19701);
xor U21852 (N_21852,N_19373,N_17872);
nor U21853 (N_21853,N_17975,N_19667);
xnor U21854 (N_21854,N_18758,N_17883);
and U21855 (N_21855,N_18719,N_18642);
or U21856 (N_21856,N_18015,N_19023);
or U21857 (N_21857,N_17818,N_18312);
xor U21858 (N_21858,N_19719,N_19057);
nand U21859 (N_21859,N_19760,N_18818);
and U21860 (N_21860,N_18342,N_19551);
or U21861 (N_21861,N_18732,N_18560);
or U21862 (N_21862,N_19725,N_19635);
nor U21863 (N_21863,N_19652,N_19744);
and U21864 (N_21864,N_19634,N_18536);
or U21865 (N_21865,N_17853,N_19375);
and U21866 (N_21866,N_18856,N_18648);
nor U21867 (N_21867,N_18163,N_17828);
and U21868 (N_21868,N_19704,N_18922);
nand U21869 (N_21869,N_17855,N_19156);
xor U21870 (N_21870,N_19877,N_18346);
xnor U21871 (N_21871,N_18489,N_18826);
nand U21872 (N_21872,N_18218,N_19011);
nor U21873 (N_21873,N_17943,N_17834);
or U21874 (N_21874,N_19980,N_17946);
and U21875 (N_21875,N_19674,N_18551);
xnor U21876 (N_21876,N_19104,N_19663);
xnor U21877 (N_21877,N_18259,N_19747);
xor U21878 (N_21878,N_19487,N_18927);
nand U21879 (N_21879,N_18030,N_17866);
and U21880 (N_21880,N_17996,N_18397);
or U21881 (N_21881,N_17731,N_18973);
nor U21882 (N_21882,N_19757,N_19350);
xnor U21883 (N_21883,N_19054,N_18914);
xnor U21884 (N_21884,N_19265,N_18229);
or U21885 (N_21885,N_18952,N_19128);
xnor U21886 (N_21886,N_17538,N_18214);
or U21887 (N_21887,N_17910,N_19080);
xnor U21888 (N_21888,N_17593,N_19651);
nand U21889 (N_21889,N_17723,N_19258);
nor U21890 (N_21890,N_18023,N_19489);
xor U21891 (N_21891,N_18088,N_19169);
or U21892 (N_21892,N_19194,N_18945);
nor U21893 (N_21893,N_19264,N_18714);
nand U21894 (N_21894,N_18636,N_17633);
and U21895 (N_21895,N_18517,N_19041);
xnor U21896 (N_21896,N_19223,N_19360);
or U21897 (N_21897,N_18829,N_18337);
xnor U21898 (N_21898,N_19446,N_18913);
nor U21899 (N_21899,N_18069,N_18091);
xnor U21900 (N_21900,N_18299,N_19318);
nand U21901 (N_21901,N_18552,N_19297);
and U21902 (N_21902,N_18945,N_19862);
and U21903 (N_21903,N_19014,N_18117);
nand U21904 (N_21904,N_17507,N_19806);
nor U21905 (N_21905,N_18056,N_18905);
and U21906 (N_21906,N_17799,N_18947);
nor U21907 (N_21907,N_18769,N_19390);
xnor U21908 (N_21908,N_18628,N_18867);
and U21909 (N_21909,N_17747,N_17757);
or U21910 (N_21910,N_18368,N_19564);
xnor U21911 (N_21911,N_18937,N_19043);
or U21912 (N_21912,N_18076,N_18972);
or U21913 (N_21913,N_18933,N_18773);
nor U21914 (N_21914,N_19275,N_19791);
nor U21915 (N_21915,N_18638,N_17758);
xor U21916 (N_21916,N_18466,N_18282);
nand U21917 (N_21917,N_19203,N_19418);
nor U21918 (N_21918,N_17974,N_18823);
and U21919 (N_21919,N_17742,N_18528);
and U21920 (N_21920,N_19727,N_17924);
or U21921 (N_21921,N_19599,N_19004);
and U21922 (N_21922,N_17956,N_19340);
or U21923 (N_21923,N_19811,N_17522);
nor U21924 (N_21924,N_17640,N_18281);
nor U21925 (N_21925,N_19870,N_17982);
nor U21926 (N_21926,N_18047,N_19334);
or U21927 (N_21927,N_18887,N_19147);
and U21928 (N_21928,N_18890,N_17700);
and U21929 (N_21929,N_19826,N_17731);
nand U21930 (N_21930,N_17567,N_19007);
xor U21931 (N_21931,N_19677,N_18059);
nor U21932 (N_21932,N_19510,N_18734);
or U21933 (N_21933,N_18259,N_19265);
nand U21934 (N_21934,N_18757,N_18632);
and U21935 (N_21935,N_19617,N_17506);
xor U21936 (N_21936,N_17563,N_19349);
nand U21937 (N_21937,N_17811,N_18429);
xor U21938 (N_21938,N_18549,N_19230);
or U21939 (N_21939,N_19737,N_19908);
nor U21940 (N_21940,N_18299,N_18323);
xor U21941 (N_21941,N_19911,N_18304);
nand U21942 (N_21942,N_18022,N_17731);
nand U21943 (N_21943,N_19594,N_19189);
or U21944 (N_21944,N_17537,N_17710);
nand U21945 (N_21945,N_18457,N_17957);
and U21946 (N_21946,N_17770,N_18980);
or U21947 (N_21947,N_18545,N_18651);
and U21948 (N_21948,N_18313,N_17502);
nor U21949 (N_21949,N_19638,N_18400);
nand U21950 (N_21950,N_18568,N_19914);
nor U21951 (N_21951,N_19346,N_19207);
nor U21952 (N_21952,N_19347,N_18690);
nor U21953 (N_21953,N_18147,N_18944);
xnor U21954 (N_21954,N_18838,N_19683);
xor U21955 (N_21955,N_19211,N_19930);
nor U21956 (N_21956,N_19822,N_18140);
and U21957 (N_21957,N_18128,N_18189);
and U21958 (N_21958,N_19236,N_17843);
nor U21959 (N_21959,N_18346,N_18313);
nor U21960 (N_21960,N_18066,N_19794);
xnor U21961 (N_21961,N_19151,N_17506);
nor U21962 (N_21962,N_18095,N_19901);
nand U21963 (N_21963,N_18228,N_18852);
and U21964 (N_21964,N_18636,N_19397);
nor U21965 (N_21965,N_17754,N_18231);
nand U21966 (N_21966,N_19346,N_18853);
or U21967 (N_21967,N_19960,N_19034);
nor U21968 (N_21968,N_18298,N_19178);
xnor U21969 (N_21969,N_18874,N_19750);
xnor U21970 (N_21970,N_19305,N_19802);
and U21971 (N_21971,N_18529,N_19761);
or U21972 (N_21972,N_18627,N_18024);
xor U21973 (N_21973,N_18848,N_18735);
xor U21974 (N_21974,N_18464,N_19536);
or U21975 (N_21975,N_19634,N_17969);
and U21976 (N_21976,N_17555,N_18368);
or U21977 (N_21977,N_18461,N_17663);
nor U21978 (N_21978,N_18150,N_19734);
and U21979 (N_21979,N_19330,N_18599);
nand U21980 (N_21980,N_17534,N_19028);
or U21981 (N_21981,N_17946,N_19173);
or U21982 (N_21982,N_18297,N_18115);
nand U21983 (N_21983,N_19735,N_19035);
or U21984 (N_21984,N_17566,N_18742);
xor U21985 (N_21985,N_17632,N_19435);
and U21986 (N_21986,N_19434,N_19314);
or U21987 (N_21987,N_19158,N_19995);
or U21988 (N_21988,N_17954,N_19390);
and U21989 (N_21989,N_18387,N_19530);
or U21990 (N_21990,N_19152,N_18825);
nor U21991 (N_21991,N_19321,N_18315);
nand U21992 (N_21992,N_19289,N_18076);
xor U21993 (N_21993,N_17796,N_18980);
and U21994 (N_21994,N_18001,N_19849);
or U21995 (N_21995,N_18511,N_19185);
xor U21996 (N_21996,N_19201,N_18555);
xor U21997 (N_21997,N_19997,N_19290);
or U21998 (N_21998,N_17599,N_17620);
xor U21999 (N_21999,N_17854,N_17853);
or U22000 (N_22000,N_19637,N_19082);
nand U22001 (N_22001,N_17799,N_19083);
nand U22002 (N_22002,N_19277,N_18141);
nand U22003 (N_22003,N_17578,N_17918);
or U22004 (N_22004,N_18913,N_18440);
nand U22005 (N_22005,N_18856,N_17656);
nand U22006 (N_22006,N_19239,N_18183);
or U22007 (N_22007,N_17803,N_19747);
nand U22008 (N_22008,N_18157,N_19063);
or U22009 (N_22009,N_18230,N_19087);
nor U22010 (N_22010,N_18557,N_19082);
xnor U22011 (N_22011,N_19570,N_18553);
nor U22012 (N_22012,N_18823,N_19180);
nor U22013 (N_22013,N_18945,N_17997);
nor U22014 (N_22014,N_17633,N_18194);
nand U22015 (N_22015,N_19668,N_18492);
and U22016 (N_22016,N_19996,N_18161);
xnor U22017 (N_22017,N_19592,N_19827);
and U22018 (N_22018,N_19007,N_17954);
and U22019 (N_22019,N_17675,N_17986);
nand U22020 (N_22020,N_17730,N_19149);
and U22021 (N_22021,N_19067,N_19069);
or U22022 (N_22022,N_18969,N_19047);
xor U22023 (N_22023,N_19591,N_18041);
or U22024 (N_22024,N_18433,N_18097);
and U22025 (N_22025,N_19589,N_18483);
nand U22026 (N_22026,N_17822,N_17579);
nor U22027 (N_22027,N_18531,N_19130);
nand U22028 (N_22028,N_19164,N_18804);
nor U22029 (N_22029,N_18956,N_18562);
nor U22030 (N_22030,N_17555,N_18689);
or U22031 (N_22031,N_17783,N_17769);
nand U22032 (N_22032,N_17710,N_18586);
nand U22033 (N_22033,N_19517,N_17800);
xor U22034 (N_22034,N_17513,N_17733);
nor U22035 (N_22035,N_19293,N_18464);
xor U22036 (N_22036,N_19562,N_19375);
xor U22037 (N_22037,N_19915,N_17693);
or U22038 (N_22038,N_18622,N_17633);
and U22039 (N_22039,N_17959,N_19456);
xnor U22040 (N_22040,N_18891,N_17717);
nor U22041 (N_22041,N_19764,N_19055);
nand U22042 (N_22042,N_18309,N_17652);
nand U22043 (N_22043,N_19938,N_17536);
xnor U22044 (N_22044,N_18251,N_18092);
and U22045 (N_22045,N_18254,N_18723);
nor U22046 (N_22046,N_18027,N_19203);
xnor U22047 (N_22047,N_18820,N_17788);
or U22048 (N_22048,N_18216,N_17636);
xor U22049 (N_22049,N_19360,N_19308);
and U22050 (N_22050,N_17648,N_19087);
and U22051 (N_22051,N_18340,N_17586);
and U22052 (N_22052,N_19845,N_17800);
or U22053 (N_22053,N_18966,N_18339);
and U22054 (N_22054,N_19796,N_18696);
xnor U22055 (N_22055,N_18821,N_17547);
nand U22056 (N_22056,N_19121,N_17512);
or U22057 (N_22057,N_18557,N_19202);
nor U22058 (N_22058,N_19587,N_19145);
and U22059 (N_22059,N_19824,N_18239);
nor U22060 (N_22060,N_19529,N_17714);
nand U22061 (N_22061,N_19825,N_19237);
xor U22062 (N_22062,N_17738,N_18124);
or U22063 (N_22063,N_18298,N_17501);
or U22064 (N_22064,N_18061,N_17547);
nand U22065 (N_22065,N_19408,N_18403);
and U22066 (N_22066,N_18865,N_17514);
and U22067 (N_22067,N_18563,N_18915);
or U22068 (N_22068,N_18808,N_19881);
and U22069 (N_22069,N_19517,N_19984);
or U22070 (N_22070,N_18812,N_19181);
or U22071 (N_22071,N_19409,N_19155);
or U22072 (N_22072,N_19955,N_19526);
or U22073 (N_22073,N_19097,N_17813);
or U22074 (N_22074,N_19150,N_19377);
and U22075 (N_22075,N_17625,N_18384);
or U22076 (N_22076,N_18292,N_17749);
nand U22077 (N_22077,N_19586,N_19150);
nor U22078 (N_22078,N_18548,N_19572);
and U22079 (N_22079,N_19892,N_18591);
nand U22080 (N_22080,N_19771,N_18928);
nor U22081 (N_22081,N_18655,N_18297);
nor U22082 (N_22082,N_18895,N_17779);
or U22083 (N_22083,N_19487,N_18279);
and U22084 (N_22084,N_18931,N_17763);
or U22085 (N_22085,N_18078,N_18271);
xnor U22086 (N_22086,N_17747,N_18500);
or U22087 (N_22087,N_17595,N_18146);
xnor U22088 (N_22088,N_18774,N_18788);
nand U22089 (N_22089,N_18370,N_18343);
and U22090 (N_22090,N_18996,N_17999);
and U22091 (N_22091,N_18149,N_19006);
nor U22092 (N_22092,N_17800,N_18332);
xnor U22093 (N_22093,N_18345,N_17817);
nand U22094 (N_22094,N_17704,N_18822);
or U22095 (N_22095,N_19596,N_18457);
nand U22096 (N_22096,N_18175,N_19795);
nor U22097 (N_22097,N_18503,N_19184);
or U22098 (N_22098,N_18403,N_18037);
nor U22099 (N_22099,N_17618,N_18242);
nor U22100 (N_22100,N_17620,N_19676);
and U22101 (N_22101,N_18887,N_19965);
or U22102 (N_22102,N_18139,N_18360);
nand U22103 (N_22103,N_17750,N_17826);
nor U22104 (N_22104,N_19168,N_18249);
or U22105 (N_22105,N_17869,N_18882);
xor U22106 (N_22106,N_18534,N_18260);
nand U22107 (N_22107,N_18704,N_18703);
and U22108 (N_22108,N_18220,N_19745);
nand U22109 (N_22109,N_17700,N_19300);
and U22110 (N_22110,N_18136,N_18371);
nand U22111 (N_22111,N_18845,N_19601);
nand U22112 (N_22112,N_17630,N_18002);
or U22113 (N_22113,N_17697,N_18854);
nor U22114 (N_22114,N_19187,N_19933);
xnor U22115 (N_22115,N_18267,N_19930);
xor U22116 (N_22116,N_17876,N_19432);
nand U22117 (N_22117,N_18094,N_18160);
nor U22118 (N_22118,N_19882,N_18081);
and U22119 (N_22119,N_19623,N_18792);
or U22120 (N_22120,N_18602,N_19230);
nand U22121 (N_22121,N_18695,N_18195);
nand U22122 (N_22122,N_19822,N_19239);
nand U22123 (N_22123,N_19042,N_18171);
nor U22124 (N_22124,N_18861,N_19689);
or U22125 (N_22125,N_19834,N_19085);
or U22126 (N_22126,N_18165,N_19743);
or U22127 (N_22127,N_18271,N_19451);
nor U22128 (N_22128,N_19376,N_19749);
xor U22129 (N_22129,N_19469,N_19075);
or U22130 (N_22130,N_18289,N_19971);
xnor U22131 (N_22131,N_18549,N_17689);
nor U22132 (N_22132,N_18152,N_19188);
nor U22133 (N_22133,N_19706,N_19694);
and U22134 (N_22134,N_18249,N_18180);
nand U22135 (N_22135,N_19161,N_19927);
nor U22136 (N_22136,N_18760,N_19410);
nand U22137 (N_22137,N_19631,N_18446);
xor U22138 (N_22138,N_18635,N_18380);
nor U22139 (N_22139,N_19011,N_18382);
or U22140 (N_22140,N_19799,N_18772);
and U22141 (N_22141,N_17830,N_18670);
nand U22142 (N_22142,N_18926,N_18573);
nand U22143 (N_22143,N_19071,N_19844);
or U22144 (N_22144,N_19490,N_17635);
xnor U22145 (N_22145,N_17860,N_17518);
xnor U22146 (N_22146,N_18844,N_17967);
nand U22147 (N_22147,N_19115,N_19797);
or U22148 (N_22148,N_17692,N_17996);
nand U22149 (N_22149,N_18051,N_19674);
nor U22150 (N_22150,N_17563,N_19482);
and U22151 (N_22151,N_17592,N_19328);
or U22152 (N_22152,N_19131,N_18958);
and U22153 (N_22153,N_18098,N_18962);
or U22154 (N_22154,N_18411,N_17507);
or U22155 (N_22155,N_18380,N_19632);
or U22156 (N_22156,N_18503,N_19378);
nand U22157 (N_22157,N_19305,N_18029);
nor U22158 (N_22158,N_19969,N_18126);
and U22159 (N_22159,N_19056,N_19212);
and U22160 (N_22160,N_19326,N_19792);
nand U22161 (N_22161,N_19389,N_19846);
and U22162 (N_22162,N_18463,N_19876);
nor U22163 (N_22163,N_18230,N_17872);
and U22164 (N_22164,N_18184,N_18357);
and U22165 (N_22165,N_18449,N_17743);
or U22166 (N_22166,N_19181,N_17663);
nor U22167 (N_22167,N_19408,N_19543);
xor U22168 (N_22168,N_18200,N_17633);
or U22169 (N_22169,N_19185,N_18168);
nor U22170 (N_22170,N_18672,N_17612);
xnor U22171 (N_22171,N_19090,N_19231);
and U22172 (N_22172,N_18010,N_19178);
nand U22173 (N_22173,N_19475,N_18277);
nand U22174 (N_22174,N_19092,N_19867);
nor U22175 (N_22175,N_18796,N_18995);
or U22176 (N_22176,N_17889,N_18628);
or U22177 (N_22177,N_19503,N_18421);
nand U22178 (N_22178,N_19407,N_17632);
xor U22179 (N_22179,N_19528,N_19913);
nor U22180 (N_22180,N_19988,N_18375);
nor U22181 (N_22181,N_18435,N_17742);
nand U22182 (N_22182,N_19892,N_17897);
or U22183 (N_22183,N_19121,N_18886);
or U22184 (N_22184,N_18691,N_18871);
and U22185 (N_22185,N_19591,N_19573);
and U22186 (N_22186,N_19444,N_19967);
nor U22187 (N_22187,N_19801,N_18783);
nor U22188 (N_22188,N_19384,N_18149);
or U22189 (N_22189,N_18134,N_18203);
xor U22190 (N_22190,N_19873,N_19325);
xnor U22191 (N_22191,N_18921,N_17979);
xor U22192 (N_22192,N_17542,N_18351);
nor U22193 (N_22193,N_19437,N_18722);
nor U22194 (N_22194,N_19344,N_19571);
or U22195 (N_22195,N_18046,N_18514);
nor U22196 (N_22196,N_19104,N_19838);
xnor U22197 (N_22197,N_18559,N_18403);
nor U22198 (N_22198,N_18788,N_17835);
nand U22199 (N_22199,N_18327,N_19372);
nand U22200 (N_22200,N_19668,N_18350);
or U22201 (N_22201,N_19651,N_18510);
nor U22202 (N_22202,N_19199,N_19848);
nand U22203 (N_22203,N_19252,N_19599);
and U22204 (N_22204,N_19681,N_18210);
and U22205 (N_22205,N_18161,N_18397);
or U22206 (N_22206,N_18395,N_18427);
xor U22207 (N_22207,N_18190,N_18462);
xor U22208 (N_22208,N_18078,N_18988);
nand U22209 (N_22209,N_19018,N_18512);
or U22210 (N_22210,N_18590,N_18915);
xnor U22211 (N_22211,N_18263,N_19576);
xnor U22212 (N_22212,N_19101,N_17713);
xnor U22213 (N_22213,N_19141,N_19418);
or U22214 (N_22214,N_18286,N_19513);
xor U22215 (N_22215,N_19167,N_19513);
or U22216 (N_22216,N_17825,N_18173);
and U22217 (N_22217,N_18202,N_19682);
xnor U22218 (N_22218,N_19716,N_18472);
xnor U22219 (N_22219,N_17807,N_19335);
nor U22220 (N_22220,N_18095,N_18123);
or U22221 (N_22221,N_19471,N_17921);
nand U22222 (N_22222,N_18502,N_17729);
nor U22223 (N_22223,N_19454,N_18938);
nand U22224 (N_22224,N_18470,N_17623);
nand U22225 (N_22225,N_18581,N_18567);
xor U22226 (N_22226,N_18188,N_19154);
or U22227 (N_22227,N_19612,N_19601);
xnor U22228 (N_22228,N_19930,N_18650);
and U22229 (N_22229,N_17995,N_19574);
or U22230 (N_22230,N_18743,N_19671);
nor U22231 (N_22231,N_19360,N_19142);
nor U22232 (N_22232,N_17882,N_17879);
nor U22233 (N_22233,N_17874,N_19207);
nor U22234 (N_22234,N_19986,N_18346);
and U22235 (N_22235,N_18233,N_17913);
or U22236 (N_22236,N_19468,N_18680);
nand U22237 (N_22237,N_17738,N_19945);
or U22238 (N_22238,N_18683,N_19751);
nor U22239 (N_22239,N_19904,N_19237);
nand U22240 (N_22240,N_18063,N_19180);
or U22241 (N_22241,N_18477,N_19799);
xor U22242 (N_22242,N_19645,N_19979);
xor U22243 (N_22243,N_18738,N_19390);
xnor U22244 (N_22244,N_18141,N_17935);
xnor U22245 (N_22245,N_19728,N_19480);
nor U22246 (N_22246,N_18464,N_18115);
nor U22247 (N_22247,N_18609,N_19600);
nand U22248 (N_22248,N_19852,N_19648);
nand U22249 (N_22249,N_18381,N_17507);
nand U22250 (N_22250,N_18649,N_18291);
or U22251 (N_22251,N_19479,N_18178);
or U22252 (N_22252,N_19811,N_19923);
nor U22253 (N_22253,N_19992,N_19101);
nor U22254 (N_22254,N_17688,N_18045);
and U22255 (N_22255,N_17977,N_18856);
and U22256 (N_22256,N_18998,N_19853);
and U22257 (N_22257,N_17821,N_19160);
or U22258 (N_22258,N_19204,N_18513);
nand U22259 (N_22259,N_18288,N_19198);
and U22260 (N_22260,N_17777,N_18247);
nand U22261 (N_22261,N_19605,N_18066);
nand U22262 (N_22262,N_18708,N_17808);
and U22263 (N_22263,N_17635,N_18745);
or U22264 (N_22264,N_17651,N_19237);
or U22265 (N_22265,N_18383,N_18574);
and U22266 (N_22266,N_19996,N_18749);
and U22267 (N_22267,N_18079,N_18600);
nand U22268 (N_22268,N_19172,N_18778);
xnor U22269 (N_22269,N_19490,N_18345);
and U22270 (N_22270,N_19136,N_18616);
or U22271 (N_22271,N_18775,N_18909);
nor U22272 (N_22272,N_19548,N_18750);
nand U22273 (N_22273,N_19693,N_18230);
xnor U22274 (N_22274,N_19391,N_18278);
or U22275 (N_22275,N_18978,N_19566);
or U22276 (N_22276,N_19177,N_19732);
and U22277 (N_22277,N_18135,N_19712);
xnor U22278 (N_22278,N_19965,N_18995);
xnor U22279 (N_22279,N_19439,N_18964);
xnor U22280 (N_22280,N_19694,N_18010);
nor U22281 (N_22281,N_19023,N_19726);
nand U22282 (N_22282,N_18948,N_18159);
and U22283 (N_22283,N_18736,N_18113);
or U22284 (N_22284,N_18510,N_18281);
xor U22285 (N_22285,N_19075,N_19545);
xor U22286 (N_22286,N_18801,N_19087);
and U22287 (N_22287,N_19141,N_18169);
xnor U22288 (N_22288,N_18075,N_18033);
xnor U22289 (N_22289,N_17969,N_19339);
nor U22290 (N_22290,N_19884,N_18872);
or U22291 (N_22291,N_18808,N_19170);
and U22292 (N_22292,N_18364,N_18678);
nor U22293 (N_22293,N_19455,N_17904);
nand U22294 (N_22294,N_19421,N_19043);
nand U22295 (N_22295,N_18681,N_19060);
and U22296 (N_22296,N_18244,N_18600);
xnor U22297 (N_22297,N_17998,N_18338);
or U22298 (N_22298,N_18288,N_19700);
nor U22299 (N_22299,N_19625,N_19772);
nor U22300 (N_22300,N_17507,N_18363);
nand U22301 (N_22301,N_19368,N_17641);
nand U22302 (N_22302,N_19576,N_18698);
or U22303 (N_22303,N_19358,N_18498);
and U22304 (N_22304,N_17926,N_18841);
nor U22305 (N_22305,N_17787,N_18997);
or U22306 (N_22306,N_19263,N_19532);
and U22307 (N_22307,N_18186,N_18876);
and U22308 (N_22308,N_19763,N_19349);
nand U22309 (N_22309,N_19118,N_19304);
and U22310 (N_22310,N_19373,N_19922);
or U22311 (N_22311,N_18418,N_18059);
or U22312 (N_22312,N_19546,N_18116);
and U22313 (N_22313,N_18510,N_18001);
xor U22314 (N_22314,N_18929,N_19503);
nand U22315 (N_22315,N_18532,N_19118);
nor U22316 (N_22316,N_19692,N_19832);
or U22317 (N_22317,N_17748,N_19625);
nand U22318 (N_22318,N_18882,N_19861);
xnor U22319 (N_22319,N_19221,N_19822);
or U22320 (N_22320,N_19413,N_19539);
and U22321 (N_22321,N_17794,N_18192);
and U22322 (N_22322,N_19087,N_18295);
nor U22323 (N_22323,N_17557,N_18141);
xor U22324 (N_22324,N_18433,N_19411);
xnor U22325 (N_22325,N_19246,N_18574);
and U22326 (N_22326,N_19449,N_18389);
and U22327 (N_22327,N_19260,N_18019);
xor U22328 (N_22328,N_18692,N_19453);
nand U22329 (N_22329,N_18777,N_19094);
or U22330 (N_22330,N_17594,N_18946);
nor U22331 (N_22331,N_18689,N_18409);
and U22332 (N_22332,N_19847,N_18219);
nor U22333 (N_22333,N_19825,N_17783);
nand U22334 (N_22334,N_19710,N_19583);
and U22335 (N_22335,N_18423,N_18737);
or U22336 (N_22336,N_19894,N_18760);
xor U22337 (N_22337,N_19556,N_18757);
xor U22338 (N_22338,N_18650,N_18591);
and U22339 (N_22339,N_19205,N_18848);
xnor U22340 (N_22340,N_17734,N_19932);
nand U22341 (N_22341,N_19250,N_19312);
and U22342 (N_22342,N_17777,N_19353);
or U22343 (N_22343,N_19960,N_19212);
xor U22344 (N_22344,N_17883,N_19881);
or U22345 (N_22345,N_18993,N_18254);
or U22346 (N_22346,N_19159,N_18798);
and U22347 (N_22347,N_19991,N_19085);
and U22348 (N_22348,N_19400,N_19982);
nor U22349 (N_22349,N_19666,N_19596);
nor U22350 (N_22350,N_18480,N_18194);
nor U22351 (N_22351,N_19496,N_19952);
nor U22352 (N_22352,N_17610,N_19796);
xnor U22353 (N_22353,N_17686,N_17509);
and U22354 (N_22354,N_18395,N_19198);
nand U22355 (N_22355,N_18940,N_17917);
nor U22356 (N_22356,N_19164,N_17541);
or U22357 (N_22357,N_17857,N_19385);
nand U22358 (N_22358,N_19579,N_18702);
nor U22359 (N_22359,N_19211,N_18951);
nand U22360 (N_22360,N_17554,N_17620);
nand U22361 (N_22361,N_17604,N_19173);
xnor U22362 (N_22362,N_18630,N_17682);
xor U22363 (N_22363,N_18741,N_18003);
nor U22364 (N_22364,N_18793,N_19226);
nand U22365 (N_22365,N_17718,N_19658);
nand U22366 (N_22366,N_17740,N_18724);
nand U22367 (N_22367,N_17578,N_19898);
or U22368 (N_22368,N_18597,N_17756);
nand U22369 (N_22369,N_19749,N_17656);
nor U22370 (N_22370,N_18989,N_18093);
nand U22371 (N_22371,N_18153,N_19788);
xor U22372 (N_22372,N_17519,N_18048);
or U22373 (N_22373,N_19197,N_18308);
nor U22374 (N_22374,N_19959,N_17763);
nor U22375 (N_22375,N_19809,N_19325);
or U22376 (N_22376,N_17801,N_18339);
xor U22377 (N_22377,N_19463,N_17779);
or U22378 (N_22378,N_18321,N_19349);
or U22379 (N_22379,N_19629,N_19580);
and U22380 (N_22380,N_17953,N_18301);
xnor U22381 (N_22381,N_17903,N_19497);
xnor U22382 (N_22382,N_19398,N_17633);
xnor U22383 (N_22383,N_19785,N_18088);
nor U22384 (N_22384,N_18258,N_19611);
nor U22385 (N_22385,N_18722,N_18188);
nor U22386 (N_22386,N_17759,N_18082);
and U22387 (N_22387,N_18181,N_19331);
nor U22388 (N_22388,N_19491,N_18513);
xnor U22389 (N_22389,N_19356,N_18164);
nand U22390 (N_22390,N_19206,N_18756);
or U22391 (N_22391,N_19184,N_18501);
nand U22392 (N_22392,N_18291,N_19636);
nor U22393 (N_22393,N_18565,N_18642);
nor U22394 (N_22394,N_19217,N_19089);
or U22395 (N_22395,N_18578,N_17525);
nor U22396 (N_22396,N_18019,N_19626);
nor U22397 (N_22397,N_18013,N_18390);
and U22398 (N_22398,N_19535,N_18338);
xor U22399 (N_22399,N_19413,N_19321);
and U22400 (N_22400,N_18856,N_17750);
or U22401 (N_22401,N_19111,N_17976);
nand U22402 (N_22402,N_19294,N_19217);
or U22403 (N_22403,N_18419,N_18508);
nor U22404 (N_22404,N_18709,N_18260);
nand U22405 (N_22405,N_19144,N_17707);
nor U22406 (N_22406,N_17685,N_18722);
nand U22407 (N_22407,N_19452,N_19014);
xnor U22408 (N_22408,N_18733,N_18787);
xor U22409 (N_22409,N_18607,N_18803);
and U22410 (N_22410,N_19615,N_17762);
or U22411 (N_22411,N_19151,N_17713);
nand U22412 (N_22412,N_17797,N_19782);
or U22413 (N_22413,N_19137,N_19366);
nor U22414 (N_22414,N_19708,N_18468);
nand U22415 (N_22415,N_17668,N_18851);
nand U22416 (N_22416,N_17665,N_19340);
nor U22417 (N_22417,N_18351,N_18901);
and U22418 (N_22418,N_19442,N_18554);
or U22419 (N_22419,N_18268,N_18438);
and U22420 (N_22420,N_19988,N_19346);
nor U22421 (N_22421,N_18589,N_19565);
or U22422 (N_22422,N_19400,N_18276);
nor U22423 (N_22423,N_19076,N_19097);
xor U22424 (N_22424,N_19871,N_19453);
nor U22425 (N_22425,N_19975,N_19188);
xor U22426 (N_22426,N_18434,N_18383);
nand U22427 (N_22427,N_19268,N_19279);
or U22428 (N_22428,N_18399,N_19818);
xnor U22429 (N_22429,N_17724,N_19495);
nand U22430 (N_22430,N_18345,N_17841);
and U22431 (N_22431,N_19193,N_19883);
nor U22432 (N_22432,N_18425,N_19566);
nor U22433 (N_22433,N_17978,N_18320);
and U22434 (N_22434,N_19774,N_17809);
nand U22435 (N_22435,N_18037,N_18433);
or U22436 (N_22436,N_17784,N_19531);
nand U22437 (N_22437,N_19810,N_17706);
xor U22438 (N_22438,N_17967,N_17808);
nand U22439 (N_22439,N_19973,N_17666);
nand U22440 (N_22440,N_18335,N_19724);
xnor U22441 (N_22441,N_19369,N_18699);
nor U22442 (N_22442,N_18335,N_19103);
nand U22443 (N_22443,N_19386,N_19089);
or U22444 (N_22444,N_19216,N_19474);
nand U22445 (N_22445,N_17828,N_17617);
nand U22446 (N_22446,N_19531,N_19764);
nor U22447 (N_22447,N_19039,N_18598);
or U22448 (N_22448,N_17700,N_18424);
xnor U22449 (N_22449,N_19069,N_17838);
nor U22450 (N_22450,N_19494,N_18038);
nor U22451 (N_22451,N_17761,N_19050);
and U22452 (N_22452,N_19389,N_18766);
xnor U22453 (N_22453,N_19691,N_18806);
or U22454 (N_22454,N_18235,N_19663);
or U22455 (N_22455,N_19305,N_17806);
xnor U22456 (N_22456,N_17550,N_18653);
xnor U22457 (N_22457,N_18957,N_19778);
nor U22458 (N_22458,N_17967,N_19196);
and U22459 (N_22459,N_19321,N_19368);
nor U22460 (N_22460,N_18323,N_19575);
nand U22461 (N_22461,N_17605,N_18418);
nor U22462 (N_22462,N_18524,N_18376);
nor U22463 (N_22463,N_17574,N_19124);
nor U22464 (N_22464,N_17833,N_18981);
xnor U22465 (N_22465,N_19132,N_17948);
and U22466 (N_22466,N_19572,N_17904);
nand U22467 (N_22467,N_17584,N_18057);
nand U22468 (N_22468,N_17794,N_19347);
xor U22469 (N_22469,N_17783,N_18044);
xor U22470 (N_22470,N_18081,N_18450);
and U22471 (N_22471,N_19313,N_19319);
nor U22472 (N_22472,N_17567,N_19274);
xor U22473 (N_22473,N_19690,N_18890);
xnor U22474 (N_22474,N_18196,N_19871);
xnor U22475 (N_22475,N_19881,N_17945);
and U22476 (N_22476,N_19179,N_18077);
and U22477 (N_22477,N_17887,N_18687);
xnor U22478 (N_22478,N_19723,N_19403);
and U22479 (N_22479,N_18809,N_17656);
or U22480 (N_22480,N_19037,N_17920);
nor U22481 (N_22481,N_17645,N_17984);
and U22482 (N_22482,N_18759,N_19533);
nand U22483 (N_22483,N_17917,N_18650);
or U22484 (N_22484,N_18469,N_19436);
or U22485 (N_22485,N_17619,N_18741);
xnor U22486 (N_22486,N_18545,N_18619);
xor U22487 (N_22487,N_18644,N_18323);
nor U22488 (N_22488,N_18541,N_19435);
xnor U22489 (N_22489,N_17821,N_19621);
xor U22490 (N_22490,N_19873,N_19134);
xor U22491 (N_22491,N_18199,N_18155);
and U22492 (N_22492,N_19083,N_18382);
nand U22493 (N_22493,N_18345,N_19567);
and U22494 (N_22494,N_18322,N_19122);
or U22495 (N_22495,N_17641,N_19711);
and U22496 (N_22496,N_17594,N_17916);
and U22497 (N_22497,N_18223,N_18133);
or U22498 (N_22498,N_18604,N_19794);
or U22499 (N_22499,N_18206,N_18848);
or U22500 (N_22500,N_20778,N_20850);
nor U22501 (N_22501,N_22341,N_22062);
nand U22502 (N_22502,N_21666,N_21094);
and U22503 (N_22503,N_20518,N_21265);
or U22504 (N_22504,N_21281,N_21180);
nand U22505 (N_22505,N_20992,N_21851);
xnor U22506 (N_22506,N_21423,N_21704);
nand U22507 (N_22507,N_20797,N_21867);
nor U22508 (N_22508,N_20431,N_21780);
xor U22509 (N_22509,N_20250,N_20294);
or U22510 (N_22510,N_22453,N_20001);
nor U22511 (N_22511,N_20826,N_20280);
nor U22512 (N_22512,N_21403,N_20696);
nand U22513 (N_22513,N_21231,N_21257);
nor U22514 (N_22514,N_21635,N_21646);
and U22515 (N_22515,N_22193,N_20028);
xor U22516 (N_22516,N_20003,N_20502);
nand U22517 (N_22517,N_21830,N_21847);
nand U22518 (N_22518,N_20589,N_22337);
nor U22519 (N_22519,N_22000,N_22447);
or U22520 (N_22520,N_20757,N_20705);
nand U22521 (N_22521,N_22104,N_21006);
nor U22522 (N_22522,N_20836,N_20307);
nand U22523 (N_22523,N_21116,N_20766);
and U22524 (N_22524,N_21648,N_21579);
nand U22525 (N_22525,N_21673,N_20122);
nor U22526 (N_22526,N_20442,N_20851);
and U22527 (N_22527,N_22041,N_21630);
or U22528 (N_22528,N_22315,N_21819);
nor U22529 (N_22529,N_22162,N_21395);
or U22530 (N_22530,N_21751,N_21814);
nand U22531 (N_22531,N_20828,N_21963);
xnor U22532 (N_22532,N_21296,N_22357);
nor U22533 (N_22533,N_21409,N_20584);
and U22534 (N_22534,N_22072,N_21383);
or U22535 (N_22535,N_20939,N_20593);
or U22536 (N_22536,N_20603,N_22141);
nor U22537 (N_22537,N_21315,N_21767);
nor U22538 (N_22538,N_20954,N_21772);
nor U22539 (N_22539,N_21389,N_20635);
and U22540 (N_22540,N_20728,N_20081);
xnor U22541 (N_22541,N_21567,N_21424);
xor U22542 (N_22542,N_20950,N_20838);
nor U22543 (N_22543,N_20904,N_20746);
nor U22544 (N_22544,N_22407,N_21922);
or U22545 (N_22545,N_20161,N_21259);
or U22546 (N_22546,N_20066,N_21360);
or U22547 (N_22547,N_21698,N_20187);
nand U22548 (N_22548,N_20205,N_22251);
nand U22549 (N_22549,N_20643,N_21081);
or U22550 (N_22550,N_22347,N_21978);
and U22551 (N_22551,N_21743,N_20934);
nand U22552 (N_22552,N_21759,N_21996);
nor U22553 (N_22553,N_20395,N_21515);
nor U22554 (N_22554,N_21888,N_20374);
and U22555 (N_22555,N_21039,N_22277);
xnor U22556 (N_22556,N_21363,N_22384);
or U22557 (N_22557,N_20360,N_20346);
nand U22558 (N_22558,N_22353,N_22165);
and U22559 (N_22559,N_20881,N_20788);
nand U22560 (N_22560,N_21926,N_21657);
nand U22561 (N_22561,N_22014,N_22432);
nand U22562 (N_22562,N_22408,N_22022);
xnor U22563 (N_22563,N_22005,N_21884);
xor U22564 (N_22564,N_21077,N_21393);
nor U22565 (N_22565,N_21909,N_21735);
xor U22566 (N_22566,N_21527,N_21840);
and U22567 (N_22567,N_21397,N_20179);
or U22568 (N_22568,N_22271,N_22234);
nor U22569 (N_22569,N_21411,N_21222);
or U22570 (N_22570,N_20648,N_20932);
xor U22571 (N_22571,N_20978,N_21069);
nand U22572 (N_22572,N_20915,N_21047);
or U22573 (N_22573,N_21367,N_20784);
nor U22574 (N_22574,N_20270,N_21004);
nor U22575 (N_22575,N_21162,N_21811);
and U22576 (N_22576,N_20988,N_21833);
nor U22577 (N_22577,N_20683,N_21054);
nand U22578 (N_22578,N_21994,N_20641);
and U22579 (N_22579,N_21087,N_20156);
or U22580 (N_22580,N_20535,N_20961);
nand U22581 (N_22581,N_21481,N_22358);
nand U22582 (N_22582,N_21025,N_20661);
nand U22583 (N_22583,N_22469,N_21053);
or U22584 (N_22584,N_20802,N_20596);
and U22585 (N_22585,N_20040,N_22138);
and U22586 (N_22586,N_21100,N_21073);
nor U22587 (N_22587,N_21384,N_22371);
xnor U22588 (N_22588,N_21332,N_20198);
or U22589 (N_22589,N_20289,N_21610);
or U22590 (N_22590,N_21234,N_22496);
nand U22591 (N_22591,N_20494,N_22285);
nand U22592 (N_22592,N_20064,N_21364);
and U22593 (N_22593,N_22451,N_22435);
and U22594 (N_22594,N_21822,N_21981);
or U22595 (N_22595,N_22151,N_22485);
nand U22596 (N_22596,N_22120,N_20631);
or U22597 (N_22597,N_20243,N_22322);
and U22598 (N_22598,N_21096,N_21179);
nand U22599 (N_22599,N_20521,N_21607);
nor U22600 (N_22600,N_21799,N_21758);
xor U22601 (N_22601,N_20142,N_21969);
xor U22602 (N_22602,N_21672,N_22342);
nand U22603 (N_22603,N_22032,N_21968);
xor U22604 (N_22604,N_20335,N_20324);
nor U22605 (N_22605,N_20195,N_20392);
xnor U22606 (N_22606,N_20771,N_22215);
and U22607 (N_22607,N_21739,N_21573);
xnor U22608 (N_22608,N_22040,N_21189);
nor U22609 (N_22609,N_21581,N_20569);
or U22610 (N_22610,N_20565,N_20126);
or U22611 (N_22611,N_20211,N_22119);
xnor U22612 (N_22612,N_20450,N_20979);
and U22613 (N_22613,N_21316,N_22255);
xor U22614 (N_22614,N_21547,N_20472);
nor U22615 (N_22615,N_21876,N_20519);
or U22616 (N_22616,N_22340,N_20279);
nand U22617 (N_22617,N_21226,N_20647);
nor U22618 (N_22618,N_21569,N_21421);
nand U22619 (N_22619,N_21408,N_21707);
and U22620 (N_22620,N_21750,N_21987);
nor U22621 (N_22621,N_20088,N_20835);
or U22622 (N_22622,N_20514,N_21908);
and U22623 (N_22623,N_22064,N_20281);
nor U22624 (N_22624,N_20624,N_20403);
xnor U22625 (N_22625,N_21262,N_21385);
xnor U22626 (N_22626,N_22129,N_21390);
and U22627 (N_22627,N_22361,N_22012);
xnor U22628 (N_22628,N_20278,N_20191);
xor U22629 (N_22629,N_21499,N_22218);
xor U22630 (N_22630,N_21260,N_21146);
xor U22631 (N_22631,N_20348,N_21827);
and U22632 (N_22632,N_22352,N_20486);
and U22633 (N_22633,N_20076,N_22377);
nor U22634 (N_22634,N_22236,N_21855);
or U22635 (N_22635,N_21119,N_22490);
or U22636 (N_22636,N_20995,N_20970);
xor U22637 (N_22637,N_21609,N_22320);
nor U22638 (N_22638,N_22063,N_22254);
and U22639 (N_22639,N_21318,N_20257);
nor U22640 (N_22640,N_21651,N_21432);
xor U22641 (N_22641,N_20220,N_22449);
nand U22642 (N_22642,N_22202,N_21614);
nor U22643 (N_22643,N_20448,N_22133);
nand U22644 (N_22644,N_21307,N_20739);
xor U22645 (N_22645,N_21034,N_21115);
nand U22646 (N_22646,N_20049,N_20980);
and U22647 (N_22647,N_20884,N_21725);
and U22648 (N_22648,N_20394,N_20332);
nor U22649 (N_22649,N_20328,N_20599);
nor U22650 (N_22650,N_20938,N_20776);
nor U22651 (N_22651,N_21960,N_21687);
or U22652 (N_22652,N_20157,N_20352);
nor U22653 (N_22653,N_20704,N_21837);
nand U22654 (N_22654,N_20758,N_21204);
or U22655 (N_22655,N_20310,N_22441);
nand U22656 (N_22656,N_21021,N_20429);
xor U22657 (N_22657,N_21308,N_21214);
nor U22658 (N_22658,N_21498,N_21902);
nor U22659 (N_22659,N_22217,N_20695);
nor U22660 (N_22660,N_21661,N_20614);
xnor U22661 (N_22661,N_20618,N_21097);
nand U22662 (N_22662,N_20342,N_20852);
nand U22663 (N_22663,N_21156,N_20206);
nand U22664 (N_22664,N_20261,N_20436);
or U22665 (N_22665,N_21040,N_22111);
nand U22666 (N_22666,N_20622,N_20558);
xor U22667 (N_22667,N_20931,N_21414);
xor U22668 (N_22668,N_20740,N_20240);
nor U22669 (N_22669,N_21330,N_22175);
or U22670 (N_22670,N_21337,N_20759);
or U22671 (N_22671,N_20796,N_22126);
or U22672 (N_22672,N_22433,N_20662);
nand U22673 (N_22673,N_20207,N_20591);
xnor U22674 (N_22674,N_20953,N_21303);
nor U22675 (N_22675,N_22195,N_20414);
or U22676 (N_22676,N_21449,N_21613);
nor U22677 (N_22677,N_20132,N_22267);
and U22678 (N_22678,N_20125,N_22429);
and U22679 (N_22679,N_20227,N_22172);
xor U22680 (N_22680,N_21061,N_20685);
nor U22681 (N_22681,N_21496,N_20571);
and U22682 (N_22682,N_20060,N_22338);
and U22683 (N_22683,N_22048,N_20137);
nand U22684 (N_22684,N_21721,N_21187);
nand U22685 (N_22685,N_20869,N_20121);
or U22686 (N_22686,N_22065,N_21241);
nand U22687 (N_22687,N_20765,N_21741);
and U22688 (N_22688,N_21931,N_20547);
xor U22689 (N_22689,N_21205,N_20466);
nor U22690 (N_22690,N_20166,N_20221);
xor U22691 (N_22691,N_21340,N_20073);
nor U22692 (N_22692,N_21599,N_21401);
nand U22693 (N_22693,N_20288,N_20609);
and U22694 (N_22694,N_20406,N_20907);
and U22695 (N_22695,N_22379,N_21011);
nand U22696 (N_22696,N_20717,N_21717);
nand U22697 (N_22697,N_20928,N_20086);
or U22698 (N_22698,N_20480,N_21010);
xnor U22699 (N_22699,N_20181,N_21768);
xnor U22700 (N_22700,N_21882,N_22246);
nor U22701 (N_22701,N_20713,N_20204);
or U22702 (N_22702,N_21055,N_20886);
nor U22703 (N_22703,N_21427,N_20655);
or U22704 (N_22704,N_21985,N_22359);
nor U22705 (N_22705,N_21636,N_21106);
or U22706 (N_22706,N_20576,N_21153);
xor U22707 (N_22707,N_21368,N_22294);
nand U22708 (N_22708,N_20427,N_21706);
xnor U22709 (N_22709,N_21667,N_20016);
or U22710 (N_22710,N_21829,N_21365);
and U22711 (N_22711,N_22436,N_20541);
and U22712 (N_22712,N_22410,N_20537);
xor U22713 (N_22713,N_21605,N_22365);
or U22714 (N_22714,N_21771,N_22248);
nor U22715 (N_22715,N_20878,N_21826);
nor U22716 (N_22716,N_22149,N_20908);
and U22717 (N_22717,N_21183,N_20079);
or U22718 (N_22718,N_20200,N_20789);
nand U22719 (N_22719,N_21023,N_21977);
nand U22720 (N_22720,N_21326,N_21689);
nand U22721 (N_22721,N_21076,N_22108);
and U22722 (N_22722,N_21731,N_21132);
nor U22723 (N_22723,N_20941,N_20699);
nand U22724 (N_22724,N_20905,N_22393);
or U22725 (N_22725,N_21877,N_21934);
xor U22726 (N_22726,N_21165,N_22397);
nor U22727 (N_22727,N_22281,N_22488);
and U22728 (N_22728,N_20634,N_20391);
and U22729 (N_22729,N_21658,N_21975);
and U22730 (N_22730,N_21677,N_22049);
nand U22731 (N_22731,N_21891,N_21377);
and U22732 (N_22732,N_20301,N_20175);
nand U22733 (N_22733,N_20610,N_20943);
or U22734 (N_22734,N_20165,N_21310);
nor U22735 (N_22735,N_20860,N_20973);
or U22736 (N_22736,N_22015,N_21450);
or U22737 (N_22737,N_21225,N_20664);
and U22738 (N_22738,N_20871,N_21186);
nor U22739 (N_22739,N_21426,N_20912);
nor U22740 (N_22740,N_20022,N_21537);
xor U22741 (N_22741,N_21353,N_22194);
nor U22742 (N_22742,N_20801,N_22421);
nor U22743 (N_22743,N_21553,N_20082);
xnor U22744 (N_22744,N_20947,N_20302);
nor U22745 (N_22745,N_21805,N_21852);
or U22746 (N_22746,N_22306,N_21092);
and U22747 (N_22747,N_20870,N_22261);
nand U22748 (N_22748,N_20291,N_21105);
nand U22749 (N_22749,N_21320,N_21169);
nor U22750 (N_22750,N_20167,N_20265);
or U22751 (N_22751,N_20174,N_20188);
nand U22752 (N_22752,N_21208,N_20775);
nor U22753 (N_22753,N_21455,N_21945);
nor U22754 (N_22754,N_20501,N_20667);
xor U22755 (N_22755,N_22031,N_21086);
or U22756 (N_22756,N_21875,N_21720);
xnor U22757 (N_22757,N_22205,N_20151);
nand U22758 (N_22758,N_21272,N_20413);
and U22759 (N_22759,N_20671,N_20859);
nand U22760 (N_22760,N_22475,N_22304);
or U22761 (N_22761,N_21293,N_20083);
xor U22762 (N_22762,N_21082,N_20632);
or U22763 (N_22763,N_21338,N_21220);
nor U22764 (N_22764,N_20652,N_22226);
nand U22765 (N_22765,N_20949,N_20298);
and U22766 (N_22766,N_20135,N_22264);
and U22767 (N_22767,N_22197,N_22472);
nor U22768 (N_22768,N_21295,N_20026);
nand U22769 (N_22769,N_21331,N_21292);
nor U22770 (N_22770,N_21901,N_20090);
and U22771 (N_22771,N_21691,N_21774);
nor U22772 (N_22772,N_22047,N_20546);
or U22773 (N_22773,N_22235,N_20714);
nor U22774 (N_22774,N_21083,N_20260);
nand U22775 (N_22775,N_22057,N_21287);
nand U22776 (N_22776,N_21064,N_20650);
xor U22777 (N_22777,N_22188,N_21201);
and U22778 (N_22778,N_21150,N_21235);
or U22779 (N_22779,N_20865,N_22019);
xnor U22780 (N_22780,N_20942,N_20715);
xor U22781 (N_22781,N_20242,N_20991);
nand U22782 (N_22782,N_20485,N_20041);
and U22783 (N_22783,N_20783,N_21356);
and U22784 (N_22784,N_20574,N_21810);
nor U22785 (N_22785,N_22450,N_20477);
or U22786 (N_22786,N_22329,N_22333);
xnor U22787 (N_22787,N_21343,N_20321);
nor U22788 (N_22788,N_21534,N_20727);
nand U22789 (N_22789,N_21905,N_21379);
nor U22790 (N_22790,N_22495,N_21964);
xor U22791 (N_22791,N_22166,N_20960);
xor U22792 (N_22792,N_21580,N_22308);
or U22793 (N_22793,N_20330,N_21709);
xnor U22794 (N_22794,N_20130,N_20363);
nand U22795 (N_22795,N_21522,N_20665);
nand U22796 (N_22796,N_21650,N_21907);
nor U22797 (N_22797,N_21932,N_21122);
and U22798 (N_22798,N_20533,N_20951);
xnor U22799 (N_22799,N_22150,N_22098);
nor U22800 (N_22800,N_21020,N_21048);
or U22801 (N_22801,N_20767,N_22257);
xnor U22802 (N_22802,N_20538,N_20756);
and U22803 (N_22803,N_20670,N_22351);
nor U22804 (N_22804,N_20411,N_22044);
and U22805 (N_22805,N_20749,N_21467);
xnor U22806 (N_22806,N_20186,N_20013);
xor U22807 (N_22807,N_21806,N_22084);
xnor U22808 (N_22808,N_20620,N_21632);
and U22809 (N_22809,N_20072,N_21892);
and U22810 (N_22810,N_22375,N_21446);
or U22811 (N_22811,N_21641,N_20234);
or U22812 (N_22812,N_20127,N_20275);
and U22813 (N_22813,N_21746,N_21182);
nand U22814 (N_22814,N_20532,N_21280);
and U22815 (N_22815,N_21211,N_22383);
nand U22816 (N_22816,N_21133,N_22157);
xor U22817 (N_22817,N_20059,N_22278);
and U22818 (N_22818,N_20336,N_21958);
or U22819 (N_22819,N_21923,N_21246);
or U22820 (N_22820,N_21928,N_20921);
nand U22821 (N_22821,N_21655,N_20500);
nand U22822 (N_22822,N_22198,N_22258);
xor U22823 (N_22823,N_22069,N_21576);
nand U22824 (N_22824,N_22113,N_21074);
or U22825 (N_22825,N_20831,N_20772);
nand U22826 (N_22826,N_22229,N_21311);
nand U22827 (N_22827,N_20792,N_21688);
or U22828 (N_22828,N_21125,N_21894);
and U22829 (N_22829,N_21361,N_20284);
or U22830 (N_22830,N_20462,N_20226);
nor U22831 (N_22831,N_21369,N_20058);
or U22832 (N_22832,N_21342,N_20663);
and U22833 (N_22833,N_21800,N_20409);
and U22834 (N_22834,N_21559,N_21407);
and U22835 (N_22835,N_20731,N_21662);
nand U22836 (N_22836,N_20868,N_20734);
nand U22837 (N_22837,N_22189,N_21459);
and U22838 (N_22838,N_22091,N_20358);
nor U22839 (N_22839,N_21637,N_22356);
or U22840 (N_22840,N_20654,N_21845);
and U22841 (N_22841,N_22011,N_21857);
and U22842 (N_22842,N_20709,N_21873);
nand U22843 (N_22843,N_21917,N_21252);
and U22844 (N_22844,N_20046,N_20613);
nand U22845 (N_22845,N_21550,N_21197);
and U22846 (N_22846,N_21198,N_20113);
or U22847 (N_22847,N_21887,N_20787);
xnor U22848 (N_22848,N_20964,N_21117);
xor U22849 (N_22849,N_20366,N_21986);
and U22850 (N_22850,N_21859,N_20827);
or U22851 (N_22851,N_22403,N_22164);
or U22852 (N_22852,N_21843,N_20504);
nand U22853 (N_22853,N_21728,N_20209);
and U22854 (N_22854,N_21608,N_21807);
nand U22855 (N_22855,N_22137,N_21157);
or U22856 (N_22856,N_20735,N_20005);
or U22857 (N_22857,N_20522,N_21711);
nor U22858 (N_22858,N_21715,N_20525);
xnor U22859 (N_22859,N_21542,N_21302);
xnor U22860 (N_22860,N_21541,N_20723);
or U22861 (N_22861,N_22415,N_20148);
xnor U22862 (N_22862,N_20420,N_20441);
or U22863 (N_22863,N_20590,N_21992);
or U22864 (N_22864,N_22125,N_21675);
xnor U22865 (N_22865,N_21993,N_20790);
and U22866 (N_22866,N_20523,N_21112);
or U22867 (N_22867,N_22391,N_21883);
nand U22868 (N_22868,N_20119,N_20594);
and U22869 (N_22869,N_21846,N_21948);
or U22870 (N_22870,N_21041,N_21686);
nor U22871 (N_22871,N_22286,N_20183);
xnor U22872 (N_22872,N_21195,N_21416);
xnor U22873 (N_22873,N_21405,N_21477);
or U22874 (N_22874,N_20182,N_20552);
nor U22875 (N_22875,N_20024,N_20550);
nand U22876 (N_22876,N_20990,N_21701);
and U22877 (N_22877,N_20638,N_21294);
nor U22878 (N_22878,N_22275,N_20455);
xor U22879 (N_22879,N_20067,N_20512);
and U22880 (N_22880,N_22094,N_21284);
xnor U22881 (N_22881,N_20861,N_20743);
nor U22882 (N_22882,N_21912,N_21591);
nand U22883 (N_22883,N_20193,N_21890);
nor U22884 (N_22884,N_20967,N_21503);
and U22885 (N_22885,N_22420,N_21139);
nor U22886 (N_22886,N_20317,N_21463);
xor U22887 (N_22887,N_20585,N_20996);
nand U22888 (N_22888,N_20432,N_21842);
or U22889 (N_22889,N_22438,N_20019);
nand U22890 (N_22890,N_20112,N_22256);
or U22891 (N_22891,N_21410,N_21752);
nor U22892 (N_22892,N_22096,N_21695);
xor U22893 (N_22893,N_21504,N_22335);
nor U22894 (N_22894,N_22050,N_21161);
nor U22895 (N_22895,N_21713,N_21063);
nand U22896 (N_22896,N_21387,N_20601);
xnor U22897 (N_22897,N_21300,N_21797);
nor U22898 (N_22898,N_20520,N_20457);
xnor U22899 (N_22899,N_20602,N_22477);
and U22900 (N_22900,N_22483,N_20323);
or U22901 (N_22901,N_20829,N_21560);
nand U22902 (N_22902,N_22176,N_21391);
nor U22903 (N_22903,N_20820,N_20966);
xor U22904 (N_22904,N_22122,N_20267);
nor U22905 (N_22905,N_21680,N_20600);
nor U22906 (N_22906,N_20233,N_20417);
or U22907 (N_22907,N_20305,N_21080);
nand U22908 (N_22908,N_20810,N_20216);
nor U22909 (N_22909,N_20421,N_21825);
nand U22910 (N_22910,N_20678,N_20936);
or U22911 (N_22911,N_21374,N_20803);
or U22912 (N_22912,N_22362,N_21848);
nand U22913 (N_22913,N_22200,N_20171);
xor U22914 (N_22914,N_21032,N_21324);
and U22915 (N_22915,N_21600,N_20946);
xor U22916 (N_22916,N_21152,N_20557);
and U22917 (N_22917,N_21177,N_20239);
xnor U22918 (N_22918,N_20843,N_20000);
or U22919 (N_22919,N_20014,N_22136);
or U22920 (N_22920,N_20164,N_21528);
and U22921 (N_22921,N_20536,N_22029);
and U22922 (N_22922,N_20093,N_20168);
or U22923 (N_22923,N_20617,N_20312);
xnor U22924 (N_22924,N_22292,N_21606);
nand U22925 (N_22925,N_22370,N_21386);
and U22926 (N_22926,N_21479,N_20693);
and U22927 (N_22927,N_21555,N_21065);
and U22928 (N_22928,N_20659,N_20228);
xnor U22929 (N_22929,N_20390,N_20848);
nand U22930 (N_22930,N_20471,N_20476);
nor U22931 (N_22931,N_21016,N_20891);
and U22932 (N_22932,N_21946,N_22457);
nor U22933 (N_22933,N_20103,N_20292);
and U22934 (N_22934,N_20959,N_20170);
and U22935 (N_22935,N_21263,N_21228);
and U22936 (N_22936,N_20386,N_22115);
and U22937 (N_22937,N_20897,N_21586);
or U22938 (N_22938,N_22238,N_21130);
and U22939 (N_22939,N_20818,N_21545);
or U22940 (N_22940,N_21627,N_20208);
nor U22941 (N_22941,N_22241,N_20733);
or U22942 (N_22942,N_21967,N_22300);
or U22943 (N_22943,N_21430,N_22380);
nand U22944 (N_22944,N_21916,N_21154);
nand U22945 (N_22945,N_22387,N_21566);
or U22946 (N_22946,N_21714,N_21557);
or U22947 (N_22947,N_20568,N_20545);
nand U22948 (N_22948,N_21131,N_21649);
or U22949 (N_22949,N_22487,N_21699);
nor U22950 (N_22950,N_20027,N_20917);
xnor U22951 (N_22951,N_21137,N_20282);
or U22952 (N_22952,N_20986,N_20008);
xnor U22953 (N_22953,N_20854,N_22430);
or U22954 (N_22954,N_22039,N_21188);
or U22955 (N_22955,N_21619,N_20134);
nor U22956 (N_22956,N_20877,N_20674);
and U22957 (N_22957,N_20458,N_21170);
or U22958 (N_22958,N_21474,N_21038);
nor U22959 (N_22959,N_21242,N_21500);
nor U22960 (N_22960,N_20384,N_20178);
nor U22961 (N_22961,N_20143,N_20098);
nor U22962 (N_22962,N_21418,N_21435);
or U22963 (N_22963,N_21483,N_22309);
and U22964 (N_22964,N_20567,N_21428);
nand U22965 (N_22965,N_22140,N_20745);
or U22966 (N_22966,N_22045,N_22132);
nand U22967 (N_22967,N_21953,N_20464);
nand U22968 (N_22968,N_21535,N_22389);
nor U22969 (N_22969,N_21596,N_22034);
or U22970 (N_22970,N_21181,N_21400);
or U22971 (N_22971,N_21863,N_22321);
nand U22972 (N_22972,N_20977,N_22299);
xor U22973 (N_22973,N_20252,N_20190);
or U22974 (N_22974,N_21584,N_21118);
xnor U22975 (N_22975,N_20308,N_20491);
xnor U22976 (N_22976,N_20892,N_21267);
nand U22977 (N_22977,N_21603,N_21289);
nand U22978 (N_22978,N_21869,N_21854);
xnor U22979 (N_22979,N_21373,N_22401);
or U22980 (N_22980,N_20553,N_20981);
and U22981 (N_22981,N_21473,N_21939);
xor U22982 (N_22982,N_21861,N_21357);
and U22983 (N_22983,N_21744,N_22276);
nand U22984 (N_22984,N_20983,N_20779);
xor U22985 (N_22985,N_21935,N_21530);
nand U22986 (N_22986,N_20454,N_21820);
xnor U22987 (N_22987,N_20325,N_20976);
or U22988 (N_22988,N_21818,N_21413);
and U22989 (N_22989,N_20903,N_22004);
and U22990 (N_22990,N_20253,N_20372);
nor U22991 (N_22991,N_22478,N_21510);
nor U22992 (N_22992,N_20586,N_20511);
and U22993 (N_22993,N_20439,N_22180);
xnor U22994 (N_22994,N_20720,N_20393);
and U22995 (N_22995,N_22268,N_22003);
and U22996 (N_22996,N_20218,N_22017);
and U22997 (N_22997,N_22066,N_22163);
or U22998 (N_22998,N_21556,N_21862);
and U22999 (N_22999,N_21109,N_22183);
or U23000 (N_23000,N_20236,N_21788);
and U23001 (N_23001,N_21464,N_20559);
nor U23002 (N_23002,N_21947,N_21312);
and U23003 (N_23003,N_20300,N_20415);
nor U23004 (N_23004,N_20068,N_20012);
or U23005 (N_23005,N_22324,N_21484);
and U23006 (N_23006,N_22160,N_20673);
or U23007 (N_23007,N_21445,N_22155);
and U23008 (N_23008,N_22244,N_21176);
nor U23009 (N_23009,N_21452,N_22154);
nand U23010 (N_23010,N_20231,N_20867);
or U23011 (N_23011,N_21172,N_21458);
xor U23012 (N_23012,N_22118,N_22075);
or U23013 (N_23013,N_20102,N_20529);
nand U23014 (N_23014,N_20587,N_20189);
nor U23015 (N_23015,N_20844,N_22325);
nor U23016 (N_23016,N_20180,N_21516);
xor U23017 (N_23017,N_21200,N_20124);
nor U23018 (N_23018,N_21417,N_21471);
nand U23019 (N_23019,N_20075,N_21778);
xnor U23020 (N_23020,N_20063,N_21955);
and U23021 (N_23021,N_22224,N_21785);
and U23022 (N_23022,N_22223,N_22060);
nor U23023 (N_23023,N_20817,N_20637);
xor U23024 (N_23024,N_20998,N_21067);
or U23025 (N_23025,N_21514,N_21533);
xnor U23026 (N_23026,N_20578,N_20682);
and U23027 (N_23027,N_21910,N_21991);
nand U23028 (N_23028,N_21942,N_21669);
xnor U23029 (N_23029,N_22135,N_20583);
and U23030 (N_23030,N_20021,N_22458);
nand U23031 (N_23031,N_21532,N_21103);
nor U23032 (N_23032,N_22272,N_21029);
or U23033 (N_23033,N_21671,N_20899);
xnor U23034 (N_23034,N_21517,N_20675);
or U23035 (N_23035,N_22148,N_21052);
nand U23036 (N_23036,N_21952,N_20377);
xnor U23037 (N_23037,N_20381,N_21285);
xor U23038 (N_23038,N_21742,N_20994);
and U23039 (N_23039,N_22112,N_20306);
xor U23040 (N_23040,N_22424,N_21050);
xor U23041 (N_23041,N_21000,N_22127);
nand U23042 (N_23042,N_20542,N_22006);
or U23043 (N_23043,N_22284,N_21468);
nor U23044 (N_23044,N_20237,N_21817);
nor U23045 (N_23045,N_22303,N_20192);
nand U23046 (N_23046,N_22214,N_20140);
or U23047 (N_23047,N_22092,N_20389);
nor U23048 (N_23048,N_20011,N_22400);
nor U23049 (N_23049,N_20139,N_20153);
xnor U23050 (N_23050,N_22426,N_20770);
nand U23051 (N_23051,N_21563,N_22225);
xor U23052 (N_23052,N_22443,N_21723);
nor U23053 (N_23053,N_21007,N_21885);
or U23054 (N_23054,N_21927,N_20623);
xor U23055 (N_23055,N_21022,N_21113);
nand U23056 (N_23056,N_22085,N_20794);
nand U23057 (N_23057,N_21679,N_21670);
or U23058 (N_23058,N_21753,N_20123);
nor U23059 (N_23059,N_21638,N_20607);
nor U23060 (N_23060,N_21142,N_21961);
or U23061 (N_23061,N_20447,N_21724);
and U23062 (N_23062,N_20326,N_20397);
and U23063 (N_23063,N_20636,N_21005);
xnor U23064 (N_23064,N_20331,N_21787);
xor U23065 (N_23065,N_22171,N_21333);
or U23066 (N_23066,N_20316,N_22083);
and U23067 (N_23067,N_22269,N_21250);
xnor U23068 (N_23068,N_22422,N_22110);
nor U23069 (N_23069,N_21433,N_21990);
and U23070 (N_23070,N_20969,N_21359);
nand U23071 (N_23071,N_20428,N_22026);
nor U23072 (N_23072,N_20782,N_21734);
nand U23073 (N_23073,N_22128,N_20702);
nor U23074 (N_23074,N_21217,N_20297);
and U23075 (N_23075,N_21678,N_22203);
nor U23076 (N_23076,N_21453,N_20461);
xnor U23077 (N_23077,N_20748,N_20010);
and U23078 (N_23078,N_21766,N_20906);
nor U23079 (N_23079,N_20919,N_20217);
xnor U23080 (N_23080,N_21973,N_20901);
or U23081 (N_23081,N_21729,N_22103);
or U23082 (N_23082,N_21959,N_22402);
nand U23083 (N_23083,N_20197,N_21617);
and U23084 (N_23084,N_20229,N_21249);
nand U23085 (N_23085,N_22059,N_20825);
nand U23086 (N_23086,N_21451,N_21104);
and U23087 (N_23087,N_21013,N_22142);
nor U23088 (N_23088,N_20379,N_22056);
nor U23089 (N_23089,N_21203,N_20730);
or U23090 (N_23090,N_21856,N_21017);
and U23091 (N_23091,N_20055,N_20097);
nand U23092 (N_23092,N_21018,N_20773);
and U23093 (N_23093,N_20684,N_21621);
nand U23094 (N_23094,N_20616,N_22456);
nand U23095 (N_23095,N_21929,N_20262);
or U23096 (N_23096,N_21511,N_22018);
and U23097 (N_23097,N_20111,N_22068);
and U23098 (N_23098,N_21223,N_21278);
or U23099 (N_23099,N_21769,N_21904);
xnor U23100 (N_23100,N_20105,N_22367);
and U23101 (N_23101,N_20923,N_20666);
and U23102 (N_23102,N_20837,N_21593);
and U23103 (N_23103,N_22093,N_20194);
nand U23104 (N_23104,N_21068,N_20184);
nand U23105 (N_23105,N_21587,N_21486);
xor U23106 (N_23106,N_21989,N_21461);
and U23107 (N_23107,N_21380,N_21878);
or U23108 (N_23108,N_21668,N_22455);
or U23109 (N_23109,N_21972,N_21941);
nand U23110 (N_23110,N_21652,N_20416);
nand U23111 (N_23111,N_20215,N_21665);
nor U23112 (N_23112,N_22168,N_20456);
nand U23113 (N_23113,N_21881,N_21794);
or U23114 (N_23114,N_20030,N_21595);
xor U23115 (N_23115,N_20688,N_20679);
and U23116 (N_23116,N_20927,N_20440);
nand U23117 (N_23117,N_22295,N_21765);
nor U23118 (N_23118,N_21521,N_21378);
xor U23119 (N_23119,N_20581,N_22009);
xnor U23120 (N_23120,N_20697,N_20469);
nand U23121 (N_23121,N_22498,N_21160);
nor U23122 (N_23122,N_20350,N_22307);
nand U23123 (N_23123,N_20753,N_21508);
and U23124 (N_23124,N_21031,N_21492);
xnor U23125 (N_23125,N_21816,N_20319);
or U23126 (N_23126,N_21136,N_21126);
xor U23127 (N_23127,N_22348,N_22181);
or U23128 (N_23128,N_20633,N_21506);
xnor U23129 (N_23129,N_20033,N_20212);
nor U23130 (N_23130,N_20318,N_20483);
xnor U23131 (N_23131,N_21440,N_22473);
nand U23132 (N_23132,N_21489,N_21355);
nand U23133 (N_23133,N_21899,N_20971);
nand U23134 (N_23134,N_22090,N_20423);
xor U23135 (N_23135,N_22042,N_20385);
nand U23136 (N_23136,N_22159,N_20645);
and U23137 (N_23137,N_21915,N_21798);
xor U23138 (N_23138,N_20929,N_22273);
nor U23139 (N_23139,N_20115,N_20626);
xor U23140 (N_23140,N_22213,N_22212);
nor U23141 (N_23141,N_22178,N_22465);
or U23142 (N_23142,N_20795,N_21618);
nor U23143 (N_23143,N_20554,N_22099);
nand U23144 (N_23144,N_20896,N_20701);
and U23145 (N_23145,N_20468,N_20196);
and U23146 (N_23146,N_20726,N_21163);
nor U23147 (N_23147,N_22283,N_21762);
or U23148 (N_23148,N_20006,N_21345);
and U23149 (N_23149,N_22187,N_22468);
or U23150 (N_23150,N_21350,N_21702);
and U23151 (N_23151,N_21736,N_20201);
nand U23152 (N_23152,N_21792,N_22071);
nand U23153 (N_23153,N_20849,N_21505);
and U23154 (N_23154,N_21870,N_21341);
and U23155 (N_23155,N_21879,N_21726);
nor U23156 (N_23156,N_21493,N_20050);
xor U23157 (N_23157,N_21328,N_22156);
and U23158 (N_23158,N_21779,N_21309);
xor U23159 (N_23159,N_22378,N_21956);
xnor U23160 (N_23160,N_20467,N_20517);
nor U23161 (N_23161,N_20224,N_21079);
nor U23162 (N_23162,N_22206,N_21549);
and U23163 (N_23163,N_22209,N_20577);
nand U23164 (N_23164,N_20378,N_20888);
and U23165 (N_23165,N_22078,N_22395);
and U23166 (N_23166,N_20922,N_20295);
or U23167 (N_23167,N_20401,N_21042);
or U23168 (N_23168,N_22480,N_20444);
nand U23169 (N_23169,N_22270,N_22470);
and U23170 (N_23170,N_20875,N_22374);
or U23171 (N_23171,N_21431,N_22196);
and U23172 (N_23172,N_21215,N_20549);
nand U23173 (N_23173,N_21821,N_20913);
and U23174 (N_23174,N_20984,N_20299);
or U23175 (N_23175,N_20592,N_20375);
nor U23176 (N_23176,N_20349,N_22484);
or U23177 (N_23177,N_21194,N_21777);
nand U23178 (N_23178,N_20354,N_20706);
xor U23179 (N_23179,N_20653,N_20449);
and U23180 (N_23180,N_20070,N_22179);
nor U23181 (N_23181,N_22302,N_20885);
nand U23182 (N_23182,N_21036,N_20092);
xor U23183 (N_23183,N_21290,N_20887);
or U23184 (N_23184,N_20649,N_22105);
nor U23185 (N_23185,N_22314,N_22208);
xor U23186 (N_23186,N_20387,N_22167);
and U23187 (N_23187,N_21676,N_21544);
or U23188 (N_23188,N_21329,N_22412);
and U23189 (N_23189,N_21664,N_20786);
nor U23190 (N_23190,N_22437,N_20213);
or U23191 (N_23191,N_21809,N_21148);
or U23192 (N_23192,N_20692,N_22282);
nor U23193 (N_23193,N_21903,N_22486);
or U23194 (N_23194,N_21275,N_20489);
and U23195 (N_23195,N_20129,N_20443);
xnor U23196 (N_23196,N_21623,N_21336);
and U23197 (N_23197,N_22334,N_20780);
or U23198 (N_23198,N_22076,N_21098);
or U23199 (N_23199,N_20370,N_21997);
xor U23200 (N_23200,N_22230,N_21168);
or U23201 (N_23201,N_22124,N_21660);
or U23202 (N_23202,N_21209,N_21588);
and U23203 (N_23203,N_20362,N_20805);
nand U23204 (N_23204,N_21149,N_20094);
nor U23205 (N_23205,N_20777,N_20061);
nand U23206 (N_23206,N_21647,N_22097);
nand U23207 (N_23207,N_21755,N_22316);
nor U23208 (N_23208,N_21072,N_20287);
xor U23209 (N_23209,N_21643,N_21334);
nand U23210 (N_23210,N_20840,N_21078);
nand U23211 (N_23211,N_21692,N_22355);
and U23212 (N_23212,N_21351,N_20277);
nor U23213 (N_23213,N_20232,N_20380);
xnor U23214 (N_23214,N_22265,N_20219);
and U23215 (N_23215,N_20724,N_21868);
nor U23216 (N_23216,N_21173,N_21317);
nor U23217 (N_23217,N_21376,N_21719);
or U23218 (N_23218,N_21980,N_21754);
or U23219 (N_23219,N_20031,N_21795);
xnor U23220 (N_23220,N_20799,N_20051);
and U23221 (N_23221,N_21441,N_21070);
nand U23222 (N_23222,N_21362,N_20290);
nand U23223 (N_23223,N_20627,N_20259);
xnor U23224 (N_23224,N_21319,N_22233);
nor U23225 (N_23225,N_22418,N_20573);
or U23226 (N_23226,N_20925,N_20089);
nand U23227 (N_23227,N_20054,N_20425);
and U23228 (N_23228,N_20555,N_21469);
and U23229 (N_23229,N_21305,N_20690);
and U23230 (N_23230,N_21045,N_21398);
nand U23231 (N_23231,N_20285,N_22087);
nor U23232 (N_23232,N_21886,N_22344);
and U23233 (N_23233,N_20710,N_21155);
nor U23234 (N_23234,N_22262,N_20725);
nand U23235 (N_23235,N_21030,N_21239);
nand U23236 (N_23236,N_20266,N_20846);
nand U23237 (N_23237,N_21261,N_21944);
nor U23238 (N_23238,N_21472,N_20677);
and U23239 (N_23239,N_20834,N_21244);
nor U23240 (N_23240,N_21654,N_22204);
or U23241 (N_23241,N_22025,N_21140);
nor U23242 (N_23242,N_21102,N_22116);
nor U23243 (N_23243,N_22388,N_21835);
or U23244 (N_23244,N_20847,N_20879);
nor U23245 (N_23245,N_22394,N_21920);
xor U23246 (N_23246,N_20152,N_22274);
or U23247 (N_23247,N_20337,N_21012);
or U23248 (N_23248,N_21612,N_22073);
and U23249 (N_23249,N_20169,N_20515);
nand U23250 (N_23250,N_20172,N_20876);
and U23251 (N_23251,N_20371,N_20141);
and U23252 (N_23252,N_20422,N_21507);
nand U23253 (N_23253,N_21954,N_20038);
or U23254 (N_23254,N_21640,N_22425);
or U23255 (N_23255,N_21488,N_20813);
or U23256 (N_23256,N_21625,N_22086);
nor U23257 (N_23257,N_20303,N_22190);
and U23258 (N_23258,N_20751,N_21202);
nor U23259 (N_23259,N_20722,N_22052);
and U23260 (N_23260,N_22428,N_21943);
nand U23261 (N_23261,N_20505,N_21003);
or U23262 (N_23262,N_20032,N_22024);
and U23263 (N_23263,N_21525,N_20644);
or U23264 (N_23264,N_20222,N_20074);
xor U23265 (N_23265,N_22088,N_22231);
xor U23266 (N_23266,N_20508,N_20883);
or U23267 (N_23267,N_21174,N_20732);
or U23268 (N_23268,N_20902,N_22413);
nor U23269 (N_23269,N_21979,N_20163);
or U23270 (N_23270,N_22173,N_20866);
or U23271 (N_23271,N_21276,N_21712);
or U23272 (N_23272,N_21594,N_22328);
nor U23273 (N_23273,N_21207,N_20327);
or U23274 (N_23274,N_20926,N_20276);
nor U23275 (N_23275,N_20862,N_21727);
nand U23276 (N_23276,N_20035,N_21685);
xor U23277 (N_23277,N_20539,N_22144);
or U23278 (N_23278,N_20646,N_22381);
xor U23279 (N_23279,N_21274,N_21167);
nor U23280 (N_23280,N_21577,N_21914);
and U23281 (N_23281,N_22385,N_22253);
or U23282 (N_23282,N_20509,N_21487);
or U23283 (N_23283,N_22219,N_22398);
nor U23284 (N_23284,N_20025,N_21193);
nand U23285 (N_23285,N_21382,N_21227);
nor U23286 (N_23286,N_20982,N_21583);
xnor U23287 (N_23287,N_21175,N_21526);
or U23288 (N_23288,N_21219,N_20272);
nor U23289 (N_23289,N_21722,N_20238);
and U23290 (N_23290,N_20890,N_22007);
xnor U23291 (N_23291,N_20721,N_20526);
or U23292 (N_23292,N_22082,N_20669);
and U23293 (N_23293,N_20945,N_20686);
nand U23294 (N_23294,N_20566,N_22288);
xnor U23295 (N_23295,N_20920,N_21348);
and U23296 (N_23296,N_21419,N_21429);
nand U23297 (N_23297,N_22499,N_22476);
nor U23298 (N_23298,N_21465,N_20419);
and U23299 (N_23299,N_21775,N_22464);
nand U23300 (N_23300,N_21190,N_21095);
nor U23301 (N_23301,N_21111,N_22399);
and U23302 (N_23302,N_21921,N_20451);
xor U23303 (N_23303,N_22170,N_20597);
nand U23304 (N_23304,N_22349,N_22109);
and U23305 (N_23305,N_21354,N_20672);
or U23306 (N_23306,N_20133,N_21572);
and U23307 (N_23307,N_21358,N_22123);
or U23308 (N_23308,N_22454,N_21645);
nor U23309 (N_23309,N_22386,N_20952);
or U23310 (N_23310,N_20263,N_22207);
nand U23311 (N_23311,N_20754,N_21066);
xnor U23312 (N_23312,N_21143,N_21043);
and U23313 (N_23313,N_22130,N_21804);
nand U23314 (N_23314,N_21490,N_21454);
and U23315 (N_23315,N_20551,N_20760);
nand U23316 (N_23316,N_20039,N_20095);
and U23317 (N_23317,N_21268,N_20460);
or U23318 (N_23318,N_21396,N_20694);
nand U23319 (N_23319,N_20580,N_20230);
and U23320 (N_23320,N_20595,N_22301);
nand U23321 (N_23321,N_21057,N_21590);
or U23322 (N_23322,N_20761,N_21447);
nor U23323 (N_23323,N_21900,N_22058);
xnor U23324 (N_23324,N_21238,N_21784);
nand U23325 (N_23325,N_22152,N_21002);
xor U23326 (N_23326,N_20225,N_21243);
and U23327 (N_23327,N_21121,N_22343);
xor U23328 (N_23328,N_20914,N_21738);
or U23329 (N_23329,N_20804,N_20488);
or U23330 (N_23330,N_21697,N_20608);
nor U23331 (N_23331,N_21849,N_21495);
nor U23332 (N_23332,N_20490,N_20473);
nor U23333 (N_23333,N_20314,N_22240);
nor U23334 (N_23334,N_21107,N_22074);
and U23335 (N_23335,N_21682,N_21135);
and U23336 (N_23336,N_22446,N_21366);
nand U23337 (N_23337,N_20598,N_20453);
xnor U23338 (N_23338,N_22461,N_20309);
and U23339 (N_23339,N_22323,N_22372);
or U23340 (N_23340,N_22250,N_20689);
or U23341 (N_23341,N_22392,N_20479);
xnor U23342 (N_23342,N_21520,N_22249);
or U23343 (N_23343,N_21585,N_21124);
xor U23344 (N_23344,N_21918,N_21936);
nor U23345 (N_23345,N_20900,N_20793);
xor U23346 (N_23346,N_21836,N_21009);
xnor U23347 (N_23347,N_21789,N_21930);
nand U23348 (N_23348,N_20147,N_20128);
or U23349 (N_23349,N_20474,N_20036);
xor U23350 (N_23350,N_22027,N_20811);
nor U23351 (N_23351,N_21014,N_22293);
and U23352 (N_23352,N_20104,N_21564);
nor U23353 (N_23353,N_22497,N_21803);
or U23354 (N_23354,N_20106,N_22013);
or U23355 (N_23355,N_20241,N_21957);
or U23356 (N_23356,N_22313,N_22185);
nor U23357 (N_23357,N_22492,N_20548);
xnor U23358 (N_23358,N_21808,N_22239);
or U23359 (N_23359,N_21834,N_21760);
nand U23360 (N_23360,N_22227,N_21075);
and U23361 (N_23361,N_21791,N_20513);
xor U23362 (N_23362,N_21620,N_21622);
and U23363 (N_23363,N_21213,N_20364);
nand U23364 (N_23364,N_21028,N_20651);
or U23365 (N_23365,N_20680,N_20893);
xnor U23366 (N_23366,N_22145,N_22366);
xnor U23367 (N_23367,N_20681,N_20402);
or U23368 (N_23368,N_20972,N_20880);
and U23369 (N_23369,N_21782,N_20071);
nand U23370 (N_23370,N_21254,N_22061);
xor U23371 (N_23371,N_20367,N_21653);
nand U23372 (N_23372,N_21552,N_21478);
nor U23373 (N_23373,N_22020,N_20698);
xor U23374 (N_23374,N_20322,N_21089);
xnor U23375 (N_23375,N_20895,N_22423);
or U23376 (N_23376,N_20345,N_22139);
xor U23377 (N_23377,N_21536,N_20855);
nand U23378 (N_23378,N_21710,N_22327);
nor U23379 (N_23379,N_20249,N_20408);
xnor U23380 (N_23380,N_21027,N_21998);
or U23381 (N_23381,N_20344,N_20320);
and U23382 (N_23382,N_21853,N_21925);
nand U23383 (N_23383,N_20563,N_21570);
nand U23384 (N_23384,N_20719,N_20034);
xor U23385 (N_23385,N_20096,N_21199);
and U23386 (N_23386,N_22177,N_20144);
nand U23387 (N_23387,N_21035,N_20839);
xor U23388 (N_23388,N_21158,N_20149);
xor U23389 (N_23389,N_20399,N_21502);
or U23390 (N_23390,N_22242,N_20729);
nor U23391 (N_23391,N_22192,N_20062);
or U23392 (N_23392,N_22010,N_21864);
or U23393 (N_23393,N_20099,N_20118);
nor U23394 (N_23394,N_21895,N_20935);
nor U23395 (N_23395,N_20497,N_20564);
and U23396 (N_23396,N_21248,N_20100);
nand U23397 (N_23397,N_20357,N_22266);
or U23398 (N_23398,N_22081,N_22016);
nand U23399 (N_23399,N_22291,N_20750);
nand U23400 (N_23400,N_21683,N_20481);
or U23401 (N_23401,N_21245,N_22216);
and U23402 (N_23402,N_20177,N_20814);
xor U23403 (N_23403,N_20109,N_20918);
xnor U23404 (N_23404,N_22199,N_21436);
xnor U23405 (N_23405,N_20069,N_21718);
nor U23406 (N_23406,N_20446,N_20863);
xor U23407 (N_23407,N_21494,N_21984);
nor U23408 (N_23408,N_21425,N_20340);
or U23409 (N_23409,N_20987,N_20044);
or U23410 (N_23410,N_20562,N_20687);
nor U23411 (N_23411,N_22289,N_22463);
nor U23412 (N_23412,N_21748,N_21529);
nand U23413 (N_23413,N_21575,N_22460);
nand U23414 (N_23414,N_22221,N_21776);
or U23415 (N_23415,N_21860,N_20045);
or U23416 (N_23416,N_21602,N_21335);
xnor U23417 (N_23417,N_20056,N_20619);
nand U23418 (N_23418,N_21733,N_21898);
xnor U23419 (N_23419,N_21370,N_20916);
nand U23420 (N_23420,N_20629,N_21858);
nand U23421 (N_23421,N_20459,N_21026);
nor U23422 (N_23422,N_21460,N_21626);
and U23423 (N_23423,N_20493,N_20334);
nor U23424 (N_23424,N_21976,N_21582);
and U23425 (N_23425,N_20579,N_21684);
or U23426 (N_23426,N_20373,N_20176);
or U23427 (N_23427,N_21159,N_20117);
nand U23428 (N_23428,N_21831,N_21044);
or U23429 (N_23429,N_20630,N_20146);
nand U23430 (N_23430,N_22143,N_20245);
or U23431 (N_23431,N_21513,N_22067);
nand U23432 (N_23432,N_20264,N_21298);
xnor U23433 (N_23433,N_21297,N_22252);
or U23434 (N_23434,N_21893,N_20223);
xnor U23435 (N_23435,N_21192,N_21802);
and U23436 (N_23436,N_21911,N_20985);
and U23437 (N_23437,N_22290,N_21060);
or U23438 (N_23438,N_21313,N_21266);
or U23439 (N_23439,N_20256,N_21347);
nor U23440 (N_23440,N_21110,N_20845);
nand U23441 (N_23441,N_22237,N_21813);
nand U23442 (N_23442,N_20544,N_21056);
and U23443 (N_23443,N_22406,N_20809);
nand U23444 (N_23444,N_20359,N_22114);
xor U23445 (N_23445,N_21444,N_21299);
xor U23446 (N_23446,N_20575,N_21574);
and U23447 (N_23447,N_21224,N_22416);
and U23448 (N_23448,N_22079,N_21538);
xnor U23449 (N_23449,N_20785,N_20410);
nand U23450 (N_23450,N_20963,N_20369);
and U23451 (N_23451,N_20424,N_20273);
xnor U23452 (N_23452,N_21974,N_20768);
or U23453 (N_23453,N_21982,N_21770);
nand U23454 (N_23454,N_20009,N_21889);
nand U23455 (N_23455,N_20807,N_21264);
xor U23456 (N_23456,N_22030,N_21790);
nor U23457 (N_23457,N_20716,N_21540);
nand U23458 (N_23458,N_20781,N_21597);
nand U23459 (N_23459,N_20628,N_22038);
and U23460 (N_23460,N_20078,N_22442);
or U23461 (N_23461,N_20924,N_22184);
and U23462 (N_23462,N_21352,N_21938);
nor U23463 (N_23463,N_20274,N_21700);
nor U23464 (N_23464,N_20311,N_21740);
nand U23465 (N_23465,N_20268,N_22474);
xnor U23466 (N_23466,N_20214,N_21663);
or U23467 (N_23467,N_22471,N_20433);
and U23468 (N_23468,N_21255,N_21321);
nor U23469 (N_23469,N_21631,N_21485);
nor U23470 (N_23470,N_21412,N_22043);
xnor U23471 (N_23471,N_20524,N_21951);
nor U23472 (N_23472,N_20368,N_20248);
nand U23473 (N_23473,N_21381,N_20065);
or U23474 (N_23474,N_20329,N_21093);
nor U23475 (N_23475,N_21099,N_20639);
nand U23476 (N_23476,N_20158,N_20660);
or U23477 (N_23477,N_22245,N_22070);
or U23478 (N_23478,N_21966,N_20930);
or U23479 (N_23479,N_21512,N_21286);
nand U23480 (N_23480,N_22444,N_21434);
or U23481 (N_23481,N_20823,N_21151);
nor U23482 (N_23482,N_20475,N_21872);
or U23483 (N_23483,N_20017,N_22033);
nand U23484 (N_23484,N_20842,N_20540);
nor U23485 (N_23485,N_20313,N_22186);
nor U23486 (N_23486,N_20791,N_20997);
or U23487 (N_23487,N_22434,N_21191);
nand U23488 (N_23488,N_21443,N_22174);
nand U23489 (N_23489,N_22182,N_22332);
and U23490 (N_23490,N_21084,N_20812);
or U23491 (N_23491,N_20404,N_20712);
xor U23492 (N_23492,N_21229,N_20138);
nand U23493 (N_23493,N_22310,N_21476);
nand U23494 (N_23494,N_20185,N_21598);
xor U23495 (N_23495,N_21783,N_21291);
xnor U23496 (N_23496,N_21773,N_21372);
and U23497 (N_23497,N_21824,N_21578);
xor U23498 (N_23498,N_21218,N_21051);
nand U23499 (N_23499,N_21144,N_22021);
nor U23500 (N_23500,N_21832,N_20763);
nand U23501 (N_23501,N_20283,N_22263);
nand U23502 (N_23502,N_20872,N_20999);
xnor U23503 (N_23503,N_20755,N_21480);
xor U23504 (N_23504,N_20499,N_22131);
and U23505 (N_23505,N_20173,N_20426);
nor U23506 (N_23506,N_21839,N_21301);
or U23507 (N_23507,N_21815,N_22493);
or U23508 (N_23508,N_21524,N_21604);
or U23509 (N_23509,N_20821,N_20484);
and U23510 (N_23510,N_21639,N_20944);
xnor U23511 (N_23511,N_21518,N_20962);
nor U23512 (N_23512,N_20437,N_22368);
or U23513 (N_23513,N_21346,N_22055);
nor U23514 (N_23514,N_20703,N_20762);
nor U23515 (N_23515,N_21253,N_21793);
xnor U23516 (N_23516,N_21940,N_22396);
nor U23517 (N_23517,N_22146,N_21874);
and U23518 (N_23518,N_22158,N_21482);
nor U23519 (N_23519,N_20808,N_20293);
and U23520 (N_23520,N_21497,N_20202);
xor U23521 (N_23521,N_22317,N_20625);
and U23522 (N_23522,N_20975,N_20077);
and U23523 (N_23523,N_21221,N_22037);
or U23524 (N_23524,N_21950,N_20815);
xor U23525 (N_23525,N_22419,N_21304);
and U23526 (N_23526,N_20769,N_21015);
or U23527 (N_23527,N_20333,N_21656);
or U23528 (N_23528,N_21256,N_22452);
xnor U23529 (N_23529,N_22481,N_21091);
xnor U23530 (N_23530,N_21866,N_22330);
nand U23531 (N_23531,N_21693,N_20611);
nand U23532 (N_23532,N_22287,N_20048);
nand U23533 (N_23533,N_21615,N_21402);
or U23534 (N_23534,N_22298,N_20434);
or U23535 (N_23535,N_21323,N_20894);
nor U23536 (N_23536,N_21786,N_20909);
and U23537 (N_23537,N_21288,N_20741);
nor U23538 (N_23538,N_21141,N_21781);
xnor U23539 (N_23539,N_20160,N_20355);
nand U23540 (N_23540,N_21988,N_20937);
or U23541 (N_23541,N_21761,N_21554);
nor U23542 (N_23542,N_20700,N_21059);
and U23543 (N_23543,N_21548,N_21546);
or U23544 (N_23544,N_21716,N_22319);
nor U23545 (N_23545,N_21539,N_20604);
or U23546 (N_23546,N_21279,N_20131);
nor U23547 (N_23547,N_20351,N_22046);
and U23548 (N_23548,N_21178,N_20210);
and U23549 (N_23549,N_21624,N_20007);
and U23550 (N_23550,N_20656,N_20736);
or U23551 (N_23551,N_20707,N_22491);
or U23552 (N_23552,N_21314,N_22054);
xor U23553 (N_23553,N_20889,N_20247);
or U23554 (N_23554,N_22445,N_20341);
nand U23555 (N_23555,N_21392,N_21206);
nand U23556 (N_23556,N_21085,N_21422);
and U23557 (N_23557,N_21764,N_22220);
nor U23558 (N_23558,N_20269,N_20606);
or U23559 (N_23559,N_21129,N_20933);
and U23560 (N_23560,N_20108,N_22489);
or U23561 (N_23561,N_20107,N_20534);
or U23562 (N_23562,N_20806,N_22363);
or U23563 (N_23563,N_21001,N_20819);
nor U23564 (N_23564,N_22318,N_20470);
nand U23565 (N_23565,N_20800,N_20612);
nand U23566 (N_23566,N_22297,N_20304);
xor U23567 (N_23567,N_21230,N_21756);
xor U23568 (N_23568,N_22414,N_21236);
nand U23569 (N_23569,N_21273,N_21058);
xor U23570 (N_23570,N_22494,N_20832);
nand U23571 (N_23571,N_20708,N_22382);
and U23572 (N_23572,N_22339,N_20052);
and U23573 (N_23573,N_21232,N_22279);
xnor U23574 (N_23574,N_20244,N_21732);
nor U23575 (N_23575,N_20376,N_22107);
and U23576 (N_23576,N_20388,N_20543);
nand U23577 (N_23577,N_22228,N_20864);
and U23578 (N_23578,N_21897,N_20155);
or U23579 (N_23579,N_20445,N_21949);
or U23580 (N_23580,N_21282,N_20853);
or U23581 (N_23581,N_21491,N_21730);
xor U23582 (N_23582,N_21470,N_20037);
nor U23583 (N_23583,N_20435,N_20091);
nor U23584 (N_23584,N_22326,N_21166);
or U23585 (N_23585,N_20235,N_20856);
nand U23586 (N_23586,N_22296,N_20940);
nor U23587 (N_23587,N_22376,N_20315);
and U23588 (N_23588,N_20816,N_21558);
and U23589 (N_23589,N_21049,N_20910);
xor U23590 (N_23590,N_21247,N_21933);
or U23591 (N_23591,N_20347,N_22036);
or U23592 (N_23592,N_20495,N_21844);
nor U23593 (N_23593,N_21128,N_20430);
or U23594 (N_23594,N_20570,N_21937);
xnor U23595 (N_23595,N_20120,N_21164);
xnor U23596 (N_23596,N_20874,N_22232);
nand U23597 (N_23597,N_20478,N_21394);
or U23598 (N_23598,N_20343,N_21210);
or U23599 (N_23599,N_20405,N_21237);
nor U23600 (N_23600,N_20718,N_20711);
xor U23601 (N_23601,N_22008,N_21616);
nor U23602 (N_23602,N_20833,N_20057);
xor U23603 (N_23603,N_20136,N_22431);
and U23604 (N_23604,N_21404,N_21138);
xor U23605 (N_23605,N_21271,N_22035);
nand U23606 (N_23606,N_20492,N_21983);
and U23607 (N_23607,N_20116,N_20015);
nand U23608 (N_23608,N_21523,N_21399);
or U23609 (N_23609,N_21850,N_20452);
xor U23610 (N_23610,N_21325,N_21568);
xnor U23611 (N_23611,N_22121,N_21277);
nor U23612 (N_23612,N_21747,N_21008);
and U23613 (N_23613,N_20203,N_22102);
xor U23614 (N_23614,N_20958,N_21457);
nor U23615 (N_23615,N_22243,N_20465);
or U23616 (N_23616,N_21216,N_22404);
nor U23617 (N_23617,N_22089,N_22153);
or U23618 (N_23618,N_20561,N_22448);
or U23619 (N_23619,N_20418,N_20114);
xnor U23620 (N_23620,N_20255,N_22345);
nor U23621 (N_23621,N_22350,N_20528);
and U23622 (N_23622,N_21101,N_20407);
xor U23623 (N_23623,N_20955,N_22390);
nand U23624 (N_23624,N_20503,N_21757);
xnor U23625 (N_23625,N_22354,N_22201);
or U23626 (N_23626,N_20527,N_22427);
and U23627 (N_23627,N_21306,N_21906);
or U23628 (N_23628,N_20676,N_21634);
nor U23629 (N_23629,N_20531,N_20642);
and U23630 (N_23630,N_20948,N_20412);
nand U23631 (N_23631,N_21812,N_22305);
xnor U23632 (N_23632,N_20199,N_21841);
nor U23633 (N_23633,N_21033,N_20029);
or U23634 (N_23634,N_22211,N_22439);
or U23635 (N_23635,N_21551,N_20020);
xnor U23636 (N_23636,N_22482,N_22411);
nand U23637 (N_23637,N_20398,N_21763);
and U23638 (N_23638,N_21592,N_21349);
nor U23639 (N_23639,N_20588,N_22440);
and U23640 (N_23640,N_21442,N_21611);
xor U23641 (N_23641,N_21196,N_21562);
nor U23642 (N_23642,N_21644,N_20356);
xnor U23643 (N_23643,N_20338,N_20150);
nand U23644 (N_23644,N_21962,N_20084);
and U23645 (N_23645,N_21745,N_21339);
or U23646 (N_23646,N_21127,N_21519);
nand U23647 (N_23647,N_21543,N_21233);
and U23648 (N_23648,N_22028,N_21046);
nand U23649 (N_23649,N_21123,N_22147);
xor U23650 (N_23650,N_20506,N_21415);
nor U23651 (N_23651,N_20824,N_20658);
nand U23652 (N_23652,N_20286,N_20254);
nand U23653 (N_23653,N_20957,N_21108);
nand U23654 (N_23654,N_22364,N_20145);
and U23655 (N_23655,N_21448,N_21737);
and U23656 (N_23656,N_20691,N_20615);
xor U23657 (N_23657,N_22479,N_21565);
or U23658 (N_23658,N_20657,N_20822);
nor U23659 (N_23659,N_20396,N_21705);
nand U23660 (N_23660,N_22369,N_20841);
nor U23661 (N_23661,N_20023,N_22023);
or U23662 (N_23662,N_22222,N_22210);
xor U23663 (N_23663,N_21114,N_21185);
nor U23664 (N_23664,N_21629,N_22312);
or U23665 (N_23665,N_21659,N_20482);
nor U23666 (N_23666,N_22053,N_22002);
nand U23667 (N_23667,N_22191,N_20246);
and U23668 (N_23668,N_20053,N_20258);
and U23669 (N_23669,N_21703,N_22311);
and U23670 (N_23670,N_20365,N_21681);
nor U23671 (N_23671,N_21406,N_21147);
xor U23672 (N_23672,N_21601,N_21388);
nand U23673 (N_23673,N_20516,N_20400);
or U23674 (N_23674,N_21375,N_20463);
nand U23675 (N_23675,N_21509,N_21965);
and U23676 (N_23676,N_20993,N_22101);
xor U23677 (N_23677,N_22280,N_20974);
nand U23678 (N_23678,N_20911,N_20764);
xnor U23679 (N_23679,N_22405,N_21371);
nand U23680 (N_23680,N_21642,N_21749);
xor U23681 (N_23681,N_21589,N_21344);
xnor U23682 (N_23682,N_20154,N_21269);
and U23683 (N_23683,N_20968,N_20857);
xnor U23684 (N_23684,N_22051,N_21212);
nand U23685 (N_23685,N_20047,N_20159);
or U23686 (N_23686,N_22161,N_22336);
and U23687 (N_23687,N_22100,N_20487);
or U23688 (N_23688,N_20858,N_21561);
nand U23689 (N_23689,N_20882,N_21439);
nor U23690 (N_23690,N_21270,N_21171);
or U23691 (N_23691,N_20271,N_21690);
xnor U23692 (N_23692,N_20339,N_21694);
nand U23693 (N_23693,N_21322,N_21466);
and U23694 (N_23694,N_21801,N_20668);
nor U23695 (N_23695,N_21674,N_22080);
nand U23696 (N_23696,N_20510,N_20752);
or U23697 (N_23697,N_20965,N_21258);
nor U23698 (N_23698,N_21970,N_21999);
or U23699 (N_23699,N_20162,N_21871);
or U23700 (N_23700,N_20560,N_22467);
and U23701 (N_23701,N_20002,N_22095);
and U23702 (N_23702,N_21120,N_20737);
nand U23703 (N_23703,N_20353,N_20621);
and U23704 (N_23704,N_21019,N_20774);
xor U23705 (N_23705,N_21896,N_20087);
xnor U23706 (N_23706,N_22466,N_21838);
nand U23707 (N_23707,N_21283,N_21184);
nand U23708 (N_23708,N_20496,N_20830);
nor U23709 (N_23709,N_22077,N_22106);
or U23710 (N_23710,N_22373,N_21456);
nor U23711 (N_23711,N_22001,N_21475);
xor U23712 (N_23712,N_21420,N_21134);
xor U23713 (N_23713,N_21971,N_21571);
nand U23714 (N_23714,N_20361,N_21145);
nand U23715 (N_23715,N_21088,N_21865);
and U23716 (N_23716,N_22259,N_22260);
nand U23717 (N_23717,N_21240,N_21024);
xor U23718 (N_23718,N_22169,N_21880);
or U23719 (N_23719,N_20382,N_20498);
or U23720 (N_23720,N_20043,N_20798);
and U23721 (N_23721,N_20004,N_21090);
and U23722 (N_23722,N_21696,N_22331);
nand U23723 (N_23723,N_21531,N_21995);
nand U23724 (N_23724,N_20989,N_21708);
nor U23725 (N_23725,N_20556,N_21919);
xor U23726 (N_23726,N_22346,N_21628);
xor U23727 (N_23727,N_20530,N_21823);
nor U23728 (N_23728,N_20640,N_20080);
and U23729 (N_23729,N_22462,N_20744);
nand U23730 (N_23730,N_21924,N_21501);
xnor U23731 (N_23731,N_21438,N_20507);
or U23732 (N_23732,N_20956,N_21913);
or U23733 (N_23733,N_20042,N_20101);
and U23734 (N_23734,N_20605,N_21633);
nand U23735 (N_23735,N_21462,N_20018);
or U23736 (N_23736,N_22117,N_21071);
or U23737 (N_23737,N_20085,N_22409);
nand U23738 (N_23738,N_21037,N_21828);
xor U23739 (N_23739,N_21062,N_22134);
xor U23740 (N_23740,N_22360,N_20296);
nor U23741 (N_23741,N_22417,N_20582);
nor U23742 (N_23742,N_22247,N_20110);
nor U23743 (N_23743,N_20898,N_20251);
nor U23744 (N_23744,N_20747,N_20438);
and U23745 (N_23745,N_21251,N_20383);
and U23746 (N_23746,N_21437,N_21327);
nand U23747 (N_23747,N_20873,N_21796);
and U23748 (N_23748,N_20742,N_20572);
nor U23749 (N_23749,N_20738,N_22459);
xnor U23750 (N_23750,N_21180,N_20957);
or U23751 (N_23751,N_21319,N_20665);
or U23752 (N_23752,N_21229,N_20055);
nor U23753 (N_23753,N_20896,N_20210);
nor U23754 (N_23754,N_20658,N_21590);
nand U23755 (N_23755,N_20292,N_20937);
nand U23756 (N_23756,N_20037,N_21438);
xnor U23757 (N_23757,N_21636,N_20760);
and U23758 (N_23758,N_22038,N_21707);
and U23759 (N_23759,N_21381,N_22010);
or U23760 (N_23760,N_20525,N_21871);
and U23761 (N_23761,N_20103,N_22041);
xor U23762 (N_23762,N_20479,N_20875);
or U23763 (N_23763,N_21069,N_22074);
xnor U23764 (N_23764,N_22335,N_21232);
nor U23765 (N_23765,N_21893,N_21264);
or U23766 (N_23766,N_20970,N_21955);
nor U23767 (N_23767,N_20482,N_20641);
nor U23768 (N_23768,N_20368,N_22334);
nand U23769 (N_23769,N_22181,N_21021);
nor U23770 (N_23770,N_21694,N_20048);
and U23771 (N_23771,N_21098,N_20596);
and U23772 (N_23772,N_21256,N_20887);
nor U23773 (N_23773,N_21689,N_21801);
nand U23774 (N_23774,N_22126,N_22193);
nor U23775 (N_23775,N_21975,N_20276);
and U23776 (N_23776,N_21850,N_21766);
and U23777 (N_23777,N_20316,N_20192);
or U23778 (N_23778,N_20458,N_21408);
and U23779 (N_23779,N_22110,N_21363);
xor U23780 (N_23780,N_20044,N_20088);
nor U23781 (N_23781,N_22492,N_22199);
and U23782 (N_23782,N_20128,N_21245);
or U23783 (N_23783,N_21774,N_22246);
nand U23784 (N_23784,N_21496,N_21634);
or U23785 (N_23785,N_20110,N_20321);
nor U23786 (N_23786,N_20223,N_20334);
and U23787 (N_23787,N_21756,N_21540);
xnor U23788 (N_23788,N_20948,N_22470);
or U23789 (N_23789,N_20252,N_20329);
nand U23790 (N_23790,N_21375,N_21091);
and U23791 (N_23791,N_21805,N_21969);
nand U23792 (N_23792,N_21413,N_22299);
and U23793 (N_23793,N_22135,N_20925);
or U23794 (N_23794,N_21436,N_20362);
nand U23795 (N_23795,N_22472,N_21407);
nand U23796 (N_23796,N_21498,N_21983);
nor U23797 (N_23797,N_22456,N_21007);
nor U23798 (N_23798,N_21015,N_20121);
nand U23799 (N_23799,N_21436,N_20976);
xor U23800 (N_23800,N_20288,N_21543);
nor U23801 (N_23801,N_20061,N_20387);
xnor U23802 (N_23802,N_21938,N_22095);
nor U23803 (N_23803,N_20150,N_22497);
nor U23804 (N_23804,N_22498,N_20471);
and U23805 (N_23805,N_21607,N_21281);
and U23806 (N_23806,N_21430,N_21477);
nand U23807 (N_23807,N_20654,N_20837);
and U23808 (N_23808,N_21380,N_21693);
or U23809 (N_23809,N_20826,N_20675);
xor U23810 (N_23810,N_21886,N_20930);
and U23811 (N_23811,N_20305,N_21737);
xnor U23812 (N_23812,N_21229,N_20192);
and U23813 (N_23813,N_21163,N_22287);
nor U23814 (N_23814,N_22370,N_21474);
and U23815 (N_23815,N_20334,N_22154);
and U23816 (N_23816,N_20709,N_22211);
nor U23817 (N_23817,N_20142,N_22195);
nor U23818 (N_23818,N_22204,N_21559);
or U23819 (N_23819,N_21815,N_21557);
and U23820 (N_23820,N_20695,N_21539);
nor U23821 (N_23821,N_21872,N_21762);
xnor U23822 (N_23822,N_22468,N_20845);
xnor U23823 (N_23823,N_20734,N_20310);
and U23824 (N_23824,N_20605,N_21655);
xnor U23825 (N_23825,N_22253,N_20130);
or U23826 (N_23826,N_20146,N_21104);
and U23827 (N_23827,N_21808,N_21044);
xor U23828 (N_23828,N_21708,N_22480);
xor U23829 (N_23829,N_21092,N_20318);
nand U23830 (N_23830,N_22390,N_21749);
xnor U23831 (N_23831,N_22156,N_21605);
nand U23832 (N_23832,N_22126,N_21125);
nor U23833 (N_23833,N_21764,N_20705);
nand U23834 (N_23834,N_22008,N_20000);
or U23835 (N_23835,N_20751,N_21198);
and U23836 (N_23836,N_21900,N_20972);
or U23837 (N_23837,N_20470,N_22075);
or U23838 (N_23838,N_21356,N_21072);
nand U23839 (N_23839,N_20620,N_20138);
nor U23840 (N_23840,N_20623,N_22030);
nand U23841 (N_23841,N_21329,N_21341);
and U23842 (N_23842,N_21564,N_20615);
nand U23843 (N_23843,N_21765,N_21820);
and U23844 (N_23844,N_21744,N_22296);
nand U23845 (N_23845,N_22084,N_21919);
nand U23846 (N_23846,N_21032,N_21841);
nor U23847 (N_23847,N_21305,N_21996);
or U23848 (N_23848,N_21613,N_22223);
xnor U23849 (N_23849,N_20404,N_21433);
or U23850 (N_23850,N_20575,N_21205);
nor U23851 (N_23851,N_21559,N_20350);
and U23852 (N_23852,N_21355,N_20147);
nor U23853 (N_23853,N_20896,N_21100);
nand U23854 (N_23854,N_20828,N_21669);
or U23855 (N_23855,N_20536,N_20248);
and U23856 (N_23856,N_20197,N_20537);
and U23857 (N_23857,N_22040,N_22005);
and U23858 (N_23858,N_22336,N_22196);
nor U23859 (N_23859,N_21698,N_20689);
xor U23860 (N_23860,N_20500,N_20358);
or U23861 (N_23861,N_20264,N_21381);
nor U23862 (N_23862,N_22005,N_21454);
nand U23863 (N_23863,N_22071,N_20406);
nor U23864 (N_23864,N_20999,N_21307);
nand U23865 (N_23865,N_21575,N_21554);
xnor U23866 (N_23866,N_22221,N_20621);
nor U23867 (N_23867,N_21965,N_20439);
xor U23868 (N_23868,N_22377,N_21734);
xnor U23869 (N_23869,N_21322,N_22169);
nor U23870 (N_23870,N_21332,N_21720);
and U23871 (N_23871,N_21672,N_20314);
or U23872 (N_23872,N_21942,N_20629);
xnor U23873 (N_23873,N_21120,N_21173);
xor U23874 (N_23874,N_22272,N_20776);
and U23875 (N_23875,N_21917,N_20263);
xor U23876 (N_23876,N_22296,N_22324);
and U23877 (N_23877,N_21563,N_20416);
nor U23878 (N_23878,N_20547,N_22291);
or U23879 (N_23879,N_20782,N_22179);
and U23880 (N_23880,N_20444,N_20165);
nand U23881 (N_23881,N_20128,N_21777);
nand U23882 (N_23882,N_21100,N_21194);
nand U23883 (N_23883,N_21204,N_22206);
nand U23884 (N_23884,N_21974,N_21317);
or U23885 (N_23885,N_20287,N_20180);
nand U23886 (N_23886,N_22140,N_20513);
and U23887 (N_23887,N_21515,N_22284);
nand U23888 (N_23888,N_22061,N_20017);
nor U23889 (N_23889,N_20865,N_22493);
xnor U23890 (N_23890,N_21869,N_22148);
nand U23891 (N_23891,N_22011,N_20090);
nand U23892 (N_23892,N_21790,N_22028);
and U23893 (N_23893,N_22417,N_20205);
nand U23894 (N_23894,N_21707,N_20835);
and U23895 (N_23895,N_21533,N_22149);
nor U23896 (N_23896,N_21562,N_21081);
nand U23897 (N_23897,N_21974,N_20521);
and U23898 (N_23898,N_22335,N_20774);
and U23899 (N_23899,N_21662,N_20047);
nand U23900 (N_23900,N_21175,N_22310);
nor U23901 (N_23901,N_21043,N_22336);
or U23902 (N_23902,N_21568,N_20877);
or U23903 (N_23903,N_22083,N_22275);
and U23904 (N_23904,N_20667,N_20201);
and U23905 (N_23905,N_21440,N_20736);
or U23906 (N_23906,N_22440,N_21377);
nor U23907 (N_23907,N_20376,N_21232);
nand U23908 (N_23908,N_20853,N_21423);
or U23909 (N_23909,N_21483,N_22365);
nand U23910 (N_23910,N_20629,N_21066);
or U23911 (N_23911,N_21812,N_20185);
or U23912 (N_23912,N_20399,N_22346);
xnor U23913 (N_23913,N_21482,N_20770);
xor U23914 (N_23914,N_20094,N_22243);
nor U23915 (N_23915,N_22361,N_22486);
xnor U23916 (N_23916,N_20035,N_20176);
or U23917 (N_23917,N_21245,N_20702);
or U23918 (N_23918,N_21738,N_21070);
or U23919 (N_23919,N_21747,N_21668);
or U23920 (N_23920,N_21232,N_21718);
xnor U23921 (N_23921,N_22337,N_21478);
or U23922 (N_23922,N_22153,N_22112);
and U23923 (N_23923,N_20367,N_21165);
and U23924 (N_23924,N_22000,N_21060);
nand U23925 (N_23925,N_20863,N_21299);
or U23926 (N_23926,N_22422,N_21566);
nor U23927 (N_23927,N_20289,N_20533);
and U23928 (N_23928,N_21126,N_22495);
xor U23929 (N_23929,N_21916,N_21227);
nor U23930 (N_23930,N_20205,N_21403);
or U23931 (N_23931,N_21163,N_22122);
nand U23932 (N_23932,N_20882,N_21933);
and U23933 (N_23933,N_21023,N_21594);
nand U23934 (N_23934,N_20120,N_20462);
and U23935 (N_23935,N_20153,N_21102);
xnor U23936 (N_23936,N_21630,N_20543);
nor U23937 (N_23937,N_21848,N_21998);
nor U23938 (N_23938,N_21304,N_21023);
nor U23939 (N_23939,N_22464,N_21062);
or U23940 (N_23940,N_20659,N_21549);
nor U23941 (N_23941,N_21507,N_22457);
or U23942 (N_23942,N_22027,N_20501);
nand U23943 (N_23943,N_20287,N_22160);
or U23944 (N_23944,N_20854,N_20456);
nand U23945 (N_23945,N_22161,N_22287);
nand U23946 (N_23946,N_21514,N_21318);
nand U23947 (N_23947,N_21215,N_20870);
nor U23948 (N_23948,N_21628,N_20833);
nor U23949 (N_23949,N_22073,N_22224);
or U23950 (N_23950,N_21344,N_22307);
nand U23951 (N_23951,N_22344,N_22099);
xnor U23952 (N_23952,N_20282,N_21658);
nand U23953 (N_23953,N_22321,N_20182);
nor U23954 (N_23954,N_20327,N_21482);
or U23955 (N_23955,N_20289,N_21366);
or U23956 (N_23956,N_20148,N_20821);
xnor U23957 (N_23957,N_20437,N_20056);
nand U23958 (N_23958,N_20999,N_20688);
nand U23959 (N_23959,N_21822,N_20286);
or U23960 (N_23960,N_22030,N_20381);
or U23961 (N_23961,N_22207,N_20685);
nor U23962 (N_23962,N_21994,N_20801);
or U23963 (N_23963,N_22129,N_22177);
or U23964 (N_23964,N_20932,N_22329);
nor U23965 (N_23965,N_20361,N_21108);
nor U23966 (N_23966,N_22194,N_20135);
nand U23967 (N_23967,N_21746,N_20048);
xor U23968 (N_23968,N_22280,N_20724);
xor U23969 (N_23969,N_22450,N_20369);
or U23970 (N_23970,N_20210,N_21613);
or U23971 (N_23971,N_22307,N_22047);
nand U23972 (N_23972,N_20989,N_20650);
or U23973 (N_23973,N_20617,N_20835);
xor U23974 (N_23974,N_20760,N_22284);
or U23975 (N_23975,N_21417,N_21551);
nand U23976 (N_23976,N_22395,N_20599);
xnor U23977 (N_23977,N_21280,N_20987);
xor U23978 (N_23978,N_22414,N_21702);
or U23979 (N_23979,N_20269,N_20976);
or U23980 (N_23980,N_20979,N_21560);
nand U23981 (N_23981,N_21855,N_22428);
or U23982 (N_23982,N_22124,N_21861);
nor U23983 (N_23983,N_22162,N_21556);
and U23984 (N_23984,N_21619,N_20896);
and U23985 (N_23985,N_22088,N_21894);
nor U23986 (N_23986,N_20217,N_21934);
and U23987 (N_23987,N_22165,N_22257);
nand U23988 (N_23988,N_20541,N_20657);
and U23989 (N_23989,N_20853,N_21415);
nand U23990 (N_23990,N_22295,N_22089);
nand U23991 (N_23991,N_20674,N_21286);
nor U23992 (N_23992,N_21094,N_21773);
xor U23993 (N_23993,N_22293,N_22272);
nand U23994 (N_23994,N_20319,N_21225);
or U23995 (N_23995,N_21650,N_22094);
nor U23996 (N_23996,N_22270,N_21138);
or U23997 (N_23997,N_20887,N_21000);
and U23998 (N_23998,N_21285,N_22446);
and U23999 (N_23999,N_21851,N_20490);
xor U24000 (N_24000,N_20711,N_21910);
nand U24001 (N_24001,N_21491,N_20368);
or U24002 (N_24002,N_21302,N_20596);
nor U24003 (N_24003,N_20839,N_21230);
and U24004 (N_24004,N_22483,N_21148);
or U24005 (N_24005,N_22432,N_20206);
nand U24006 (N_24006,N_22163,N_20627);
xnor U24007 (N_24007,N_21396,N_20454);
nor U24008 (N_24008,N_22013,N_21514);
nor U24009 (N_24009,N_20589,N_21909);
nor U24010 (N_24010,N_20098,N_22263);
or U24011 (N_24011,N_21341,N_20310);
xnor U24012 (N_24012,N_21025,N_20455);
or U24013 (N_24013,N_20057,N_21857);
and U24014 (N_24014,N_21747,N_20881);
nand U24015 (N_24015,N_21119,N_21925);
nand U24016 (N_24016,N_22409,N_21783);
xnor U24017 (N_24017,N_22068,N_20978);
nor U24018 (N_24018,N_22371,N_21950);
nand U24019 (N_24019,N_20516,N_21169);
nand U24020 (N_24020,N_21564,N_21665);
nor U24021 (N_24021,N_21370,N_21056);
xnor U24022 (N_24022,N_22036,N_22312);
and U24023 (N_24023,N_21032,N_20980);
or U24024 (N_24024,N_20923,N_21494);
xnor U24025 (N_24025,N_21295,N_22068);
xor U24026 (N_24026,N_21809,N_21250);
and U24027 (N_24027,N_21146,N_20947);
nor U24028 (N_24028,N_21889,N_21718);
or U24029 (N_24029,N_20860,N_21940);
xnor U24030 (N_24030,N_21489,N_21167);
nor U24031 (N_24031,N_21429,N_21043);
nand U24032 (N_24032,N_20163,N_22255);
or U24033 (N_24033,N_22003,N_21467);
xnor U24034 (N_24034,N_22169,N_22048);
or U24035 (N_24035,N_20479,N_20599);
and U24036 (N_24036,N_20675,N_22276);
xnor U24037 (N_24037,N_22074,N_20241);
nand U24038 (N_24038,N_21239,N_21814);
nor U24039 (N_24039,N_21384,N_21036);
nor U24040 (N_24040,N_20508,N_20223);
nor U24041 (N_24041,N_20660,N_20279);
or U24042 (N_24042,N_21768,N_21333);
or U24043 (N_24043,N_22018,N_22425);
or U24044 (N_24044,N_21614,N_20790);
xor U24045 (N_24045,N_20987,N_21655);
and U24046 (N_24046,N_21004,N_20285);
and U24047 (N_24047,N_20645,N_20868);
and U24048 (N_24048,N_21556,N_21175);
or U24049 (N_24049,N_20591,N_20910);
and U24050 (N_24050,N_21409,N_21132);
and U24051 (N_24051,N_21905,N_21646);
or U24052 (N_24052,N_20486,N_21269);
xnor U24053 (N_24053,N_21230,N_21367);
or U24054 (N_24054,N_21316,N_22044);
or U24055 (N_24055,N_21742,N_20256);
xor U24056 (N_24056,N_20457,N_20260);
nand U24057 (N_24057,N_21929,N_21791);
xnor U24058 (N_24058,N_21392,N_21439);
or U24059 (N_24059,N_21004,N_22216);
or U24060 (N_24060,N_21953,N_21115);
and U24061 (N_24061,N_21298,N_21359);
and U24062 (N_24062,N_22218,N_21751);
xor U24063 (N_24063,N_21870,N_21741);
or U24064 (N_24064,N_20831,N_20386);
xnor U24065 (N_24065,N_21162,N_22154);
and U24066 (N_24066,N_22276,N_21539);
or U24067 (N_24067,N_20032,N_22240);
nor U24068 (N_24068,N_20191,N_21745);
nor U24069 (N_24069,N_21921,N_20828);
and U24070 (N_24070,N_21985,N_20525);
nor U24071 (N_24071,N_20039,N_20096);
or U24072 (N_24072,N_21444,N_21857);
or U24073 (N_24073,N_22008,N_21512);
nor U24074 (N_24074,N_21190,N_20053);
or U24075 (N_24075,N_22024,N_20659);
or U24076 (N_24076,N_20712,N_20255);
nand U24077 (N_24077,N_21183,N_20923);
xor U24078 (N_24078,N_20229,N_20034);
or U24079 (N_24079,N_21062,N_20955);
nor U24080 (N_24080,N_22146,N_21740);
xnor U24081 (N_24081,N_21862,N_20542);
nand U24082 (N_24082,N_20264,N_20460);
xnor U24083 (N_24083,N_20102,N_21996);
or U24084 (N_24084,N_22122,N_21403);
or U24085 (N_24085,N_20741,N_21209);
nor U24086 (N_24086,N_20623,N_20928);
xnor U24087 (N_24087,N_22210,N_20776);
nand U24088 (N_24088,N_21267,N_21324);
and U24089 (N_24089,N_20169,N_20755);
nand U24090 (N_24090,N_20094,N_21685);
and U24091 (N_24091,N_22220,N_20586);
nor U24092 (N_24092,N_21185,N_22060);
xnor U24093 (N_24093,N_22144,N_20259);
xnor U24094 (N_24094,N_20639,N_21168);
and U24095 (N_24095,N_21194,N_21302);
and U24096 (N_24096,N_22012,N_22168);
xnor U24097 (N_24097,N_22085,N_20904);
and U24098 (N_24098,N_21626,N_20844);
xor U24099 (N_24099,N_22213,N_22210);
xor U24100 (N_24100,N_20604,N_20735);
and U24101 (N_24101,N_21258,N_21836);
nand U24102 (N_24102,N_20174,N_20099);
or U24103 (N_24103,N_20418,N_21185);
and U24104 (N_24104,N_21828,N_20223);
or U24105 (N_24105,N_21534,N_21316);
xnor U24106 (N_24106,N_21692,N_21449);
nand U24107 (N_24107,N_22409,N_21138);
or U24108 (N_24108,N_21080,N_20883);
nor U24109 (N_24109,N_21232,N_21183);
xnor U24110 (N_24110,N_20767,N_22321);
xor U24111 (N_24111,N_22488,N_22331);
xor U24112 (N_24112,N_21592,N_22111);
or U24113 (N_24113,N_21325,N_21342);
or U24114 (N_24114,N_20543,N_20994);
and U24115 (N_24115,N_21489,N_22057);
nor U24116 (N_24116,N_21998,N_20911);
and U24117 (N_24117,N_21909,N_20454);
and U24118 (N_24118,N_21414,N_22421);
nor U24119 (N_24119,N_22090,N_21730);
nand U24120 (N_24120,N_22189,N_22163);
xor U24121 (N_24121,N_20608,N_21664);
or U24122 (N_24122,N_22414,N_20113);
and U24123 (N_24123,N_20444,N_20418);
and U24124 (N_24124,N_21295,N_22469);
or U24125 (N_24125,N_20599,N_21576);
nand U24126 (N_24126,N_22181,N_20734);
nand U24127 (N_24127,N_21610,N_21238);
or U24128 (N_24128,N_21245,N_21841);
and U24129 (N_24129,N_21921,N_21022);
nand U24130 (N_24130,N_21610,N_20403);
nand U24131 (N_24131,N_22451,N_20061);
and U24132 (N_24132,N_22259,N_21673);
and U24133 (N_24133,N_21130,N_20667);
xor U24134 (N_24134,N_20800,N_21465);
nor U24135 (N_24135,N_21090,N_20902);
nor U24136 (N_24136,N_21192,N_22378);
xor U24137 (N_24137,N_20033,N_21776);
and U24138 (N_24138,N_22027,N_20634);
nor U24139 (N_24139,N_21475,N_20002);
or U24140 (N_24140,N_21478,N_21144);
xnor U24141 (N_24141,N_20561,N_21945);
nor U24142 (N_24142,N_20564,N_20176);
xnor U24143 (N_24143,N_20172,N_20445);
and U24144 (N_24144,N_20922,N_20864);
xor U24145 (N_24145,N_22076,N_20160);
or U24146 (N_24146,N_20748,N_22132);
xnor U24147 (N_24147,N_20943,N_21054);
nand U24148 (N_24148,N_20080,N_22480);
or U24149 (N_24149,N_22457,N_22368);
and U24150 (N_24150,N_20308,N_21143);
xnor U24151 (N_24151,N_21165,N_21267);
and U24152 (N_24152,N_20190,N_20449);
nand U24153 (N_24153,N_22394,N_21155);
and U24154 (N_24154,N_20971,N_20542);
xnor U24155 (N_24155,N_20227,N_21848);
and U24156 (N_24156,N_20555,N_22188);
and U24157 (N_24157,N_20687,N_22179);
xnor U24158 (N_24158,N_21906,N_21686);
xnor U24159 (N_24159,N_21211,N_21393);
nand U24160 (N_24160,N_21388,N_21594);
nand U24161 (N_24161,N_21240,N_21488);
nor U24162 (N_24162,N_20926,N_22190);
or U24163 (N_24163,N_20725,N_20406);
xor U24164 (N_24164,N_20577,N_21404);
xor U24165 (N_24165,N_21457,N_20804);
and U24166 (N_24166,N_21092,N_22291);
and U24167 (N_24167,N_21117,N_21398);
and U24168 (N_24168,N_20222,N_21180);
or U24169 (N_24169,N_22056,N_21743);
nand U24170 (N_24170,N_22436,N_20643);
nand U24171 (N_24171,N_21843,N_21702);
xnor U24172 (N_24172,N_21666,N_22152);
and U24173 (N_24173,N_22333,N_22326);
or U24174 (N_24174,N_21202,N_22280);
xor U24175 (N_24175,N_20987,N_21717);
nand U24176 (N_24176,N_22457,N_21300);
or U24177 (N_24177,N_21787,N_22488);
or U24178 (N_24178,N_20849,N_21261);
nor U24179 (N_24179,N_21812,N_20364);
or U24180 (N_24180,N_21884,N_20693);
or U24181 (N_24181,N_20293,N_20496);
and U24182 (N_24182,N_21259,N_20098);
and U24183 (N_24183,N_20399,N_21382);
and U24184 (N_24184,N_22409,N_20657);
xor U24185 (N_24185,N_22036,N_22446);
nor U24186 (N_24186,N_22345,N_20529);
xnor U24187 (N_24187,N_20538,N_22254);
xor U24188 (N_24188,N_20585,N_20776);
nor U24189 (N_24189,N_20529,N_21745);
or U24190 (N_24190,N_20103,N_21834);
nand U24191 (N_24191,N_22067,N_20554);
xnor U24192 (N_24192,N_21525,N_20653);
and U24193 (N_24193,N_20139,N_21785);
nand U24194 (N_24194,N_20130,N_22428);
nand U24195 (N_24195,N_21697,N_20043);
nand U24196 (N_24196,N_20465,N_22489);
or U24197 (N_24197,N_22461,N_21226);
nor U24198 (N_24198,N_21165,N_22114);
nor U24199 (N_24199,N_21484,N_20837);
nor U24200 (N_24200,N_21574,N_20539);
xnor U24201 (N_24201,N_21410,N_20296);
nor U24202 (N_24202,N_21480,N_21977);
or U24203 (N_24203,N_21351,N_20255);
nand U24204 (N_24204,N_22213,N_20417);
nor U24205 (N_24205,N_21229,N_20610);
and U24206 (N_24206,N_21632,N_20573);
nor U24207 (N_24207,N_22338,N_20388);
xor U24208 (N_24208,N_21494,N_21804);
xnor U24209 (N_24209,N_21127,N_22475);
xnor U24210 (N_24210,N_21478,N_22068);
or U24211 (N_24211,N_22139,N_20592);
nand U24212 (N_24212,N_22267,N_21668);
or U24213 (N_24213,N_20498,N_21036);
nor U24214 (N_24214,N_20452,N_21768);
and U24215 (N_24215,N_20061,N_20603);
nor U24216 (N_24216,N_20985,N_21156);
or U24217 (N_24217,N_20150,N_20617);
xnor U24218 (N_24218,N_21099,N_22309);
or U24219 (N_24219,N_20955,N_20069);
and U24220 (N_24220,N_22307,N_22334);
nand U24221 (N_24221,N_20900,N_20364);
xor U24222 (N_24222,N_21107,N_22389);
nand U24223 (N_24223,N_21497,N_20016);
nor U24224 (N_24224,N_21447,N_20585);
or U24225 (N_24225,N_20345,N_21078);
xnor U24226 (N_24226,N_21546,N_20430);
and U24227 (N_24227,N_20667,N_20177);
and U24228 (N_24228,N_21941,N_21039);
and U24229 (N_24229,N_20449,N_21706);
nand U24230 (N_24230,N_20207,N_20940);
and U24231 (N_24231,N_21050,N_20938);
nand U24232 (N_24232,N_20350,N_21712);
and U24233 (N_24233,N_22224,N_20424);
or U24234 (N_24234,N_20787,N_21404);
and U24235 (N_24235,N_20806,N_20853);
or U24236 (N_24236,N_22012,N_22094);
or U24237 (N_24237,N_22193,N_21374);
nor U24238 (N_24238,N_22028,N_20689);
nand U24239 (N_24239,N_20304,N_21710);
and U24240 (N_24240,N_20987,N_21759);
or U24241 (N_24241,N_21972,N_21313);
or U24242 (N_24242,N_21005,N_20616);
nand U24243 (N_24243,N_21724,N_20160);
xnor U24244 (N_24244,N_21191,N_21236);
nand U24245 (N_24245,N_20483,N_20012);
xnor U24246 (N_24246,N_20432,N_22480);
nand U24247 (N_24247,N_21788,N_20924);
nand U24248 (N_24248,N_20723,N_20659);
nand U24249 (N_24249,N_21569,N_21318);
nor U24250 (N_24250,N_20219,N_21344);
and U24251 (N_24251,N_21715,N_21170);
nor U24252 (N_24252,N_20644,N_22291);
and U24253 (N_24253,N_20453,N_21416);
nor U24254 (N_24254,N_21232,N_21563);
and U24255 (N_24255,N_21032,N_20984);
xor U24256 (N_24256,N_21461,N_20194);
xor U24257 (N_24257,N_20947,N_21480);
nor U24258 (N_24258,N_22428,N_20560);
or U24259 (N_24259,N_21865,N_22139);
and U24260 (N_24260,N_20024,N_21820);
nor U24261 (N_24261,N_20494,N_21844);
xor U24262 (N_24262,N_20826,N_20219);
xor U24263 (N_24263,N_22047,N_20407);
and U24264 (N_24264,N_20709,N_20448);
xnor U24265 (N_24265,N_21400,N_20500);
or U24266 (N_24266,N_20174,N_21768);
or U24267 (N_24267,N_21485,N_21138);
nand U24268 (N_24268,N_21572,N_20406);
xor U24269 (N_24269,N_20046,N_22205);
or U24270 (N_24270,N_20037,N_22183);
and U24271 (N_24271,N_21935,N_20056);
nand U24272 (N_24272,N_20181,N_20827);
nand U24273 (N_24273,N_21963,N_20710);
and U24274 (N_24274,N_20529,N_21769);
or U24275 (N_24275,N_20177,N_22278);
xnor U24276 (N_24276,N_20907,N_21463);
nor U24277 (N_24277,N_20477,N_20781);
or U24278 (N_24278,N_21634,N_20198);
xor U24279 (N_24279,N_20189,N_20216);
or U24280 (N_24280,N_22458,N_21998);
nand U24281 (N_24281,N_20317,N_20961);
nor U24282 (N_24282,N_22021,N_20028);
nand U24283 (N_24283,N_21911,N_22341);
or U24284 (N_24284,N_20217,N_20893);
nor U24285 (N_24285,N_20565,N_21150);
nand U24286 (N_24286,N_20113,N_21807);
nor U24287 (N_24287,N_20045,N_20934);
nand U24288 (N_24288,N_22004,N_20989);
or U24289 (N_24289,N_20026,N_22088);
nor U24290 (N_24290,N_20855,N_20910);
or U24291 (N_24291,N_20021,N_22401);
xor U24292 (N_24292,N_20475,N_20308);
and U24293 (N_24293,N_20642,N_22243);
nor U24294 (N_24294,N_21970,N_21376);
nor U24295 (N_24295,N_21766,N_21762);
and U24296 (N_24296,N_21392,N_20427);
nor U24297 (N_24297,N_21572,N_21277);
nand U24298 (N_24298,N_22424,N_22354);
and U24299 (N_24299,N_21331,N_20946);
nor U24300 (N_24300,N_20078,N_22087);
and U24301 (N_24301,N_20206,N_21006);
nand U24302 (N_24302,N_21193,N_22056);
xor U24303 (N_24303,N_22330,N_20791);
and U24304 (N_24304,N_20718,N_21314);
nand U24305 (N_24305,N_21321,N_20929);
or U24306 (N_24306,N_22328,N_22473);
xor U24307 (N_24307,N_22460,N_20930);
and U24308 (N_24308,N_20770,N_22253);
and U24309 (N_24309,N_20984,N_20674);
nand U24310 (N_24310,N_21001,N_20762);
or U24311 (N_24311,N_22410,N_21279);
xnor U24312 (N_24312,N_20626,N_21764);
xnor U24313 (N_24313,N_21130,N_22193);
nand U24314 (N_24314,N_20976,N_20785);
xor U24315 (N_24315,N_20005,N_21858);
nor U24316 (N_24316,N_20229,N_21423);
xor U24317 (N_24317,N_21582,N_20188);
or U24318 (N_24318,N_20567,N_20591);
xnor U24319 (N_24319,N_20645,N_20997);
and U24320 (N_24320,N_22027,N_21568);
and U24321 (N_24321,N_20497,N_20781);
and U24322 (N_24322,N_21715,N_20972);
nor U24323 (N_24323,N_21582,N_20292);
nand U24324 (N_24324,N_20700,N_21770);
or U24325 (N_24325,N_21803,N_22013);
and U24326 (N_24326,N_20995,N_20556);
or U24327 (N_24327,N_20294,N_20054);
or U24328 (N_24328,N_20240,N_20808);
and U24329 (N_24329,N_21293,N_20815);
or U24330 (N_24330,N_21277,N_20657);
nor U24331 (N_24331,N_20366,N_20580);
xnor U24332 (N_24332,N_20639,N_21447);
xnor U24333 (N_24333,N_20389,N_22287);
or U24334 (N_24334,N_21825,N_22227);
and U24335 (N_24335,N_20668,N_21333);
nand U24336 (N_24336,N_21123,N_21944);
nor U24337 (N_24337,N_21201,N_20559);
and U24338 (N_24338,N_20648,N_20766);
xor U24339 (N_24339,N_20158,N_20770);
nor U24340 (N_24340,N_20383,N_20371);
nand U24341 (N_24341,N_21842,N_21556);
nand U24342 (N_24342,N_22229,N_20611);
xor U24343 (N_24343,N_21619,N_22407);
nand U24344 (N_24344,N_20818,N_20090);
or U24345 (N_24345,N_20883,N_20185);
nand U24346 (N_24346,N_20272,N_22240);
nor U24347 (N_24347,N_21455,N_21781);
or U24348 (N_24348,N_21249,N_21661);
nand U24349 (N_24349,N_22327,N_20386);
or U24350 (N_24350,N_21307,N_22279);
xor U24351 (N_24351,N_22234,N_22123);
nand U24352 (N_24352,N_21405,N_21297);
xor U24353 (N_24353,N_21386,N_21538);
nand U24354 (N_24354,N_21990,N_21793);
and U24355 (N_24355,N_20295,N_20619);
nand U24356 (N_24356,N_21137,N_21290);
and U24357 (N_24357,N_21354,N_22162);
and U24358 (N_24358,N_21922,N_20754);
or U24359 (N_24359,N_22402,N_21902);
or U24360 (N_24360,N_22434,N_22330);
nor U24361 (N_24361,N_21391,N_21690);
nand U24362 (N_24362,N_20096,N_20612);
nand U24363 (N_24363,N_21643,N_22119);
nor U24364 (N_24364,N_20813,N_21234);
or U24365 (N_24365,N_20545,N_22312);
or U24366 (N_24366,N_20736,N_20095);
nand U24367 (N_24367,N_21271,N_20861);
or U24368 (N_24368,N_22332,N_20448);
and U24369 (N_24369,N_21666,N_21996);
or U24370 (N_24370,N_20907,N_21722);
and U24371 (N_24371,N_20089,N_20700);
nor U24372 (N_24372,N_20058,N_20766);
xor U24373 (N_24373,N_22161,N_21763);
nor U24374 (N_24374,N_21020,N_22324);
or U24375 (N_24375,N_20024,N_20720);
nand U24376 (N_24376,N_22317,N_21591);
xor U24377 (N_24377,N_20043,N_21993);
nor U24378 (N_24378,N_20628,N_21095);
nand U24379 (N_24379,N_20199,N_22466);
nand U24380 (N_24380,N_21576,N_21648);
xor U24381 (N_24381,N_21201,N_21332);
nor U24382 (N_24382,N_22351,N_20468);
and U24383 (N_24383,N_20249,N_20859);
or U24384 (N_24384,N_20945,N_20406);
nor U24385 (N_24385,N_20281,N_20221);
and U24386 (N_24386,N_21608,N_20479);
or U24387 (N_24387,N_21095,N_21662);
nand U24388 (N_24388,N_20129,N_21809);
or U24389 (N_24389,N_21643,N_20347);
nand U24390 (N_24390,N_20953,N_20593);
and U24391 (N_24391,N_20490,N_22197);
and U24392 (N_24392,N_20288,N_20776);
nand U24393 (N_24393,N_21275,N_22454);
or U24394 (N_24394,N_20586,N_21451);
and U24395 (N_24395,N_22104,N_21712);
nor U24396 (N_24396,N_20547,N_20477);
xnor U24397 (N_24397,N_20737,N_21122);
or U24398 (N_24398,N_21004,N_21896);
nand U24399 (N_24399,N_21289,N_21776);
and U24400 (N_24400,N_20713,N_21436);
nand U24401 (N_24401,N_20861,N_22192);
nand U24402 (N_24402,N_20205,N_21788);
xor U24403 (N_24403,N_21547,N_22056);
or U24404 (N_24404,N_22443,N_21719);
nor U24405 (N_24405,N_20677,N_21053);
or U24406 (N_24406,N_20044,N_20930);
xnor U24407 (N_24407,N_20521,N_20846);
and U24408 (N_24408,N_20900,N_21792);
nor U24409 (N_24409,N_21377,N_20521);
nand U24410 (N_24410,N_21807,N_22348);
or U24411 (N_24411,N_22109,N_21584);
xnor U24412 (N_24412,N_22114,N_22220);
nor U24413 (N_24413,N_22313,N_20120);
xor U24414 (N_24414,N_22045,N_20730);
nor U24415 (N_24415,N_22215,N_22401);
nor U24416 (N_24416,N_21439,N_20869);
or U24417 (N_24417,N_22116,N_20146);
xnor U24418 (N_24418,N_21042,N_20873);
and U24419 (N_24419,N_22407,N_21639);
or U24420 (N_24420,N_22163,N_21079);
nand U24421 (N_24421,N_20563,N_21468);
or U24422 (N_24422,N_20673,N_21766);
nand U24423 (N_24423,N_20439,N_21664);
xnor U24424 (N_24424,N_22395,N_21567);
nand U24425 (N_24425,N_20476,N_21347);
and U24426 (N_24426,N_21045,N_21798);
and U24427 (N_24427,N_20457,N_22454);
xor U24428 (N_24428,N_20750,N_21009);
nor U24429 (N_24429,N_22063,N_22163);
or U24430 (N_24430,N_22368,N_20156);
nor U24431 (N_24431,N_21649,N_21273);
nand U24432 (N_24432,N_20785,N_21439);
or U24433 (N_24433,N_22302,N_21638);
nand U24434 (N_24434,N_22154,N_22078);
xnor U24435 (N_24435,N_22179,N_21367);
nor U24436 (N_24436,N_21624,N_21931);
and U24437 (N_24437,N_20610,N_21461);
xor U24438 (N_24438,N_20526,N_20447);
and U24439 (N_24439,N_21550,N_22224);
or U24440 (N_24440,N_21021,N_20054);
or U24441 (N_24441,N_21324,N_22349);
and U24442 (N_24442,N_20452,N_21700);
nand U24443 (N_24443,N_22160,N_20664);
nor U24444 (N_24444,N_20611,N_21579);
nor U24445 (N_24445,N_20314,N_21475);
xor U24446 (N_24446,N_21711,N_20484);
nor U24447 (N_24447,N_20776,N_21040);
or U24448 (N_24448,N_21075,N_22377);
nand U24449 (N_24449,N_21463,N_21841);
or U24450 (N_24450,N_21780,N_21271);
and U24451 (N_24451,N_20629,N_22008);
nand U24452 (N_24452,N_22143,N_20795);
and U24453 (N_24453,N_21824,N_21149);
nor U24454 (N_24454,N_22436,N_22347);
and U24455 (N_24455,N_20324,N_22165);
or U24456 (N_24456,N_22437,N_22248);
nor U24457 (N_24457,N_20527,N_20292);
nor U24458 (N_24458,N_22153,N_20165);
nor U24459 (N_24459,N_20278,N_20699);
nand U24460 (N_24460,N_20105,N_20901);
or U24461 (N_24461,N_20445,N_20558);
or U24462 (N_24462,N_20094,N_21613);
nand U24463 (N_24463,N_20061,N_21861);
nor U24464 (N_24464,N_21490,N_21367);
xor U24465 (N_24465,N_22109,N_20864);
nor U24466 (N_24466,N_21178,N_20077);
or U24467 (N_24467,N_20640,N_20892);
xnor U24468 (N_24468,N_20628,N_22296);
xor U24469 (N_24469,N_21234,N_20585);
or U24470 (N_24470,N_21857,N_22420);
xor U24471 (N_24471,N_22126,N_20826);
and U24472 (N_24472,N_22252,N_20517);
nor U24473 (N_24473,N_20175,N_20110);
and U24474 (N_24474,N_20023,N_20195);
nand U24475 (N_24475,N_20215,N_22101);
nand U24476 (N_24476,N_20738,N_20046);
nand U24477 (N_24477,N_20904,N_21304);
or U24478 (N_24478,N_22032,N_20854);
or U24479 (N_24479,N_20071,N_22023);
and U24480 (N_24480,N_20483,N_20046);
nor U24481 (N_24481,N_20023,N_20227);
nand U24482 (N_24482,N_21111,N_20452);
xnor U24483 (N_24483,N_21926,N_20658);
nor U24484 (N_24484,N_21040,N_20550);
nor U24485 (N_24485,N_22134,N_20471);
nand U24486 (N_24486,N_21414,N_21734);
or U24487 (N_24487,N_20427,N_22226);
or U24488 (N_24488,N_22039,N_20686);
xor U24489 (N_24489,N_21920,N_21756);
or U24490 (N_24490,N_20696,N_21321);
or U24491 (N_24491,N_21962,N_21657);
nor U24492 (N_24492,N_22294,N_20058);
and U24493 (N_24493,N_20179,N_21141);
and U24494 (N_24494,N_20755,N_21416);
nand U24495 (N_24495,N_21616,N_20570);
xor U24496 (N_24496,N_21150,N_20950);
xor U24497 (N_24497,N_20884,N_20802);
nor U24498 (N_24498,N_20771,N_20153);
or U24499 (N_24499,N_21436,N_22277);
nor U24500 (N_24500,N_21922,N_22280);
nor U24501 (N_24501,N_21296,N_20225);
and U24502 (N_24502,N_21674,N_21253);
or U24503 (N_24503,N_22328,N_21118);
xnor U24504 (N_24504,N_20726,N_20588);
and U24505 (N_24505,N_20120,N_20563);
xnor U24506 (N_24506,N_20762,N_21906);
nor U24507 (N_24507,N_22166,N_21672);
and U24508 (N_24508,N_20545,N_22323);
and U24509 (N_24509,N_20313,N_20210);
or U24510 (N_24510,N_20882,N_20302);
nor U24511 (N_24511,N_22055,N_21455);
xor U24512 (N_24512,N_20322,N_21876);
xnor U24513 (N_24513,N_22296,N_20385);
or U24514 (N_24514,N_20084,N_21391);
and U24515 (N_24515,N_20039,N_20555);
and U24516 (N_24516,N_22080,N_22246);
nor U24517 (N_24517,N_20507,N_21129);
nand U24518 (N_24518,N_20830,N_21039);
xnor U24519 (N_24519,N_20537,N_21784);
nand U24520 (N_24520,N_22388,N_20064);
nand U24521 (N_24521,N_22181,N_21405);
nand U24522 (N_24522,N_21615,N_21698);
nand U24523 (N_24523,N_21465,N_21860);
xnor U24524 (N_24524,N_21306,N_20068);
xor U24525 (N_24525,N_20168,N_20201);
and U24526 (N_24526,N_22280,N_22036);
or U24527 (N_24527,N_21808,N_20759);
or U24528 (N_24528,N_20948,N_21045);
nand U24529 (N_24529,N_22364,N_21598);
nor U24530 (N_24530,N_20962,N_21348);
nor U24531 (N_24531,N_20060,N_22238);
nand U24532 (N_24532,N_21632,N_21300);
and U24533 (N_24533,N_22033,N_21936);
or U24534 (N_24534,N_22134,N_20509);
nor U24535 (N_24535,N_20508,N_22320);
and U24536 (N_24536,N_22271,N_21553);
or U24537 (N_24537,N_20382,N_21142);
nand U24538 (N_24538,N_20213,N_22051);
xnor U24539 (N_24539,N_21365,N_21017);
or U24540 (N_24540,N_20252,N_20636);
xor U24541 (N_24541,N_21470,N_22007);
nand U24542 (N_24542,N_20672,N_21842);
nand U24543 (N_24543,N_21770,N_21995);
and U24544 (N_24544,N_21781,N_20682);
nand U24545 (N_24545,N_20991,N_21190);
xor U24546 (N_24546,N_22220,N_22495);
xnor U24547 (N_24547,N_21561,N_21206);
nor U24548 (N_24548,N_21385,N_21526);
nor U24549 (N_24549,N_20791,N_21620);
nor U24550 (N_24550,N_20383,N_21244);
nand U24551 (N_24551,N_21276,N_20225);
nand U24552 (N_24552,N_22462,N_20301);
and U24553 (N_24553,N_21879,N_21320);
xnor U24554 (N_24554,N_21103,N_21556);
or U24555 (N_24555,N_20800,N_21064);
nor U24556 (N_24556,N_22302,N_20906);
xnor U24557 (N_24557,N_22356,N_21903);
xnor U24558 (N_24558,N_20048,N_21404);
or U24559 (N_24559,N_21311,N_22417);
nor U24560 (N_24560,N_20166,N_22456);
nor U24561 (N_24561,N_21343,N_21085);
nand U24562 (N_24562,N_20838,N_21933);
and U24563 (N_24563,N_20331,N_21334);
and U24564 (N_24564,N_20722,N_21781);
nor U24565 (N_24565,N_22080,N_21037);
xnor U24566 (N_24566,N_20257,N_20916);
nand U24567 (N_24567,N_20422,N_20875);
nor U24568 (N_24568,N_20472,N_21149);
or U24569 (N_24569,N_21055,N_21936);
nand U24570 (N_24570,N_20356,N_20331);
nand U24571 (N_24571,N_21514,N_20561);
and U24572 (N_24572,N_21263,N_21572);
nand U24573 (N_24573,N_21194,N_22188);
nor U24574 (N_24574,N_21182,N_21254);
nor U24575 (N_24575,N_22195,N_20275);
nand U24576 (N_24576,N_21241,N_22405);
nand U24577 (N_24577,N_20688,N_21731);
nand U24578 (N_24578,N_21121,N_20296);
and U24579 (N_24579,N_21851,N_22444);
and U24580 (N_24580,N_22164,N_20565);
xor U24581 (N_24581,N_21915,N_20276);
nand U24582 (N_24582,N_20933,N_21118);
or U24583 (N_24583,N_22472,N_21605);
xor U24584 (N_24584,N_21753,N_21867);
and U24585 (N_24585,N_22063,N_20255);
xnor U24586 (N_24586,N_20642,N_20582);
and U24587 (N_24587,N_21391,N_20183);
and U24588 (N_24588,N_20722,N_20679);
nand U24589 (N_24589,N_20034,N_22245);
or U24590 (N_24590,N_21097,N_21326);
or U24591 (N_24591,N_20582,N_21657);
and U24592 (N_24592,N_21249,N_21068);
or U24593 (N_24593,N_22023,N_21691);
xnor U24594 (N_24594,N_21412,N_20151);
nand U24595 (N_24595,N_20601,N_20593);
nand U24596 (N_24596,N_21146,N_22265);
or U24597 (N_24597,N_21655,N_20678);
or U24598 (N_24598,N_21944,N_21260);
nor U24599 (N_24599,N_22193,N_20512);
and U24600 (N_24600,N_20171,N_21005);
xor U24601 (N_24601,N_21257,N_21044);
or U24602 (N_24602,N_22268,N_20370);
nor U24603 (N_24603,N_20683,N_21699);
and U24604 (N_24604,N_20031,N_21404);
xor U24605 (N_24605,N_20722,N_22346);
or U24606 (N_24606,N_21620,N_21358);
nor U24607 (N_24607,N_22296,N_22190);
nor U24608 (N_24608,N_21886,N_22305);
xnor U24609 (N_24609,N_21886,N_22354);
xor U24610 (N_24610,N_22454,N_21701);
nor U24611 (N_24611,N_20027,N_22068);
nor U24612 (N_24612,N_20751,N_20294);
and U24613 (N_24613,N_21062,N_20354);
or U24614 (N_24614,N_20514,N_22149);
nand U24615 (N_24615,N_20305,N_21978);
and U24616 (N_24616,N_20384,N_21698);
and U24617 (N_24617,N_21540,N_22155);
and U24618 (N_24618,N_20651,N_20911);
xor U24619 (N_24619,N_22090,N_21657);
or U24620 (N_24620,N_20197,N_20851);
and U24621 (N_24621,N_21234,N_21572);
xor U24622 (N_24622,N_21432,N_22347);
xnor U24623 (N_24623,N_21797,N_21869);
or U24624 (N_24624,N_20022,N_21608);
xnor U24625 (N_24625,N_21556,N_20336);
and U24626 (N_24626,N_21831,N_20241);
nor U24627 (N_24627,N_21395,N_20747);
xor U24628 (N_24628,N_21755,N_20004);
nor U24629 (N_24629,N_20530,N_21657);
nand U24630 (N_24630,N_21534,N_22306);
or U24631 (N_24631,N_22409,N_20590);
and U24632 (N_24632,N_21201,N_20800);
nor U24633 (N_24633,N_20593,N_21289);
nand U24634 (N_24634,N_20952,N_21262);
nor U24635 (N_24635,N_20960,N_20428);
nor U24636 (N_24636,N_21488,N_21034);
nor U24637 (N_24637,N_20254,N_20259);
nand U24638 (N_24638,N_21586,N_21460);
xnor U24639 (N_24639,N_22088,N_20945);
or U24640 (N_24640,N_21747,N_20017);
or U24641 (N_24641,N_21809,N_20243);
xor U24642 (N_24642,N_22048,N_22175);
and U24643 (N_24643,N_22439,N_21656);
or U24644 (N_24644,N_21198,N_21619);
nor U24645 (N_24645,N_20068,N_21406);
xnor U24646 (N_24646,N_20810,N_20194);
xor U24647 (N_24647,N_22106,N_21985);
nand U24648 (N_24648,N_21957,N_20220);
xnor U24649 (N_24649,N_21082,N_21652);
xnor U24650 (N_24650,N_21459,N_20294);
nor U24651 (N_24651,N_21862,N_20739);
or U24652 (N_24652,N_21129,N_22298);
nor U24653 (N_24653,N_21839,N_20260);
and U24654 (N_24654,N_22308,N_20193);
nor U24655 (N_24655,N_21847,N_21688);
nand U24656 (N_24656,N_21131,N_20678);
xnor U24657 (N_24657,N_21940,N_22292);
and U24658 (N_24658,N_21125,N_20096);
nand U24659 (N_24659,N_20467,N_20253);
or U24660 (N_24660,N_21589,N_21724);
xor U24661 (N_24661,N_22324,N_20957);
or U24662 (N_24662,N_21007,N_20687);
xor U24663 (N_24663,N_21692,N_22291);
xor U24664 (N_24664,N_22128,N_20724);
xnor U24665 (N_24665,N_21284,N_22025);
and U24666 (N_24666,N_21458,N_20065);
xor U24667 (N_24667,N_21130,N_21374);
nand U24668 (N_24668,N_21219,N_21963);
nor U24669 (N_24669,N_22428,N_21332);
xor U24670 (N_24670,N_20733,N_20309);
xor U24671 (N_24671,N_20419,N_22266);
and U24672 (N_24672,N_22283,N_21614);
nor U24673 (N_24673,N_21147,N_21168);
or U24674 (N_24674,N_22269,N_21555);
nand U24675 (N_24675,N_20277,N_20296);
nand U24676 (N_24676,N_21988,N_20056);
nor U24677 (N_24677,N_20739,N_20734);
or U24678 (N_24678,N_22064,N_20463);
xor U24679 (N_24679,N_20679,N_21916);
nor U24680 (N_24680,N_20499,N_22214);
or U24681 (N_24681,N_21352,N_22333);
xor U24682 (N_24682,N_20653,N_20510);
or U24683 (N_24683,N_21192,N_20848);
nor U24684 (N_24684,N_22125,N_20321);
and U24685 (N_24685,N_21203,N_22228);
or U24686 (N_24686,N_20131,N_20495);
and U24687 (N_24687,N_20953,N_22388);
nor U24688 (N_24688,N_22215,N_21162);
and U24689 (N_24689,N_20913,N_21350);
and U24690 (N_24690,N_21574,N_21426);
xnor U24691 (N_24691,N_22026,N_21282);
nand U24692 (N_24692,N_20113,N_20066);
and U24693 (N_24693,N_22386,N_22475);
nor U24694 (N_24694,N_20599,N_21572);
nand U24695 (N_24695,N_20963,N_20196);
xor U24696 (N_24696,N_20571,N_22039);
and U24697 (N_24697,N_22166,N_20147);
nor U24698 (N_24698,N_20377,N_20524);
and U24699 (N_24699,N_21707,N_20475);
and U24700 (N_24700,N_22360,N_20437);
and U24701 (N_24701,N_21072,N_21095);
and U24702 (N_24702,N_22001,N_21046);
or U24703 (N_24703,N_20420,N_20962);
and U24704 (N_24704,N_20723,N_21721);
xnor U24705 (N_24705,N_21723,N_21541);
nor U24706 (N_24706,N_20826,N_20365);
nor U24707 (N_24707,N_21098,N_20317);
nor U24708 (N_24708,N_21387,N_22456);
and U24709 (N_24709,N_20240,N_22246);
and U24710 (N_24710,N_20706,N_20087);
nor U24711 (N_24711,N_20289,N_20281);
nor U24712 (N_24712,N_21499,N_22237);
and U24713 (N_24713,N_21280,N_21781);
nor U24714 (N_24714,N_21426,N_22026);
or U24715 (N_24715,N_20133,N_21525);
xnor U24716 (N_24716,N_21521,N_21718);
nand U24717 (N_24717,N_20178,N_20506);
or U24718 (N_24718,N_20644,N_21998);
nor U24719 (N_24719,N_22358,N_21484);
xor U24720 (N_24720,N_22430,N_21733);
and U24721 (N_24721,N_20216,N_20827);
nand U24722 (N_24722,N_21198,N_21733);
and U24723 (N_24723,N_21856,N_20128);
xnor U24724 (N_24724,N_20811,N_22367);
and U24725 (N_24725,N_21207,N_20167);
nor U24726 (N_24726,N_21218,N_21109);
or U24727 (N_24727,N_20247,N_20573);
nor U24728 (N_24728,N_21199,N_22486);
nand U24729 (N_24729,N_22206,N_21968);
nor U24730 (N_24730,N_21458,N_21133);
nor U24731 (N_24731,N_20656,N_22393);
or U24732 (N_24732,N_21479,N_21130);
nand U24733 (N_24733,N_20116,N_20566);
nor U24734 (N_24734,N_22247,N_20405);
nor U24735 (N_24735,N_21818,N_20613);
xnor U24736 (N_24736,N_21563,N_21605);
or U24737 (N_24737,N_20961,N_20738);
xor U24738 (N_24738,N_21607,N_22035);
or U24739 (N_24739,N_22302,N_21331);
xnor U24740 (N_24740,N_22091,N_21144);
or U24741 (N_24741,N_21753,N_20726);
or U24742 (N_24742,N_20666,N_21174);
nor U24743 (N_24743,N_21027,N_21959);
nor U24744 (N_24744,N_22223,N_20209);
nor U24745 (N_24745,N_20960,N_20552);
and U24746 (N_24746,N_21594,N_22365);
xor U24747 (N_24747,N_21266,N_21902);
nand U24748 (N_24748,N_20830,N_21353);
nor U24749 (N_24749,N_21450,N_21214);
nor U24750 (N_24750,N_22085,N_20780);
nor U24751 (N_24751,N_22106,N_21948);
or U24752 (N_24752,N_20880,N_20757);
nand U24753 (N_24753,N_21550,N_22441);
and U24754 (N_24754,N_21248,N_20219);
and U24755 (N_24755,N_21116,N_20688);
or U24756 (N_24756,N_21934,N_20999);
or U24757 (N_24757,N_21130,N_20612);
and U24758 (N_24758,N_20826,N_20309);
nor U24759 (N_24759,N_21734,N_22391);
nand U24760 (N_24760,N_20478,N_20750);
nor U24761 (N_24761,N_21411,N_20995);
nand U24762 (N_24762,N_20396,N_21833);
nor U24763 (N_24763,N_22066,N_21327);
or U24764 (N_24764,N_22473,N_22067);
nand U24765 (N_24765,N_21456,N_21720);
xnor U24766 (N_24766,N_20367,N_21716);
xnor U24767 (N_24767,N_21996,N_22126);
nor U24768 (N_24768,N_20476,N_20979);
and U24769 (N_24769,N_20556,N_21077);
nor U24770 (N_24770,N_20714,N_21276);
nand U24771 (N_24771,N_21092,N_20879);
nor U24772 (N_24772,N_20517,N_22326);
and U24773 (N_24773,N_22409,N_21444);
or U24774 (N_24774,N_21384,N_20616);
xnor U24775 (N_24775,N_20738,N_20718);
nor U24776 (N_24776,N_20924,N_21480);
and U24777 (N_24777,N_20608,N_20075);
nor U24778 (N_24778,N_20661,N_20879);
nand U24779 (N_24779,N_20045,N_21574);
or U24780 (N_24780,N_20041,N_20417);
or U24781 (N_24781,N_22495,N_20993);
and U24782 (N_24782,N_21068,N_20494);
and U24783 (N_24783,N_22472,N_21711);
nand U24784 (N_24784,N_20068,N_21842);
nand U24785 (N_24785,N_20984,N_22353);
and U24786 (N_24786,N_20283,N_20255);
and U24787 (N_24787,N_20768,N_21739);
or U24788 (N_24788,N_20410,N_20766);
xnor U24789 (N_24789,N_22041,N_22019);
nand U24790 (N_24790,N_22215,N_21937);
or U24791 (N_24791,N_20323,N_22094);
xnor U24792 (N_24792,N_22256,N_21071);
nand U24793 (N_24793,N_22361,N_21413);
xnor U24794 (N_24794,N_21655,N_21051);
xnor U24795 (N_24795,N_20670,N_20495);
nor U24796 (N_24796,N_20853,N_21490);
xor U24797 (N_24797,N_21831,N_20902);
nand U24798 (N_24798,N_21255,N_22355);
xnor U24799 (N_24799,N_20246,N_22459);
xor U24800 (N_24800,N_21900,N_21134);
xor U24801 (N_24801,N_20483,N_21308);
and U24802 (N_24802,N_22100,N_21904);
nor U24803 (N_24803,N_21803,N_20633);
and U24804 (N_24804,N_22304,N_21379);
nor U24805 (N_24805,N_22093,N_21876);
and U24806 (N_24806,N_21168,N_21497);
xor U24807 (N_24807,N_21344,N_20462);
nor U24808 (N_24808,N_21141,N_20086);
nor U24809 (N_24809,N_20886,N_20701);
xnor U24810 (N_24810,N_21488,N_21973);
and U24811 (N_24811,N_22261,N_20846);
or U24812 (N_24812,N_21199,N_22471);
nand U24813 (N_24813,N_21296,N_20964);
nand U24814 (N_24814,N_21554,N_20234);
and U24815 (N_24815,N_20379,N_20381);
xnor U24816 (N_24816,N_21079,N_22236);
and U24817 (N_24817,N_21148,N_21304);
xnor U24818 (N_24818,N_21708,N_22388);
or U24819 (N_24819,N_21382,N_20775);
and U24820 (N_24820,N_20660,N_21268);
nor U24821 (N_24821,N_21303,N_21965);
nand U24822 (N_24822,N_22144,N_21133);
and U24823 (N_24823,N_20284,N_21974);
xnor U24824 (N_24824,N_21171,N_21403);
or U24825 (N_24825,N_20136,N_21498);
or U24826 (N_24826,N_21705,N_22336);
or U24827 (N_24827,N_20315,N_21210);
xnor U24828 (N_24828,N_21983,N_22102);
xnor U24829 (N_24829,N_21318,N_22118);
nand U24830 (N_24830,N_22287,N_20253);
xor U24831 (N_24831,N_20805,N_20309);
nand U24832 (N_24832,N_20839,N_20427);
and U24833 (N_24833,N_20775,N_21517);
nor U24834 (N_24834,N_20387,N_22312);
xor U24835 (N_24835,N_22025,N_20570);
nor U24836 (N_24836,N_21145,N_20007);
xnor U24837 (N_24837,N_20386,N_21335);
and U24838 (N_24838,N_22396,N_20544);
or U24839 (N_24839,N_21290,N_20659);
xor U24840 (N_24840,N_22093,N_20451);
nand U24841 (N_24841,N_20277,N_22040);
xnor U24842 (N_24842,N_22289,N_21454);
nand U24843 (N_24843,N_21168,N_21850);
nor U24844 (N_24844,N_20023,N_21550);
nor U24845 (N_24845,N_21472,N_20922);
nor U24846 (N_24846,N_20906,N_21879);
and U24847 (N_24847,N_22352,N_21556);
xor U24848 (N_24848,N_21497,N_21334);
xor U24849 (N_24849,N_22427,N_20740);
xor U24850 (N_24850,N_22236,N_22266);
or U24851 (N_24851,N_22411,N_22326);
xnor U24852 (N_24852,N_20883,N_21377);
xnor U24853 (N_24853,N_20018,N_21829);
nor U24854 (N_24854,N_20752,N_20229);
xor U24855 (N_24855,N_20279,N_21401);
and U24856 (N_24856,N_21565,N_22373);
and U24857 (N_24857,N_20448,N_20938);
or U24858 (N_24858,N_20037,N_22407);
nor U24859 (N_24859,N_20041,N_22479);
nor U24860 (N_24860,N_22158,N_22352);
or U24861 (N_24861,N_21858,N_20374);
nand U24862 (N_24862,N_20907,N_20998);
or U24863 (N_24863,N_20030,N_22260);
xor U24864 (N_24864,N_20677,N_20900);
or U24865 (N_24865,N_21445,N_22222);
or U24866 (N_24866,N_22257,N_21141);
xor U24867 (N_24867,N_20553,N_20665);
nand U24868 (N_24868,N_21558,N_22020);
or U24869 (N_24869,N_21568,N_20724);
nor U24870 (N_24870,N_21207,N_20533);
nor U24871 (N_24871,N_20135,N_20080);
xor U24872 (N_24872,N_22130,N_21343);
or U24873 (N_24873,N_20661,N_22116);
xor U24874 (N_24874,N_22001,N_21869);
xnor U24875 (N_24875,N_22450,N_20620);
nor U24876 (N_24876,N_21954,N_21098);
and U24877 (N_24877,N_20572,N_20384);
nor U24878 (N_24878,N_21233,N_20662);
nor U24879 (N_24879,N_21050,N_22238);
or U24880 (N_24880,N_20297,N_21723);
nor U24881 (N_24881,N_20259,N_20852);
and U24882 (N_24882,N_20035,N_22361);
nor U24883 (N_24883,N_21928,N_21136);
and U24884 (N_24884,N_20974,N_20066);
xnor U24885 (N_24885,N_20512,N_20515);
nor U24886 (N_24886,N_20128,N_20803);
or U24887 (N_24887,N_21974,N_21985);
or U24888 (N_24888,N_20360,N_22327);
xnor U24889 (N_24889,N_20638,N_21806);
nand U24890 (N_24890,N_20182,N_22124);
nor U24891 (N_24891,N_22413,N_21844);
nor U24892 (N_24892,N_21143,N_21195);
or U24893 (N_24893,N_20665,N_20397);
nor U24894 (N_24894,N_20960,N_20003);
nor U24895 (N_24895,N_20672,N_21537);
nand U24896 (N_24896,N_21553,N_20240);
or U24897 (N_24897,N_20809,N_21454);
nor U24898 (N_24898,N_21669,N_20130);
nand U24899 (N_24899,N_22033,N_21618);
xor U24900 (N_24900,N_22124,N_21505);
or U24901 (N_24901,N_21485,N_22266);
and U24902 (N_24902,N_22414,N_20324);
and U24903 (N_24903,N_21159,N_22196);
nand U24904 (N_24904,N_20053,N_22229);
and U24905 (N_24905,N_21105,N_20899);
nand U24906 (N_24906,N_21983,N_20066);
or U24907 (N_24907,N_21690,N_20149);
or U24908 (N_24908,N_22343,N_21220);
nor U24909 (N_24909,N_21189,N_21373);
nor U24910 (N_24910,N_20764,N_20895);
nand U24911 (N_24911,N_21134,N_21282);
or U24912 (N_24912,N_20758,N_20505);
nand U24913 (N_24913,N_20532,N_20351);
or U24914 (N_24914,N_21076,N_20044);
nor U24915 (N_24915,N_21858,N_20726);
xnor U24916 (N_24916,N_20053,N_20020);
xor U24917 (N_24917,N_21802,N_20731);
or U24918 (N_24918,N_22443,N_21271);
and U24919 (N_24919,N_21777,N_21928);
and U24920 (N_24920,N_20953,N_22116);
and U24921 (N_24921,N_20620,N_21820);
xor U24922 (N_24922,N_21473,N_20433);
and U24923 (N_24923,N_21008,N_21305);
xor U24924 (N_24924,N_20170,N_21321);
nand U24925 (N_24925,N_22116,N_22451);
nand U24926 (N_24926,N_21813,N_20388);
nor U24927 (N_24927,N_20470,N_21177);
nor U24928 (N_24928,N_21887,N_21127);
or U24929 (N_24929,N_21296,N_20496);
nand U24930 (N_24930,N_20842,N_20444);
nor U24931 (N_24931,N_21856,N_20246);
nand U24932 (N_24932,N_20176,N_20392);
or U24933 (N_24933,N_21027,N_21157);
nor U24934 (N_24934,N_21628,N_21771);
or U24935 (N_24935,N_21914,N_21002);
xor U24936 (N_24936,N_20352,N_21899);
and U24937 (N_24937,N_21700,N_21170);
nor U24938 (N_24938,N_20507,N_20776);
nand U24939 (N_24939,N_22106,N_20440);
nand U24940 (N_24940,N_20564,N_21856);
xor U24941 (N_24941,N_20492,N_21348);
or U24942 (N_24942,N_21068,N_22273);
and U24943 (N_24943,N_21387,N_21946);
and U24944 (N_24944,N_21269,N_20654);
and U24945 (N_24945,N_21427,N_21663);
nor U24946 (N_24946,N_20426,N_20208);
nand U24947 (N_24947,N_21952,N_21135);
or U24948 (N_24948,N_20161,N_20864);
or U24949 (N_24949,N_20575,N_21879);
and U24950 (N_24950,N_21799,N_22240);
nand U24951 (N_24951,N_20759,N_21200);
or U24952 (N_24952,N_20152,N_21480);
and U24953 (N_24953,N_22137,N_20768);
nor U24954 (N_24954,N_21846,N_22081);
xnor U24955 (N_24955,N_22145,N_20188);
xor U24956 (N_24956,N_20193,N_21912);
and U24957 (N_24957,N_21194,N_22312);
nand U24958 (N_24958,N_22341,N_22405);
xnor U24959 (N_24959,N_21556,N_21413);
xor U24960 (N_24960,N_22240,N_20067);
or U24961 (N_24961,N_21647,N_21338);
and U24962 (N_24962,N_21880,N_21753);
nor U24963 (N_24963,N_21211,N_21827);
or U24964 (N_24964,N_21427,N_22314);
or U24965 (N_24965,N_20726,N_22215);
and U24966 (N_24966,N_20180,N_20503);
or U24967 (N_24967,N_20431,N_21431);
or U24968 (N_24968,N_20865,N_22397);
nand U24969 (N_24969,N_20222,N_22445);
and U24970 (N_24970,N_20809,N_21195);
xor U24971 (N_24971,N_21818,N_20630);
nor U24972 (N_24972,N_21117,N_20606);
and U24973 (N_24973,N_20864,N_21530);
nor U24974 (N_24974,N_21751,N_20110);
nor U24975 (N_24975,N_22298,N_21038);
or U24976 (N_24976,N_21576,N_22089);
nor U24977 (N_24977,N_20514,N_20015);
and U24978 (N_24978,N_20347,N_21171);
xor U24979 (N_24979,N_20435,N_20943);
xor U24980 (N_24980,N_20417,N_22238);
nand U24981 (N_24981,N_20836,N_21162);
or U24982 (N_24982,N_21152,N_22345);
nand U24983 (N_24983,N_20977,N_21904);
nor U24984 (N_24984,N_21872,N_22273);
xnor U24985 (N_24985,N_20023,N_20855);
nor U24986 (N_24986,N_20590,N_21083);
and U24987 (N_24987,N_21023,N_20215);
or U24988 (N_24988,N_22253,N_21146);
xor U24989 (N_24989,N_22106,N_20549);
nor U24990 (N_24990,N_22496,N_20301);
nor U24991 (N_24991,N_22472,N_20218);
xor U24992 (N_24992,N_22264,N_21647);
or U24993 (N_24993,N_22268,N_21871);
nand U24994 (N_24994,N_21424,N_20131);
nor U24995 (N_24995,N_20850,N_21893);
and U24996 (N_24996,N_20622,N_21674);
and U24997 (N_24997,N_20697,N_21302);
and U24998 (N_24998,N_20881,N_20408);
nand U24999 (N_24999,N_21814,N_20050);
nand UO_0 (O_0,N_23770,N_24377);
nor UO_1 (O_1,N_23856,N_23278);
nand UO_2 (O_2,N_24344,N_23103);
nand UO_3 (O_3,N_22823,N_23041);
or UO_4 (O_4,N_23849,N_23197);
and UO_5 (O_5,N_23642,N_22624);
xnor UO_6 (O_6,N_24396,N_23218);
nor UO_7 (O_7,N_24689,N_23579);
xnor UO_8 (O_8,N_23824,N_24244);
xnor UO_9 (O_9,N_24728,N_23787);
nor UO_10 (O_10,N_23006,N_23040);
xnor UO_11 (O_11,N_23811,N_23998);
or UO_12 (O_12,N_23556,N_23424);
xor UO_13 (O_13,N_23241,N_23349);
xnor UO_14 (O_14,N_24658,N_23653);
and UO_15 (O_15,N_24670,N_23479);
or UO_16 (O_16,N_23359,N_23171);
nand UO_17 (O_17,N_23011,N_24767);
nor UO_18 (O_18,N_22978,N_23298);
xor UO_19 (O_19,N_23082,N_22924);
or UO_20 (O_20,N_24167,N_23932);
xor UO_21 (O_21,N_24856,N_24332);
nor UO_22 (O_22,N_24092,N_24574);
and UO_23 (O_23,N_22903,N_23522);
nor UO_24 (O_24,N_24623,N_23220);
nand UO_25 (O_25,N_22586,N_22791);
xnor UO_26 (O_26,N_24541,N_24605);
xnor UO_27 (O_27,N_22936,N_24366);
xnor UO_28 (O_28,N_22737,N_23416);
or UO_29 (O_29,N_23099,N_24241);
nand UO_30 (O_30,N_23555,N_23979);
xnor UO_31 (O_31,N_24812,N_23108);
and UO_32 (O_32,N_24188,N_23543);
nor UO_33 (O_33,N_24341,N_23832);
xor UO_34 (O_34,N_24773,N_23509);
or UO_35 (O_35,N_24679,N_24888);
and UO_36 (O_36,N_23842,N_24403);
or UO_37 (O_37,N_23230,N_24229);
or UO_38 (O_38,N_24149,N_24480);
and UO_39 (O_39,N_23274,N_24277);
nand UO_40 (O_40,N_24998,N_23153);
and UO_41 (O_41,N_23833,N_24506);
nor UO_42 (O_42,N_23978,N_23352);
or UO_43 (O_43,N_22644,N_23635);
and UO_44 (O_44,N_22617,N_23880);
and UO_45 (O_45,N_24422,N_23384);
and UO_46 (O_46,N_22975,N_24462);
xnor UO_47 (O_47,N_24004,N_24761);
xnor UO_48 (O_48,N_23098,N_24395);
or UO_49 (O_49,N_24068,N_24599);
and UO_50 (O_50,N_24710,N_24905);
or UO_51 (O_51,N_23261,N_22837);
and UO_52 (O_52,N_23752,N_24939);
and UO_53 (O_53,N_24521,N_23378);
nor UO_54 (O_54,N_22935,N_24629);
and UO_55 (O_55,N_22818,N_23212);
nor UO_56 (O_56,N_23367,N_23091);
and UO_57 (O_57,N_22859,N_24170);
nand UO_58 (O_58,N_23597,N_22509);
xnor UO_59 (O_59,N_22807,N_24391);
nand UO_60 (O_60,N_24006,N_23994);
xnor UO_61 (O_61,N_24460,N_22681);
and UO_62 (O_62,N_23004,N_24636);
nand UO_63 (O_63,N_24774,N_23682);
and UO_64 (O_64,N_23474,N_23810);
nand UO_65 (O_65,N_24001,N_24340);
and UO_66 (O_66,N_23596,N_24483);
xor UO_67 (O_67,N_24284,N_22609);
or UO_68 (O_68,N_23411,N_23694);
nor UO_69 (O_69,N_24858,N_22566);
or UO_70 (O_70,N_24977,N_23496);
nor UO_71 (O_71,N_24876,N_23264);
nand UO_72 (O_72,N_23311,N_24474);
nor UO_73 (O_73,N_22684,N_23090);
nand UO_74 (O_74,N_23183,N_23545);
xor UO_75 (O_75,N_23105,N_23174);
nor UO_76 (O_76,N_24989,N_23113);
nand UO_77 (O_77,N_23990,N_22635);
and UO_78 (O_78,N_23354,N_22941);
and UO_79 (O_79,N_24193,N_24999);
xnor UO_80 (O_80,N_23506,N_22541);
and UO_81 (O_81,N_22694,N_24690);
or UO_82 (O_82,N_24975,N_23460);
or UO_83 (O_83,N_23982,N_22639);
or UO_84 (O_84,N_24631,N_24606);
nand UO_85 (O_85,N_24920,N_23455);
and UO_86 (O_86,N_23695,N_23085);
nand UO_87 (O_87,N_22579,N_22551);
and UO_88 (O_88,N_24681,N_23343);
nor UO_89 (O_89,N_22977,N_23494);
nor UO_90 (O_90,N_22567,N_24881);
or UO_91 (O_91,N_24090,N_22890);
and UO_92 (O_92,N_22649,N_23247);
or UO_93 (O_93,N_24398,N_24443);
nor UO_94 (O_94,N_24890,N_22519);
nor UO_95 (O_95,N_22795,N_22862);
nor UO_96 (O_96,N_23737,N_24650);
nand UO_97 (O_97,N_22674,N_22619);
and UO_98 (O_98,N_22904,N_23609);
nand UO_99 (O_99,N_23818,N_24447);
xnor UO_100 (O_100,N_24732,N_22664);
nor UO_101 (O_101,N_23662,N_23145);
or UO_102 (O_102,N_22683,N_23129);
nand UO_103 (O_103,N_23079,N_23563);
xor UO_104 (O_104,N_22638,N_23876);
and UO_105 (O_105,N_24757,N_24417);
xor UO_106 (O_106,N_23947,N_23054);
nand UO_107 (O_107,N_23371,N_23203);
and UO_108 (O_108,N_24694,N_23143);
or UO_109 (O_109,N_24766,N_24855);
or UO_110 (O_110,N_23330,N_24162);
xnor UO_111 (O_111,N_22958,N_23120);
or UO_112 (O_112,N_24067,N_23826);
and UO_113 (O_113,N_23659,N_23062);
nand UO_114 (O_114,N_24116,N_22914);
and UO_115 (O_115,N_23589,N_24972);
nand UO_116 (O_116,N_23528,N_24568);
and UO_117 (O_117,N_22938,N_22558);
or UO_118 (O_118,N_22928,N_23484);
nor UO_119 (O_119,N_22946,N_23841);
xor UO_120 (O_120,N_22610,N_23689);
nand UO_121 (O_121,N_22532,N_23732);
nand UO_122 (O_122,N_23630,N_24492);
and UO_123 (O_123,N_22881,N_23946);
or UO_124 (O_124,N_23191,N_24719);
nand UO_125 (O_125,N_24850,N_24826);
nor UO_126 (O_126,N_22848,N_24497);
or UO_127 (O_127,N_23291,N_24263);
xnor UO_128 (O_128,N_24563,N_22725);
nor UO_129 (O_129,N_24079,N_22696);
nand UO_130 (O_130,N_23450,N_23179);
nand UO_131 (O_131,N_23785,N_24820);
and UO_132 (O_132,N_23781,N_24020);
xnor UO_133 (O_133,N_23290,N_22648);
and UO_134 (O_134,N_24307,N_23008);
or UO_135 (O_135,N_22621,N_23444);
and UO_136 (O_136,N_24048,N_22962);
and UO_137 (O_137,N_23495,N_23933);
xnor UO_138 (O_138,N_22563,N_23764);
nand UO_139 (O_139,N_24660,N_23071);
nand UO_140 (O_140,N_24343,N_24313);
and UO_141 (O_141,N_24464,N_24893);
or UO_142 (O_142,N_24355,N_22597);
or UO_143 (O_143,N_22716,N_22929);
xnor UO_144 (O_144,N_22502,N_24583);
nor UO_145 (O_145,N_24573,N_24183);
and UO_146 (O_146,N_24723,N_22593);
xnor UO_147 (O_147,N_24538,N_23934);
nor UO_148 (O_148,N_24220,N_23139);
or UO_149 (O_149,N_24592,N_24873);
and UO_150 (O_150,N_22741,N_23049);
and UO_151 (O_151,N_23704,N_23156);
or UO_152 (O_152,N_23162,N_22671);
nand UO_153 (O_153,N_22759,N_23281);
xor UO_154 (O_154,N_23043,N_24647);
xor UO_155 (O_155,N_24037,N_22607);
or UO_156 (O_156,N_22965,N_23313);
or UO_157 (O_157,N_24379,N_22629);
xor UO_158 (O_158,N_23333,N_23688);
xnor UO_159 (O_159,N_22789,N_22806);
nor UO_160 (O_160,N_24708,N_23462);
nand UO_161 (O_161,N_24891,N_22829);
nand UO_162 (O_162,N_22544,N_24451);
xor UO_163 (O_163,N_22626,N_24080);
nor UO_164 (O_164,N_24010,N_23061);
and UO_165 (O_165,N_23692,N_24519);
xnor UO_166 (O_166,N_22940,N_24196);
and UO_167 (O_167,N_24936,N_24966);
and UO_168 (O_168,N_23756,N_23340);
xnor UO_169 (O_169,N_24834,N_22800);
or UO_170 (O_170,N_24027,N_22662);
or UO_171 (O_171,N_24946,N_23951);
nand UO_172 (O_172,N_23121,N_22745);
and UO_173 (O_173,N_24415,N_22944);
and UO_174 (O_174,N_22739,N_22992);
or UO_175 (O_175,N_24074,N_23211);
xor UO_176 (O_176,N_23564,N_24338);
nor UO_177 (O_177,N_22732,N_24018);
nor UO_178 (O_178,N_23167,N_23341);
nor UO_179 (O_179,N_24425,N_23257);
or UO_180 (O_180,N_24087,N_24522);
and UO_181 (O_181,N_24954,N_23468);
nand UO_182 (O_182,N_24853,N_23165);
or UO_183 (O_183,N_23164,N_23458);
or UO_184 (O_184,N_22836,N_24223);
nand UO_185 (O_185,N_23716,N_23332);
or UO_186 (O_186,N_23467,N_24556);
or UO_187 (O_187,N_24019,N_22699);
nor UO_188 (O_188,N_23489,N_24144);
xor UO_189 (O_189,N_23173,N_23652);
xor UO_190 (O_190,N_23956,N_22564);
nor UO_191 (O_191,N_23622,N_24476);
xor UO_192 (O_192,N_22604,N_24983);
or UO_193 (O_193,N_23913,N_23485);
nand UO_194 (O_194,N_24127,N_23339);
and UO_195 (O_195,N_24084,N_22568);
or UO_196 (O_196,N_22529,N_22548);
xor UO_197 (O_197,N_23205,N_23225);
and UO_198 (O_198,N_23393,N_24827);
nand UO_199 (O_199,N_23569,N_23063);
nor UO_200 (O_200,N_24300,N_23052);
nor UO_201 (O_201,N_23272,N_23927);
xor UO_202 (O_202,N_23314,N_23295);
nor UO_203 (O_203,N_22655,N_23745);
xnor UO_204 (O_204,N_22953,N_23287);
or UO_205 (O_205,N_22917,N_23395);
and UO_206 (O_206,N_23065,N_24712);
nand UO_207 (O_207,N_22501,N_24974);
or UO_208 (O_208,N_22679,N_23407);
xnor UO_209 (O_209,N_23426,N_24184);
nor UO_210 (O_210,N_23408,N_23806);
and UO_211 (O_211,N_22668,N_23971);
nor UO_212 (O_212,N_23730,N_23476);
and UO_213 (O_213,N_24158,N_23267);
nand UO_214 (O_214,N_24316,N_23862);
xor UO_215 (O_215,N_23464,N_23789);
nand UO_216 (O_216,N_23221,N_24166);
or UO_217 (O_217,N_24976,N_23375);
or UO_218 (O_218,N_23196,N_24231);
nand UO_219 (O_219,N_24691,N_24958);
nand UO_220 (O_220,N_23975,N_24380);
nor UO_221 (O_221,N_24400,N_23388);
or UO_222 (O_222,N_23723,N_23967);
nand UO_223 (O_223,N_24979,N_24782);
and UO_224 (O_224,N_23533,N_22792);
nor UO_225 (O_225,N_24202,N_22550);
and UO_226 (O_226,N_23326,N_24108);
and UO_227 (O_227,N_23850,N_23719);
or UO_228 (O_228,N_24580,N_22933);
and UO_229 (O_229,N_23970,N_24938);
and UO_230 (O_230,N_23707,N_24684);
and UO_231 (O_231,N_22991,N_22980);
or UO_232 (O_232,N_24654,N_23943);
nand UO_233 (O_233,N_23442,N_23751);
nand UO_234 (O_234,N_22738,N_24045);
and UO_235 (O_235,N_24327,N_23915);
xor UO_236 (O_236,N_24516,N_24866);
or UO_237 (O_237,N_24121,N_22869);
nor UO_238 (O_238,N_23318,N_24867);
xnor UO_239 (O_239,N_24981,N_24361);
nor UO_240 (O_240,N_23920,N_23319);
and UO_241 (O_241,N_23800,N_24887);
and UO_242 (O_242,N_23775,N_23557);
nand UO_243 (O_243,N_22811,N_23096);
xnor UO_244 (O_244,N_23023,N_23661);
or UO_245 (O_245,N_24000,N_23387);
or UO_246 (O_246,N_22750,N_23588);
and UO_247 (O_247,N_24402,N_23030);
xnor UO_248 (O_248,N_24477,N_23860);
or UO_249 (O_249,N_23537,N_24992);
or UO_250 (O_250,N_24478,N_22814);
or UO_251 (O_251,N_24346,N_23396);
or UO_252 (O_252,N_23398,N_22822);
nand UO_253 (O_253,N_24434,N_23586);
or UO_254 (O_254,N_23991,N_24830);
and UO_255 (O_255,N_23936,N_24482);
and UO_256 (O_256,N_23320,N_22802);
nand UO_257 (O_257,N_23536,N_23507);
nand UO_258 (O_258,N_24816,N_23151);
xor UO_259 (O_259,N_23392,N_23526);
and UO_260 (O_260,N_24256,N_22786);
xor UO_261 (O_261,N_22983,N_23422);
xnor UO_262 (O_262,N_24206,N_24135);
xnor UO_263 (O_263,N_23572,N_23500);
and UO_264 (O_264,N_23648,N_23779);
and UO_265 (O_265,N_23819,N_22594);
nand UO_266 (O_266,N_24214,N_23578);
or UO_267 (O_267,N_24302,N_24505);
and UO_268 (O_268,N_24960,N_24209);
nor UO_269 (O_269,N_22880,N_23149);
and UO_270 (O_270,N_22994,N_23198);
nor UO_271 (O_271,N_24248,N_24513);
nand UO_272 (O_272,N_23034,N_22600);
and UO_273 (O_273,N_24661,N_24065);
xnor UO_274 (O_274,N_23118,N_22727);
or UO_275 (O_275,N_24311,N_24738);
nor UO_276 (O_276,N_23406,N_24616);
and UO_277 (O_277,N_24584,N_23997);
or UO_278 (O_278,N_24445,N_24169);
or UO_279 (O_279,N_23187,N_24285);
nor UO_280 (O_280,N_24937,N_24755);
nor UO_281 (O_281,N_23604,N_22968);
nor UO_282 (O_282,N_24825,N_24034);
nand UO_283 (O_283,N_22539,N_24680);
xor UO_284 (O_284,N_24924,N_24515);
and UO_285 (O_285,N_24995,N_23611);
and UO_286 (O_286,N_24106,N_23836);
xor UO_287 (O_287,N_24228,N_24931);
xor UO_288 (O_288,N_22872,N_22740);
or UO_289 (O_289,N_24264,N_22522);
and UO_290 (O_290,N_23042,N_23448);
xor UO_291 (O_291,N_23447,N_23093);
nor UO_292 (O_292,N_23702,N_24002);
xor UO_293 (O_293,N_23577,N_23996);
nand UO_294 (O_294,N_23344,N_23914);
nor UO_295 (O_295,N_24315,N_24390);
or UO_296 (O_296,N_23571,N_23134);
and UO_297 (O_297,N_24435,N_24544);
or UO_298 (O_298,N_24458,N_23618);
nor UO_299 (O_299,N_24536,N_22653);
nor UO_300 (O_300,N_23415,N_24633);
or UO_301 (O_301,N_23879,N_23930);
nand UO_302 (O_302,N_23977,N_23993);
xor UO_303 (O_303,N_24734,N_23888);
nand UO_304 (O_304,N_24286,N_22521);
xor UO_305 (O_305,N_22752,N_22838);
xnor UO_306 (O_306,N_23954,N_24024);
nor UO_307 (O_307,N_24044,N_22860);
or UO_308 (O_308,N_24347,N_23686);
or UO_309 (O_309,N_23935,N_23399);
and UO_310 (O_310,N_23805,N_23923);
and UO_311 (O_311,N_22855,N_23172);
or UO_312 (O_312,N_24198,N_22794);
xor UO_313 (O_313,N_24383,N_23092);
nor UO_314 (O_314,N_23962,N_22678);
or UO_315 (O_315,N_23434,N_24810);
xnor UO_316 (O_316,N_23182,N_24288);
and UO_317 (O_317,N_24414,N_23358);
nand UO_318 (O_318,N_24789,N_22540);
nand UO_319 (O_319,N_22816,N_22996);
or UO_320 (O_320,N_22592,N_22570);
or UO_321 (O_321,N_23405,N_24225);
and UO_322 (O_322,N_23866,N_23275);
nand UO_323 (O_323,N_24570,N_24715);
nor UO_324 (O_324,N_24357,N_22585);
nand UO_325 (O_325,N_23132,N_23863);
nor UO_326 (O_326,N_22891,N_23992);
xor UO_327 (O_327,N_23282,N_23964);
nand UO_328 (O_328,N_24015,N_22731);
nor UO_329 (O_329,N_24275,N_24164);
or UO_330 (O_330,N_22711,N_24230);
or UO_331 (O_331,N_24746,N_23931);
nor UO_332 (O_332,N_23083,N_24870);
nand UO_333 (O_333,N_23871,N_23624);
nand UO_334 (O_334,N_23020,N_24322);
or UO_335 (O_335,N_24351,N_24781);
or UO_336 (O_336,N_24175,N_23246);
nand UO_337 (O_337,N_22784,N_24587);
xnor UO_338 (O_338,N_23877,N_22511);
nor UO_339 (O_339,N_24655,N_24649);
nor UO_340 (O_340,N_24103,N_24790);
or UO_341 (O_341,N_24571,N_22864);
nor UO_342 (O_342,N_24779,N_24449);
nand UO_343 (O_343,N_24145,N_24711);
nand UO_344 (O_344,N_23312,N_23503);
or UO_345 (O_345,N_24189,N_23763);
and UO_346 (O_346,N_24635,N_23657);
xnor UO_347 (O_347,N_23180,N_24008);
nand UO_348 (O_348,N_24486,N_23420);
nor UO_349 (O_349,N_22552,N_22921);
nor UO_350 (O_350,N_24261,N_22504);
nand UO_351 (O_351,N_22841,N_23905);
nand UO_352 (O_352,N_24013,N_23066);
xor UO_353 (O_353,N_22916,N_23908);
and UO_354 (O_354,N_22961,N_23687);
nand UO_355 (O_355,N_23893,N_23409);
nor UO_356 (O_356,N_23605,N_23838);
or UO_357 (O_357,N_24877,N_24806);
or UO_358 (O_358,N_24171,N_24575);
nor UO_359 (O_359,N_22850,N_24663);
nand UO_360 (O_360,N_22866,N_22553);
or UO_361 (O_361,N_23987,N_24671);
and UO_362 (O_362,N_24259,N_24055);
nor UO_363 (O_363,N_24572,N_23660);
and UO_364 (O_364,N_22754,N_24283);
nand UO_365 (O_365,N_22615,N_24542);
and UO_366 (O_366,N_24369,N_23304);
or UO_367 (O_367,N_22598,N_22700);
nand UO_368 (O_368,N_24303,N_24243);
nor UO_369 (O_369,N_24823,N_24182);
and UO_370 (O_370,N_24883,N_22643);
nand UO_371 (O_371,N_24266,N_24579);
nor UO_372 (O_372,N_24685,N_24569);
nor UO_373 (O_373,N_23360,N_24201);
and UO_374 (O_374,N_23874,N_22680);
nor UO_375 (O_375,N_24421,N_23427);
and UO_376 (O_376,N_23795,N_23302);
nor UO_377 (O_377,N_22882,N_24123);
and UO_378 (O_378,N_22858,N_22787);
nor UO_379 (O_379,N_23204,N_24620);
nand UO_380 (O_380,N_23046,N_22525);
nor UO_381 (O_381,N_22883,N_23729);
and UO_382 (O_382,N_23135,N_22561);
and UO_383 (O_383,N_24921,N_22954);
and UO_384 (O_384,N_22581,N_24385);
or UO_385 (O_385,N_23575,N_24423);
nor UO_386 (O_386,N_23086,N_23678);
and UO_387 (O_387,N_24107,N_23498);
nor UO_388 (O_388,N_24269,N_23133);
nor UO_389 (O_389,N_23804,N_24955);
xnor UO_390 (O_390,N_24951,N_23002);
or UO_391 (O_391,N_23338,N_23109);
nor UO_392 (O_392,N_24354,N_23827);
xor UO_393 (O_393,N_24485,N_22813);
xnor UO_394 (O_394,N_22950,N_24797);
xnor UO_395 (O_395,N_23847,N_23148);
or UO_396 (O_396,N_22575,N_23906);
and UO_397 (O_397,N_23194,N_22557);
or UO_398 (O_398,N_24762,N_22707);
nor UO_399 (O_399,N_24612,N_24317);
nor UO_400 (O_400,N_23403,N_22785);
or UO_401 (O_401,N_23346,N_24880);
nand UO_402 (O_402,N_23234,N_24701);
nor UO_403 (O_403,N_22960,N_24982);
nand UO_404 (O_404,N_23674,N_23268);
nand UO_405 (O_405,N_22934,N_24996);
nor UO_406 (O_406,N_23816,N_24526);
xnor UO_407 (O_407,N_23676,N_23757);
xnor UO_408 (O_408,N_23316,N_24438);
nor UO_409 (O_409,N_23336,N_24086);
and UO_410 (O_410,N_24114,N_23390);
nor UO_411 (O_411,N_22507,N_23525);
or UO_412 (O_412,N_23381,N_22761);
or UO_413 (O_413,N_23620,N_23834);
and UO_414 (O_414,N_22966,N_23155);
and UO_415 (O_415,N_24586,N_24078);
nor UO_416 (O_416,N_24021,N_24441);
or UO_417 (O_417,N_24785,N_24987);
nor UO_418 (O_418,N_24181,N_23169);
nand UO_419 (O_419,N_23175,N_24707);
nor UO_420 (O_420,N_24993,N_23972);
or UO_421 (O_421,N_23273,N_23839);
nor UO_422 (O_422,N_23513,N_23848);
and UO_423 (O_423,N_24963,N_22835);
xor UO_424 (O_424,N_23025,N_23514);
nand UO_425 (O_425,N_23955,N_24662);
xnor UO_426 (O_426,N_24499,N_22777);
or UO_427 (O_427,N_24838,N_24319);
and UO_428 (O_428,N_24949,N_24057);
nand UO_429 (O_429,N_22815,N_24363);
and UO_430 (O_430,N_24187,N_24942);
and UO_431 (O_431,N_24430,N_23735);
and UO_432 (O_432,N_23315,N_22780);
nor UO_433 (O_433,N_23331,N_22714);
or UO_434 (O_434,N_23033,N_23741);
and UO_435 (O_435,N_23902,N_24540);
nand UO_436 (O_436,N_24058,N_23727);
xor UO_437 (O_437,N_24863,N_24336);
and UO_438 (O_438,N_23961,N_24023);
or UO_439 (O_439,N_22849,N_24577);
or UO_440 (O_440,N_22827,N_22969);
nand UO_441 (O_441,N_23433,N_24677);
or UO_442 (O_442,N_24743,N_23058);
and UO_443 (O_443,N_22695,N_23898);
nand UO_444 (O_444,N_24518,N_24788);
and UO_445 (O_445,N_22633,N_24535);
and UO_446 (O_446,N_23413,N_22863);
xor UO_447 (O_447,N_22620,N_24155);
and UO_448 (O_448,N_24576,N_24604);
and UO_449 (O_449,N_23711,N_23665);
nor UO_450 (O_450,N_23709,N_24444);
and UO_451 (O_451,N_23361,N_24043);
nand UO_452 (O_452,N_22893,N_22717);
or UO_453 (O_453,N_24919,N_23168);
xnor UO_454 (O_454,N_24598,N_24875);
xnor UO_455 (O_455,N_23896,N_23457);
xor UO_456 (O_456,N_23808,N_24927);
or UO_457 (O_457,N_23483,N_23591);
or UO_458 (O_458,N_24765,N_23101);
or UO_459 (O_459,N_23492,N_23250);
and UO_460 (O_460,N_22758,N_23161);
nand UO_461 (O_461,N_23843,N_22907);
nand UO_462 (O_462,N_24173,N_24520);
or UO_463 (O_463,N_24213,N_23201);
xor UO_464 (O_464,N_23032,N_23292);
nand UO_465 (O_465,N_22673,N_23724);
xnor UO_466 (O_466,N_23229,N_22796);
xor UO_467 (O_467,N_24308,N_23215);
nor UO_468 (O_468,N_24368,N_24532);
nand UO_469 (O_469,N_23088,N_24097);
nor UO_470 (O_470,N_23505,N_24190);
and UO_471 (O_471,N_24846,N_24533);
xor UO_472 (O_472,N_24388,N_22772);
nand UO_473 (O_473,N_22832,N_22797);
and UO_474 (O_474,N_24410,N_23573);
and UO_475 (O_475,N_22756,N_24642);
and UO_476 (O_476,N_23718,N_22747);
and UO_477 (O_477,N_24272,N_23114);
nor UO_478 (O_478,N_22920,N_24722);
and UO_479 (O_479,N_23015,N_23431);
nor UO_480 (O_480,N_22526,N_23750);
nor UO_481 (O_481,N_24896,N_22776);
nand UO_482 (O_482,N_23176,N_24622);
nor UO_483 (O_483,N_23562,N_23646);
nor UO_484 (O_484,N_24778,N_22595);
nand UO_485 (O_485,N_23232,N_24617);
nand UO_486 (O_486,N_23958,N_23253);
or UO_487 (O_487,N_23631,N_22778);
nor UO_488 (O_488,N_24626,N_23645);
and UO_489 (O_489,N_24236,N_22712);
xnor UO_490 (O_490,N_23073,N_24066);
and UO_491 (O_491,N_23087,N_24412);
or UO_492 (O_492,N_23080,N_23369);
nor UO_493 (O_493,N_22757,N_23502);
nand UO_494 (O_494,N_24122,N_24358);
or UO_495 (O_495,N_23809,N_23216);
and UO_496 (O_496,N_22908,N_24798);
nor UO_497 (O_497,N_22697,N_24208);
nor UO_498 (O_498,N_24038,N_24433);
xnor UO_499 (O_499,N_23649,N_24833);
nor UO_500 (O_500,N_24278,N_23837);
xnor UO_501 (O_501,N_23929,N_23158);
nand UO_502 (O_502,N_23580,N_24212);
and UO_503 (O_503,N_24558,N_22985);
or UO_504 (O_504,N_24291,N_22826);
nand UO_505 (O_505,N_22533,N_24716);
and UO_506 (O_506,N_24686,N_23710);
nand UO_507 (O_507,N_24648,N_22582);
nand UO_508 (O_508,N_24903,N_24758);
nand UO_509 (O_509,N_22952,N_24967);
nand UO_510 (O_510,N_22942,N_24393);
and UO_511 (O_511,N_23026,N_23259);
nand UO_512 (O_512,N_23891,N_24935);
or UO_513 (O_513,N_24703,N_23650);
or UO_514 (O_514,N_24036,N_23345);
or UO_515 (O_515,N_23651,N_23031);
nand UO_516 (O_516,N_24783,N_23401);
or UO_517 (O_517,N_23470,N_23598);
or UO_518 (O_518,N_24726,N_23235);
nor UO_519 (O_519,N_23869,N_24900);
and UO_520 (O_520,N_22972,N_23984);
nor UO_521 (O_521,N_24384,N_23739);
or UO_522 (O_522,N_23391,N_23705);
nor UO_523 (O_523,N_22693,N_24721);
nor UO_524 (O_524,N_24298,N_24469);
nand UO_525 (O_525,N_24280,N_23747);
xnor UO_526 (O_526,N_24968,N_24934);
and UO_527 (O_527,N_24795,N_23497);
and UO_528 (O_528,N_24442,N_24320);
nor UO_529 (O_529,N_23262,N_24374);
xnor UO_530 (O_530,N_24614,N_22669);
and UO_531 (O_531,N_24709,N_23112);
or UO_532 (O_532,N_24233,N_24751);
or UO_533 (O_533,N_22889,N_23632);
or UO_534 (O_534,N_22887,N_23472);
or UO_535 (O_535,N_24871,N_23144);
nor UO_536 (O_536,N_24537,N_22899);
and UO_537 (O_537,N_24821,N_23084);
nand UO_538 (O_538,N_24744,N_23224);
nand UO_539 (O_539,N_23919,N_22765);
or UO_540 (O_540,N_24401,N_23067);
nor UO_541 (O_541,N_24985,N_23193);
nor UO_542 (O_542,N_23097,N_23553);
xnor UO_543 (O_543,N_22622,N_24892);
xnor UO_544 (O_544,N_24644,N_24052);
and UO_545 (O_545,N_23603,N_24672);
xor UO_546 (O_546,N_23774,N_23949);
nor UO_547 (O_547,N_23491,N_23535);
xnor UO_548 (O_548,N_22660,N_22516);
nor UO_549 (O_549,N_24050,N_24547);
nor UO_550 (O_550,N_22506,N_23542);
or UO_551 (O_551,N_22995,N_22825);
xnor UO_552 (O_552,N_23177,N_23122);
nand UO_553 (O_553,N_23188,N_23094);
or UO_554 (O_554,N_23321,N_23452);
nand UO_555 (O_555,N_24367,N_22583);
nand UO_556 (O_556,N_24695,N_23960);
or UO_557 (O_557,N_24740,N_24091);
xnor UO_558 (O_558,N_23899,N_24796);
and UO_559 (O_559,N_24141,N_23897);
and UO_560 (O_560,N_24119,N_23515);
nand UO_561 (O_561,N_24407,N_23146);
nor UO_562 (O_562,N_23907,N_24382);
nand UO_563 (O_563,N_22744,N_24026);
nor UO_564 (O_564,N_24450,N_23223);
nand UO_565 (O_565,N_23310,N_24907);
or UO_566 (O_566,N_24980,N_22888);
nor UO_567 (O_567,N_23035,N_24468);
and UO_568 (O_568,N_23377,N_23477);
nor UO_569 (O_569,N_23803,N_24714);
and UO_570 (O_570,N_22868,N_24697);
and UO_571 (O_571,N_23019,N_22923);
nor UO_572 (O_572,N_24372,N_23673);
and UO_573 (O_573,N_22790,N_23892);
nand UO_574 (O_574,N_24754,N_23983);
nor UO_575 (O_575,N_24780,N_24845);
nor UO_576 (O_576,N_23296,N_22951);
and UO_577 (O_577,N_24392,N_24353);
and UO_578 (O_578,N_22735,N_22879);
nand UO_579 (O_579,N_23001,N_23743);
nand UO_580 (O_580,N_22931,N_22805);
nand UO_581 (O_581,N_24705,N_23758);
or UO_582 (O_582,N_22909,N_23095);
and UO_583 (O_583,N_22748,N_22867);
nor UO_584 (O_584,N_22876,N_24249);
xor UO_585 (O_585,N_23668,N_23059);
nor UO_586 (O_586,N_24242,N_23070);
or UO_587 (O_587,N_24828,N_24111);
nand UO_588 (O_588,N_22554,N_24381);
nand UO_589 (O_589,N_23851,N_23547);
or UO_590 (O_590,N_23701,N_24739);
and UO_591 (O_591,N_23768,N_23853);
nand UO_592 (O_592,N_23950,N_23685);
xor UO_593 (O_593,N_23374,N_22718);
xor UO_594 (O_594,N_23742,N_24318);
nand UO_595 (O_595,N_22763,N_22611);
or UO_596 (O_596,N_23921,N_22625);
xor UO_597 (O_597,N_23269,N_23844);
and UO_598 (O_598,N_24467,N_24759);
or UO_599 (O_599,N_22537,N_24459);
xor UO_600 (O_600,N_24096,N_23952);
xnor UO_601 (O_601,N_22779,N_23623);
nor UO_602 (O_602,N_24800,N_23255);
and UO_603 (O_603,N_22808,N_24262);
xnor UO_604 (O_604,N_22656,N_23213);
nand UO_605 (O_605,N_22781,N_24165);
nor UO_606 (O_606,N_24325,N_24137);
xnor UO_607 (O_607,N_24267,N_22569);
and UO_608 (O_608,N_23446,N_22602);
and UO_609 (O_609,N_23738,N_22710);
and UO_610 (O_610,N_22746,N_23550);
and UO_611 (O_611,N_23802,N_23807);
and UO_612 (O_612,N_24088,N_22896);
or UO_613 (O_613,N_24056,N_23000);
xnor UO_614 (O_614,N_23696,N_24994);
or UO_615 (O_615,N_24502,N_23428);
nand UO_616 (O_616,N_24548,N_23538);
or UO_617 (O_617,N_24257,N_23968);
xor UO_618 (O_618,N_22831,N_23325);
and UO_619 (O_619,N_22877,N_23190);
nor UO_620 (O_620,N_24582,N_24207);
and UO_621 (O_621,N_24912,N_24488);
and UO_622 (O_622,N_24546,N_24003);
nor UO_623 (O_623,N_24869,N_22675);
or UO_624 (O_624,N_24424,N_24473);
nand UO_625 (O_625,N_24105,N_22902);
or UO_626 (O_626,N_23508,N_23466);
xnor UO_627 (O_627,N_24523,N_22535);
xor UO_628 (O_628,N_23684,N_23568);
nor UO_629 (O_629,N_23610,N_23909);
nand UO_630 (O_630,N_22599,N_23691);
or UO_631 (O_631,N_23429,N_24894);
nor UO_632 (O_632,N_23671,N_24857);
nand UO_633 (O_633,N_22546,N_24882);
xnor UO_634 (O_634,N_24926,N_23233);
or UO_635 (O_635,N_24948,N_23865);
nor UO_636 (O_636,N_23022,N_23587);
nand UO_637 (O_637,N_24032,N_23613);
and UO_638 (O_638,N_22628,N_22528);
and UO_639 (O_639,N_23355,N_24060);
xor UO_640 (O_640,N_23380,N_22783);
and UO_641 (O_641,N_22724,N_23731);
nand UO_642 (O_642,N_24925,N_23207);
and UO_643 (O_643,N_23890,N_23773);
and UO_644 (O_644,N_23252,N_23534);
or UO_645 (O_645,N_23048,N_23106);
nor UO_646 (O_646,N_24791,N_24693);
nor UO_647 (O_647,N_24234,N_24487);
or UO_648 (O_648,N_23142,N_23111);
or UO_649 (O_649,N_24072,N_24222);
xor UO_650 (O_650,N_23130,N_23616);
and UO_651 (O_651,N_24504,N_24534);
nand UO_652 (O_652,N_23110,N_24470);
and UO_653 (O_653,N_23038,N_24495);
or UO_654 (O_654,N_22726,N_22665);
or UO_655 (O_655,N_24841,N_24324);
or UO_656 (O_656,N_23518,N_23200);
and UO_657 (O_657,N_22865,N_24501);
or UO_658 (O_658,N_24033,N_23353);
xnor UO_659 (O_659,N_22556,N_22852);
nand UO_660 (O_660,N_24988,N_23647);
nand UO_661 (O_661,N_23459,N_23107);
or UO_662 (O_662,N_23576,N_24039);
xnor UO_663 (O_663,N_23208,N_23337);
nor UO_664 (O_664,N_24205,N_24772);
or UO_665 (O_665,N_24260,N_22703);
nor UO_666 (O_666,N_22733,N_24294);
nand UO_667 (O_667,N_23771,N_22676);
and UO_668 (O_668,N_22720,N_24352);
and UO_669 (O_669,N_23131,N_22809);
nand UO_670 (O_670,N_22884,N_23516);
nor UO_671 (O_671,N_22913,N_22686);
xor UO_672 (O_672,N_23733,N_22774);
or UO_673 (O_673,N_24930,N_24130);
and UO_674 (O_674,N_22512,N_24717);
and UO_675 (O_675,N_23565,N_22788);
nor UO_676 (O_676,N_23840,N_22947);
and UO_677 (O_677,N_22998,N_23527);
nor UO_678 (O_678,N_24192,N_24878);
and UO_679 (O_679,N_22565,N_24077);
xnor UO_680 (O_680,N_23210,N_24142);
nand UO_681 (O_681,N_24132,N_24978);
and UO_682 (O_682,N_24418,N_23926);
nand UO_683 (O_683,N_23895,N_24042);
nor UO_684 (O_684,N_22630,N_22721);
nor UO_685 (O_685,N_23055,N_22659);
or UO_686 (O_686,N_23297,N_23010);
and UO_687 (O_687,N_24140,N_24297);
and UO_688 (O_688,N_24879,N_22873);
nand UO_689 (O_689,N_24564,N_23417);
and UO_690 (O_690,N_24131,N_24808);
nand UO_691 (O_691,N_24742,N_22989);
and UO_692 (O_692,N_24652,N_24238);
and UO_693 (O_693,N_22894,N_22736);
nand UO_694 (O_694,N_22905,N_24735);
nand UO_695 (O_695,N_24157,N_24562);
nor UO_696 (O_696,N_24898,N_23617);
xor UO_697 (O_697,N_23453,N_23793);
and UO_698 (O_698,N_24046,N_23219);
nor UO_699 (O_699,N_23185,N_24362);
xor UO_700 (O_700,N_23619,N_23266);
nor UO_701 (O_701,N_23289,N_24553);
nor UO_702 (O_702,N_22510,N_23823);
nor UO_703 (O_703,N_24475,N_23740);
or UO_704 (O_704,N_24640,N_22616);
or UO_705 (O_705,N_23790,N_24718);
nor UO_706 (O_706,N_22542,N_23940);
xnor UO_707 (O_707,N_22910,N_22821);
and UO_708 (O_708,N_22636,N_24837);
or UO_709 (O_709,N_23157,N_23288);
nor UO_710 (O_710,N_23600,N_22817);
xnor UO_711 (O_711,N_24491,N_24752);
or UO_712 (O_712,N_22590,N_24786);
xnor UO_713 (O_713,N_24945,N_22839);
xor UO_714 (O_714,N_23366,N_24730);
xnor UO_715 (O_715,N_24787,N_23965);
nor UO_716 (O_716,N_23602,N_24962);
nor UO_717 (O_717,N_24842,N_23656);
nand UO_718 (O_718,N_23217,N_24054);
nor UO_719 (O_719,N_24289,N_24489);
xnor UO_720 (O_720,N_22854,N_24254);
nor UO_721 (O_721,N_24397,N_24203);
xor UO_722 (O_722,N_23138,N_23959);
nand UO_723 (O_723,N_22973,N_23986);
nor UO_724 (O_724,N_24862,N_24112);
xnor UO_725 (O_725,N_22637,N_23548);
nor UO_726 (O_726,N_23301,N_24557);
nand UO_727 (O_727,N_23386,N_24217);
or UO_728 (O_728,N_24022,N_23988);
and UO_729 (O_729,N_23722,N_22861);
or UO_730 (O_730,N_24364,N_24524);
nor UO_731 (O_731,N_24997,N_22538);
or UO_732 (O_732,N_24479,N_24543);
or UO_733 (O_733,N_24404,N_23308);
nor UO_734 (O_734,N_24665,N_23828);
nor UO_735 (O_735,N_24457,N_23703);
and UO_736 (O_736,N_24959,N_24641);
and UO_737 (O_737,N_24688,N_23634);
nand UO_738 (O_738,N_23400,N_24093);
nand UO_739 (O_739,N_23150,N_22729);
nand UO_740 (O_740,N_24897,N_24657);
and UO_741 (O_741,N_24664,N_23394);
or UO_742 (O_742,N_23294,N_24159);
xor UO_743 (O_743,N_24593,N_24824);
or UO_744 (O_744,N_23835,N_24645);
and UO_745 (O_745,N_22606,N_23402);
nor UO_746 (O_746,N_23830,N_23435);
nand UO_747 (O_747,N_23858,N_24419);
nand UO_748 (O_748,N_23539,N_22885);
or UO_749 (O_749,N_23242,N_23822);
or UO_750 (O_750,N_24101,N_23126);
or UO_751 (O_751,N_24176,N_22704);
nand UO_752 (O_752,N_24452,N_24376);
nand UO_753 (O_753,N_24178,N_22524);
xor UO_754 (O_754,N_24625,N_24909);
or UO_755 (O_755,N_24219,N_24095);
xor UO_756 (O_756,N_23432,N_24822);
xor UO_757 (O_757,N_24168,N_24699);
xnor UO_758 (O_758,N_23766,N_24607);
and UO_759 (O_759,N_23347,N_22828);
and UO_760 (O_760,N_24818,N_23251);
xor UO_761 (O_761,N_23989,N_23532);
nand UO_762 (O_762,N_23801,N_22981);
nor UO_763 (O_763,N_23436,N_22767);
xnor UO_764 (O_764,N_24813,N_22949);
nor UO_765 (O_765,N_24776,N_22749);
nor UO_766 (O_766,N_24763,N_23356);
xor UO_767 (O_767,N_24104,N_24760);
and UO_768 (O_768,N_23490,N_24472);
nand UO_769 (O_769,N_24731,N_23948);
and UO_770 (O_770,N_23236,N_24359);
nand UO_771 (O_771,N_24062,N_23601);
xor UO_772 (O_772,N_24794,N_22559);
or UO_773 (O_773,N_23584,N_22640);
nor UO_774 (O_774,N_23831,N_22770);
or UO_775 (O_775,N_23626,N_24836);
and UO_776 (O_776,N_24864,N_24792);
xor UO_777 (O_777,N_23005,N_23260);
nor UO_778 (O_778,N_23357,N_23013);
and UO_779 (O_779,N_24128,N_23638);
or UO_780 (O_780,N_24426,N_23814);
nor UO_781 (O_781,N_23451,N_22911);
nor UO_782 (O_782,N_23654,N_23794);
and UO_783 (O_783,N_23581,N_23720);
or UO_784 (O_784,N_23231,N_22875);
and UO_785 (O_785,N_24348,N_23846);
xnor UO_786 (O_786,N_24851,N_22742);
xor UO_787 (O_787,N_23199,N_24565);
and UO_788 (O_788,N_23655,N_24059);
nand UO_789 (O_789,N_24941,N_23627);
xor UO_790 (O_790,N_24394,N_24683);
nand UO_791 (O_791,N_24560,N_22661);
or UO_792 (O_792,N_23945,N_24621);
xnor UO_793 (O_793,N_24312,N_24848);
xor UO_794 (O_794,N_23797,N_24530);
or UO_795 (O_795,N_24618,N_24063);
or UO_796 (O_796,N_24832,N_24186);
xor UO_797 (O_797,N_24700,N_24180);
and UO_798 (O_798,N_23753,N_24608);
xnor UO_799 (O_799,N_24990,N_23937);
and UO_800 (O_800,N_22897,N_22743);
nor UO_801 (O_801,N_24287,N_23437);
nand UO_802 (O_802,N_22764,N_23540);
xnor UO_803 (O_803,N_23963,N_22932);
or UO_804 (O_804,N_24859,N_24639);
and UO_805 (O_805,N_23570,N_24292);
nand UO_806 (O_806,N_23881,N_22906);
nand UO_807 (O_807,N_24333,N_22688);
xor UO_808 (O_808,N_23640,N_24713);
xor UO_809 (O_809,N_22534,N_22536);
or UO_810 (O_810,N_24545,N_24041);
xor UO_811 (O_811,N_24904,N_23772);
and UO_812 (O_812,N_23027,N_22820);
or UO_813 (O_813,N_22870,N_23867);
or UO_814 (O_814,N_22775,N_24197);
xor UO_815 (O_815,N_24456,N_23700);
nor UO_816 (O_816,N_24854,N_24129);
nand UO_817 (O_817,N_23412,N_23957);
and UO_818 (O_818,N_24124,N_22967);
nand UO_819 (O_819,N_24591,N_23209);
xor UO_820 (O_820,N_24463,N_24339);
nor UO_821 (O_821,N_24769,N_24016);
and UO_822 (O_822,N_24793,N_23641);
xor UO_823 (O_823,N_23309,N_23152);
or UO_824 (O_824,N_24295,N_24437);
xor UO_825 (O_825,N_23690,N_24215);
xnor UO_826 (O_826,N_24809,N_24191);
nor UO_827 (O_827,N_23551,N_23762);
xor UO_828 (O_828,N_24973,N_24011);
nand UO_829 (O_829,N_24747,N_23263);
and UO_830 (O_830,N_24446,N_24031);
nor UO_831 (O_831,N_23749,N_22596);
or UO_832 (O_832,N_24017,N_24682);
nand UO_833 (O_833,N_24517,N_22587);
nand UO_834 (O_834,N_22919,N_24305);
nor UO_835 (O_835,N_24440,N_22627);
or UO_836 (O_836,N_24630,N_22571);
xnor UO_837 (O_837,N_24172,N_23903);
and UO_838 (O_838,N_23894,N_24012);
nand UO_839 (O_839,N_24005,N_24678);
or UO_840 (O_840,N_23170,N_23531);
and UO_841 (O_841,N_22666,N_24009);
or UO_842 (O_842,N_23350,N_24561);
or UO_843 (O_843,N_23999,N_24290);
and UO_844 (O_844,N_24724,N_22987);
or UO_845 (O_845,N_24118,N_23342);
nand UO_846 (O_846,N_23222,N_24578);
or UO_847 (O_847,N_24194,N_24329);
nand UO_848 (O_848,N_23119,N_23681);
or UO_849 (O_849,N_23449,N_23524);
nor UO_850 (O_850,N_24195,N_24432);
nor UO_851 (O_851,N_23478,N_23076);
and UO_852 (O_852,N_22613,N_24179);
nand UO_853 (O_853,N_22672,N_24030);
nand UO_854 (O_854,N_24335,N_24799);
or UO_855 (O_855,N_22922,N_23419);
nor UO_856 (O_856,N_24409,N_23329);
nor UO_857 (O_857,N_23324,N_23666);
nand UO_858 (O_858,N_23721,N_24251);
or UO_859 (O_859,N_23878,N_24160);
or UO_860 (O_860,N_23036,N_23379);
nand UO_861 (O_861,N_23754,N_23636);
nor UO_862 (O_862,N_22670,N_22708);
nand UO_863 (O_863,N_22623,N_22614);
nor UO_864 (O_864,N_23248,N_22728);
xor UO_865 (O_865,N_23300,N_24296);
xnor UO_866 (O_866,N_23683,N_22514);
xor UO_867 (O_867,N_22824,N_23117);
and UO_868 (O_868,N_24839,N_23658);
xor UO_869 (O_869,N_24613,N_23372);
nor UO_870 (O_870,N_24885,N_24865);
and UO_871 (O_871,N_23100,N_22857);
or UO_872 (O_872,N_24309,N_24588);
or UO_873 (O_873,N_23159,N_23184);
and UO_874 (O_874,N_24861,N_23480);
nor UO_875 (O_875,N_22874,N_22979);
nand UO_876 (O_876,N_23081,N_24330);
and UO_877 (O_877,N_24073,N_23546);
and UO_878 (O_878,N_22833,N_24991);
nor UO_879 (O_879,N_23736,N_22945);
or UO_880 (O_880,N_23595,N_22988);
nor UO_881 (O_881,N_22588,N_22810);
or UO_882 (O_882,N_24461,N_24246);
nor UO_883 (O_883,N_22650,N_24378);
or UO_884 (O_884,N_24831,N_22631);
or UO_885 (O_885,N_24943,N_24455);
nor UO_886 (O_886,N_24136,N_22646);
nor UO_887 (O_887,N_24306,N_22605);
or UO_888 (O_888,N_23717,N_24247);
nand UO_889 (O_889,N_24070,N_23410);
or UO_890 (O_890,N_22657,N_22574);
or UO_891 (O_891,N_24692,N_23003);
nor UO_892 (O_892,N_22549,N_24085);
xnor UO_893 (O_893,N_24386,N_23529);
nand UO_894 (O_894,N_23074,N_23285);
nor UO_895 (O_895,N_22576,N_24115);
or UO_896 (O_896,N_24232,N_22722);
xor UO_897 (O_897,N_22957,N_24471);
xnor UO_898 (O_898,N_23567,N_22578);
or UO_899 (O_899,N_23916,N_24185);
and UO_900 (O_900,N_24293,N_23728);
nand UO_901 (O_901,N_24049,N_22793);
nor UO_902 (O_902,N_23277,N_22976);
nor UO_903 (O_903,N_22918,N_23376);
and UO_904 (O_904,N_22577,N_22804);
or UO_905 (O_905,N_24040,N_24610);
or UO_906 (O_906,N_23373,N_23163);
and UO_907 (O_907,N_23249,N_23397);
or UO_908 (O_908,N_24600,N_23461);
xnor UO_909 (O_909,N_24304,N_24273);
nand UO_910 (O_910,N_24109,N_24961);
xnor UO_911 (O_911,N_23922,N_22687);
nor UO_912 (O_912,N_22766,N_23748);
or UO_913 (O_913,N_23755,N_23882);
nor UO_914 (O_914,N_22997,N_23389);
nor UO_915 (O_915,N_23585,N_24706);
or UO_916 (O_916,N_23792,N_24270);
or UO_917 (O_917,N_23521,N_24595);
nor UO_918 (O_918,N_23693,N_24134);
or UO_919 (O_919,N_22948,N_24634);
nand UO_920 (O_920,N_23900,N_23544);
xnor UO_921 (O_921,N_22986,N_24431);
or UO_922 (O_922,N_24147,N_23075);
and UO_923 (O_923,N_23510,N_24053);
or UO_924 (O_924,N_24342,N_24720);
and UO_925 (O_925,N_23024,N_24148);
or UO_926 (O_926,N_23872,N_23614);
nor UO_927 (O_927,N_22503,N_24956);
xor UO_928 (O_928,N_23166,N_24696);
nor UO_929 (O_929,N_24551,N_24125);
or UO_930 (O_930,N_23192,N_24624);
xor UO_931 (O_931,N_24736,N_24807);
nand UO_932 (O_932,N_23769,N_23323);
nor UO_933 (O_933,N_23599,N_22842);
nand UO_934 (O_934,N_22589,N_24874);
xnor UO_935 (O_935,N_24727,N_22982);
nand UO_936 (O_936,N_22753,N_23561);
nor UO_937 (O_937,N_23439,N_24947);
or UO_938 (O_938,N_23064,N_22799);
nor UO_939 (O_939,N_24550,N_23317);
nand UO_940 (O_940,N_22762,N_22645);
or UO_941 (O_941,N_23784,N_22963);
nor UO_942 (O_942,N_23549,N_24775);
and UO_943 (O_943,N_24153,N_24667);
or UO_944 (O_944,N_24083,N_23160);
and UO_945 (O_945,N_23825,N_24139);
nand UO_946 (O_946,N_23414,N_23469);
nand UO_947 (O_947,N_24200,N_23966);
nor UO_948 (O_948,N_24815,N_24035);
and UO_949 (O_949,N_24872,N_23817);
nor UO_950 (O_950,N_23829,N_23441);
nor UO_951 (O_951,N_24659,N_24218);
xor UO_952 (O_952,N_24704,N_23712);
nor UO_953 (O_953,N_24113,N_24555);
or UO_954 (O_954,N_24323,N_24416);
nand UO_955 (O_955,N_22618,N_23418);
or UO_956 (O_956,N_24539,N_23590);
or UO_957 (O_957,N_24370,N_24817);
nand UO_958 (O_958,N_22654,N_22573);
xnor UO_959 (O_959,N_23786,N_23214);
and UO_960 (O_960,N_22798,N_24916);
nor UO_961 (O_961,N_24609,N_24453);
nand UO_962 (O_962,N_23136,N_23780);
nor UO_963 (O_963,N_24064,N_23115);
and UO_964 (O_964,N_22959,N_23016);
nand UO_965 (O_965,N_22773,N_24334);
nand UO_966 (O_966,N_23942,N_24389);
nand UO_967 (O_967,N_23625,N_22878);
and UO_968 (O_968,N_24337,N_24802);
nand UO_969 (O_969,N_22701,N_24227);
nor UO_970 (O_970,N_23045,N_24500);
xnor UO_971 (O_971,N_23629,N_23364);
nand UO_972 (O_972,N_22974,N_24895);
nor UO_973 (O_973,N_22689,N_23454);
or UO_974 (O_974,N_24061,N_23473);
xor UO_975 (O_975,N_22846,N_24514);
nand UO_976 (O_976,N_22572,N_24527);
xor UO_977 (O_977,N_22999,N_24922);
or UO_978 (O_978,N_23995,N_24923);
nor UO_979 (O_979,N_23560,N_24886);
and UO_980 (O_980,N_24849,N_24764);
and UO_981 (O_981,N_24884,N_24408);
xor UO_982 (O_982,N_24098,N_24529);
and UO_983 (O_983,N_23976,N_23014);
and UO_984 (O_984,N_23465,N_23280);
xnor UO_985 (O_985,N_22652,N_22608);
or UO_986 (O_986,N_23680,N_24814);
or UO_987 (O_987,N_24750,N_22943);
xnor UO_988 (O_988,N_23859,N_23286);
and UO_989 (O_989,N_23007,N_23029);
or UO_990 (O_990,N_24510,N_24299);
xor UO_991 (O_991,N_24911,N_24559);
nand UO_992 (O_992,N_23541,N_23512);
or UO_993 (O_993,N_24745,N_24581);
and UO_994 (O_994,N_24174,N_23488);
and UO_995 (O_995,N_24399,N_23669);
nor UO_996 (O_996,N_22751,N_24902);
and UO_997 (O_997,N_24258,N_24590);
nor UO_998 (O_998,N_22634,N_24226);
and UO_999 (O_999,N_24076,N_24901);
or UO_1000 (O_1000,N_24152,N_23382);
xor UO_1001 (O_1001,N_23924,N_24094);
or UO_1002 (O_1002,N_24025,N_22898);
nor UO_1003 (O_1003,N_24150,N_23607);
nand UO_1004 (O_1004,N_24950,N_22601);
and UO_1005 (O_1005,N_22886,N_23582);
nor UO_1006 (O_1006,N_23404,N_24089);
nand UO_1007 (O_1007,N_22769,N_24161);
nand UO_1008 (O_1008,N_24669,N_23044);
xnor UO_1009 (O_1009,N_22518,N_24615);
and UO_1010 (O_1010,N_24216,N_22971);
nand UO_1011 (O_1011,N_23973,N_23938);
nand UO_1012 (O_1012,N_23368,N_23917);
nor UO_1013 (O_1013,N_22677,N_24429);
nand UO_1014 (O_1014,N_23885,N_24525);
and UO_1015 (O_1015,N_23334,N_22990);
and UO_1016 (O_1016,N_24047,N_24651);
or UO_1017 (O_1017,N_24448,N_24503);
nand UO_1018 (O_1018,N_24268,N_22845);
and UO_1019 (O_1019,N_24733,N_24597);
and UO_1020 (O_1020,N_23918,N_24146);
or UO_1021 (O_1021,N_22768,N_24151);
nand UO_1022 (O_1022,N_23069,N_22555);
nand UO_1023 (O_1023,N_24314,N_22505);
nor UO_1024 (O_1024,N_24940,N_22706);
and UO_1025 (O_1025,N_23475,N_22782);
xor UO_1026 (O_1026,N_23939,N_23592);
xnor UO_1027 (O_1027,N_24585,N_23519);
nand UO_1028 (O_1028,N_24611,N_23925);
and UO_1029 (O_1029,N_24075,N_24804);
nand UO_1030 (O_1030,N_23821,N_24619);
and UO_1031 (O_1031,N_23910,N_23504);
nor UO_1032 (O_1032,N_23815,N_23128);
nor UO_1033 (O_1033,N_23195,N_24970);
xor UO_1034 (O_1034,N_23886,N_23471);
or UO_1035 (O_1035,N_23363,N_22562);
xor UO_1036 (O_1036,N_24932,N_24199);
xnor UO_1037 (O_1037,N_23178,N_23487);
nand UO_1038 (O_1038,N_23305,N_22803);
or UO_1039 (O_1039,N_23639,N_22702);
xor UO_1040 (O_1040,N_23425,N_24117);
nor UO_1041 (O_1041,N_22734,N_23270);
or UO_1042 (O_1042,N_23137,N_24632);
xor UO_1043 (O_1043,N_22760,N_23140);
nor UO_1044 (O_1044,N_24454,N_24420);
and UO_1045 (O_1045,N_23708,N_24250);
nand UO_1046 (O_1046,N_22691,N_23237);
nor UO_1047 (O_1047,N_24081,N_22755);
or UO_1048 (O_1048,N_22508,N_23864);
xnor UO_1049 (O_1049,N_23440,N_24952);
and UO_1050 (O_1050,N_23104,N_23969);
or UO_1051 (O_1051,N_24552,N_23953);
and UO_1052 (O_1052,N_23370,N_23782);
nor UO_1053 (O_1053,N_24596,N_23243);
or UO_1054 (O_1054,N_22834,N_24373);
nor UO_1055 (O_1055,N_24110,N_23227);
or UO_1056 (O_1056,N_23812,N_24594);
and UO_1057 (O_1057,N_24933,N_24906);
nor UO_1058 (O_1058,N_23078,N_23244);
and UO_1059 (O_1059,N_23284,N_24628);
nor UO_1060 (O_1060,N_24281,N_23445);
nor UO_1061 (O_1061,N_24120,N_24549);
or UO_1062 (O_1062,N_22801,N_24413);
nor UO_1063 (O_1063,N_23855,N_24847);
xor UO_1064 (O_1064,N_24387,N_24484);
nor UO_1065 (O_1065,N_23637,N_23271);
or UO_1066 (O_1066,N_22682,N_24224);
or UO_1067 (O_1067,N_24638,N_22719);
nor UO_1068 (O_1068,N_23443,N_24014);
nand UO_1069 (O_1069,N_23486,N_23511);
nand UO_1070 (O_1070,N_23181,N_23226);
nor UO_1071 (O_1071,N_23186,N_23240);
xor UO_1072 (O_1072,N_23047,N_24805);
and UO_1073 (O_1073,N_22840,N_23706);
or UO_1074 (O_1074,N_24301,N_24509);
and UO_1075 (O_1075,N_23985,N_24749);
and UO_1076 (O_1076,N_23697,N_23463);
or UO_1077 (O_1077,N_24674,N_23672);
xor UO_1078 (O_1078,N_22591,N_23348);
nand UO_1079 (O_1079,N_22930,N_24554);
or UO_1080 (O_1080,N_24493,N_23012);
nand UO_1081 (O_1081,N_24007,N_24481);
xor UO_1082 (O_1082,N_22642,N_24255);
and UO_1083 (O_1083,N_23820,N_23628);
nand UO_1084 (O_1084,N_23777,N_24852);
xor UO_1085 (O_1085,N_23633,N_24528);
and UO_1086 (O_1086,N_22685,N_22647);
xor UO_1087 (O_1087,N_23053,N_22771);
xnor UO_1088 (O_1088,N_24803,N_24868);
or UO_1089 (O_1089,N_24156,N_24365);
nand UO_1090 (O_1090,N_23776,N_23520);
xor UO_1091 (O_1091,N_23854,N_22844);
xnor UO_1092 (O_1092,N_24310,N_23765);
nor UO_1093 (O_1093,N_24819,N_23189);
xnor UO_1094 (O_1094,N_24725,N_22500);
xor UO_1095 (O_1095,N_24784,N_23228);
nand UO_1096 (O_1096,N_22692,N_24567);
and UO_1097 (O_1097,N_23530,N_22520);
xnor UO_1098 (O_1098,N_23238,N_24252);
or UO_1099 (O_1099,N_23760,N_22530);
nor UO_1100 (O_1100,N_23493,N_22723);
or UO_1101 (O_1101,N_23327,N_23077);
or UO_1102 (O_1102,N_23928,N_23385);
nand UO_1103 (O_1103,N_23699,N_24126);
xor UO_1104 (O_1104,N_23206,N_24102);
xor UO_1105 (O_1105,N_24843,N_23593);
and UO_1106 (O_1106,N_23021,N_24777);
and UO_1107 (O_1107,N_23102,N_22912);
and UO_1108 (O_1108,N_22939,N_24964);
and UO_1109 (O_1109,N_24666,N_23726);
and UO_1110 (O_1110,N_24082,N_24771);
nor UO_1111 (O_1111,N_22964,N_24643);
xnor UO_1112 (O_1112,N_24498,N_24729);
or UO_1113 (O_1113,N_24844,N_24512);
xnor UO_1114 (O_1114,N_23068,N_23254);
nor UO_1115 (O_1115,N_22926,N_23421);
nor UO_1116 (O_1116,N_23845,N_22851);
and UO_1117 (O_1117,N_24914,N_22819);
nor UO_1118 (O_1118,N_24239,N_24737);
xor UO_1119 (O_1119,N_23981,N_23725);
or UO_1120 (O_1120,N_23667,N_23675);
xnor UO_1121 (O_1121,N_22641,N_24811);
nand UO_1122 (O_1122,N_23328,N_23857);
xor UO_1123 (O_1123,N_24860,N_24511);
nor UO_1124 (O_1124,N_23481,N_23594);
nand UO_1125 (O_1125,N_24411,N_22955);
xor UO_1126 (O_1126,N_23056,N_24237);
xnor UO_1127 (O_1127,N_23127,N_23744);
nor UO_1128 (O_1128,N_24356,N_23875);
xor UO_1129 (O_1129,N_24375,N_23123);
xnor UO_1130 (O_1130,N_24829,N_24350);
nor UO_1131 (O_1131,N_23799,N_24687);
or UO_1132 (O_1132,N_24138,N_24235);
nand UO_1133 (O_1133,N_24245,N_23303);
nor UO_1134 (O_1134,N_24835,N_23456);
nand UO_1135 (O_1135,N_23430,N_22812);
nand UO_1136 (O_1136,N_24918,N_24768);
nand UO_1137 (O_1137,N_23276,N_22713);
nor UO_1138 (O_1138,N_22513,N_24276);
nor UO_1139 (O_1139,N_24971,N_24428);
nand UO_1140 (O_1140,N_23239,N_22603);
xnor UO_1141 (O_1141,N_22900,N_24071);
nand UO_1142 (O_1142,N_22690,N_24154);
nand UO_1143 (O_1143,N_23245,N_24753);
and UO_1144 (O_1144,N_24163,N_22843);
xnor UO_1145 (O_1145,N_23335,N_23734);
nand UO_1146 (O_1146,N_24405,N_22715);
and UO_1147 (O_1147,N_23499,N_24439);
and UO_1148 (O_1148,N_23664,N_23698);
and UO_1149 (O_1149,N_24210,N_24840);
nor UO_1150 (O_1150,N_22993,N_23154);
nor UO_1151 (O_1151,N_23523,N_24889);
nand UO_1152 (O_1152,N_23559,N_23778);
nand UO_1153 (O_1153,N_22937,N_24627);
nand UO_1154 (O_1154,N_23050,N_24702);
nand UO_1155 (O_1155,N_24676,N_22667);
nand UO_1156 (O_1156,N_22915,N_23852);
nor UO_1157 (O_1157,N_22612,N_24603);
or UO_1158 (O_1158,N_22545,N_24371);
nor UO_1159 (O_1159,N_23009,N_24928);
nor UO_1160 (O_1160,N_22651,N_23884);
or UO_1161 (O_1161,N_24331,N_23615);
xor UO_1162 (O_1162,N_24770,N_24675);
xor UO_1163 (O_1163,N_22517,N_24673);
nor UO_1164 (O_1164,N_23279,N_23307);
and UO_1165 (O_1165,N_24957,N_24756);
and UO_1166 (O_1166,N_23060,N_24741);
nand UO_1167 (O_1167,N_24698,N_23116);
xnor UO_1168 (O_1168,N_24899,N_23791);
nand UO_1169 (O_1169,N_23873,N_23039);
xor UO_1170 (O_1170,N_23679,N_24913);
and UO_1171 (O_1171,N_23798,N_24490);
nand UO_1172 (O_1172,N_24531,N_23608);
or UO_1173 (O_1173,N_23256,N_23941);
or UO_1174 (O_1174,N_23438,N_22892);
xnor UO_1175 (O_1175,N_22901,N_23974);
nand UO_1176 (O_1176,N_23713,N_24143);
xor UO_1177 (O_1177,N_22632,N_23583);
and UO_1178 (O_1178,N_23362,N_23606);
or UO_1179 (O_1179,N_23868,N_23887);
and UO_1180 (O_1180,N_23783,N_24969);
xor UO_1181 (O_1181,N_23554,N_23566);
nand UO_1182 (O_1182,N_22856,N_22984);
xor UO_1183 (O_1183,N_23746,N_23028);
nand UO_1184 (O_1184,N_24279,N_22709);
xor UO_1185 (O_1185,N_24100,N_24986);
xnor UO_1186 (O_1186,N_22853,N_23643);
and UO_1187 (O_1187,N_24221,N_24984);
or UO_1188 (O_1188,N_24637,N_23258);
or UO_1189 (O_1189,N_23911,N_24265);
nor UO_1190 (O_1190,N_23944,N_23293);
nor UO_1191 (O_1191,N_24801,N_22970);
nor UO_1192 (O_1192,N_24908,N_23283);
xor UO_1193 (O_1193,N_22515,N_24133);
nand UO_1194 (O_1194,N_22927,N_22956);
or UO_1195 (O_1195,N_23306,N_24360);
and UO_1196 (O_1196,N_24496,N_24321);
or UO_1197 (O_1197,N_24508,N_23072);
and UO_1198 (O_1198,N_23761,N_24406);
nor UO_1199 (O_1199,N_24099,N_23788);
or UO_1200 (O_1200,N_23051,N_24602);
or UO_1201 (O_1201,N_24965,N_24566);
or UO_1202 (O_1202,N_22531,N_23980);
and UO_1203 (O_1203,N_23265,N_22698);
and UO_1204 (O_1204,N_24507,N_23365);
nand UO_1205 (O_1205,N_24646,N_24944);
and UO_1206 (O_1206,N_22663,N_24436);
nor UO_1207 (O_1207,N_22658,N_23057);
and UO_1208 (O_1208,N_24177,N_24748);
or UO_1209 (O_1209,N_23714,N_22543);
xnor UO_1210 (O_1210,N_23644,N_23677);
or UO_1211 (O_1211,N_23351,N_24653);
and UO_1212 (O_1212,N_23423,N_24668);
nor UO_1213 (O_1213,N_23621,N_23759);
and UO_1214 (O_1214,N_23322,N_23558);
or UO_1215 (O_1215,N_24028,N_23147);
or UO_1216 (O_1216,N_23861,N_23202);
nor UO_1217 (O_1217,N_23501,N_22705);
nand UO_1218 (O_1218,N_23141,N_24953);
nor UO_1219 (O_1219,N_24282,N_24915);
or UO_1220 (O_1220,N_23796,N_23574);
nor UO_1221 (O_1221,N_23552,N_23017);
nor UO_1222 (O_1222,N_23517,N_24601);
xor UO_1223 (O_1223,N_23912,N_24274);
or UO_1224 (O_1224,N_23037,N_24349);
nor UO_1225 (O_1225,N_23767,N_23124);
or UO_1226 (O_1226,N_24253,N_24204);
nor UO_1227 (O_1227,N_24929,N_22871);
or UO_1228 (O_1228,N_22730,N_23670);
nor UO_1229 (O_1229,N_23663,N_24029);
or UO_1230 (O_1230,N_24271,N_23125);
xnor UO_1231 (O_1231,N_24910,N_23089);
nor UO_1232 (O_1232,N_24051,N_23383);
nand UO_1233 (O_1233,N_24211,N_23883);
or UO_1234 (O_1234,N_24345,N_22527);
nor UO_1235 (O_1235,N_24656,N_23901);
nor UO_1236 (O_1236,N_24326,N_24465);
nand UO_1237 (O_1237,N_23904,N_22895);
xor UO_1238 (O_1238,N_23813,N_23482);
nor UO_1239 (O_1239,N_24069,N_24917);
nand UO_1240 (O_1240,N_24328,N_22584);
nand UO_1241 (O_1241,N_23889,N_23299);
xnor UO_1242 (O_1242,N_23612,N_22523);
xor UO_1243 (O_1243,N_23870,N_22925);
or UO_1244 (O_1244,N_22580,N_22560);
and UO_1245 (O_1245,N_24466,N_24240);
and UO_1246 (O_1246,N_22547,N_24427);
nand UO_1247 (O_1247,N_22830,N_23018);
nor UO_1248 (O_1248,N_22847,N_24589);
and UO_1249 (O_1249,N_24494,N_23715);
or UO_1250 (O_1250,N_24856,N_22649);
nand UO_1251 (O_1251,N_24276,N_22939);
xnor UO_1252 (O_1252,N_24013,N_23286);
xnor UO_1253 (O_1253,N_23612,N_24631);
xor UO_1254 (O_1254,N_24700,N_24085);
nor UO_1255 (O_1255,N_23215,N_23184);
or UO_1256 (O_1256,N_23313,N_23193);
nand UO_1257 (O_1257,N_23741,N_24055);
nor UO_1258 (O_1258,N_24447,N_24057);
nor UO_1259 (O_1259,N_23975,N_24110);
and UO_1260 (O_1260,N_22681,N_23700);
and UO_1261 (O_1261,N_24813,N_23714);
xnor UO_1262 (O_1262,N_24419,N_23152);
nor UO_1263 (O_1263,N_23109,N_23104);
xnor UO_1264 (O_1264,N_24391,N_24203);
and UO_1265 (O_1265,N_22841,N_22529);
and UO_1266 (O_1266,N_22934,N_24109);
and UO_1267 (O_1267,N_24554,N_23823);
xor UO_1268 (O_1268,N_23163,N_24680);
and UO_1269 (O_1269,N_23666,N_23164);
nor UO_1270 (O_1270,N_24464,N_24264);
nand UO_1271 (O_1271,N_24131,N_23532);
or UO_1272 (O_1272,N_24951,N_23056);
nand UO_1273 (O_1273,N_22611,N_24175);
nand UO_1274 (O_1274,N_23956,N_23656);
and UO_1275 (O_1275,N_23213,N_23237);
or UO_1276 (O_1276,N_24262,N_23245);
nor UO_1277 (O_1277,N_23337,N_22835);
and UO_1278 (O_1278,N_24201,N_24273);
nor UO_1279 (O_1279,N_22671,N_24568);
nor UO_1280 (O_1280,N_23553,N_22751);
and UO_1281 (O_1281,N_24329,N_23147);
nor UO_1282 (O_1282,N_24782,N_23322);
xor UO_1283 (O_1283,N_24561,N_24831);
xor UO_1284 (O_1284,N_24650,N_24610);
and UO_1285 (O_1285,N_22543,N_23316);
nor UO_1286 (O_1286,N_23730,N_24361);
nand UO_1287 (O_1287,N_24896,N_22520);
and UO_1288 (O_1288,N_23897,N_24458);
nor UO_1289 (O_1289,N_24841,N_23488);
and UO_1290 (O_1290,N_23070,N_24578);
nand UO_1291 (O_1291,N_23797,N_22732);
nand UO_1292 (O_1292,N_22881,N_22655);
or UO_1293 (O_1293,N_24121,N_22951);
xnor UO_1294 (O_1294,N_24351,N_24694);
or UO_1295 (O_1295,N_23272,N_23605);
and UO_1296 (O_1296,N_23789,N_24055);
xnor UO_1297 (O_1297,N_23611,N_23982);
and UO_1298 (O_1298,N_23654,N_23318);
nor UO_1299 (O_1299,N_22659,N_23126);
or UO_1300 (O_1300,N_22524,N_23453);
xor UO_1301 (O_1301,N_24255,N_23610);
nand UO_1302 (O_1302,N_23638,N_24297);
nand UO_1303 (O_1303,N_23401,N_24465);
nor UO_1304 (O_1304,N_23457,N_24988);
nor UO_1305 (O_1305,N_24167,N_24647);
or UO_1306 (O_1306,N_23177,N_24221);
or UO_1307 (O_1307,N_23726,N_24941);
and UO_1308 (O_1308,N_23858,N_24799);
nand UO_1309 (O_1309,N_24973,N_23902);
nor UO_1310 (O_1310,N_23215,N_23009);
nand UO_1311 (O_1311,N_24973,N_24978);
xor UO_1312 (O_1312,N_23491,N_22622);
and UO_1313 (O_1313,N_24544,N_22647);
nor UO_1314 (O_1314,N_24880,N_24524);
nor UO_1315 (O_1315,N_23185,N_23529);
nor UO_1316 (O_1316,N_23847,N_22880);
or UO_1317 (O_1317,N_24731,N_22940);
and UO_1318 (O_1318,N_24356,N_23151);
nor UO_1319 (O_1319,N_24287,N_23959);
nand UO_1320 (O_1320,N_24509,N_24627);
nor UO_1321 (O_1321,N_22772,N_23084);
and UO_1322 (O_1322,N_24664,N_24871);
and UO_1323 (O_1323,N_22663,N_24178);
nor UO_1324 (O_1324,N_22806,N_24315);
and UO_1325 (O_1325,N_22502,N_22949);
xnor UO_1326 (O_1326,N_24579,N_24395);
xor UO_1327 (O_1327,N_23850,N_23464);
nand UO_1328 (O_1328,N_24873,N_23492);
or UO_1329 (O_1329,N_24066,N_24671);
or UO_1330 (O_1330,N_24225,N_23761);
nor UO_1331 (O_1331,N_22592,N_24685);
nor UO_1332 (O_1332,N_23353,N_24695);
nand UO_1333 (O_1333,N_23377,N_23525);
xor UO_1334 (O_1334,N_24338,N_22679);
nand UO_1335 (O_1335,N_23189,N_24079);
or UO_1336 (O_1336,N_22950,N_23827);
nor UO_1337 (O_1337,N_24126,N_24099);
and UO_1338 (O_1338,N_24882,N_24725);
nor UO_1339 (O_1339,N_23588,N_24150);
nor UO_1340 (O_1340,N_23665,N_24705);
nand UO_1341 (O_1341,N_23766,N_23417);
or UO_1342 (O_1342,N_22570,N_23533);
and UO_1343 (O_1343,N_24185,N_22582);
or UO_1344 (O_1344,N_23106,N_24259);
or UO_1345 (O_1345,N_22740,N_22924);
xnor UO_1346 (O_1346,N_23682,N_23944);
nand UO_1347 (O_1347,N_23182,N_22558);
nor UO_1348 (O_1348,N_23925,N_23401);
nand UO_1349 (O_1349,N_23436,N_23553);
nand UO_1350 (O_1350,N_22952,N_24332);
nand UO_1351 (O_1351,N_24955,N_22861);
nor UO_1352 (O_1352,N_22771,N_23643);
xnor UO_1353 (O_1353,N_24762,N_23265);
nand UO_1354 (O_1354,N_22763,N_22937);
xnor UO_1355 (O_1355,N_22820,N_23367);
xnor UO_1356 (O_1356,N_24549,N_24656);
nor UO_1357 (O_1357,N_24531,N_23168);
xor UO_1358 (O_1358,N_24989,N_23634);
or UO_1359 (O_1359,N_24316,N_24234);
or UO_1360 (O_1360,N_23756,N_23481);
nand UO_1361 (O_1361,N_23305,N_24032);
nand UO_1362 (O_1362,N_23970,N_23616);
and UO_1363 (O_1363,N_23187,N_23574);
nand UO_1364 (O_1364,N_24759,N_24299);
nand UO_1365 (O_1365,N_24981,N_24169);
nand UO_1366 (O_1366,N_22894,N_24395);
nand UO_1367 (O_1367,N_24447,N_24662);
or UO_1368 (O_1368,N_22566,N_22512);
xor UO_1369 (O_1369,N_23166,N_23071);
or UO_1370 (O_1370,N_24866,N_23532);
nand UO_1371 (O_1371,N_23465,N_22650);
nand UO_1372 (O_1372,N_23943,N_24878);
nor UO_1373 (O_1373,N_24356,N_24278);
nand UO_1374 (O_1374,N_24005,N_23000);
xnor UO_1375 (O_1375,N_24496,N_24051);
xor UO_1376 (O_1376,N_22619,N_24151);
xnor UO_1377 (O_1377,N_23954,N_24060);
nand UO_1378 (O_1378,N_23143,N_22848);
xnor UO_1379 (O_1379,N_22563,N_22620);
nor UO_1380 (O_1380,N_22702,N_23557);
xor UO_1381 (O_1381,N_24459,N_24891);
nor UO_1382 (O_1382,N_24901,N_23922);
nand UO_1383 (O_1383,N_22901,N_24149);
or UO_1384 (O_1384,N_23032,N_24197);
and UO_1385 (O_1385,N_22837,N_22972);
xor UO_1386 (O_1386,N_23590,N_24370);
xor UO_1387 (O_1387,N_22674,N_24268);
nand UO_1388 (O_1388,N_23468,N_22744);
nand UO_1389 (O_1389,N_22800,N_22753);
or UO_1390 (O_1390,N_24511,N_24504);
or UO_1391 (O_1391,N_23615,N_24529);
and UO_1392 (O_1392,N_22549,N_24750);
and UO_1393 (O_1393,N_24126,N_22977);
nand UO_1394 (O_1394,N_23523,N_23822);
and UO_1395 (O_1395,N_22703,N_23513);
and UO_1396 (O_1396,N_23003,N_23710);
xor UO_1397 (O_1397,N_23041,N_23435);
or UO_1398 (O_1398,N_24391,N_22916);
and UO_1399 (O_1399,N_22689,N_24623);
nor UO_1400 (O_1400,N_23304,N_22937);
and UO_1401 (O_1401,N_24933,N_24087);
xnor UO_1402 (O_1402,N_24976,N_24178);
or UO_1403 (O_1403,N_24503,N_23623);
and UO_1404 (O_1404,N_24728,N_24636);
or UO_1405 (O_1405,N_24321,N_23260);
and UO_1406 (O_1406,N_24774,N_24223);
or UO_1407 (O_1407,N_23596,N_23731);
nor UO_1408 (O_1408,N_24677,N_23816);
nor UO_1409 (O_1409,N_23905,N_23245);
and UO_1410 (O_1410,N_23378,N_22628);
xor UO_1411 (O_1411,N_22728,N_23858);
nor UO_1412 (O_1412,N_24954,N_23461);
nor UO_1413 (O_1413,N_24293,N_23177);
nor UO_1414 (O_1414,N_22722,N_23193);
or UO_1415 (O_1415,N_24497,N_23235);
nand UO_1416 (O_1416,N_24543,N_24872);
nand UO_1417 (O_1417,N_23593,N_23203);
nand UO_1418 (O_1418,N_23635,N_24181);
or UO_1419 (O_1419,N_23954,N_23390);
and UO_1420 (O_1420,N_24608,N_24438);
and UO_1421 (O_1421,N_23188,N_24674);
xnor UO_1422 (O_1422,N_23567,N_24199);
nor UO_1423 (O_1423,N_22543,N_24198);
nand UO_1424 (O_1424,N_24108,N_22987);
and UO_1425 (O_1425,N_24360,N_24111);
or UO_1426 (O_1426,N_23522,N_24776);
and UO_1427 (O_1427,N_23260,N_22671);
or UO_1428 (O_1428,N_24532,N_22824);
xor UO_1429 (O_1429,N_23998,N_24389);
xnor UO_1430 (O_1430,N_23221,N_24425);
and UO_1431 (O_1431,N_22622,N_24871);
and UO_1432 (O_1432,N_23687,N_24329);
xnor UO_1433 (O_1433,N_24812,N_22529);
nand UO_1434 (O_1434,N_22999,N_22891);
and UO_1435 (O_1435,N_24407,N_24289);
xor UO_1436 (O_1436,N_24631,N_23244);
nand UO_1437 (O_1437,N_24488,N_23916);
and UO_1438 (O_1438,N_24636,N_24281);
nand UO_1439 (O_1439,N_22577,N_23832);
and UO_1440 (O_1440,N_24263,N_24015);
nand UO_1441 (O_1441,N_24665,N_23766);
xnor UO_1442 (O_1442,N_23373,N_24145);
or UO_1443 (O_1443,N_23173,N_24189);
and UO_1444 (O_1444,N_24107,N_22593);
xnor UO_1445 (O_1445,N_23581,N_22896);
xnor UO_1446 (O_1446,N_22956,N_23825);
and UO_1447 (O_1447,N_24136,N_24972);
and UO_1448 (O_1448,N_23503,N_23465);
and UO_1449 (O_1449,N_24909,N_22785);
or UO_1450 (O_1450,N_23397,N_23813);
nor UO_1451 (O_1451,N_24452,N_24077);
xnor UO_1452 (O_1452,N_23960,N_23904);
and UO_1453 (O_1453,N_24284,N_23016);
nor UO_1454 (O_1454,N_24072,N_24002);
and UO_1455 (O_1455,N_23207,N_24250);
nor UO_1456 (O_1456,N_23209,N_23810);
nand UO_1457 (O_1457,N_24334,N_22762);
nor UO_1458 (O_1458,N_23376,N_23981);
and UO_1459 (O_1459,N_23072,N_23277);
nor UO_1460 (O_1460,N_22993,N_24481);
xor UO_1461 (O_1461,N_23721,N_23770);
and UO_1462 (O_1462,N_24097,N_24489);
or UO_1463 (O_1463,N_23284,N_22630);
nor UO_1464 (O_1464,N_23134,N_23805);
or UO_1465 (O_1465,N_22838,N_23254);
xor UO_1466 (O_1466,N_23098,N_24935);
nor UO_1467 (O_1467,N_22947,N_24492);
xnor UO_1468 (O_1468,N_24421,N_23265);
xnor UO_1469 (O_1469,N_23686,N_23913);
nor UO_1470 (O_1470,N_22687,N_24990);
nand UO_1471 (O_1471,N_23803,N_24553);
or UO_1472 (O_1472,N_23721,N_24067);
nor UO_1473 (O_1473,N_24294,N_24135);
nand UO_1474 (O_1474,N_23845,N_23259);
nor UO_1475 (O_1475,N_23765,N_24957);
nor UO_1476 (O_1476,N_24378,N_24369);
nor UO_1477 (O_1477,N_23282,N_24937);
xnor UO_1478 (O_1478,N_24182,N_24022);
nand UO_1479 (O_1479,N_24858,N_24449);
and UO_1480 (O_1480,N_22968,N_24384);
nand UO_1481 (O_1481,N_24037,N_24457);
and UO_1482 (O_1482,N_24002,N_24465);
or UO_1483 (O_1483,N_24390,N_22886);
nor UO_1484 (O_1484,N_24648,N_22796);
nor UO_1485 (O_1485,N_24805,N_22548);
and UO_1486 (O_1486,N_24945,N_23297);
nor UO_1487 (O_1487,N_23536,N_22802);
xor UO_1488 (O_1488,N_24936,N_22767);
xnor UO_1489 (O_1489,N_23747,N_24227);
and UO_1490 (O_1490,N_24659,N_24031);
xor UO_1491 (O_1491,N_23053,N_24486);
and UO_1492 (O_1492,N_22931,N_23109);
nand UO_1493 (O_1493,N_22941,N_24986);
and UO_1494 (O_1494,N_23003,N_24298);
or UO_1495 (O_1495,N_24020,N_24001);
nand UO_1496 (O_1496,N_22756,N_22503);
and UO_1497 (O_1497,N_24087,N_23170);
xnor UO_1498 (O_1498,N_24081,N_22580);
nor UO_1499 (O_1499,N_22597,N_23962);
nor UO_1500 (O_1500,N_23582,N_22556);
or UO_1501 (O_1501,N_24134,N_24765);
nand UO_1502 (O_1502,N_23372,N_24136);
and UO_1503 (O_1503,N_24741,N_24213);
or UO_1504 (O_1504,N_23137,N_24020);
xor UO_1505 (O_1505,N_23600,N_22990);
xor UO_1506 (O_1506,N_23400,N_23687);
and UO_1507 (O_1507,N_23469,N_22585);
nor UO_1508 (O_1508,N_24749,N_23586);
or UO_1509 (O_1509,N_23004,N_24083);
and UO_1510 (O_1510,N_23992,N_23949);
nand UO_1511 (O_1511,N_23215,N_24842);
and UO_1512 (O_1512,N_24160,N_22934);
and UO_1513 (O_1513,N_24250,N_23783);
or UO_1514 (O_1514,N_24478,N_23197);
nand UO_1515 (O_1515,N_24601,N_22537);
nand UO_1516 (O_1516,N_23169,N_22508);
and UO_1517 (O_1517,N_23362,N_23006);
and UO_1518 (O_1518,N_22533,N_23183);
nor UO_1519 (O_1519,N_24864,N_24145);
nor UO_1520 (O_1520,N_22584,N_24184);
nand UO_1521 (O_1521,N_24444,N_23011);
xor UO_1522 (O_1522,N_22503,N_22858);
or UO_1523 (O_1523,N_24833,N_22919);
and UO_1524 (O_1524,N_22558,N_23427);
nor UO_1525 (O_1525,N_23800,N_23893);
xor UO_1526 (O_1526,N_23083,N_23031);
nor UO_1527 (O_1527,N_22890,N_23978);
or UO_1528 (O_1528,N_23427,N_24362);
xor UO_1529 (O_1529,N_24998,N_23577);
or UO_1530 (O_1530,N_23662,N_23487);
or UO_1531 (O_1531,N_24898,N_24672);
and UO_1532 (O_1532,N_22885,N_23832);
nand UO_1533 (O_1533,N_22944,N_23610);
nand UO_1534 (O_1534,N_22617,N_24016);
nand UO_1535 (O_1535,N_23976,N_23409);
xor UO_1536 (O_1536,N_23876,N_22616);
nor UO_1537 (O_1537,N_24171,N_22739);
and UO_1538 (O_1538,N_24788,N_24631);
nor UO_1539 (O_1539,N_23697,N_24526);
or UO_1540 (O_1540,N_24656,N_24878);
nor UO_1541 (O_1541,N_24111,N_24973);
xnor UO_1542 (O_1542,N_23956,N_24649);
or UO_1543 (O_1543,N_24987,N_24372);
and UO_1544 (O_1544,N_23094,N_23198);
nand UO_1545 (O_1545,N_24440,N_24729);
nor UO_1546 (O_1546,N_22668,N_22544);
nand UO_1547 (O_1547,N_24155,N_24926);
or UO_1548 (O_1548,N_23166,N_24858);
nand UO_1549 (O_1549,N_23331,N_22529);
nor UO_1550 (O_1550,N_22572,N_23996);
or UO_1551 (O_1551,N_22531,N_23185);
or UO_1552 (O_1552,N_24300,N_23611);
nor UO_1553 (O_1553,N_23078,N_24667);
nor UO_1554 (O_1554,N_22980,N_23551);
and UO_1555 (O_1555,N_24543,N_24806);
nor UO_1556 (O_1556,N_22750,N_23084);
or UO_1557 (O_1557,N_23872,N_23376);
and UO_1558 (O_1558,N_23535,N_24689);
xor UO_1559 (O_1559,N_24830,N_24727);
or UO_1560 (O_1560,N_23395,N_23872);
nor UO_1561 (O_1561,N_24003,N_24307);
nand UO_1562 (O_1562,N_24487,N_24813);
or UO_1563 (O_1563,N_22501,N_24283);
nor UO_1564 (O_1564,N_23562,N_23543);
xor UO_1565 (O_1565,N_24440,N_23515);
and UO_1566 (O_1566,N_22880,N_24361);
or UO_1567 (O_1567,N_23544,N_23342);
or UO_1568 (O_1568,N_23002,N_24587);
or UO_1569 (O_1569,N_24476,N_24954);
xnor UO_1570 (O_1570,N_24671,N_24895);
xnor UO_1571 (O_1571,N_24848,N_23955);
and UO_1572 (O_1572,N_23470,N_23092);
xnor UO_1573 (O_1573,N_24405,N_24295);
and UO_1574 (O_1574,N_24735,N_24838);
nor UO_1575 (O_1575,N_24248,N_23909);
nand UO_1576 (O_1576,N_22681,N_24566);
nor UO_1577 (O_1577,N_24941,N_24946);
nor UO_1578 (O_1578,N_22535,N_23157);
nand UO_1579 (O_1579,N_23079,N_24331);
nand UO_1580 (O_1580,N_24249,N_24147);
nand UO_1581 (O_1581,N_24357,N_24928);
xnor UO_1582 (O_1582,N_22774,N_23051);
or UO_1583 (O_1583,N_24538,N_24167);
or UO_1584 (O_1584,N_24854,N_22891);
xnor UO_1585 (O_1585,N_24973,N_24286);
nand UO_1586 (O_1586,N_24262,N_24253);
and UO_1587 (O_1587,N_22748,N_24273);
xnor UO_1588 (O_1588,N_23976,N_22981);
or UO_1589 (O_1589,N_23132,N_23202);
and UO_1590 (O_1590,N_24215,N_24193);
or UO_1591 (O_1591,N_23033,N_24273);
or UO_1592 (O_1592,N_23261,N_24001);
or UO_1593 (O_1593,N_23069,N_24528);
or UO_1594 (O_1594,N_22500,N_24553);
and UO_1595 (O_1595,N_23385,N_24805);
and UO_1596 (O_1596,N_23005,N_23744);
xor UO_1597 (O_1597,N_24990,N_22915);
or UO_1598 (O_1598,N_24093,N_24371);
xor UO_1599 (O_1599,N_22767,N_24860);
nand UO_1600 (O_1600,N_24577,N_22692);
nor UO_1601 (O_1601,N_23029,N_24887);
and UO_1602 (O_1602,N_22942,N_22872);
nor UO_1603 (O_1603,N_23507,N_22814);
xor UO_1604 (O_1604,N_22559,N_24578);
or UO_1605 (O_1605,N_24316,N_23509);
or UO_1606 (O_1606,N_23931,N_24556);
nand UO_1607 (O_1607,N_22898,N_24149);
or UO_1608 (O_1608,N_22697,N_23735);
or UO_1609 (O_1609,N_23340,N_24848);
and UO_1610 (O_1610,N_22648,N_22775);
or UO_1611 (O_1611,N_22995,N_24233);
and UO_1612 (O_1612,N_23236,N_23556);
or UO_1613 (O_1613,N_23180,N_24468);
nor UO_1614 (O_1614,N_23131,N_22691);
nor UO_1615 (O_1615,N_23199,N_22994);
nand UO_1616 (O_1616,N_24468,N_24207);
or UO_1617 (O_1617,N_23998,N_23727);
and UO_1618 (O_1618,N_22704,N_24580);
and UO_1619 (O_1619,N_24046,N_22643);
nand UO_1620 (O_1620,N_24772,N_24074);
or UO_1621 (O_1621,N_24317,N_24299);
nand UO_1622 (O_1622,N_22970,N_24988);
and UO_1623 (O_1623,N_24170,N_24607);
or UO_1624 (O_1624,N_24480,N_23647);
nor UO_1625 (O_1625,N_24437,N_24944);
and UO_1626 (O_1626,N_24175,N_23454);
and UO_1627 (O_1627,N_22901,N_22876);
or UO_1628 (O_1628,N_24495,N_24395);
or UO_1629 (O_1629,N_22972,N_23153);
or UO_1630 (O_1630,N_24536,N_23378);
xor UO_1631 (O_1631,N_23478,N_24894);
nor UO_1632 (O_1632,N_23898,N_23839);
nand UO_1633 (O_1633,N_24007,N_22962);
nor UO_1634 (O_1634,N_23155,N_22746);
nand UO_1635 (O_1635,N_24226,N_24102);
or UO_1636 (O_1636,N_23848,N_24408);
and UO_1637 (O_1637,N_22615,N_24459);
nor UO_1638 (O_1638,N_22984,N_24566);
nand UO_1639 (O_1639,N_22630,N_23402);
xor UO_1640 (O_1640,N_24483,N_23773);
xnor UO_1641 (O_1641,N_23275,N_22632);
nor UO_1642 (O_1642,N_24957,N_24853);
and UO_1643 (O_1643,N_23512,N_22586);
or UO_1644 (O_1644,N_23020,N_23681);
xnor UO_1645 (O_1645,N_23638,N_24730);
nor UO_1646 (O_1646,N_24803,N_24873);
nor UO_1647 (O_1647,N_23693,N_23291);
nand UO_1648 (O_1648,N_24123,N_23147);
xnor UO_1649 (O_1649,N_23602,N_23388);
xor UO_1650 (O_1650,N_24182,N_24947);
nor UO_1651 (O_1651,N_24626,N_24612);
nand UO_1652 (O_1652,N_23208,N_23635);
nand UO_1653 (O_1653,N_24108,N_22753);
xnor UO_1654 (O_1654,N_23238,N_24622);
or UO_1655 (O_1655,N_22797,N_24090);
nand UO_1656 (O_1656,N_24430,N_23381);
nor UO_1657 (O_1657,N_23970,N_22596);
or UO_1658 (O_1658,N_24465,N_24285);
or UO_1659 (O_1659,N_24849,N_24473);
and UO_1660 (O_1660,N_24023,N_22852);
and UO_1661 (O_1661,N_23744,N_24538);
xnor UO_1662 (O_1662,N_23382,N_24068);
or UO_1663 (O_1663,N_22937,N_23184);
xor UO_1664 (O_1664,N_23150,N_22814);
xnor UO_1665 (O_1665,N_23387,N_24500);
and UO_1666 (O_1666,N_24486,N_23401);
and UO_1667 (O_1667,N_24227,N_23354);
xnor UO_1668 (O_1668,N_24042,N_24479);
nor UO_1669 (O_1669,N_23643,N_23950);
or UO_1670 (O_1670,N_23226,N_24079);
and UO_1671 (O_1671,N_22840,N_22744);
or UO_1672 (O_1672,N_22947,N_24230);
and UO_1673 (O_1673,N_23279,N_24999);
or UO_1674 (O_1674,N_22662,N_23788);
and UO_1675 (O_1675,N_23455,N_24900);
and UO_1676 (O_1676,N_23098,N_23031);
or UO_1677 (O_1677,N_23137,N_24116);
nand UO_1678 (O_1678,N_24700,N_24618);
xnor UO_1679 (O_1679,N_22833,N_23605);
nor UO_1680 (O_1680,N_22690,N_22796);
or UO_1681 (O_1681,N_23481,N_23363);
and UO_1682 (O_1682,N_24157,N_24758);
or UO_1683 (O_1683,N_23679,N_24609);
nor UO_1684 (O_1684,N_23297,N_22708);
and UO_1685 (O_1685,N_22713,N_23580);
nor UO_1686 (O_1686,N_24851,N_24916);
and UO_1687 (O_1687,N_23771,N_24058);
or UO_1688 (O_1688,N_23431,N_24973);
or UO_1689 (O_1689,N_23612,N_23032);
nand UO_1690 (O_1690,N_24510,N_23629);
xnor UO_1691 (O_1691,N_23892,N_24576);
or UO_1692 (O_1692,N_22522,N_23756);
or UO_1693 (O_1693,N_22817,N_24260);
xnor UO_1694 (O_1694,N_24794,N_22849);
and UO_1695 (O_1695,N_23204,N_22891);
nand UO_1696 (O_1696,N_24317,N_24891);
nor UO_1697 (O_1697,N_24921,N_22665);
xor UO_1698 (O_1698,N_24185,N_24680);
or UO_1699 (O_1699,N_24292,N_23663);
nand UO_1700 (O_1700,N_24692,N_23587);
nor UO_1701 (O_1701,N_23216,N_24200);
and UO_1702 (O_1702,N_24729,N_24771);
nor UO_1703 (O_1703,N_22733,N_24966);
nor UO_1704 (O_1704,N_22755,N_24109);
or UO_1705 (O_1705,N_24177,N_23806);
nand UO_1706 (O_1706,N_23010,N_23779);
and UO_1707 (O_1707,N_22727,N_24759);
nand UO_1708 (O_1708,N_24475,N_22679);
nor UO_1709 (O_1709,N_24979,N_23557);
or UO_1710 (O_1710,N_23958,N_23417);
nand UO_1711 (O_1711,N_23266,N_24176);
nand UO_1712 (O_1712,N_24446,N_23948);
or UO_1713 (O_1713,N_23265,N_22761);
nor UO_1714 (O_1714,N_22902,N_24991);
or UO_1715 (O_1715,N_22510,N_24117);
or UO_1716 (O_1716,N_24489,N_24958);
and UO_1717 (O_1717,N_24968,N_23395);
nor UO_1718 (O_1718,N_23294,N_24714);
nand UO_1719 (O_1719,N_22557,N_22949);
nor UO_1720 (O_1720,N_24245,N_24866);
or UO_1721 (O_1721,N_24058,N_23302);
or UO_1722 (O_1722,N_22652,N_23802);
nor UO_1723 (O_1723,N_23871,N_23410);
nor UO_1724 (O_1724,N_24352,N_23209);
xor UO_1725 (O_1725,N_24734,N_24545);
nand UO_1726 (O_1726,N_22930,N_24621);
or UO_1727 (O_1727,N_24504,N_22617);
and UO_1728 (O_1728,N_22722,N_24625);
nor UO_1729 (O_1729,N_22786,N_23125);
nor UO_1730 (O_1730,N_24818,N_24473);
nor UO_1731 (O_1731,N_24875,N_22774);
nand UO_1732 (O_1732,N_22956,N_22832);
or UO_1733 (O_1733,N_24024,N_23158);
nand UO_1734 (O_1734,N_23472,N_22823);
or UO_1735 (O_1735,N_22527,N_22727);
or UO_1736 (O_1736,N_23239,N_23346);
and UO_1737 (O_1737,N_24683,N_24414);
and UO_1738 (O_1738,N_24752,N_24142);
nor UO_1739 (O_1739,N_23301,N_23614);
nand UO_1740 (O_1740,N_24929,N_24304);
and UO_1741 (O_1741,N_23561,N_23588);
and UO_1742 (O_1742,N_23157,N_24130);
and UO_1743 (O_1743,N_24231,N_23991);
nand UO_1744 (O_1744,N_24856,N_24594);
nor UO_1745 (O_1745,N_24442,N_23329);
or UO_1746 (O_1746,N_23871,N_23185);
nor UO_1747 (O_1747,N_22583,N_22846);
and UO_1748 (O_1748,N_24834,N_23984);
nand UO_1749 (O_1749,N_22955,N_23164);
xor UO_1750 (O_1750,N_24630,N_24754);
nor UO_1751 (O_1751,N_23056,N_24939);
and UO_1752 (O_1752,N_22973,N_23190);
xnor UO_1753 (O_1753,N_23980,N_23549);
xnor UO_1754 (O_1754,N_22554,N_24977);
and UO_1755 (O_1755,N_24568,N_24513);
nand UO_1756 (O_1756,N_24943,N_23548);
nor UO_1757 (O_1757,N_23524,N_23761);
or UO_1758 (O_1758,N_24361,N_22543);
xnor UO_1759 (O_1759,N_22628,N_22674);
or UO_1760 (O_1760,N_24974,N_23395);
xnor UO_1761 (O_1761,N_24191,N_24338);
xnor UO_1762 (O_1762,N_24157,N_23542);
or UO_1763 (O_1763,N_22744,N_24451);
and UO_1764 (O_1764,N_22925,N_23927);
nand UO_1765 (O_1765,N_22734,N_23503);
nand UO_1766 (O_1766,N_22508,N_23114);
xor UO_1767 (O_1767,N_23636,N_22969);
xnor UO_1768 (O_1768,N_24621,N_23875);
nor UO_1769 (O_1769,N_23798,N_23678);
nor UO_1770 (O_1770,N_24627,N_22515);
and UO_1771 (O_1771,N_23270,N_23140);
nor UO_1772 (O_1772,N_24900,N_23071);
or UO_1773 (O_1773,N_23937,N_22968);
and UO_1774 (O_1774,N_23636,N_23114);
nand UO_1775 (O_1775,N_23684,N_24707);
and UO_1776 (O_1776,N_24354,N_23996);
and UO_1777 (O_1777,N_24911,N_23864);
nor UO_1778 (O_1778,N_24970,N_22619);
and UO_1779 (O_1779,N_22963,N_23523);
and UO_1780 (O_1780,N_24279,N_24797);
or UO_1781 (O_1781,N_23187,N_23976);
or UO_1782 (O_1782,N_24481,N_22930);
nand UO_1783 (O_1783,N_24923,N_23908);
nor UO_1784 (O_1784,N_22935,N_23477);
nor UO_1785 (O_1785,N_23078,N_24080);
or UO_1786 (O_1786,N_23900,N_23315);
nand UO_1787 (O_1787,N_22577,N_23464);
and UO_1788 (O_1788,N_23121,N_24231);
xor UO_1789 (O_1789,N_24585,N_23128);
or UO_1790 (O_1790,N_23370,N_24391);
nor UO_1791 (O_1791,N_23020,N_23273);
and UO_1792 (O_1792,N_24567,N_22959);
xnor UO_1793 (O_1793,N_23796,N_24325);
or UO_1794 (O_1794,N_24344,N_24364);
or UO_1795 (O_1795,N_24357,N_22704);
xnor UO_1796 (O_1796,N_24401,N_22906);
nor UO_1797 (O_1797,N_23275,N_23195);
nor UO_1798 (O_1798,N_23527,N_23729);
nand UO_1799 (O_1799,N_24447,N_23135);
and UO_1800 (O_1800,N_22521,N_23731);
xnor UO_1801 (O_1801,N_23979,N_23491);
or UO_1802 (O_1802,N_22904,N_24818);
xor UO_1803 (O_1803,N_24534,N_22567);
and UO_1804 (O_1804,N_22748,N_23008);
and UO_1805 (O_1805,N_24817,N_24593);
xnor UO_1806 (O_1806,N_23221,N_24999);
nand UO_1807 (O_1807,N_24568,N_24356);
and UO_1808 (O_1808,N_24041,N_23521);
nand UO_1809 (O_1809,N_23950,N_23489);
nand UO_1810 (O_1810,N_24770,N_24521);
nor UO_1811 (O_1811,N_22521,N_24453);
xor UO_1812 (O_1812,N_24685,N_23067);
xor UO_1813 (O_1813,N_23414,N_24073);
or UO_1814 (O_1814,N_24318,N_22722);
or UO_1815 (O_1815,N_24859,N_24550);
nor UO_1816 (O_1816,N_23293,N_23460);
nand UO_1817 (O_1817,N_24799,N_24235);
nand UO_1818 (O_1818,N_22968,N_24627);
xor UO_1819 (O_1819,N_23350,N_24518);
and UO_1820 (O_1820,N_23545,N_24410);
and UO_1821 (O_1821,N_22729,N_23801);
nor UO_1822 (O_1822,N_22644,N_23969);
xor UO_1823 (O_1823,N_24532,N_23676);
and UO_1824 (O_1824,N_22508,N_24414);
xor UO_1825 (O_1825,N_23710,N_23633);
nor UO_1826 (O_1826,N_22786,N_23700);
nor UO_1827 (O_1827,N_24470,N_23213);
nor UO_1828 (O_1828,N_23212,N_24865);
xor UO_1829 (O_1829,N_24477,N_24879);
nand UO_1830 (O_1830,N_23462,N_23642);
or UO_1831 (O_1831,N_24120,N_24800);
nor UO_1832 (O_1832,N_23977,N_24329);
xnor UO_1833 (O_1833,N_24832,N_24883);
and UO_1834 (O_1834,N_24616,N_24780);
nand UO_1835 (O_1835,N_24438,N_23831);
or UO_1836 (O_1836,N_24465,N_24734);
or UO_1837 (O_1837,N_23203,N_24938);
and UO_1838 (O_1838,N_23716,N_24332);
xor UO_1839 (O_1839,N_23504,N_24314);
and UO_1840 (O_1840,N_24326,N_23349);
xnor UO_1841 (O_1841,N_23008,N_24594);
nor UO_1842 (O_1842,N_24050,N_23713);
xnor UO_1843 (O_1843,N_24233,N_23428);
and UO_1844 (O_1844,N_23622,N_22534);
nor UO_1845 (O_1845,N_24114,N_23431);
or UO_1846 (O_1846,N_24778,N_24685);
and UO_1847 (O_1847,N_23370,N_24279);
nor UO_1848 (O_1848,N_22882,N_24928);
nand UO_1849 (O_1849,N_23364,N_24487);
nor UO_1850 (O_1850,N_24077,N_23828);
nand UO_1851 (O_1851,N_23876,N_24850);
or UO_1852 (O_1852,N_23915,N_22871);
nand UO_1853 (O_1853,N_24928,N_23192);
nor UO_1854 (O_1854,N_23004,N_24825);
or UO_1855 (O_1855,N_23281,N_22611);
or UO_1856 (O_1856,N_24220,N_24782);
xor UO_1857 (O_1857,N_23149,N_24885);
nor UO_1858 (O_1858,N_24291,N_24791);
and UO_1859 (O_1859,N_23757,N_24719);
nand UO_1860 (O_1860,N_23581,N_24189);
or UO_1861 (O_1861,N_24696,N_23275);
and UO_1862 (O_1862,N_24621,N_23068);
xor UO_1863 (O_1863,N_24257,N_24290);
and UO_1864 (O_1864,N_22987,N_24055);
and UO_1865 (O_1865,N_23749,N_23996);
nor UO_1866 (O_1866,N_24190,N_24327);
nand UO_1867 (O_1867,N_23390,N_23945);
or UO_1868 (O_1868,N_24945,N_22526);
nand UO_1869 (O_1869,N_23669,N_24266);
xnor UO_1870 (O_1870,N_23783,N_23515);
and UO_1871 (O_1871,N_23571,N_22746);
and UO_1872 (O_1872,N_24809,N_23555);
nand UO_1873 (O_1873,N_24416,N_22532);
and UO_1874 (O_1874,N_23536,N_24697);
or UO_1875 (O_1875,N_24076,N_22688);
nand UO_1876 (O_1876,N_23349,N_24376);
nor UO_1877 (O_1877,N_23095,N_24069);
nand UO_1878 (O_1878,N_24128,N_22653);
nand UO_1879 (O_1879,N_24327,N_23504);
xnor UO_1880 (O_1880,N_24182,N_23872);
and UO_1881 (O_1881,N_23655,N_22962);
nand UO_1882 (O_1882,N_23624,N_24892);
and UO_1883 (O_1883,N_22826,N_22975);
or UO_1884 (O_1884,N_23208,N_22507);
nor UO_1885 (O_1885,N_24006,N_23244);
nor UO_1886 (O_1886,N_22625,N_23664);
nand UO_1887 (O_1887,N_22645,N_24265);
nor UO_1888 (O_1888,N_24135,N_24197);
xnor UO_1889 (O_1889,N_23006,N_23048);
and UO_1890 (O_1890,N_22831,N_23872);
nor UO_1891 (O_1891,N_23520,N_24622);
xor UO_1892 (O_1892,N_22991,N_22867);
nor UO_1893 (O_1893,N_24607,N_24338);
nand UO_1894 (O_1894,N_22639,N_24900);
nor UO_1895 (O_1895,N_24775,N_23892);
and UO_1896 (O_1896,N_23696,N_23961);
nand UO_1897 (O_1897,N_23629,N_23125);
nand UO_1898 (O_1898,N_24382,N_23169);
or UO_1899 (O_1899,N_23259,N_23832);
nor UO_1900 (O_1900,N_22850,N_23995);
and UO_1901 (O_1901,N_23364,N_22741);
nand UO_1902 (O_1902,N_24404,N_23286);
nand UO_1903 (O_1903,N_23391,N_24621);
nand UO_1904 (O_1904,N_24626,N_24009);
and UO_1905 (O_1905,N_22553,N_24290);
and UO_1906 (O_1906,N_24949,N_24925);
or UO_1907 (O_1907,N_24925,N_23900);
nor UO_1908 (O_1908,N_23134,N_23757);
or UO_1909 (O_1909,N_22862,N_22955);
nor UO_1910 (O_1910,N_22557,N_23529);
and UO_1911 (O_1911,N_24287,N_23779);
nor UO_1912 (O_1912,N_24189,N_23841);
and UO_1913 (O_1913,N_23475,N_24205);
and UO_1914 (O_1914,N_24451,N_23694);
or UO_1915 (O_1915,N_23069,N_23412);
and UO_1916 (O_1916,N_22799,N_23584);
and UO_1917 (O_1917,N_23117,N_24897);
and UO_1918 (O_1918,N_24612,N_24331);
nand UO_1919 (O_1919,N_23772,N_24472);
xnor UO_1920 (O_1920,N_24956,N_22592);
nor UO_1921 (O_1921,N_23604,N_22896);
xor UO_1922 (O_1922,N_23138,N_23296);
or UO_1923 (O_1923,N_23274,N_24815);
nand UO_1924 (O_1924,N_23754,N_23231);
and UO_1925 (O_1925,N_24341,N_23163);
xnor UO_1926 (O_1926,N_24817,N_22555);
or UO_1927 (O_1927,N_23511,N_23869);
nor UO_1928 (O_1928,N_24805,N_22629);
xnor UO_1929 (O_1929,N_22738,N_24270);
or UO_1930 (O_1930,N_24028,N_23698);
nand UO_1931 (O_1931,N_24557,N_24208);
or UO_1932 (O_1932,N_24914,N_22726);
nor UO_1933 (O_1933,N_23035,N_22677);
and UO_1934 (O_1934,N_24826,N_22979);
nor UO_1935 (O_1935,N_23327,N_22813);
or UO_1936 (O_1936,N_22697,N_22534);
and UO_1937 (O_1937,N_23484,N_24847);
or UO_1938 (O_1938,N_24890,N_24351);
nor UO_1939 (O_1939,N_24206,N_24628);
and UO_1940 (O_1940,N_24117,N_23824);
and UO_1941 (O_1941,N_23582,N_24910);
or UO_1942 (O_1942,N_23578,N_23496);
and UO_1943 (O_1943,N_23485,N_22674);
nand UO_1944 (O_1944,N_23663,N_24266);
nand UO_1945 (O_1945,N_23325,N_22656);
nand UO_1946 (O_1946,N_24015,N_24480);
or UO_1947 (O_1947,N_22626,N_22590);
or UO_1948 (O_1948,N_24744,N_24795);
xnor UO_1949 (O_1949,N_23738,N_24166);
or UO_1950 (O_1950,N_24276,N_23953);
nor UO_1951 (O_1951,N_22532,N_24625);
nor UO_1952 (O_1952,N_23538,N_24336);
or UO_1953 (O_1953,N_24520,N_24406);
nor UO_1954 (O_1954,N_23630,N_24976);
and UO_1955 (O_1955,N_23981,N_24128);
xor UO_1956 (O_1956,N_23086,N_24111);
xor UO_1957 (O_1957,N_24975,N_23621);
xor UO_1958 (O_1958,N_23872,N_22915);
nor UO_1959 (O_1959,N_24378,N_23755);
xor UO_1960 (O_1960,N_22545,N_24406);
or UO_1961 (O_1961,N_23960,N_24100);
nand UO_1962 (O_1962,N_23700,N_24396);
or UO_1963 (O_1963,N_22671,N_23452);
nor UO_1964 (O_1964,N_24572,N_22785);
nor UO_1965 (O_1965,N_22816,N_23103);
nor UO_1966 (O_1966,N_24759,N_22847);
xor UO_1967 (O_1967,N_24486,N_24157);
and UO_1968 (O_1968,N_23841,N_24044);
or UO_1969 (O_1969,N_23037,N_22553);
xnor UO_1970 (O_1970,N_23002,N_22866);
nand UO_1971 (O_1971,N_24514,N_24493);
and UO_1972 (O_1972,N_23157,N_24595);
nand UO_1973 (O_1973,N_23552,N_24578);
and UO_1974 (O_1974,N_22508,N_24385);
xor UO_1975 (O_1975,N_23791,N_24684);
or UO_1976 (O_1976,N_23605,N_23134);
nand UO_1977 (O_1977,N_23074,N_23994);
nand UO_1978 (O_1978,N_23156,N_24430);
and UO_1979 (O_1979,N_23956,N_24726);
nand UO_1980 (O_1980,N_24223,N_23259);
xnor UO_1981 (O_1981,N_23871,N_24667);
or UO_1982 (O_1982,N_22992,N_22507);
and UO_1983 (O_1983,N_22504,N_23090);
or UO_1984 (O_1984,N_24763,N_24425);
xor UO_1985 (O_1985,N_24888,N_22774);
nand UO_1986 (O_1986,N_23909,N_22545);
nor UO_1987 (O_1987,N_22738,N_24075);
nor UO_1988 (O_1988,N_24064,N_24116);
or UO_1989 (O_1989,N_24135,N_22615);
or UO_1990 (O_1990,N_23887,N_24987);
nor UO_1991 (O_1991,N_24590,N_22502);
nor UO_1992 (O_1992,N_23657,N_24304);
xnor UO_1993 (O_1993,N_22778,N_24973);
xor UO_1994 (O_1994,N_24447,N_23952);
and UO_1995 (O_1995,N_23090,N_23629);
and UO_1996 (O_1996,N_24074,N_24262);
and UO_1997 (O_1997,N_22930,N_24376);
nor UO_1998 (O_1998,N_23698,N_24585);
xor UO_1999 (O_1999,N_24062,N_23843);
nand UO_2000 (O_2000,N_23777,N_23441);
or UO_2001 (O_2001,N_24186,N_23832);
and UO_2002 (O_2002,N_23516,N_22999);
or UO_2003 (O_2003,N_23681,N_23533);
or UO_2004 (O_2004,N_24344,N_22960);
nor UO_2005 (O_2005,N_23475,N_24522);
or UO_2006 (O_2006,N_24079,N_24181);
or UO_2007 (O_2007,N_23271,N_23814);
xnor UO_2008 (O_2008,N_22663,N_23124);
and UO_2009 (O_2009,N_23123,N_23118);
nor UO_2010 (O_2010,N_22765,N_23679);
nand UO_2011 (O_2011,N_23843,N_24714);
and UO_2012 (O_2012,N_23170,N_24072);
and UO_2013 (O_2013,N_24162,N_22694);
nand UO_2014 (O_2014,N_24686,N_24965);
or UO_2015 (O_2015,N_23291,N_24949);
nand UO_2016 (O_2016,N_23059,N_23406);
or UO_2017 (O_2017,N_23377,N_23102);
xnor UO_2018 (O_2018,N_23219,N_22623);
and UO_2019 (O_2019,N_22894,N_24609);
or UO_2020 (O_2020,N_23454,N_24330);
nand UO_2021 (O_2021,N_22847,N_23334);
or UO_2022 (O_2022,N_22703,N_24323);
and UO_2023 (O_2023,N_24293,N_24489);
xor UO_2024 (O_2024,N_24279,N_24540);
xnor UO_2025 (O_2025,N_24783,N_24141);
nor UO_2026 (O_2026,N_24900,N_22837);
or UO_2027 (O_2027,N_24752,N_24096);
nor UO_2028 (O_2028,N_23938,N_24238);
nor UO_2029 (O_2029,N_24967,N_23442);
and UO_2030 (O_2030,N_22885,N_22814);
or UO_2031 (O_2031,N_24157,N_23726);
nor UO_2032 (O_2032,N_24190,N_23207);
and UO_2033 (O_2033,N_24614,N_24518);
nor UO_2034 (O_2034,N_24818,N_22556);
nor UO_2035 (O_2035,N_23716,N_23350);
xor UO_2036 (O_2036,N_23038,N_23046);
or UO_2037 (O_2037,N_22545,N_24198);
or UO_2038 (O_2038,N_24131,N_22560);
xnor UO_2039 (O_2039,N_23017,N_24925);
and UO_2040 (O_2040,N_24782,N_24226);
xnor UO_2041 (O_2041,N_23370,N_22500);
nand UO_2042 (O_2042,N_24396,N_24229);
nor UO_2043 (O_2043,N_24237,N_23411);
and UO_2044 (O_2044,N_24721,N_24921);
nand UO_2045 (O_2045,N_23689,N_22525);
and UO_2046 (O_2046,N_23621,N_24973);
nor UO_2047 (O_2047,N_23528,N_23531);
and UO_2048 (O_2048,N_23048,N_24058);
nand UO_2049 (O_2049,N_22587,N_22625);
or UO_2050 (O_2050,N_23639,N_23217);
nor UO_2051 (O_2051,N_22863,N_23140);
or UO_2052 (O_2052,N_23808,N_24036);
or UO_2053 (O_2053,N_23993,N_22698);
or UO_2054 (O_2054,N_23599,N_24620);
nand UO_2055 (O_2055,N_22916,N_22594);
or UO_2056 (O_2056,N_23754,N_23100);
and UO_2057 (O_2057,N_24857,N_23870);
xnor UO_2058 (O_2058,N_24545,N_22843);
nand UO_2059 (O_2059,N_23055,N_22836);
nand UO_2060 (O_2060,N_23069,N_24456);
and UO_2061 (O_2061,N_23706,N_24769);
or UO_2062 (O_2062,N_24995,N_23876);
nand UO_2063 (O_2063,N_23640,N_24684);
and UO_2064 (O_2064,N_23465,N_23861);
or UO_2065 (O_2065,N_22710,N_22966);
nand UO_2066 (O_2066,N_23110,N_24072);
and UO_2067 (O_2067,N_24255,N_24334);
nand UO_2068 (O_2068,N_24055,N_24359);
nor UO_2069 (O_2069,N_24366,N_23816);
nand UO_2070 (O_2070,N_24482,N_23136);
nor UO_2071 (O_2071,N_24792,N_22852);
and UO_2072 (O_2072,N_24360,N_23266);
or UO_2073 (O_2073,N_24351,N_23951);
nor UO_2074 (O_2074,N_23279,N_24116);
or UO_2075 (O_2075,N_24104,N_24861);
and UO_2076 (O_2076,N_23664,N_22824);
or UO_2077 (O_2077,N_24015,N_22876);
nand UO_2078 (O_2078,N_24272,N_24855);
nand UO_2079 (O_2079,N_23845,N_24029);
and UO_2080 (O_2080,N_24302,N_22847);
or UO_2081 (O_2081,N_23453,N_24243);
xnor UO_2082 (O_2082,N_23601,N_23104);
or UO_2083 (O_2083,N_23758,N_24591);
nand UO_2084 (O_2084,N_24125,N_24360);
or UO_2085 (O_2085,N_24929,N_24312);
xnor UO_2086 (O_2086,N_22780,N_23844);
and UO_2087 (O_2087,N_22506,N_23202);
xor UO_2088 (O_2088,N_22888,N_23159);
and UO_2089 (O_2089,N_22762,N_24174);
or UO_2090 (O_2090,N_23937,N_22733);
nand UO_2091 (O_2091,N_23202,N_24432);
nor UO_2092 (O_2092,N_23612,N_23901);
or UO_2093 (O_2093,N_24694,N_24039);
nand UO_2094 (O_2094,N_23924,N_23710);
nand UO_2095 (O_2095,N_24292,N_23730);
xnor UO_2096 (O_2096,N_24150,N_22924);
nand UO_2097 (O_2097,N_22807,N_23119);
xor UO_2098 (O_2098,N_22764,N_22729);
xnor UO_2099 (O_2099,N_24183,N_23413);
or UO_2100 (O_2100,N_23905,N_22586);
nor UO_2101 (O_2101,N_23983,N_23595);
xor UO_2102 (O_2102,N_22550,N_24582);
or UO_2103 (O_2103,N_24761,N_23403);
and UO_2104 (O_2104,N_23986,N_23442);
xor UO_2105 (O_2105,N_24885,N_22605);
xor UO_2106 (O_2106,N_23909,N_24036);
nor UO_2107 (O_2107,N_24277,N_24114);
and UO_2108 (O_2108,N_23950,N_24916);
xnor UO_2109 (O_2109,N_24911,N_22703);
and UO_2110 (O_2110,N_24861,N_24953);
or UO_2111 (O_2111,N_23753,N_22609);
nor UO_2112 (O_2112,N_24044,N_22663);
nor UO_2113 (O_2113,N_22708,N_23065);
and UO_2114 (O_2114,N_24106,N_24891);
and UO_2115 (O_2115,N_23608,N_24066);
nor UO_2116 (O_2116,N_24746,N_23483);
and UO_2117 (O_2117,N_24735,N_24162);
nor UO_2118 (O_2118,N_24727,N_24958);
and UO_2119 (O_2119,N_23067,N_23852);
nand UO_2120 (O_2120,N_22982,N_24870);
xor UO_2121 (O_2121,N_23050,N_24848);
nand UO_2122 (O_2122,N_23577,N_22793);
nor UO_2123 (O_2123,N_24455,N_23763);
and UO_2124 (O_2124,N_24976,N_23189);
xor UO_2125 (O_2125,N_23264,N_23524);
or UO_2126 (O_2126,N_24048,N_23896);
and UO_2127 (O_2127,N_23633,N_24683);
and UO_2128 (O_2128,N_24673,N_24064);
or UO_2129 (O_2129,N_24001,N_22723);
nand UO_2130 (O_2130,N_22741,N_22902);
xnor UO_2131 (O_2131,N_24078,N_23030);
and UO_2132 (O_2132,N_24674,N_24557);
or UO_2133 (O_2133,N_23350,N_24732);
nand UO_2134 (O_2134,N_23567,N_24079);
xor UO_2135 (O_2135,N_24014,N_24459);
xor UO_2136 (O_2136,N_24923,N_23600);
and UO_2137 (O_2137,N_22511,N_24903);
nand UO_2138 (O_2138,N_23217,N_23988);
xnor UO_2139 (O_2139,N_23129,N_24057);
and UO_2140 (O_2140,N_24731,N_24393);
nor UO_2141 (O_2141,N_22898,N_22654);
and UO_2142 (O_2142,N_22924,N_23656);
xor UO_2143 (O_2143,N_24141,N_23225);
nand UO_2144 (O_2144,N_24286,N_22925);
nand UO_2145 (O_2145,N_23783,N_23895);
or UO_2146 (O_2146,N_23753,N_24095);
nor UO_2147 (O_2147,N_22921,N_23061);
xnor UO_2148 (O_2148,N_22912,N_22576);
xor UO_2149 (O_2149,N_24915,N_23334);
and UO_2150 (O_2150,N_22621,N_23273);
nand UO_2151 (O_2151,N_23919,N_24129);
nor UO_2152 (O_2152,N_23333,N_24158);
or UO_2153 (O_2153,N_22723,N_24928);
xnor UO_2154 (O_2154,N_23453,N_23157);
xnor UO_2155 (O_2155,N_24742,N_23887);
nand UO_2156 (O_2156,N_24772,N_22917);
nor UO_2157 (O_2157,N_23912,N_23495);
and UO_2158 (O_2158,N_24951,N_22731);
and UO_2159 (O_2159,N_23020,N_23570);
xor UO_2160 (O_2160,N_24256,N_24349);
nand UO_2161 (O_2161,N_23416,N_23848);
and UO_2162 (O_2162,N_23998,N_23180);
and UO_2163 (O_2163,N_22767,N_23610);
nand UO_2164 (O_2164,N_23408,N_22595);
nor UO_2165 (O_2165,N_24819,N_24494);
and UO_2166 (O_2166,N_22646,N_23023);
nor UO_2167 (O_2167,N_23689,N_22641);
xnor UO_2168 (O_2168,N_24005,N_24344);
nor UO_2169 (O_2169,N_24556,N_22955);
nor UO_2170 (O_2170,N_24187,N_24273);
nand UO_2171 (O_2171,N_23681,N_24477);
nand UO_2172 (O_2172,N_23803,N_22789);
nand UO_2173 (O_2173,N_24268,N_24598);
and UO_2174 (O_2174,N_22866,N_23850);
nor UO_2175 (O_2175,N_23621,N_24503);
nand UO_2176 (O_2176,N_24513,N_22569);
nand UO_2177 (O_2177,N_23575,N_24987);
and UO_2178 (O_2178,N_24659,N_23574);
xnor UO_2179 (O_2179,N_23689,N_23789);
or UO_2180 (O_2180,N_24038,N_24859);
and UO_2181 (O_2181,N_23234,N_24806);
and UO_2182 (O_2182,N_23902,N_24779);
or UO_2183 (O_2183,N_24743,N_24129);
or UO_2184 (O_2184,N_24303,N_22562);
or UO_2185 (O_2185,N_24034,N_23482);
nor UO_2186 (O_2186,N_23794,N_22617);
or UO_2187 (O_2187,N_23121,N_24488);
xor UO_2188 (O_2188,N_24678,N_24095);
or UO_2189 (O_2189,N_24827,N_23555);
xnor UO_2190 (O_2190,N_23275,N_24457);
nand UO_2191 (O_2191,N_24190,N_22935);
or UO_2192 (O_2192,N_23786,N_24800);
nor UO_2193 (O_2193,N_23071,N_23347);
or UO_2194 (O_2194,N_22996,N_22862);
and UO_2195 (O_2195,N_24692,N_23814);
and UO_2196 (O_2196,N_22853,N_23936);
nand UO_2197 (O_2197,N_22726,N_23667);
nand UO_2198 (O_2198,N_23060,N_23347);
nor UO_2199 (O_2199,N_22945,N_22920);
or UO_2200 (O_2200,N_24412,N_23633);
or UO_2201 (O_2201,N_22822,N_24546);
nor UO_2202 (O_2202,N_23385,N_23842);
and UO_2203 (O_2203,N_24742,N_22949);
and UO_2204 (O_2204,N_24764,N_23184);
and UO_2205 (O_2205,N_24785,N_24047);
nand UO_2206 (O_2206,N_23604,N_24026);
xor UO_2207 (O_2207,N_23329,N_22604);
and UO_2208 (O_2208,N_23243,N_22601);
nor UO_2209 (O_2209,N_22680,N_23321);
and UO_2210 (O_2210,N_24873,N_22913);
or UO_2211 (O_2211,N_24235,N_24686);
and UO_2212 (O_2212,N_23642,N_24763);
nor UO_2213 (O_2213,N_24042,N_24877);
nand UO_2214 (O_2214,N_23641,N_23374);
xnor UO_2215 (O_2215,N_24575,N_22548);
or UO_2216 (O_2216,N_24290,N_23376);
nor UO_2217 (O_2217,N_24034,N_24055);
nand UO_2218 (O_2218,N_24159,N_22689);
or UO_2219 (O_2219,N_24306,N_23162);
or UO_2220 (O_2220,N_24574,N_24759);
nor UO_2221 (O_2221,N_22784,N_22734);
or UO_2222 (O_2222,N_23513,N_23452);
nor UO_2223 (O_2223,N_24313,N_23050);
nand UO_2224 (O_2224,N_23466,N_24970);
nand UO_2225 (O_2225,N_23862,N_24506);
nor UO_2226 (O_2226,N_24112,N_23803);
nand UO_2227 (O_2227,N_24985,N_22938);
xnor UO_2228 (O_2228,N_22521,N_24518);
or UO_2229 (O_2229,N_23903,N_24842);
or UO_2230 (O_2230,N_22749,N_23936);
xnor UO_2231 (O_2231,N_23242,N_22847);
xnor UO_2232 (O_2232,N_22548,N_24566);
xnor UO_2233 (O_2233,N_24954,N_22959);
nor UO_2234 (O_2234,N_23335,N_23996);
nor UO_2235 (O_2235,N_24580,N_23400);
or UO_2236 (O_2236,N_23661,N_23532);
or UO_2237 (O_2237,N_23121,N_24670);
nor UO_2238 (O_2238,N_24257,N_23894);
or UO_2239 (O_2239,N_23103,N_22523);
xnor UO_2240 (O_2240,N_24807,N_22560);
and UO_2241 (O_2241,N_23919,N_22788);
and UO_2242 (O_2242,N_24128,N_24146);
nand UO_2243 (O_2243,N_24174,N_24425);
and UO_2244 (O_2244,N_22690,N_23850);
nand UO_2245 (O_2245,N_22565,N_24620);
nand UO_2246 (O_2246,N_24644,N_24404);
xnor UO_2247 (O_2247,N_22917,N_22557);
or UO_2248 (O_2248,N_24735,N_24909);
and UO_2249 (O_2249,N_22736,N_24948);
nand UO_2250 (O_2250,N_24562,N_22861);
or UO_2251 (O_2251,N_22772,N_24836);
or UO_2252 (O_2252,N_24294,N_23135);
and UO_2253 (O_2253,N_22580,N_22582);
nor UO_2254 (O_2254,N_23871,N_23704);
or UO_2255 (O_2255,N_24598,N_23285);
xnor UO_2256 (O_2256,N_24985,N_22906);
nand UO_2257 (O_2257,N_22627,N_22588);
or UO_2258 (O_2258,N_22534,N_23022);
nor UO_2259 (O_2259,N_23856,N_22832);
nand UO_2260 (O_2260,N_22578,N_23635);
xnor UO_2261 (O_2261,N_24429,N_22699);
nor UO_2262 (O_2262,N_22578,N_24399);
nor UO_2263 (O_2263,N_22688,N_24074);
nand UO_2264 (O_2264,N_23989,N_24420);
and UO_2265 (O_2265,N_24345,N_22677);
nor UO_2266 (O_2266,N_24666,N_23685);
nand UO_2267 (O_2267,N_24424,N_23703);
and UO_2268 (O_2268,N_22776,N_24655);
and UO_2269 (O_2269,N_23181,N_24943);
nor UO_2270 (O_2270,N_23434,N_23421);
xor UO_2271 (O_2271,N_23103,N_22792);
nor UO_2272 (O_2272,N_24140,N_23589);
and UO_2273 (O_2273,N_24034,N_23605);
and UO_2274 (O_2274,N_23072,N_24101);
and UO_2275 (O_2275,N_24472,N_24730);
or UO_2276 (O_2276,N_24087,N_23216);
nor UO_2277 (O_2277,N_23827,N_23950);
nor UO_2278 (O_2278,N_22898,N_24592);
xor UO_2279 (O_2279,N_24451,N_23433);
xnor UO_2280 (O_2280,N_24642,N_23497);
and UO_2281 (O_2281,N_24261,N_24836);
xnor UO_2282 (O_2282,N_24936,N_24902);
and UO_2283 (O_2283,N_22723,N_24614);
xor UO_2284 (O_2284,N_23813,N_24895);
and UO_2285 (O_2285,N_23064,N_24128);
xor UO_2286 (O_2286,N_24498,N_22770);
nand UO_2287 (O_2287,N_23473,N_24313);
nor UO_2288 (O_2288,N_23824,N_22523);
xor UO_2289 (O_2289,N_23986,N_23726);
nor UO_2290 (O_2290,N_24985,N_22687);
and UO_2291 (O_2291,N_24096,N_24334);
nor UO_2292 (O_2292,N_24074,N_24057);
nand UO_2293 (O_2293,N_23348,N_24453);
nor UO_2294 (O_2294,N_24559,N_23347);
xor UO_2295 (O_2295,N_24800,N_24113);
xor UO_2296 (O_2296,N_24857,N_23110);
or UO_2297 (O_2297,N_23865,N_23445);
or UO_2298 (O_2298,N_22974,N_22957);
and UO_2299 (O_2299,N_22695,N_23494);
xor UO_2300 (O_2300,N_22888,N_23308);
nand UO_2301 (O_2301,N_22828,N_23820);
or UO_2302 (O_2302,N_24370,N_23563);
nand UO_2303 (O_2303,N_24879,N_24334);
nand UO_2304 (O_2304,N_24134,N_23777);
nor UO_2305 (O_2305,N_24155,N_24323);
xor UO_2306 (O_2306,N_22766,N_24932);
nor UO_2307 (O_2307,N_24275,N_24817);
nand UO_2308 (O_2308,N_22890,N_24859);
or UO_2309 (O_2309,N_24124,N_24140);
xnor UO_2310 (O_2310,N_23979,N_23729);
nor UO_2311 (O_2311,N_24943,N_23047);
nand UO_2312 (O_2312,N_24042,N_24104);
nor UO_2313 (O_2313,N_22790,N_23121);
xnor UO_2314 (O_2314,N_24750,N_23086);
nor UO_2315 (O_2315,N_22786,N_22503);
nor UO_2316 (O_2316,N_23864,N_23601);
or UO_2317 (O_2317,N_22827,N_22510);
xor UO_2318 (O_2318,N_22507,N_23906);
and UO_2319 (O_2319,N_22762,N_23727);
and UO_2320 (O_2320,N_22738,N_23123);
nor UO_2321 (O_2321,N_24234,N_23096);
and UO_2322 (O_2322,N_23423,N_22546);
nand UO_2323 (O_2323,N_24296,N_24722);
or UO_2324 (O_2324,N_23440,N_24280);
or UO_2325 (O_2325,N_22788,N_23500);
nand UO_2326 (O_2326,N_23409,N_23733);
nand UO_2327 (O_2327,N_22995,N_24421);
or UO_2328 (O_2328,N_24736,N_23305);
nor UO_2329 (O_2329,N_23572,N_24867);
nand UO_2330 (O_2330,N_24813,N_23063);
xor UO_2331 (O_2331,N_23724,N_23060);
nand UO_2332 (O_2332,N_24244,N_22885);
xnor UO_2333 (O_2333,N_23166,N_22948);
nor UO_2334 (O_2334,N_24103,N_23579);
nor UO_2335 (O_2335,N_23288,N_23393);
and UO_2336 (O_2336,N_24127,N_22504);
xnor UO_2337 (O_2337,N_23232,N_23416);
and UO_2338 (O_2338,N_22912,N_22703);
nand UO_2339 (O_2339,N_23536,N_22898);
or UO_2340 (O_2340,N_24765,N_22592);
or UO_2341 (O_2341,N_22658,N_23140);
and UO_2342 (O_2342,N_24811,N_23852);
nand UO_2343 (O_2343,N_23378,N_22507);
or UO_2344 (O_2344,N_23846,N_23448);
or UO_2345 (O_2345,N_22892,N_23792);
nor UO_2346 (O_2346,N_23368,N_24852);
or UO_2347 (O_2347,N_24610,N_22564);
and UO_2348 (O_2348,N_24197,N_24503);
or UO_2349 (O_2349,N_23961,N_24187);
and UO_2350 (O_2350,N_23151,N_23193);
nor UO_2351 (O_2351,N_24198,N_22567);
nor UO_2352 (O_2352,N_23263,N_24728);
xnor UO_2353 (O_2353,N_24090,N_24686);
nor UO_2354 (O_2354,N_22658,N_22825);
xor UO_2355 (O_2355,N_23974,N_23279);
and UO_2356 (O_2356,N_23518,N_24627);
or UO_2357 (O_2357,N_24049,N_24118);
or UO_2358 (O_2358,N_23154,N_24547);
nand UO_2359 (O_2359,N_23760,N_23318);
nand UO_2360 (O_2360,N_24211,N_23793);
xor UO_2361 (O_2361,N_23920,N_23990);
or UO_2362 (O_2362,N_24097,N_24877);
nand UO_2363 (O_2363,N_23024,N_23667);
or UO_2364 (O_2364,N_23099,N_22565);
xor UO_2365 (O_2365,N_24767,N_22678);
and UO_2366 (O_2366,N_22875,N_23767);
and UO_2367 (O_2367,N_23246,N_23592);
nor UO_2368 (O_2368,N_22772,N_24956);
nand UO_2369 (O_2369,N_23528,N_23082);
or UO_2370 (O_2370,N_23162,N_24839);
and UO_2371 (O_2371,N_23097,N_23650);
nand UO_2372 (O_2372,N_23506,N_24047);
or UO_2373 (O_2373,N_23199,N_23752);
xnor UO_2374 (O_2374,N_24180,N_23973);
or UO_2375 (O_2375,N_23937,N_23689);
xor UO_2376 (O_2376,N_23703,N_24352);
and UO_2377 (O_2377,N_23982,N_24545);
nor UO_2378 (O_2378,N_24115,N_22665);
xnor UO_2379 (O_2379,N_22871,N_23587);
xnor UO_2380 (O_2380,N_23778,N_23175);
and UO_2381 (O_2381,N_24906,N_24734);
nor UO_2382 (O_2382,N_23395,N_23151);
nor UO_2383 (O_2383,N_24069,N_24052);
nand UO_2384 (O_2384,N_23403,N_23549);
or UO_2385 (O_2385,N_22815,N_24135);
xnor UO_2386 (O_2386,N_24398,N_22814);
nor UO_2387 (O_2387,N_24242,N_23826);
and UO_2388 (O_2388,N_23428,N_24916);
nor UO_2389 (O_2389,N_22609,N_24974);
or UO_2390 (O_2390,N_22848,N_24668);
nor UO_2391 (O_2391,N_23596,N_22791);
and UO_2392 (O_2392,N_24111,N_24146);
xor UO_2393 (O_2393,N_23961,N_24251);
xnor UO_2394 (O_2394,N_24118,N_24307);
or UO_2395 (O_2395,N_23853,N_22726);
nor UO_2396 (O_2396,N_24309,N_24412);
or UO_2397 (O_2397,N_24315,N_23109);
nor UO_2398 (O_2398,N_22663,N_22774);
or UO_2399 (O_2399,N_24630,N_23429);
nand UO_2400 (O_2400,N_22950,N_23990);
or UO_2401 (O_2401,N_24228,N_23142);
nor UO_2402 (O_2402,N_23991,N_24382);
nor UO_2403 (O_2403,N_24589,N_24799);
nor UO_2404 (O_2404,N_23849,N_23069);
xnor UO_2405 (O_2405,N_22638,N_23065);
nand UO_2406 (O_2406,N_24958,N_24949);
xor UO_2407 (O_2407,N_24621,N_24107);
nand UO_2408 (O_2408,N_24754,N_24687);
or UO_2409 (O_2409,N_23677,N_24969);
or UO_2410 (O_2410,N_22984,N_24503);
nand UO_2411 (O_2411,N_23260,N_24864);
nor UO_2412 (O_2412,N_24712,N_24020);
nor UO_2413 (O_2413,N_23309,N_24606);
nand UO_2414 (O_2414,N_22951,N_23014);
xnor UO_2415 (O_2415,N_23519,N_24790);
and UO_2416 (O_2416,N_24829,N_24700);
nand UO_2417 (O_2417,N_23598,N_24584);
nor UO_2418 (O_2418,N_24211,N_23873);
xnor UO_2419 (O_2419,N_24276,N_23159);
nand UO_2420 (O_2420,N_23480,N_24408);
or UO_2421 (O_2421,N_23483,N_23764);
xor UO_2422 (O_2422,N_24885,N_24604);
or UO_2423 (O_2423,N_24377,N_23966);
or UO_2424 (O_2424,N_23099,N_23635);
xor UO_2425 (O_2425,N_22958,N_24247);
xor UO_2426 (O_2426,N_22818,N_22752);
and UO_2427 (O_2427,N_24295,N_24583);
nor UO_2428 (O_2428,N_24421,N_24619);
nand UO_2429 (O_2429,N_22653,N_23220);
nor UO_2430 (O_2430,N_23212,N_23038);
nor UO_2431 (O_2431,N_23993,N_23865);
and UO_2432 (O_2432,N_22555,N_24002);
and UO_2433 (O_2433,N_23699,N_23564);
and UO_2434 (O_2434,N_24079,N_23181);
or UO_2435 (O_2435,N_23760,N_24352);
xnor UO_2436 (O_2436,N_24051,N_23094);
and UO_2437 (O_2437,N_23429,N_23526);
and UO_2438 (O_2438,N_23425,N_22836);
xor UO_2439 (O_2439,N_22908,N_24242);
nand UO_2440 (O_2440,N_23720,N_24678);
or UO_2441 (O_2441,N_23456,N_24063);
and UO_2442 (O_2442,N_24109,N_24181);
nand UO_2443 (O_2443,N_22792,N_23765);
nor UO_2444 (O_2444,N_23720,N_24769);
nor UO_2445 (O_2445,N_24280,N_24317);
nor UO_2446 (O_2446,N_24941,N_23191);
nand UO_2447 (O_2447,N_22688,N_24683);
or UO_2448 (O_2448,N_24849,N_24154);
xnor UO_2449 (O_2449,N_23871,N_23792);
nand UO_2450 (O_2450,N_23320,N_24198);
and UO_2451 (O_2451,N_24519,N_23430);
nor UO_2452 (O_2452,N_22526,N_24545);
xnor UO_2453 (O_2453,N_24700,N_23463);
nor UO_2454 (O_2454,N_23793,N_23100);
and UO_2455 (O_2455,N_24387,N_22757);
nor UO_2456 (O_2456,N_24618,N_22509);
nor UO_2457 (O_2457,N_24631,N_22803);
or UO_2458 (O_2458,N_24900,N_24084);
nor UO_2459 (O_2459,N_24330,N_24703);
and UO_2460 (O_2460,N_23102,N_23311);
and UO_2461 (O_2461,N_24865,N_24296);
nor UO_2462 (O_2462,N_23735,N_24008);
nor UO_2463 (O_2463,N_23164,N_24280);
and UO_2464 (O_2464,N_22637,N_24983);
nand UO_2465 (O_2465,N_24693,N_22944);
and UO_2466 (O_2466,N_22765,N_24210);
nor UO_2467 (O_2467,N_24384,N_23420);
nor UO_2468 (O_2468,N_22736,N_22649);
and UO_2469 (O_2469,N_22698,N_22753);
nand UO_2470 (O_2470,N_23773,N_24062);
or UO_2471 (O_2471,N_23760,N_24011);
xor UO_2472 (O_2472,N_22896,N_23011);
nand UO_2473 (O_2473,N_24444,N_23674);
xnor UO_2474 (O_2474,N_24250,N_22774);
xor UO_2475 (O_2475,N_23532,N_24091);
nand UO_2476 (O_2476,N_24998,N_24085);
nand UO_2477 (O_2477,N_23294,N_22850);
and UO_2478 (O_2478,N_22696,N_22574);
or UO_2479 (O_2479,N_24515,N_22519);
or UO_2480 (O_2480,N_23977,N_22675);
nor UO_2481 (O_2481,N_24765,N_23009);
nor UO_2482 (O_2482,N_24654,N_23040);
nand UO_2483 (O_2483,N_24574,N_24154);
or UO_2484 (O_2484,N_24856,N_24347);
xor UO_2485 (O_2485,N_24201,N_23489);
and UO_2486 (O_2486,N_24285,N_24958);
xnor UO_2487 (O_2487,N_22776,N_23049);
nor UO_2488 (O_2488,N_23885,N_23606);
and UO_2489 (O_2489,N_22914,N_24321);
nand UO_2490 (O_2490,N_22953,N_24769);
or UO_2491 (O_2491,N_23954,N_23837);
nor UO_2492 (O_2492,N_23252,N_24083);
nor UO_2493 (O_2493,N_23517,N_23247);
xnor UO_2494 (O_2494,N_24970,N_24184);
or UO_2495 (O_2495,N_22550,N_22724);
and UO_2496 (O_2496,N_22738,N_24172);
nor UO_2497 (O_2497,N_24018,N_23281);
and UO_2498 (O_2498,N_24753,N_22709);
nand UO_2499 (O_2499,N_24416,N_23647);
nand UO_2500 (O_2500,N_24090,N_24450);
and UO_2501 (O_2501,N_24764,N_23422);
or UO_2502 (O_2502,N_24304,N_23004);
nand UO_2503 (O_2503,N_24918,N_23585);
or UO_2504 (O_2504,N_23935,N_24995);
and UO_2505 (O_2505,N_24860,N_22806);
nor UO_2506 (O_2506,N_23556,N_24908);
nand UO_2507 (O_2507,N_23012,N_22994);
or UO_2508 (O_2508,N_23008,N_24070);
and UO_2509 (O_2509,N_24121,N_23683);
nand UO_2510 (O_2510,N_24151,N_24903);
or UO_2511 (O_2511,N_23261,N_23076);
nor UO_2512 (O_2512,N_22871,N_23711);
xor UO_2513 (O_2513,N_23128,N_23024);
xor UO_2514 (O_2514,N_24842,N_24408);
and UO_2515 (O_2515,N_23965,N_22693);
or UO_2516 (O_2516,N_22824,N_23254);
and UO_2517 (O_2517,N_24055,N_23968);
nor UO_2518 (O_2518,N_23206,N_24945);
nor UO_2519 (O_2519,N_23503,N_24085);
nor UO_2520 (O_2520,N_23806,N_22598);
or UO_2521 (O_2521,N_23532,N_24907);
nor UO_2522 (O_2522,N_24242,N_22935);
xnor UO_2523 (O_2523,N_24536,N_22849);
and UO_2524 (O_2524,N_24311,N_23183);
or UO_2525 (O_2525,N_24331,N_24311);
and UO_2526 (O_2526,N_24845,N_24920);
nor UO_2527 (O_2527,N_22913,N_24292);
or UO_2528 (O_2528,N_23130,N_24266);
or UO_2529 (O_2529,N_24990,N_24797);
or UO_2530 (O_2530,N_23775,N_22524);
nor UO_2531 (O_2531,N_22860,N_22621);
and UO_2532 (O_2532,N_23859,N_24303);
xnor UO_2533 (O_2533,N_24386,N_24303);
xnor UO_2534 (O_2534,N_23288,N_23443);
and UO_2535 (O_2535,N_23338,N_22561);
nand UO_2536 (O_2536,N_24093,N_22676);
or UO_2537 (O_2537,N_23634,N_24138);
xor UO_2538 (O_2538,N_23624,N_24009);
or UO_2539 (O_2539,N_24779,N_24608);
nand UO_2540 (O_2540,N_23922,N_24804);
nand UO_2541 (O_2541,N_23495,N_24668);
and UO_2542 (O_2542,N_24769,N_23989);
nor UO_2543 (O_2543,N_24485,N_23384);
xnor UO_2544 (O_2544,N_24994,N_23255);
nor UO_2545 (O_2545,N_23340,N_23466);
or UO_2546 (O_2546,N_24084,N_23610);
and UO_2547 (O_2547,N_24080,N_24799);
xnor UO_2548 (O_2548,N_22693,N_23879);
nand UO_2549 (O_2549,N_23638,N_24329);
nor UO_2550 (O_2550,N_24106,N_23346);
xnor UO_2551 (O_2551,N_24936,N_22529);
xor UO_2552 (O_2552,N_22606,N_24602);
xnor UO_2553 (O_2553,N_23425,N_24750);
nor UO_2554 (O_2554,N_23007,N_24842);
and UO_2555 (O_2555,N_24156,N_24743);
or UO_2556 (O_2556,N_23892,N_24212);
xnor UO_2557 (O_2557,N_23368,N_23707);
nor UO_2558 (O_2558,N_23031,N_24748);
nand UO_2559 (O_2559,N_23327,N_24849);
nor UO_2560 (O_2560,N_24269,N_23023);
and UO_2561 (O_2561,N_23734,N_22910);
nand UO_2562 (O_2562,N_24900,N_24742);
nor UO_2563 (O_2563,N_24230,N_23652);
nand UO_2564 (O_2564,N_23119,N_23125);
nand UO_2565 (O_2565,N_23997,N_24972);
nor UO_2566 (O_2566,N_24113,N_23669);
and UO_2567 (O_2567,N_23673,N_23842);
and UO_2568 (O_2568,N_24897,N_24051);
xnor UO_2569 (O_2569,N_24522,N_23702);
nand UO_2570 (O_2570,N_24104,N_22906);
nor UO_2571 (O_2571,N_24738,N_23278);
xor UO_2572 (O_2572,N_23519,N_24216);
nor UO_2573 (O_2573,N_24986,N_23716);
nand UO_2574 (O_2574,N_23959,N_23883);
and UO_2575 (O_2575,N_23634,N_23959);
and UO_2576 (O_2576,N_23015,N_24887);
nand UO_2577 (O_2577,N_24391,N_23173);
xor UO_2578 (O_2578,N_24693,N_23587);
or UO_2579 (O_2579,N_24491,N_24844);
nand UO_2580 (O_2580,N_24976,N_24240);
nor UO_2581 (O_2581,N_24444,N_23818);
and UO_2582 (O_2582,N_24984,N_23870);
nand UO_2583 (O_2583,N_22603,N_22703);
or UO_2584 (O_2584,N_23274,N_22764);
nand UO_2585 (O_2585,N_24584,N_24371);
nor UO_2586 (O_2586,N_23016,N_24527);
xor UO_2587 (O_2587,N_24569,N_23052);
or UO_2588 (O_2588,N_23306,N_22555);
or UO_2589 (O_2589,N_24764,N_23778);
and UO_2590 (O_2590,N_23477,N_24425);
or UO_2591 (O_2591,N_24607,N_23286);
nor UO_2592 (O_2592,N_24261,N_22603);
nand UO_2593 (O_2593,N_23737,N_22597);
or UO_2594 (O_2594,N_22647,N_23555);
xor UO_2595 (O_2595,N_24514,N_22656);
and UO_2596 (O_2596,N_24883,N_24352);
or UO_2597 (O_2597,N_24905,N_23429);
and UO_2598 (O_2598,N_24891,N_23920);
and UO_2599 (O_2599,N_24523,N_23634);
nand UO_2600 (O_2600,N_22678,N_24595);
and UO_2601 (O_2601,N_24080,N_22708);
or UO_2602 (O_2602,N_23547,N_23696);
and UO_2603 (O_2603,N_23958,N_22671);
or UO_2604 (O_2604,N_22812,N_23140);
or UO_2605 (O_2605,N_24985,N_23473);
nor UO_2606 (O_2606,N_23697,N_24530);
and UO_2607 (O_2607,N_23038,N_24596);
or UO_2608 (O_2608,N_22680,N_24566);
or UO_2609 (O_2609,N_24810,N_24376);
xor UO_2610 (O_2610,N_23048,N_24256);
xnor UO_2611 (O_2611,N_22897,N_22790);
or UO_2612 (O_2612,N_23199,N_22856);
and UO_2613 (O_2613,N_23878,N_23787);
nand UO_2614 (O_2614,N_24244,N_22755);
or UO_2615 (O_2615,N_22920,N_22717);
xnor UO_2616 (O_2616,N_22912,N_24032);
or UO_2617 (O_2617,N_24798,N_24182);
or UO_2618 (O_2618,N_23449,N_24279);
xnor UO_2619 (O_2619,N_23479,N_24416);
nand UO_2620 (O_2620,N_24019,N_23170);
xor UO_2621 (O_2621,N_24661,N_23409);
nand UO_2622 (O_2622,N_23703,N_22775);
nor UO_2623 (O_2623,N_24241,N_23113);
or UO_2624 (O_2624,N_23105,N_24032);
nand UO_2625 (O_2625,N_23279,N_23504);
and UO_2626 (O_2626,N_23815,N_24009);
nand UO_2627 (O_2627,N_23416,N_22506);
or UO_2628 (O_2628,N_22624,N_24959);
nor UO_2629 (O_2629,N_24604,N_24876);
xor UO_2630 (O_2630,N_23532,N_23377);
nor UO_2631 (O_2631,N_22782,N_23790);
or UO_2632 (O_2632,N_24823,N_24958);
or UO_2633 (O_2633,N_23746,N_24017);
xnor UO_2634 (O_2634,N_24085,N_22759);
nand UO_2635 (O_2635,N_22568,N_24460);
nor UO_2636 (O_2636,N_22520,N_22904);
xnor UO_2637 (O_2637,N_22971,N_23967);
nor UO_2638 (O_2638,N_24644,N_23359);
or UO_2639 (O_2639,N_24135,N_24662);
xnor UO_2640 (O_2640,N_23406,N_24099);
xor UO_2641 (O_2641,N_24855,N_24943);
nor UO_2642 (O_2642,N_22967,N_23787);
nand UO_2643 (O_2643,N_23020,N_24335);
xor UO_2644 (O_2644,N_23790,N_22645);
xnor UO_2645 (O_2645,N_23405,N_22517);
nor UO_2646 (O_2646,N_24444,N_23273);
xor UO_2647 (O_2647,N_23375,N_24590);
or UO_2648 (O_2648,N_23541,N_24349);
nand UO_2649 (O_2649,N_22599,N_23131);
or UO_2650 (O_2650,N_22639,N_23454);
and UO_2651 (O_2651,N_24412,N_24066);
or UO_2652 (O_2652,N_24613,N_23084);
and UO_2653 (O_2653,N_24637,N_24702);
nor UO_2654 (O_2654,N_23013,N_23311);
or UO_2655 (O_2655,N_24537,N_22729);
and UO_2656 (O_2656,N_23369,N_24230);
nor UO_2657 (O_2657,N_22991,N_24401);
xnor UO_2658 (O_2658,N_23959,N_23010);
nand UO_2659 (O_2659,N_23168,N_23433);
and UO_2660 (O_2660,N_23624,N_23153);
nor UO_2661 (O_2661,N_24825,N_24865);
or UO_2662 (O_2662,N_22866,N_23508);
nor UO_2663 (O_2663,N_24508,N_24635);
and UO_2664 (O_2664,N_22910,N_24538);
and UO_2665 (O_2665,N_22841,N_24063);
nor UO_2666 (O_2666,N_24880,N_24206);
or UO_2667 (O_2667,N_24898,N_24281);
nand UO_2668 (O_2668,N_24194,N_24652);
nand UO_2669 (O_2669,N_23520,N_22837);
nand UO_2670 (O_2670,N_22654,N_24443);
nand UO_2671 (O_2671,N_23560,N_22807);
or UO_2672 (O_2672,N_23430,N_23642);
xor UO_2673 (O_2673,N_24463,N_22948);
xor UO_2674 (O_2674,N_24331,N_24752);
or UO_2675 (O_2675,N_24380,N_23368);
xor UO_2676 (O_2676,N_24615,N_24981);
or UO_2677 (O_2677,N_23124,N_24779);
nor UO_2678 (O_2678,N_23515,N_23548);
or UO_2679 (O_2679,N_24671,N_22852);
and UO_2680 (O_2680,N_23481,N_24083);
and UO_2681 (O_2681,N_24271,N_24124);
nor UO_2682 (O_2682,N_23082,N_24756);
or UO_2683 (O_2683,N_24327,N_22500);
and UO_2684 (O_2684,N_22648,N_22610);
or UO_2685 (O_2685,N_23729,N_24106);
xnor UO_2686 (O_2686,N_24121,N_23598);
nand UO_2687 (O_2687,N_23891,N_24757);
or UO_2688 (O_2688,N_23226,N_23943);
xor UO_2689 (O_2689,N_22533,N_23021);
or UO_2690 (O_2690,N_22647,N_24664);
xor UO_2691 (O_2691,N_24760,N_24220);
or UO_2692 (O_2692,N_24419,N_23226);
xnor UO_2693 (O_2693,N_24640,N_23298);
and UO_2694 (O_2694,N_24667,N_23355);
nand UO_2695 (O_2695,N_22793,N_23967);
and UO_2696 (O_2696,N_24191,N_23757);
xnor UO_2697 (O_2697,N_22928,N_23235);
or UO_2698 (O_2698,N_22638,N_23030);
nor UO_2699 (O_2699,N_23296,N_23331);
nor UO_2700 (O_2700,N_24053,N_22823);
and UO_2701 (O_2701,N_22611,N_24527);
and UO_2702 (O_2702,N_24634,N_24519);
nor UO_2703 (O_2703,N_23083,N_24633);
and UO_2704 (O_2704,N_24551,N_22844);
nor UO_2705 (O_2705,N_24612,N_23781);
and UO_2706 (O_2706,N_24808,N_23978);
nor UO_2707 (O_2707,N_24119,N_23157);
xor UO_2708 (O_2708,N_22765,N_24039);
xnor UO_2709 (O_2709,N_24790,N_22625);
xnor UO_2710 (O_2710,N_22532,N_23607);
nor UO_2711 (O_2711,N_23298,N_22843);
nand UO_2712 (O_2712,N_24400,N_23684);
and UO_2713 (O_2713,N_24683,N_24027);
nand UO_2714 (O_2714,N_22653,N_22605);
nor UO_2715 (O_2715,N_24106,N_23266);
or UO_2716 (O_2716,N_23916,N_24102);
or UO_2717 (O_2717,N_22541,N_23443);
xor UO_2718 (O_2718,N_23406,N_22731);
and UO_2719 (O_2719,N_24537,N_24637);
xor UO_2720 (O_2720,N_24896,N_22600);
nand UO_2721 (O_2721,N_22691,N_23482);
xnor UO_2722 (O_2722,N_23970,N_24749);
nor UO_2723 (O_2723,N_24694,N_23432);
and UO_2724 (O_2724,N_24990,N_23488);
or UO_2725 (O_2725,N_22589,N_23876);
and UO_2726 (O_2726,N_23954,N_24512);
nor UO_2727 (O_2727,N_23153,N_23682);
xnor UO_2728 (O_2728,N_23127,N_24101);
nor UO_2729 (O_2729,N_24995,N_23413);
nand UO_2730 (O_2730,N_23551,N_23553);
or UO_2731 (O_2731,N_22520,N_24042);
nor UO_2732 (O_2732,N_22768,N_24591);
or UO_2733 (O_2733,N_23309,N_24308);
and UO_2734 (O_2734,N_23954,N_23860);
nand UO_2735 (O_2735,N_22662,N_23549);
nand UO_2736 (O_2736,N_24748,N_23384);
nor UO_2737 (O_2737,N_23274,N_23396);
or UO_2738 (O_2738,N_23982,N_23162);
xnor UO_2739 (O_2739,N_24587,N_23901);
nor UO_2740 (O_2740,N_24247,N_24239);
nand UO_2741 (O_2741,N_24910,N_22642);
nand UO_2742 (O_2742,N_24908,N_23432);
or UO_2743 (O_2743,N_23549,N_23155);
nand UO_2744 (O_2744,N_23572,N_24515);
or UO_2745 (O_2745,N_23493,N_24126);
or UO_2746 (O_2746,N_23544,N_23926);
xnor UO_2747 (O_2747,N_22544,N_23011);
xor UO_2748 (O_2748,N_24511,N_22894);
xnor UO_2749 (O_2749,N_22607,N_22760);
and UO_2750 (O_2750,N_23609,N_23189);
xor UO_2751 (O_2751,N_23024,N_22686);
or UO_2752 (O_2752,N_22798,N_22751);
and UO_2753 (O_2753,N_22974,N_24012);
xnor UO_2754 (O_2754,N_24179,N_24013);
nand UO_2755 (O_2755,N_24502,N_24741);
or UO_2756 (O_2756,N_24759,N_23686);
xor UO_2757 (O_2757,N_23340,N_24995);
xor UO_2758 (O_2758,N_24581,N_24637);
xnor UO_2759 (O_2759,N_24464,N_23652);
nor UO_2760 (O_2760,N_24734,N_22679);
nand UO_2761 (O_2761,N_23874,N_24140);
xnor UO_2762 (O_2762,N_24387,N_22893);
nor UO_2763 (O_2763,N_22648,N_22558);
and UO_2764 (O_2764,N_23390,N_22749);
and UO_2765 (O_2765,N_23808,N_23659);
xor UO_2766 (O_2766,N_23180,N_22839);
nor UO_2767 (O_2767,N_23062,N_24513);
nor UO_2768 (O_2768,N_22767,N_23409);
nor UO_2769 (O_2769,N_24662,N_23845);
or UO_2770 (O_2770,N_22786,N_24149);
nand UO_2771 (O_2771,N_24245,N_24009);
and UO_2772 (O_2772,N_24577,N_24190);
or UO_2773 (O_2773,N_24517,N_24938);
xnor UO_2774 (O_2774,N_23033,N_24868);
or UO_2775 (O_2775,N_22580,N_24776);
or UO_2776 (O_2776,N_24036,N_24459);
nor UO_2777 (O_2777,N_24567,N_22749);
xor UO_2778 (O_2778,N_23164,N_22649);
nand UO_2779 (O_2779,N_23004,N_23441);
nor UO_2780 (O_2780,N_24062,N_22966);
xor UO_2781 (O_2781,N_24969,N_24653);
or UO_2782 (O_2782,N_22637,N_23498);
nor UO_2783 (O_2783,N_24657,N_22907);
nor UO_2784 (O_2784,N_24212,N_23006);
or UO_2785 (O_2785,N_24891,N_24881);
xnor UO_2786 (O_2786,N_22897,N_23605);
nor UO_2787 (O_2787,N_23153,N_22553);
and UO_2788 (O_2788,N_22840,N_23470);
xor UO_2789 (O_2789,N_22735,N_23484);
or UO_2790 (O_2790,N_24115,N_24883);
or UO_2791 (O_2791,N_22739,N_24580);
xnor UO_2792 (O_2792,N_22660,N_24198);
and UO_2793 (O_2793,N_22578,N_22589);
nor UO_2794 (O_2794,N_24922,N_23158);
and UO_2795 (O_2795,N_23614,N_23946);
xnor UO_2796 (O_2796,N_23775,N_23959);
xor UO_2797 (O_2797,N_23660,N_24642);
or UO_2798 (O_2798,N_22637,N_23196);
nand UO_2799 (O_2799,N_22669,N_23254);
nand UO_2800 (O_2800,N_24507,N_23605);
or UO_2801 (O_2801,N_24649,N_23946);
or UO_2802 (O_2802,N_23186,N_23717);
nor UO_2803 (O_2803,N_23299,N_24029);
xor UO_2804 (O_2804,N_24284,N_24527);
nor UO_2805 (O_2805,N_24552,N_23795);
or UO_2806 (O_2806,N_23272,N_23494);
nand UO_2807 (O_2807,N_23057,N_24272);
nor UO_2808 (O_2808,N_23893,N_22619);
nand UO_2809 (O_2809,N_24985,N_22774);
or UO_2810 (O_2810,N_24322,N_23368);
xnor UO_2811 (O_2811,N_24464,N_22901);
and UO_2812 (O_2812,N_23786,N_23876);
xor UO_2813 (O_2813,N_23476,N_23155);
xor UO_2814 (O_2814,N_23593,N_24340);
nand UO_2815 (O_2815,N_24373,N_24125);
and UO_2816 (O_2816,N_23378,N_23607);
nor UO_2817 (O_2817,N_22954,N_23486);
and UO_2818 (O_2818,N_23124,N_24996);
xnor UO_2819 (O_2819,N_22618,N_22727);
or UO_2820 (O_2820,N_22622,N_22763);
nor UO_2821 (O_2821,N_24868,N_23556);
and UO_2822 (O_2822,N_22625,N_22557);
or UO_2823 (O_2823,N_22614,N_23880);
nand UO_2824 (O_2824,N_22906,N_23297);
xnor UO_2825 (O_2825,N_24788,N_24258);
or UO_2826 (O_2826,N_23251,N_23846);
nor UO_2827 (O_2827,N_23415,N_22692);
xor UO_2828 (O_2828,N_24225,N_22535);
nor UO_2829 (O_2829,N_23448,N_23523);
nand UO_2830 (O_2830,N_23703,N_23217);
or UO_2831 (O_2831,N_22555,N_22548);
and UO_2832 (O_2832,N_24177,N_24630);
nand UO_2833 (O_2833,N_23544,N_24229);
or UO_2834 (O_2834,N_23630,N_24737);
nand UO_2835 (O_2835,N_22952,N_22923);
nand UO_2836 (O_2836,N_24934,N_22750);
xor UO_2837 (O_2837,N_23717,N_23693);
or UO_2838 (O_2838,N_24500,N_24787);
and UO_2839 (O_2839,N_23736,N_22871);
xnor UO_2840 (O_2840,N_22733,N_22771);
and UO_2841 (O_2841,N_24369,N_24463);
or UO_2842 (O_2842,N_24637,N_22632);
nand UO_2843 (O_2843,N_23742,N_23752);
and UO_2844 (O_2844,N_23543,N_22673);
nor UO_2845 (O_2845,N_22888,N_23253);
or UO_2846 (O_2846,N_24012,N_22864);
or UO_2847 (O_2847,N_23868,N_23435);
nand UO_2848 (O_2848,N_23432,N_23189);
nand UO_2849 (O_2849,N_23675,N_24957);
nor UO_2850 (O_2850,N_22500,N_23368);
or UO_2851 (O_2851,N_23433,N_24511);
nor UO_2852 (O_2852,N_24487,N_24165);
or UO_2853 (O_2853,N_23551,N_22685);
nor UO_2854 (O_2854,N_23941,N_24647);
and UO_2855 (O_2855,N_23784,N_23916);
nand UO_2856 (O_2856,N_24061,N_23079);
nor UO_2857 (O_2857,N_24643,N_24030);
nand UO_2858 (O_2858,N_24214,N_24313);
nor UO_2859 (O_2859,N_22861,N_24583);
nor UO_2860 (O_2860,N_22922,N_22726);
or UO_2861 (O_2861,N_23832,N_23874);
xor UO_2862 (O_2862,N_22677,N_24092);
nor UO_2863 (O_2863,N_24994,N_24310);
or UO_2864 (O_2864,N_23559,N_24866);
xnor UO_2865 (O_2865,N_24757,N_24302);
and UO_2866 (O_2866,N_23634,N_22862);
or UO_2867 (O_2867,N_22885,N_24793);
nand UO_2868 (O_2868,N_24096,N_24085);
nand UO_2869 (O_2869,N_22565,N_23778);
or UO_2870 (O_2870,N_24495,N_23266);
xnor UO_2871 (O_2871,N_23060,N_22580);
nand UO_2872 (O_2872,N_23108,N_24325);
nor UO_2873 (O_2873,N_22788,N_24484);
and UO_2874 (O_2874,N_23872,N_23193);
nand UO_2875 (O_2875,N_24816,N_23750);
and UO_2876 (O_2876,N_24835,N_23673);
xnor UO_2877 (O_2877,N_23909,N_23262);
xor UO_2878 (O_2878,N_24902,N_22813);
nor UO_2879 (O_2879,N_23003,N_24996);
nand UO_2880 (O_2880,N_22680,N_24662);
xor UO_2881 (O_2881,N_22679,N_24142);
or UO_2882 (O_2882,N_24040,N_22896);
nor UO_2883 (O_2883,N_24491,N_22646);
xor UO_2884 (O_2884,N_24668,N_23367);
nand UO_2885 (O_2885,N_24102,N_24983);
and UO_2886 (O_2886,N_24455,N_24626);
nor UO_2887 (O_2887,N_22768,N_24996);
nor UO_2888 (O_2888,N_24033,N_23561);
xor UO_2889 (O_2889,N_23845,N_24163);
or UO_2890 (O_2890,N_24662,N_24799);
nand UO_2891 (O_2891,N_22737,N_24650);
nor UO_2892 (O_2892,N_23475,N_24028);
or UO_2893 (O_2893,N_23232,N_22586);
nor UO_2894 (O_2894,N_23669,N_22928);
or UO_2895 (O_2895,N_22703,N_22535);
xnor UO_2896 (O_2896,N_24930,N_24348);
or UO_2897 (O_2897,N_23897,N_24202);
xnor UO_2898 (O_2898,N_23804,N_23584);
or UO_2899 (O_2899,N_22992,N_24027);
or UO_2900 (O_2900,N_23357,N_23383);
xnor UO_2901 (O_2901,N_22812,N_23657);
or UO_2902 (O_2902,N_23098,N_23554);
or UO_2903 (O_2903,N_23063,N_22575);
xor UO_2904 (O_2904,N_24430,N_22679);
and UO_2905 (O_2905,N_24893,N_23614);
nand UO_2906 (O_2906,N_22806,N_24079);
nor UO_2907 (O_2907,N_22794,N_22525);
or UO_2908 (O_2908,N_23805,N_24780);
and UO_2909 (O_2909,N_24349,N_23384);
and UO_2910 (O_2910,N_22604,N_22509);
nor UO_2911 (O_2911,N_24424,N_23467);
and UO_2912 (O_2912,N_23581,N_24619);
or UO_2913 (O_2913,N_24034,N_24618);
or UO_2914 (O_2914,N_22993,N_23762);
nand UO_2915 (O_2915,N_22715,N_24366);
and UO_2916 (O_2916,N_22764,N_24340);
or UO_2917 (O_2917,N_23068,N_24436);
xor UO_2918 (O_2918,N_23149,N_23533);
nor UO_2919 (O_2919,N_22653,N_24223);
xor UO_2920 (O_2920,N_23647,N_23280);
xnor UO_2921 (O_2921,N_22518,N_24264);
and UO_2922 (O_2922,N_23024,N_22666);
nand UO_2923 (O_2923,N_23218,N_24305);
nand UO_2924 (O_2924,N_23151,N_24808);
or UO_2925 (O_2925,N_23175,N_23054);
and UO_2926 (O_2926,N_24972,N_24432);
or UO_2927 (O_2927,N_22964,N_24165);
nand UO_2928 (O_2928,N_23697,N_23914);
or UO_2929 (O_2929,N_23711,N_24164);
nor UO_2930 (O_2930,N_22936,N_23255);
nand UO_2931 (O_2931,N_23835,N_23007);
or UO_2932 (O_2932,N_24590,N_24720);
nor UO_2933 (O_2933,N_23746,N_22888);
or UO_2934 (O_2934,N_23848,N_24595);
nor UO_2935 (O_2935,N_23384,N_24941);
xnor UO_2936 (O_2936,N_23817,N_23018);
and UO_2937 (O_2937,N_24943,N_23152);
or UO_2938 (O_2938,N_24843,N_22966);
nand UO_2939 (O_2939,N_23082,N_22903);
nor UO_2940 (O_2940,N_23227,N_23879);
or UO_2941 (O_2941,N_24818,N_23634);
or UO_2942 (O_2942,N_24623,N_23885);
xor UO_2943 (O_2943,N_22562,N_23242);
nand UO_2944 (O_2944,N_24751,N_24826);
xnor UO_2945 (O_2945,N_23189,N_24108);
nand UO_2946 (O_2946,N_22699,N_24024);
xnor UO_2947 (O_2947,N_24573,N_24776);
nand UO_2948 (O_2948,N_23844,N_24354);
and UO_2949 (O_2949,N_23571,N_23445);
nand UO_2950 (O_2950,N_23404,N_23321);
nor UO_2951 (O_2951,N_24894,N_24379);
nor UO_2952 (O_2952,N_23391,N_24055);
and UO_2953 (O_2953,N_23815,N_23813);
nor UO_2954 (O_2954,N_24032,N_24674);
nand UO_2955 (O_2955,N_22970,N_24989);
nor UO_2956 (O_2956,N_23551,N_24523);
nor UO_2957 (O_2957,N_24122,N_22721);
and UO_2958 (O_2958,N_23247,N_24333);
or UO_2959 (O_2959,N_24868,N_24601);
xor UO_2960 (O_2960,N_22607,N_24958);
and UO_2961 (O_2961,N_24694,N_22983);
or UO_2962 (O_2962,N_22902,N_22835);
or UO_2963 (O_2963,N_24186,N_24165);
nor UO_2964 (O_2964,N_24883,N_22684);
and UO_2965 (O_2965,N_22714,N_22544);
nand UO_2966 (O_2966,N_24049,N_22862);
or UO_2967 (O_2967,N_22873,N_23812);
and UO_2968 (O_2968,N_24890,N_22923);
nand UO_2969 (O_2969,N_23983,N_22978);
or UO_2970 (O_2970,N_23976,N_24624);
or UO_2971 (O_2971,N_22838,N_24083);
nand UO_2972 (O_2972,N_23043,N_24640);
and UO_2973 (O_2973,N_23334,N_23281);
nor UO_2974 (O_2974,N_23136,N_22604);
xor UO_2975 (O_2975,N_24457,N_23592);
xor UO_2976 (O_2976,N_22989,N_23681);
nor UO_2977 (O_2977,N_23620,N_24252);
and UO_2978 (O_2978,N_23884,N_22540);
and UO_2979 (O_2979,N_23303,N_23993);
and UO_2980 (O_2980,N_22969,N_24747);
xnor UO_2981 (O_2981,N_24646,N_23428);
nor UO_2982 (O_2982,N_24360,N_22833);
nand UO_2983 (O_2983,N_24416,N_24361);
nor UO_2984 (O_2984,N_23837,N_24511);
nand UO_2985 (O_2985,N_23924,N_24777);
nand UO_2986 (O_2986,N_24647,N_23519);
or UO_2987 (O_2987,N_23833,N_24818);
and UO_2988 (O_2988,N_23132,N_24417);
and UO_2989 (O_2989,N_24052,N_24303);
and UO_2990 (O_2990,N_24956,N_22700);
or UO_2991 (O_2991,N_23737,N_24354);
nand UO_2992 (O_2992,N_23046,N_23998);
or UO_2993 (O_2993,N_22596,N_23177);
xor UO_2994 (O_2994,N_23041,N_23415);
nand UO_2995 (O_2995,N_22560,N_24437);
or UO_2996 (O_2996,N_23586,N_24468);
or UO_2997 (O_2997,N_24680,N_23244);
nand UO_2998 (O_2998,N_22772,N_22725);
xnor UO_2999 (O_2999,N_23736,N_24287);
endmodule