module basic_1500_15000_2000_100_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_627,In_1478);
and U1 (N_1,In_1037,In_413);
xor U2 (N_2,In_223,In_472);
or U3 (N_3,In_130,In_96);
nand U4 (N_4,In_250,In_1175);
nor U5 (N_5,In_441,In_1185);
or U6 (N_6,In_801,In_649);
nand U7 (N_7,In_145,In_277);
xor U8 (N_8,In_976,In_437);
nor U9 (N_9,In_1274,In_464);
and U10 (N_10,In_1191,In_754);
nand U11 (N_11,In_99,In_789);
or U12 (N_12,In_896,In_1266);
xor U13 (N_13,In_1058,In_870);
nand U14 (N_14,In_770,In_575);
xor U15 (N_15,In_655,In_879);
nor U16 (N_16,In_348,In_772);
and U17 (N_17,In_798,In_443);
nor U18 (N_18,In_763,In_1038);
nor U19 (N_19,In_1407,In_1155);
xnor U20 (N_20,In_1219,In_1171);
and U21 (N_21,In_1265,In_1145);
nor U22 (N_22,In_1320,In_5);
nand U23 (N_23,In_502,In_1119);
nand U24 (N_24,In_50,In_714);
xor U25 (N_25,In_745,In_1138);
or U26 (N_26,In_1014,In_1246);
and U27 (N_27,In_567,In_1143);
and U28 (N_28,In_1243,In_213);
xor U29 (N_29,In_670,In_1497);
nand U30 (N_30,In_146,In_538);
xnor U31 (N_31,In_768,In_604);
nand U32 (N_32,In_946,In_967);
or U33 (N_33,In_1203,In_292);
xor U34 (N_34,In_1477,In_760);
xnor U35 (N_35,In_1031,In_124);
nor U36 (N_36,In_382,In_1140);
nand U37 (N_37,In_607,In_855);
and U38 (N_38,In_358,In_926);
nand U39 (N_39,In_1162,In_1224);
xnor U40 (N_40,In_203,In_812);
nor U41 (N_41,In_242,In_1349);
nor U42 (N_42,In_364,In_1028);
or U43 (N_43,In_1110,In_1082);
nor U44 (N_44,In_1022,In_305);
and U45 (N_45,In_174,In_692);
nor U46 (N_46,In_1357,In_532);
nand U47 (N_47,In_934,In_577);
and U48 (N_48,In_1342,In_304);
and U49 (N_49,In_620,In_546);
nor U50 (N_50,In_14,In_1396);
nor U51 (N_51,In_524,In_238);
or U52 (N_52,In_1465,In_561);
nand U53 (N_53,In_426,In_679);
xor U54 (N_54,In_1331,In_404);
nand U55 (N_55,In_433,In_738);
xnor U56 (N_56,In_52,In_401);
or U57 (N_57,In_222,In_1011);
nor U58 (N_58,In_1451,In_514);
and U59 (N_59,In_576,In_438);
and U60 (N_60,In_637,In_1315);
xnor U61 (N_61,In_536,In_200);
or U62 (N_62,In_547,In_1294);
or U63 (N_63,In_42,In_945);
xnor U64 (N_64,In_1118,In_179);
nand U65 (N_65,In_1321,In_1216);
nand U66 (N_66,In_137,In_1098);
or U67 (N_67,In_809,In_58);
nor U68 (N_68,In_446,In_995);
xnor U69 (N_69,In_1130,In_837);
nor U70 (N_70,In_376,In_975);
xor U71 (N_71,In_746,In_984);
nor U72 (N_72,In_700,In_865);
nor U73 (N_73,In_1067,In_689);
nand U74 (N_74,In_1328,In_10);
and U75 (N_75,In_299,In_962);
nor U76 (N_76,In_970,In_1431);
nand U77 (N_77,In_190,In_1239);
and U78 (N_78,In_1471,In_839);
nand U79 (N_79,In_1009,In_506);
xor U80 (N_80,In_317,In_1256);
or U81 (N_81,In_990,In_497);
and U82 (N_82,In_580,In_1042);
xor U83 (N_83,In_1277,In_733);
xnor U84 (N_84,In_362,In_1382);
nor U85 (N_85,In_1247,In_306);
nand U86 (N_86,In_1302,In_69);
nor U87 (N_87,In_259,In_925);
nor U88 (N_88,In_1488,In_862);
nand U89 (N_89,In_492,In_796);
nand U90 (N_90,In_272,In_462);
nand U91 (N_91,In_1435,In_94);
nor U92 (N_92,In_1201,In_1189);
nor U93 (N_93,In_297,In_1026);
xnor U94 (N_94,In_429,In_373);
xnor U95 (N_95,In_683,In_942);
xor U96 (N_96,In_1156,In_947);
xor U97 (N_97,In_1368,In_626);
nor U98 (N_98,In_1270,In_716);
nand U99 (N_99,In_394,In_24);
xnor U100 (N_100,In_147,In_1012);
nand U101 (N_101,In_1196,In_1350);
xnor U102 (N_102,In_728,In_933);
and U103 (N_103,In_350,In_1437);
nor U104 (N_104,In_49,In_958);
and U105 (N_105,In_873,In_465);
and U106 (N_106,In_1370,In_522);
nand U107 (N_107,In_311,In_13);
or U108 (N_108,In_530,In_1071);
xor U109 (N_109,In_140,In_936);
nand U110 (N_110,In_1013,In_1269);
and U111 (N_111,In_647,In_374);
xor U112 (N_112,In_539,In_1141);
xnor U113 (N_113,In_248,In_509);
and U114 (N_114,In_432,In_62);
nand U115 (N_115,In_483,In_390);
nand U116 (N_116,In_428,In_739);
or U117 (N_117,In_1324,In_95);
or U118 (N_118,In_1411,In_1292);
nor U119 (N_119,In_1223,In_159);
and U120 (N_120,In_398,In_1379);
or U121 (N_121,In_357,In_788);
nor U122 (N_122,In_955,In_1049);
nor U123 (N_123,In_1153,In_675);
and U124 (N_124,In_210,In_1148);
xor U125 (N_125,In_65,In_690);
or U126 (N_126,In_252,In_534);
nor U127 (N_127,In_445,In_882);
nor U128 (N_128,In_653,In_1054);
and U129 (N_129,In_225,In_339);
and U130 (N_130,In_1306,In_249);
and U131 (N_131,In_1418,In_761);
xor U132 (N_132,In_1151,In_1221);
and U133 (N_133,In_327,In_1027);
nor U134 (N_134,In_821,In_110);
nand U135 (N_135,In_168,In_199);
nand U136 (N_136,In_512,In_152);
nand U137 (N_137,In_485,In_1000);
xor U138 (N_138,In_558,In_1227);
and U139 (N_139,In_722,In_459);
and U140 (N_140,In_351,In_1424);
or U141 (N_141,In_279,In_618);
or U142 (N_142,In_1260,In_667);
or U143 (N_143,In_1047,In_1298);
and U144 (N_144,In_609,In_544);
xnor U145 (N_145,In_1263,In_1436);
or U146 (N_146,In_1187,In_1008);
nand U147 (N_147,In_1441,In_887);
nand U148 (N_148,In_616,In_499);
xor U149 (N_149,In_1493,In_321);
or U150 (N_150,In_380,In_25);
and U151 (N_151,In_2,In_818);
xnor U152 (N_152,In_102,In_1128);
xor U153 (N_153,In_681,In_540);
nand U154 (N_154,In_1399,In_469);
nor U155 (N_155,In_864,N_35);
and U156 (N_156,In_125,In_1245);
xnor U157 (N_157,In_517,In_1050);
xnor U158 (N_158,In_765,N_110);
and U159 (N_159,In_1457,In_1254);
xnor U160 (N_160,In_347,In_400);
nand U161 (N_161,In_1236,In_831);
nand U162 (N_162,In_1135,In_1157);
xnor U163 (N_163,In_399,In_844);
and U164 (N_164,In_1182,In_164);
nor U165 (N_165,In_769,In_212);
nand U166 (N_166,In_287,In_412);
or U167 (N_167,In_682,In_1417);
and U168 (N_168,In_78,In_84);
nor U169 (N_169,In_254,In_633);
nor U170 (N_170,In_1100,In_599);
or U171 (N_171,In_278,In_944);
xnor U172 (N_172,In_1466,In_204);
xor U173 (N_173,In_919,In_44);
or U174 (N_174,In_309,In_845);
nand U175 (N_175,In_859,In_1132);
xor U176 (N_176,In_82,In_268);
nor U177 (N_177,In_730,In_912);
and U178 (N_178,In_1099,In_478);
and U179 (N_179,In_80,In_435);
or U180 (N_180,In_1429,N_40);
or U181 (N_181,In_1366,In_732);
or U182 (N_182,In_1462,In_424);
xor U183 (N_183,In_537,N_61);
nor U184 (N_184,In_704,In_1329);
or U185 (N_185,In_1,In_552);
or U186 (N_186,In_1248,In_587);
nor U187 (N_187,In_1194,In_126);
or U188 (N_188,In_201,In_1210);
and U189 (N_189,In_11,In_487);
xnor U190 (N_190,In_123,In_1020);
and U191 (N_191,In_451,In_1018);
nor U192 (N_192,In_233,In_907);
and U193 (N_193,In_508,In_1147);
nand U194 (N_194,In_308,In_416);
and U195 (N_195,In_1229,In_629);
and U196 (N_196,In_332,In_785);
or U197 (N_197,In_51,In_1311);
xor U198 (N_198,N_99,In_331);
and U199 (N_199,In_1035,In_260);
nor U200 (N_200,In_151,In_1161);
or U201 (N_201,In_677,N_5);
nand U202 (N_202,In_221,In_1276);
or U203 (N_203,In_1183,In_1262);
and U204 (N_204,In_330,In_353);
xor U205 (N_205,In_301,In_721);
nor U206 (N_206,N_46,In_1259);
nand U207 (N_207,In_1186,N_12);
and U208 (N_208,In_171,In_453);
xor U209 (N_209,In_661,In_12);
and U210 (N_210,In_414,In_1450);
nor U211 (N_211,In_849,In_405);
nor U212 (N_212,In_1356,In_216);
nand U213 (N_213,In_914,In_109);
nand U214 (N_214,In_39,In_1234);
or U215 (N_215,N_50,In_479);
and U216 (N_216,N_8,In_560);
nor U217 (N_217,In_729,In_290);
or U218 (N_218,In_239,In_615);
nand U219 (N_219,In_1006,In_3);
xnor U220 (N_220,In_814,In_286);
xor U221 (N_221,In_697,In_568);
xnor U222 (N_222,In_163,In_215);
and U223 (N_223,In_1036,In_1412);
nor U224 (N_224,In_442,In_1237);
xnor U225 (N_225,In_193,In_158);
or U226 (N_226,In_100,In_601);
nor U227 (N_227,In_325,In_1101);
nand U228 (N_228,In_1285,In_1453);
and U229 (N_229,N_105,In_1233);
xnor U230 (N_230,In_1215,In_1257);
xnor U231 (N_231,In_195,In_759);
xor U232 (N_232,In_585,In_527);
or U233 (N_233,In_68,In_1440);
and U234 (N_234,In_1409,In_1218);
and U235 (N_235,In_869,In_143);
nor U236 (N_236,In_863,In_1154);
or U237 (N_237,In_194,In_594);
and U238 (N_238,In_103,In_592);
xnor U239 (N_239,In_652,In_1363);
and U240 (N_240,In_846,In_1498);
xor U241 (N_241,In_897,In_1388);
and U242 (N_242,In_756,In_209);
xor U243 (N_243,In_1106,In_64);
nor U244 (N_244,In_191,In_1422);
nand U245 (N_245,In_1184,In_1133);
xor U246 (N_246,In_1373,In_1202);
nor U247 (N_247,In_1177,In_1113);
nand U248 (N_248,In_346,In_617);
and U249 (N_249,In_750,In_375);
xnor U250 (N_250,In_885,In_511);
nor U251 (N_251,In_1069,N_109);
xor U252 (N_252,In_335,In_1492);
and U253 (N_253,In_372,N_57);
nand U254 (N_254,In_356,N_93);
xnor U255 (N_255,In_18,In_1024);
or U256 (N_256,In_598,In_1286);
nand U257 (N_257,In_890,In_224);
xnor U258 (N_258,In_1353,N_6);
or U259 (N_259,In_1343,In_55);
nand U260 (N_260,In_491,In_937);
and U261 (N_261,In_656,In_296);
xnor U262 (N_262,In_645,In_853);
nor U263 (N_263,In_1438,In_395);
and U264 (N_264,In_240,In_642);
nor U265 (N_265,In_996,N_38);
xor U266 (N_266,In_156,N_116);
and U267 (N_267,In_977,In_461);
nor U268 (N_268,N_102,In_1092);
nand U269 (N_269,In_1044,In_822);
nor U270 (N_270,In_834,In_71);
xor U271 (N_271,In_963,In_564);
nor U272 (N_272,N_83,In_1332);
and U273 (N_273,In_313,In_940);
or U274 (N_274,In_1371,In_444);
nor U275 (N_275,N_28,In_53);
nand U276 (N_276,In_1459,In_993);
xor U277 (N_277,In_127,N_19);
and U278 (N_278,In_906,In_255);
and U279 (N_279,In_85,In_207);
and U280 (N_280,In_605,In_563);
and U281 (N_281,In_198,In_1387);
or U282 (N_282,N_143,In_1169);
xor U283 (N_283,In_1125,In_323);
nor U284 (N_284,In_1220,In_368);
and U285 (N_285,In_408,In_884);
nor U286 (N_286,In_603,In_1079);
nand U287 (N_287,In_498,In_1433);
nand U288 (N_288,In_1444,N_113);
xnor U289 (N_289,In_500,In_340);
nor U290 (N_290,In_136,In_1160);
xor U291 (N_291,In_234,In_32);
nor U292 (N_292,In_40,In_134);
xnor U293 (N_293,N_25,In_1204);
nand U294 (N_294,In_1144,In_753);
xor U295 (N_295,In_959,N_104);
xnor U296 (N_296,In_186,In_261);
nor U297 (N_297,In_867,In_930);
or U298 (N_298,In_630,In_988);
xor U299 (N_299,In_928,In_1439);
nor U300 (N_300,In_1307,In_917);
or U301 (N_301,In_470,In_1163);
xor U302 (N_302,In_1374,In_289);
nand U303 (N_303,N_53,In_932);
xor U304 (N_304,In_157,N_154);
nor U305 (N_305,N_33,In_1089);
or U306 (N_306,In_1383,In_1405);
or U307 (N_307,In_861,N_79);
or U308 (N_308,In_1358,In_1129);
xor U309 (N_309,In_265,N_26);
nand U310 (N_310,In_87,In_1005);
nor U311 (N_311,In_160,In_76);
nor U312 (N_312,In_1333,In_232);
nor U313 (N_313,In_611,In_1390);
xor U314 (N_314,In_725,In_229);
or U315 (N_315,In_16,N_220);
and U316 (N_316,In_982,In_1272);
nand U317 (N_317,In_1217,In_1490);
xor U318 (N_318,In_957,N_76);
or U319 (N_319,N_64,In_904);
and U320 (N_320,In_883,In_167);
or U321 (N_321,N_158,In_1048);
or U322 (N_322,In_1468,In_1190);
xor U323 (N_323,N_234,In_920);
and U324 (N_324,In_385,In_447);
and U325 (N_325,In_584,In_314);
or U326 (N_326,In_91,N_289);
nor U327 (N_327,In_1059,In_606);
nor U328 (N_328,In_613,In_1423);
nand U329 (N_329,In_566,In_826);
xnor U330 (N_330,In_1040,In_218);
xor U331 (N_331,In_46,In_892);
xnor U332 (N_332,In_1164,In_354);
nand U333 (N_333,In_1283,N_0);
or U334 (N_334,In_574,In_836);
and U335 (N_335,In_623,In_392);
and U336 (N_336,In_467,In_381);
nor U337 (N_337,In_949,In_1318);
nor U338 (N_338,In_344,In_83);
and U339 (N_339,N_272,In_1323);
nor U340 (N_340,In_257,In_1380);
or U341 (N_341,In_359,In_1317);
nand U342 (N_342,In_31,In_1126);
or U343 (N_343,N_27,In_1404);
xnor U344 (N_344,In_666,N_72);
nand U345 (N_345,In_1420,In_956);
and U346 (N_346,In_468,In_1086);
nand U347 (N_347,N_167,In_695);
xnor U348 (N_348,In_111,N_292);
or U349 (N_349,In_815,In_253);
or U350 (N_350,In_280,In_685);
and U351 (N_351,In_1304,In_523);
and U352 (N_352,N_125,In_803);
xor U353 (N_353,In_1485,N_248);
nor U354 (N_354,In_196,In_1445);
xor U355 (N_355,In_1075,In_625);
or U356 (N_356,In_315,In_115);
and U357 (N_357,In_295,N_282);
or U358 (N_358,In_1394,In_411);
nand U359 (N_359,In_266,N_199);
or U360 (N_360,In_1428,In_1046);
nor U361 (N_361,N_49,In_952);
or U362 (N_362,N_148,In_1240);
or U363 (N_363,In_1021,In_1327);
nor U364 (N_364,In_237,In_555);
nor U365 (N_365,In_579,In_1090);
nor U366 (N_366,In_1192,N_163);
or U367 (N_367,In_651,In_545);
and U368 (N_368,In_1063,N_181);
and U369 (N_369,In_67,In_370);
nand U370 (N_370,In_342,In_1346);
and U371 (N_371,In_457,In_397);
nor U372 (N_372,In_894,N_74);
xnor U373 (N_373,In_1461,N_258);
nand U374 (N_374,N_3,N_160);
or U375 (N_375,In_663,In_1108);
nor U376 (N_376,In_774,In_966);
nor U377 (N_377,In_1473,In_101);
and U378 (N_378,N_131,In_646);
and U379 (N_379,In_777,In_1377);
or U380 (N_380,In_1214,In_1258);
nand U381 (N_381,In_969,In_740);
or U382 (N_382,In_107,N_187);
xor U383 (N_383,In_1088,N_58);
nor U384 (N_384,N_255,N_197);
and U385 (N_385,In_366,In_337);
nor U386 (N_386,N_173,In_1337);
or U387 (N_387,In_987,In_379);
xor U388 (N_388,N_278,In_1188);
nor U389 (N_389,N_284,In_981);
nor U390 (N_390,In_256,In_182);
or U391 (N_391,In_294,In_1389);
xor U392 (N_392,In_570,In_709);
xor U393 (N_393,N_151,In_66);
or U394 (N_394,In_431,In_737);
or U395 (N_395,In_1280,N_20);
nor U396 (N_396,In_703,In_891);
nand U397 (N_397,N_186,In_1312);
nand U398 (N_398,In_1206,N_21);
nor U399 (N_399,In_1268,In_450);
xnor U400 (N_400,In_1310,In_718);
nand U401 (N_401,In_1146,N_200);
and U402 (N_402,In_1273,In_1087);
or U403 (N_403,In_923,In_303);
or U404 (N_404,In_406,N_269);
or U405 (N_405,In_1193,In_1016);
xnor U406 (N_406,In_322,In_471);
or U407 (N_407,In_734,In_1454);
nand U408 (N_408,In_515,N_106);
xor U409 (N_409,N_70,In_1308);
nor U410 (N_410,In_535,In_841);
nor U411 (N_411,In_320,In_968);
or U412 (N_412,In_596,N_101);
and U413 (N_413,N_133,N_190);
nor U414 (N_414,N_22,N_217);
and U415 (N_415,In_565,In_489);
xnor U416 (N_416,In_1297,In_501);
or U417 (N_417,In_36,In_771);
nand U418 (N_418,N_214,In_1425);
and U419 (N_419,In_1180,N_254);
or U420 (N_420,In_744,N_202);
or U421 (N_421,In_185,N_162);
xnor U422 (N_422,In_1003,In_54);
and U423 (N_423,N_123,In_717);
nor U424 (N_424,In_755,In_1107);
nor U425 (N_425,In_835,N_257);
and U426 (N_426,In_1326,N_166);
xnor U427 (N_427,N_140,In_241);
nand U428 (N_428,N_276,N_211);
nor U429 (N_429,In_757,In_1406);
or U430 (N_430,In_989,In_449);
xor U431 (N_431,In_929,N_298);
nor U432 (N_432,In_211,In_578);
xor U433 (N_433,N_229,N_67);
xor U434 (N_434,N_219,In_686);
or U435 (N_435,In_983,In_691);
xor U436 (N_436,N_10,In_1004);
and U437 (N_437,In_422,In_271);
and U438 (N_438,In_1096,N_31);
xor U439 (N_439,In_155,In_1137);
nand U440 (N_440,N_77,In_954);
xor U441 (N_441,In_59,N_207);
or U442 (N_442,N_85,In_490);
or U443 (N_443,In_758,In_1172);
nor U444 (N_444,In_162,In_1261);
nand U445 (N_445,In_410,N_126);
nand U446 (N_446,In_458,N_124);
or U447 (N_447,In_843,In_766);
or U448 (N_448,N_231,In_17);
nand U449 (N_449,In_939,N_156);
nor U450 (N_450,N_139,In_148);
xnor U451 (N_451,In_773,In_1480);
xor U452 (N_452,N_54,In_262);
xor U453 (N_453,In_284,In_840);
and U454 (N_454,N_382,In_1056);
xor U455 (N_455,N_182,In_1120);
nor U456 (N_456,In_1034,In_908);
xnor U457 (N_457,In_1470,In_1205);
or U458 (N_458,N_407,In_1112);
nor U459 (N_459,In_345,N_185);
and U460 (N_460,In_219,In_1010);
nand U461 (N_461,N_392,N_121);
nor U462 (N_462,In_231,In_736);
or U463 (N_463,In_267,N_100);
and U464 (N_464,In_581,In_1482);
xor U465 (N_465,In_4,In_726);
and U466 (N_466,N_130,In_371);
xor U467 (N_467,In_850,In_886);
or U468 (N_468,N_178,N_297);
nor U469 (N_469,In_747,N_411);
or U470 (N_470,N_119,N_300);
nand U471 (N_471,In_664,N_424);
and U472 (N_472,N_302,In_1076);
or U473 (N_473,In_889,N_445);
xnor U474 (N_474,In_1097,In_189);
nor U475 (N_475,In_326,In_273);
or U476 (N_476,N_283,N_349);
or U477 (N_477,N_414,In_635);
or U478 (N_478,In_1002,In_192);
xnor U479 (N_479,In_142,In_562);
xnor U480 (N_480,In_1474,N_409);
and U481 (N_481,N_313,N_84);
xnor U482 (N_482,In_455,In_312);
and U483 (N_483,In_1052,N_175);
and U484 (N_484,In_992,N_111);
or U485 (N_485,In_1365,N_440);
and U486 (N_486,In_531,In_694);
or U487 (N_487,In_79,In_1222);
nand U488 (N_488,In_693,In_1072);
and U489 (N_489,In_1401,N_344);
nand U490 (N_490,In_1299,N_137);
nand U491 (N_491,In_1226,In_98);
xor U492 (N_492,In_1230,In_909);
xor U493 (N_493,In_648,N_357);
xor U494 (N_494,N_335,In_1065);
nand U495 (N_495,In_1181,N_203);
nand U496 (N_496,In_622,In_1322);
or U497 (N_497,In_288,N_425);
nand U498 (N_498,In_1166,In_550);
and U499 (N_499,N_29,N_381);
or U500 (N_500,N_419,In_1400);
nor U501 (N_501,In_776,N_37);
or U502 (N_502,N_235,In_866);
and U503 (N_503,N_205,N_368);
xor U504 (N_504,In_1469,In_60);
nor U505 (N_505,N_144,N_358);
or U506 (N_506,In_1345,In_659);
nand U507 (N_507,In_494,N_7);
nor U508 (N_508,In_1378,In_533);
xnor U509 (N_509,In_1413,In_794);
nand U510 (N_510,N_324,In_131);
xnor U511 (N_511,In_1167,In_246);
and U512 (N_512,N_14,In_1476);
nand U513 (N_513,N_299,N_45);
and U514 (N_514,N_92,In_593);
xor U515 (N_515,N_448,In_1385);
nor U516 (N_516,N_371,In_724);
nor U517 (N_517,N_15,N_96);
nor U518 (N_518,In_1200,In_1085);
nor U519 (N_519,In_1364,N_59);
nor U520 (N_520,N_449,N_183);
and U521 (N_521,In_1442,In_169);
nand U522 (N_522,In_513,In_153);
or U523 (N_523,In_980,In_943);
nor U524 (N_524,In_847,N_41);
and U525 (N_525,In_779,In_800);
and U526 (N_526,In_951,In_1017);
or U527 (N_527,In_1293,N_295);
and U528 (N_528,N_417,In_516);
or U529 (N_529,In_504,N_318);
or U530 (N_530,N_321,In_264);
nor U531 (N_531,In_106,In_1352);
nand U532 (N_532,In_720,In_178);
or U533 (N_533,N_347,In_918);
and U534 (N_534,In_1355,N_290);
nand U535 (N_535,In_972,In_1287);
and U536 (N_536,In_402,N_285);
and U537 (N_537,In_463,In_460);
nor U538 (N_538,N_326,In_1339);
and U539 (N_539,N_17,N_446);
and U540 (N_540,In_161,N_340);
xor U541 (N_541,In_244,In_654);
and U542 (N_542,In_1041,In_1178);
nand U543 (N_543,In_466,In_133);
and U544 (N_544,N_169,In_89);
nand U545 (N_545,In_641,In_452);
and U546 (N_546,In_1074,In_1131);
or U547 (N_547,N_224,N_405);
nand U548 (N_548,N_350,In_1449);
nor U549 (N_549,In_1430,N_44);
or U550 (N_550,In_1296,N_252);
nor U551 (N_551,N_98,N_441);
and U552 (N_552,In_588,In_556);
xnor U553 (N_553,In_678,In_660);
nor U554 (N_554,In_1252,In_1284);
nor U555 (N_555,In_1251,In_114);
nand U556 (N_556,In_1419,In_8);
nand U557 (N_557,N_9,N_384);
xnor U558 (N_558,In_324,In_1491);
or U559 (N_559,In_665,In_120);
and U560 (N_560,N_395,In_1124);
nor U561 (N_561,N_442,N_34);
xnor U562 (N_562,In_1197,In_365);
and U563 (N_563,In_1061,N_142);
and U564 (N_564,N_212,In_1025);
or U565 (N_565,In_363,N_421);
and U566 (N_566,N_13,N_150);
xor U567 (N_567,In_672,In_688);
nor U568 (N_568,N_329,In_913);
nand U569 (N_569,In_571,N_206);
or U570 (N_570,In_696,In_1139);
and U571 (N_571,N_11,N_422);
nor U572 (N_572,In_220,N_361);
and U573 (N_573,In_1170,In_281);
and U574 (N_574,In_20,In_1499);
or U575 (N_575,In_334,N_262);
nor U576 (N_576,In_804,In_628);
xor U577 (N_577,In_662,In_391);
xor U578 (N_578,N_427,In_668);
and U579 (N_579,In_1174,N_374);
nor U580 (N_580,In_230,N_331);
and U581 (N_581,N_103,In_727);
and U582 (N_582,In_899,N_179);
and U583 (N_583,In_784,N_223);
xor U584 (N_584,N_86,N_393);
or U585 (N_585,In_961,N_65);
and U586 (N_586,In_787,In_790);
or U587 (N_587,N_259,In_1053);
xnor U588 (N_588,In_1077,N_386);
and U589 (N_589,In_1463,N_24);
nand U590 (N_590,In_177,In_1235);
nor U591 (N_591,In_283,N_408);
nor U592 (N_592,In_1334,In_1208);
nor U593 (N_593,In_960,In_1057);
nor U594 (N_594,In_456,N_152);
nand U595 (N_595,In_1452,In_104);
nand U596 (N_596,In_1142,In_1338);
nand U597 (N_597,In_1319,In_731);
or U598 (N_598,N_341,In_333);
xnor U599 (N_599,In_893,In_1291);
or U600 (N_600,In_113,In_338);
nand U601 (N_601,N_237,In_56);
xnor U602 (N_602,In_999,In_829);
and U603 (N_603,In_842,In_1149);
or U604 (N_604,N_95,N_564);
and U605 (N_605,In_518,N_330);
nor U606 (N_606,N_582,N_410);
nand U607 (N_607,N_469,N_420);
xnor U608 (N_608,N_592,In_877);
and U609 (N_609,In_1384,N_328);
and U610 (N_610,N_505,In_418);
or U611 (N_611,N_577,N_492);
nor U612 (N_612,In_1496,In_1117);
nand U613 (N_613,N_241,N_136);
and U614 (N_614,In_848,In_486);
or U615 (N_615,In_118,N_204);
and U616 (N_616,N_373,N_2);
nor U617 (N_617,N_588,N_171);
nand U618 (N_618,In_741,N_394);
nor U619 (N_619,In_713,N_317);
nand U620 (N_620,In_202,In_170);
nand U621 (N_621,N_168,In_644);
and U622 (N_622,In_1391,N_43);
xor U623 (N_623,N_482,In_434);
nand U624 (N_624,In_1303,N_322);
nor U625 (N_625,N_399,N_107);
nand U626 (N_626,In_409,In_436);
or U627 (N_627,In_910,N_337);
xor U628 (N_628,In_903,N_251);
or U629 (N_629,In_529,N_62);
or U630 (N_630,In_1198,N_336);
nand U631 (N_631,N_574,N_451);
and U632 (N_632,In_1238,N_397);
xnor U633 (N_633,N_120,In_819);
and U634 (N_634,In_1340,N_380);
or U635 (N_635,In_505,N_429);
xnor U636 (N_636,In_23,N_560);
nand U637 (N_637,In_602,In_541);
xor U638 (N_638,In_791,In_1114);
nor U639 (N_639,In_1443,In_205);
xor U640 (N_640,In_986,N_516);
or U641 (N_641,N_475,N_597);
nor U642 (N_642,N_80,In_638);
and U643 (N_643,In_235,In_77);
xnor U644 (N_644,In_927,N_134);
nor U645 (N_645,In_63,N_52);
and U646 (N_646,N_471,In_214);
nor U647 (N_647,In_780,In_128);
nor U648 (N_648,N_477,N_286);
and U649 (N_649,N_293,In_132);
or U650 (N_650,In_1458,In_1483);
nor U651 (N_651,In_1015,In_1475);
xor U652 (N_652,In_482,In_582);
and U653 (N_653,In_1278,N_294);
nor U654 (N_654,N_453,In_1372);
nor U655 (N_655,N_288,In_634);
xor U656 (N_656,In_476,N_507);
or U657 (N_657,In_586,N_550);
or U658 (N_658,In_1487,N_332);
nand U659 (N_659,In_614,N_319);
xnor U660 (N_660,N_572,In_1421);
nor U661 (N_661,In_387,N_503);
nor U662 (N_662,N_312,In_857);
or U663 (N_663,In_888,N_226);
nand U664 (N_664,In_473,N_543);
nor U665 (N_665,In_673,In_360);
or U666 (N_666,N_348,In_439);
xor U667 (N_667,N_296,N_228);
nand U668 (N_668,N_236,N_465);
nor U669 (N_669,In_705,In_856);
or U670 (N_670,N_534,N_436);
and U671 (N_671,In_105,N_159);
nand U672 (N_672,N_464,N_221);
xnor U673 (N_673,In_48,N_510);
nand U674 (N_674,In_1001,N_108);
nand U675 (N_675,In_1393,In_175);
nand U676 (N_676,N_55,In_1348);
and U677 (N_677,In_336,N_60);
xor U678 (N_678,In_298,In_658);
nor U679 (N_679,In_526,N_239);
xnor U680 (N_680,In_1225,N_443);
and U681 (N_681,In_425,In_971);
or U682 (N_682,N_489,N_486);
or U683 (N_683,In_1055,In_838);
and U684 (N_684,N_56,N_47);
nor U685 (N_685,In_1414,N_304);
and U686 (N_686,In_97,N_215);
nand U687 (N_687,N_172,In_361);
xor U688 (N_688,In_1078,In_871);
nor U689 (N_689,N_468,N_352);
xor U690 (N_690,In_1242,N_565);
and U691 (N_691,In_528,N_595);
nor U692 (N_692,N_458,N_218);
and U693 (N_693,In_129,N_135);
xnor U694 (N_694,In_1410,In_824);
or U695 (N_695,N_127,In_825);
xor U696 (N_696,N_539,In_150);
xor U697 (N_697,N_314,N_391);
nor U698 (N_698,N_71,In_1432);
and U699 (N_699,In_270,In_417);
xor U700 (N_700,In_1325,N_490);
nor U701 (N_701,N_78,In_236);
nor U702 (N_702,N_379,In_901);
nand U703 (N_703,In_1207,In_1427);
xor U704 (N_704,In_764,N_434);
xnor U705 (N_705,In_868,In_180);
nand U706 (N_706,In_573,In_600);
xor U707 (N_707,N_263,N_457);
xnor U708 (N_708,In_1068,N_568);
and U709 (N_709,N_562,N_359);
and U710 (N_710,In_448,In_187);
nand U711 (N_711,N_456,N_261);
or U712 (N_712,N_94,In_81);
nand U713 (N_713,N_147,N_481);
and U714 (N_714,N_174,In_285);
and U715 (N_715,In_503,In_383);
or U716 (N_716,In_572,In_138);
xnor U717 (N_717,N_558,N_478);
or U718 (N_718,In_795,In_310);
and U719 (N_719,N_557,N_476);
or U720 (N_720,In_1282,N_460);
nor U721 (N_721,N_117,N_524);
xnor U722 (N_722,N_118,N_227);
xnor U723 (N_723,N_508,In_1073);
nor U724 (N_724,In_521,In_316);
xor U725 (N_725,In_166,In_34);
or U726 (N_726,In_355,In_1103);
or U727 (N_727,In_496,N_91);
xnor U728 (N_728,In_396,N_366);
nor U729 (N_729,In_141,In_1376);
or U730 (N_730,In_165,In_1116);
nor U731 (N_731,N_497,N_245);
nor U732 (N_732,In_699,In_1105);
nor U733 (N_733,In_712,N_271);
xor U734 (N_734,In_1228,In_1173);
or U735 (N_735,N_404,In_7);
or U736 (N_736,N_51,In_258);
nand U737 (N_737,In_1043,In_1019);
nor U738 (N_738,N_428,N_511);
and U739 (N_739,In_608,N_195);
and U740 (N_740,N_177,In_495);
nand U741 (N_741,N_356,In_245);
nor U742 (N_742,N_63,In_872);
and U743 (N_743,In_1250,In_57);
or U744 (N_744,N_584,In_589);
nand U745 (N_745,N_243,In_1123);
nor U746 (N_746,In_419,N_447);
or U747 (N_747,In_493,N_498);
and U748 (N_748,In_657,N_523);
nand U749 (N_749,In_1158,In_15);
or U750 (N_750,N_438,N_192);
xnor U751 (N_751,In_384,N_700);
or U752 (N_752,In_1104,In_1361);
and U753 (N_753,In_1347,In_911);
nor U754 (N_754,N_705,N_485);
and U755 (N_755,N_570,In_631);
nor U756 (N_756,N_184,N_716);
nor U757 (N_757,In_792,N_369);
or U758 (N_758,In_1415,In_33);
or U759 (N_759,In_950,In_293);
or U760 (N_760,N_728,N_496);
or U761 (N_761,In_1212,N_741);
xor U762 (N_762,N_260,In_964);
or U763 (N_763,In_6,In_1039);
or U764 (N_764,In_820,N_273);
nand U765 (N_765,In_1448,In_749);
or U766 (N_766,In_119,N_439);
xnor U767 (N_767,In_61,In_998);
xor U768 (N_768,In_377,N_216);
xnor U769 (N_769,N_115,In_1300);
and U770 (N_770,In_480,In_403);
xor U771 (N_771,N_462,In_329);
nand U772 (N_772,In_1109,In_1279);
nor U773 (N_773,N_583,N_546);
xnor U774 (N_774,In_21,In_1249);
nand U775 (N_775,In_276,N_387);
nor U776 (N_776,In_29,In_369);
and U777 (N_777,In_1314,N_266);
nor U778 (N_778,In_197,In_590);
or U779 (N_779,In_1115,N_670);
xnor U780 (N_780,N_18,In_1484);
nand U781 (N_781,N_697,In_420);
nand U782 (N_782,In_302,In_621);
and U783 (N_783,In_1359,In_474);
xnor U784 (N_784,N_594,N_351);
xor U785 (N_785,N_372,N_668);
or U786 (N_786,N_157,In_854);
and U787 (N_787,In_743,N_474);
xnor U788 (N_788,N_122,In_1176);
nand U789 (N_789,N_89,N_194);
xnor U790 (N_790,N_579,N_416);
nand U791 (N_791,In_1398,In_1486);
and U792 (N_792,N_242,N_87);
xor U793 (N_793,N_694,N_246);
nand U794 (N_794,N_338,In_1335);
and U795 (N_795,N_180,N_711);
nor U796 (N_796,In_639,N_640);
nor U797 (N_797,N_688,In_902);
nand U798 (N_798,In_86,N_355);
nor U799 (N_799,N_655,In_507);
nand U800 (N_800,In_139,N_375);
nand U801 (N_801,N_571,N_402);
nand U802 (N_802,In_542,N_730);
nor U803 (N_803,In_965,N_639);
and U804 (N_804,N_567,N_590);
xnor U805 (N_805,N_138,N_406);
or U806 (N_806,N_365,N_624);
nand U807 (N_807,In_488,In_1447);
or U808 (N_808,N_225,In_941);
xor U809 (N_809,In_226,In_181);
xnor U810 (N_810,In_393,N_256);
nor U811 (N_811,In_415,N_522);
xnor U812 (N_812,In_778,N_311);
or U813 (N_813,In_806,N_529);
nand U814 (N_814,N_545,N_551);
nand U815 (N_815,N_170,N_415);
xor U816 (N_816,N_712,In_1402);
xnor U817 (N_817,N_502,N_327);
nand U818 (N_818,N_210,N_535);
and U819 (N_819,N_605,In_172);
or U820 (N_820,In_708,N_735);
and U821 (N_821,In_676,N_42);
nand U822 (N_822,In_1397,In_610);
nor U823 (N_823,In_135,N_708);
nand U824 (N_824,In_88,In_208);
and U825 (N_825,N_193,N_721);
and U826 (N_826,N_649,In_1386);
and U827 (N_827,N_473,N_240);
or U828 (N_828,N_686,In_386);
and U829 (N_829,N_112,N_548);
nand U830 (N_830,N_631,N_275);
nor U831 (N_831,N_702,N_155);
nor U832 (N_832,N_176,N_608);
and U833 (N_833,N_343,N_648);
nand U834 (N_834,N_746,N_547);
nor U835 (N_835,In_1408,In_243);
xor U836 (N_836,In_1060,In_73);
nor U837 (N_837,N_606,In_924);
nand U838 (N_838,In_711,N_306);
nor U839 (N_839,N_603,N_513);
nor U840 (N_840,N_723,N_491);
xnor U841 (N_841,N_334,In_799);
xor U842 (N_842,N_559,N_437);
nor U843 (N_843,N_611,In_551);
nor U844 (N_844,N_209,In_74);
xnor U845 (N_845,N_201,In_328);
nand U846 (N_846,In_810,In_828);
xor U847 (N_847,In_108,In_1489);
or U848 (N_848,In_1267,N_743);
xor U849 (N_849,In_37,N_724);
nand U850 (N_850,In_1066,N_353);
nand U851 (N_851,In_1091,In_1255);
nand U852 (N_852,In_1121,N_636);
and U853 (N_853,In_898,N_691);
and U854 (N_854,N_736,N_250);
or U855 (N_855,In_811,N_274);
or U856 (N_856,N_674,In_624);
or U857 (N_857,In_525,N_706);
or U858 (N_858,N_709,In_782);
xor U859 (N_859,N_470,N_360);
nor U860 (N_860,In_953,N_575);
nand U861 (N_861,In_921,In_26);
and U862 (N_862,N_740,N_198);
nand U863 (N_863,N_450,N_390);
and U864 (N_864,N_363,In_1367);
and U865 (N_865,In_875,N_149);
nor U866 (N_866,In_206,N_75);
and U867 (N_867,N_161,In_1045);
and U868 (N_868,In_735,N_690);
nor U869 (N_869,N_333,In_851);
and U870 (N_870,N_388,In_687);
nand U871 (N_871,In_775,N_310);
xor U872 (N_872,N_315,N_720);
xnor U873 (N_873,N_82,In_742);
xnor U874 (N_874,In_1195,N_556);
nor U875 (N_875,In_510,N_146);
xnor U876 (N_876,N_610,N_585);
and U877 (N_877,In_72,N_270);
and U878 (N_878,N_400,N_521);
nor U879 (N_879,N_675,N_653);
and U880 (N_880,In_922,N_693);
xnor U881 (N_881,N_666,In_1159);
nor U882 (N_882,In_1081,N_472);
or U883 (N_883,In_994,In_1375);
nand U884 (N_884,N_738,In_973);
or U885 (N_885,N_418,In_519);
and U886 (N_886,N_561,In_1336);
xor U887 (N_887,In_122,In_430);
xor U888 (N_888,N_628,In_751);
and U889 (N_889,In_807,In_974);
nand U890 (N_890,N_196,In_1360);
nor U891 (N_891,N_431,N_596);
nor U892 (N_892,N_483,In_274);
xnor U893 (N_893,In_802,In_251);
or U894 (N_894,N_660,In_559);
xor U895 (N_895,N_656,N_309);
nand U896 (N_896,N_707,In_116);
xnor U897 (N_897,In_43,N_710);
nand U898 (N_898,In_880,N_377);
xor U899 (N_899,In_985,N_526);
or U900 (N_900,N_872,N_542);
or U901 (N_901,In_640,N_851);
and U902 (N_902,In_75,In_1083);
nand U903 (N_903,In_797,N_345);
and U904 (N_904,In_144,In_475);
or U905 (N_905,N_525,N_619);
nor U906 (N_906,In_1051,N_808);
xnor U907 (N_907,N_650,N_621);
xnor U908 (N_908,In_1032,In_269);
nand U909 (N_909,N_385,N_862);
xor U910 (N_910,N_222,In_300);
or U911 (N_911,In_915,N_683);
nand U912 (N_912,N_701,In_1392);
xnor U913 (N_913,N_714,N_806);
and U914 (N_914,N_658,N_748);
nor U915 (N_915,N_541,N_634);
xnor U916 (N_916,In_1456,N_892);
nand U917 (N_917,In_388,N_812);
nand U918 (N_918,N_835,In_1023);
nand U919 (N_919,N_613,N_871);
and U920 (N_920,N_843,In_341);
nor U921 (N_921,N_652,N_520);
and U922 (N_922,N_672,N_553);
xnor U923 (N_923,N_833,In_1301);
xor U924 (N_924,In_112,In_1122);
nor U925 (N_925,In_227,N_795);
nand U926 (N_926,In_1330,N_889);
or U927 (N_927,N_888,N_616);
or U928 (N_928,N_452,N_620);
and U929 (N_929,N_780,In_1275);
nor U930 (N_930,N_249,In_1455);
nor U931 (N_931,N_635,In_307);
and U932 (N_932,N_129,N_680);
nor U933 (N_933,N_466,N_776);
nor U934 (N_934,N_869,N_687);
nand U935 (N_935,N_73,N_853);
and U936 (N_936,N_758,N_495);
or U937 (N_937,N_845,In_979);
xnor U938 (N_938,N_796,N_576);
xor U939 (N_939,N_817,N_778);
and U940 (N_940,N_659,N_822);
nand U941 (N_941,N_825,N_868);
nand U942 (N_942,In_70,In_876);
nand U943 (N_943,In_1395,In_1152);
nand U944 (N_944,N_876,N_164);
nand U945 (N_945,N_749,In_1309);
or U946 (N_946,N_626,In_762);
nand U947 (N_947,In_569,N_818);
nor U948 (N_948,N_580,N_747);
xnor U949 (N_949,N_770,In_440);
nor U950 (N_950,N_618,In_793);
nand U951 (N_951,In_217,N_753);
nor U952 (N_952,N_791,N_264);
and U953 (N_953,N_423,In_1232);
xnor U954 (N_954,In_832,N_877);
or U955 (N_955,N_90,In_38);
nor U956 (N_956,In_684,N_213);
nor U957 (N_957,In_948,N_819);
xnor U958 (N_958,In_1127,N_848);
nand U959 (N_959,N_854,In_22);
nor U960 (N_960,In_895,N_287);
nand U961 (N_961,In_719,N_739);
nand U962 (N_962,In_548,N_760);
nand U963 (N_963,N_633,In_767);
and U964 (N_964,N_141,N_790);
or U965 (N_965,N_362,N_737);
nor U966 (N_966,In_916,N_698);
xnor U967 (N_967,In_671,N_779);
or U968 (N_968,N_540,N_757);
nand U969 (N_969,N_695,In_454);
nor U970 (N_970,N_828,N_763);
nor U971 (N_971,N_681,In_748);
nand U972 (N_972,N_880,N_518);
nor U973 (N_973,In_1134,N_677);
nor U974 (N_974,In_28,N_667);
or U975 (N_975,In_30,In_1241);
and U976 (N_976,N_435,N_622);
xnor U977 (N_977,N_530,In_557);
nor U978 (N_978,In_1479,N_364);
and U979 (N_979,N_527,N_774);
xor U980 (N_980,N_744,In_852);
and U981 (N_981,N_555,N_661);
nor U982 (N_982,In_1481,In_1460);
or U983 (N_983,N_426,N_253);
and U984 (N_984,N_320,N_1);
xor U985 (N_985,N_480,N_789);
xnor U986 (N_986,N_268,N_751);
and U987 (N_987,N_882,N_600);
and U988 (N_988,N_30,N_517);
and U989 (N_989,In_1084,N_145);
nand U990 (N_990,In_1464,In_1070);
xor U991 (N_991,N_831,In_650);
nor U992 (N_992,In_183,N_623);
xor U993 (N_993,N_625,N_897);
nor U994 (N_994,N_786,In_783);
xnor U995 (N_995,N_303,N_852);
xnor U996 (N_996,In_935,In_813);
nor U997 (N_997,N_874,N_591);
nand U998 (N_998,In_1381,In_680);
and U999 (N_999,In_484,N_644);
xnor U1000 (N_1000,In_636,N_488);
nand U1001 (N_1001,N_813,In_1179);
and U1002 (N_1002,N_792,N_859);
and U1003 (N_1003,In_1281,In_349);
xor U1004 (N_1004,N_756,In_1033);
or U1005 (N_1005,N_857,N_589);
nor U1006 (N_1006,N_685,In_19);
nor U1007 (N_1007,N_726,N_811);
nor U1008 (N_1008,N_367,In_1213);
and U1009 (N_1009,In_1426,N_48);
nor U1010 (N_1010,In_978,In_881);
nor U1011 (N_1011,N_403,N_866);
nor U1012 (N_1012,N_731,N_759);
xor U1013 (N_1013,In_991,In_1080);
nor U1014 (N_1014,N_401,In_833);
nor U1015 (N_1015,N_769,N_132);
nand U1016 (N_1016,N_484,N_875);
or U1017 (N_1017,In_858,N_609);
nand U1018 (N_1018,N_601,In_1416);
and U1019 (N_1019,In_1295,In_1102);
and U1020 (N_1020,N_750,N_396);
nor U1021 (N_1021,N_834,In_247);
nand U1022 (N_1022,N_602,N_279);
xnor U1023 (N_1023,N_493,N_815);
or U1024 (N_1024,In_1362,N_895);
nand U1025 (N_1025,N_827,N_614);
nor U1026 (N_1026,In_45,N_814);
nor U1027 (N_1027,N_784,N_768);
or U1028 (N_1028,N_837,In_263);
or U1029 (N_1029,N_578,N_842);
and U1030 (N_1030,In_1029,In_121);
nand U1031 (N_1031,N_467,N_598);
and U1032 (N_1032,In_1313,In_184);
nor U1033 (N_1033,In_90,N_745);
nand U1034 (N_1034,In_1095,N_499);
or U1035 (N_1035,N_208,N_487);
or U1036 (N_1036,In_674,N_604);
nor U1037 (N_1037,N_370,N_841);
or U1038 (N_1038,N_870,N_504);
xnor U1039 (N_1039,N_461,N_891);
nand U1040 (N_1040,N_627,In_698);
or U1041 (N_1041,N_673,In_1165);
or U1042 (N_1042,In_149,N_800);
or U1043 (N_1043,N_821,N_849);
nor U1044 (N_1044,N_787,N_713);
nand U1045 (N_1045,In_706,N_325);
nor U1046 (N_1046,N_865,N_662);
nor U1047 (N_1047,In_817,In_931);
or U1048 (N_1048,In_343,N_479);
nor U1049 (N_1049,N_642,N_573);
nor U1050 (N_1050,N_927,N_16);
nor U1051 (N_1051,In_900,N_1024);
xnor U1052 (N_1052,In_715,N_931);
nor U1053 (N_1053,N_32,In_830);
nand U1054 (N_1054,N_900,N_918);
xnor U1055 (N_1055,N_963,N_802);
nand U1056 (N_1056,N_727,In_291);
xnor U1057 (N_1057,N_765,N_761);
nand U1058 (N_1058,N_494,In_1494);
nor U1059 (N_1059,N_1011,N_905);
or U1060 (N_1060,N_860,N_973);
nand U1061 (N_1061,N_908,N_902);
or U1062 (N_1062,N_969,N_432);
nand U1063 (N_1063,N_785,N_189);
or U1064 (N_1064,N_794,N_979);
and U1065 (N_1065,In_878,N_956);
nand U1066 (N_1066,N_816,N_939);
or U1067 (N_1067,N_699,N_989);
and U1068 (N_1068,N_247,N_719);
or U1069 (N_1069,N_920,In_27);
nand U1070 (N_1070,N_966,N_342);
nand U1071 (N_1071,N_637,In_1467);
nand U1072 (N_1072,N_982,In_643);
nor U1073 (N_1073,In_188,N_732);
nor U1074 (N_1074,N_647,N_890);
or U1075 (N_1075,N_907,N_1025);
and U1076 (N_1076,In_1064,In_619);
nor U1077 (N_1077,N_663,In_701);
nor U1078 (N_1078,N_904,N_1027);
and U1079 (N_1079,N_722,N_641);
and U1080 (N_1080,N_867,N_994);
nor U1081 (N_1081,N_389,N_896);
nor U1082 (N_1082,N_893,N_544);
xnor U1083 (N_1083,N_941,N_948);
nor U1084 (N_1084,In_1316,N_501);
or U1085 (N_1085,N_928,N_1018);
nand U1086 (N_1086,N_915,In_597);
or U1087 (N_1087,N_783,N_68);
xor U1088 (N_1088,N_968,In_378);
nor U1089 (N_1089,In_275,N_910);
and U1090 (N_1090,N_1004,In_481);
nand U1091 (N_1091,N_188,N_1034);
and U1092 (N_1092,In_1344,N_657);
nor U1093 (N_1093,In_543,N_519);
xnor U1094 (N_1094,N_798,N_970);
nand U1095 (N_1095,N_459,N_376);
nor U1096 (N_1096,N_820,N_569);
nand U1097 (N_1097,N_554,N_514);
or U1098 (N_1098,N_836,N_788);
nand U1099 (N_1099,N_455,N_913);
and U1100 (N_1100,In_228,N_899);
xor U1101 (N_1101,N_630,N_1047);
nor U1102 (N_1102,N_413,N_629);
nand U1103 (N_1103,N_267,N_1016);
or U1104 (N_1104,In_805,N_1046);
and U1105 (N_1105,N_66,N_917);
or U1106 (N_1106,N_232,N_301);
and U1107 (N_1107,N_946,N_654);
or U1108 (N_1108,N_885,In_860);
nor U1109 (N_1109,N_307,N_1033);
and U1110 (N_1110,N_901,In_938);
nand U1111 (N_1111,N_531,In_1093);
nand U1112 (N_1112,N_651,In_92);
nor U1113 (N_1113,In_1150,N_230);
and U1114 (N_1114,N_991,N_799);
nand U1115 (N_1115,N_914,In_47);
nand U1116 (N_1116,In_117,N_265);
nand U1117 (N_1117,N_536,N_940);
xor U1118 (N_1118,N_684,N_669);
nand U1119 (N_1119,N_772,In_319);
xor U1120 (N_1120,N_988,In_781);
or U1121 (N_1121,In_41,N_679);
nand U1122 (N_1122,N_323,N_1028);
xnor U1123 (N_1123,In_520,In_1271);
nand U1124 (N_1124,N_433,N_990);
and U1125 (N_1125,N_678,In_1264);
and U1126 (N_1126,N_826,N_960);
xnor U1127 (N_1127,N_858,N_974);
nor U1128 (N_1128,N_921,N_587);
and U1129 (N_1129,In_1231,N_88);
nand U1130 (N_1130,N_775,N_277);
or U1131 (N_1131,N_552,N_563);
or U1132 (N_1132,In_632,In_1062);
or U1133 (N_1133,N_771,N_830);
nand U1134 (N_1134,In_407,N_949);
or U1135 (N_1135,N_692,N_1012);
xor U1136 (N_1136,In_669,N_916);
or U1137 (N_1137,N_165,In_1136);
and U1138 (N_1138,N_873,N_114);
nand U1139 (N_1139,N_581,N_840);
xor U1140 (N_1140,N_1013,N_906);
and U1141 (N_1141,In_554,N_1044);
xnor U1142 (N_1142,In_1472,N_883);
nor U1143 (N_1143,N_955,N_1015);
xnor U1144 (N_1144,N_944,In_1199);
or U1145 (N_1145,N_958,In_0);
xnor U1146 (N_1146,N_506,N_951);
and U1147 (N_1147,N_980,N_346);
or U1148 (N_1148,In_93,N_953);
or U1149 (N_1149,In_1030,N_764);
nand U1150 (N_1150,N_599,N_887);
xnor U1151 (N_1151,N_926,N_823);
xnor U1152 (N_1152,In_786,N_1041);
xnor U1153 (N_1153,N_878,N_664);
nand U1154 (N_1154,N_954,N_929);
nand U1155 (N_1155,N_999,N_1001);
or U1156 (N_1156,N_793,N_898);
nand U1157 (N_1157,In_549,In_1168);
and U1158 (N_1158,N_1010,N_935);
nand U1159 (N_1159,N_972,N_1035);
or U1160 (N_1160,N_824,N_704);
and U1161 (N_1161,N_538,N_128);
nand U1162 (N_1162,N_942,N_566);
nor U1163 (N_1163,N_923,N_838);
nand U1164 (N_1164,N_1039,In_1209);
xnor U1165 (N_1165,N_646,In_9);
or U1166 (N_1166,N_444,N_925);
nor U1167 (N_1167,N_932,N_632);
nand U1168 (N_1168,In_1403,N_463);
xnor U1169 (N_1169,N_612,N_992);
and U1170 (N_1170,N_959,N_952);
nor U1171 (N_1171,N_801,In_427);
nor U1172 (N_1172,N_729,N_909);
and U1173 (N_1173,N_1021,N_1049);
xnor U1174 (N_1174,N_809,N_919);
nor U1175 (N_1175,N_981,N_844);
or U1176 (N_1176,N_781,N_153);
nand U1177 (N_1177,N_607,N_804);
xnor U1178 (N_1178,N_755,In_816);
xnor U1179 (N_1179,N_412,In_1007);
and U1180 (N_1180,N_500,N_856);
or U1181 (N_1181,N_855,In_997);
and U1182 (N_1182,N_1008,N_617);
and U1183 (N_1183,N_1048,N_725);
nand U1184 (N_1184,N_975,N_515);
xnor U1185 (N_1185,N_879,N_339);
xor U1186 (N_1186,N_803,N_280);
or U1187 (N_1187,In_553,In_1211);
or U1188 (N_1188,In_1253,N_638);
nand U1189 (N_1189,In_1446,N_937);
nor U1190 (N_1190,In_1369,N_933);
nor U1191 (N_1191,N_81,In_1354);
nand U1192 (N_1192,N_665,N_4);
nor U1193 (N_1193,N_762,In_282);
or U1194 (N_1194,In_612,N_528);
or U1195 (N_1195,In_389,In_710);
nand U1196 (N_1196,N_593,N_986);
nor U1197 (N_1197,N_233,N_615);
or U1198 (N_1198,N_983,N_1007);
or U1199 (N_1199,N_671,N_586);
nand U1200 (N_1200,N_864,In_352);
nor U1201 (N_1201,N_1144,N_1171);
xnor U1202 (N_1202,In_35,N_1086);
or U1203 (N_1203,In_702,N_1196);
xnor U1204 (N_1204,N_832,N_1193);
and U1205 (N_1205,N_957,N_782);
xnor U1206 (N_1206,N_1064,N_1189);
nand U1207 (N_1207,N_1073,In_318);
nor U1208 (N_1208,N_1059,N_912);
nor U1209 (N_1209,N_1124,N_1162);
nor U1210 (N_1210,In_1305,N_1136);
xnor U1211 (N_1211,N_777,N_1150);
xor U1212 (N_1212,N_1062,N_1095);
nand U1213 (N_1213,N_1134,N_1178);
xor U1214 (N_1214,N_1186,N_676);
xnor U1215 (N_1215,N_1109,N_1123);
and U1216 (N_1216,N_1111,N_1002);
or U1217 (N_1217,N_1022,N_847);
nor U1218 (N_1218,N_1056,In_477);
nand U1219 (N_1219,N_752,N_850);
or U1220 (N_1220,N_976,N_1194);
and U1221 (N_1221,N_1187,N_1172);
nand U1222 (N_1222,N_717,N_1169);
or U1223 (N_1223,N_903,N_1076);
or U1224 (N_1224,N_1102,N_805);
nand U1225 (N_1225,N_1094,N_1067);
or U1226 (N_1226,N_1131,N_911);
nor U1227 (N_1227,N_1098,N_884);
nand U1228 (N_1228,N_1063,N_378);
nand U1229 (N_1229,N_1106,In_1434);
nor U1230 (N_1230,N_947,N_773);
xnor U1231 (N_1231,N_1032,N_1148);
nor U1232 (N_1232,N_1164,N_1085);
nor U1233 (N_1233,N_1151,N_863);
xnor U1234 (N_1234,In_154,N_1199);
xor U1235 (N_1235,N_1158,N_291);
and U1236 (N_1236,N_1177,N_1129);
xnor U1237 (N_1237,N_1092,N_829);
nor U1238 (N_1238,N_924,N_1184);
nor U1239 (N_1239,N_537,N_1080);
nand U1240 (N_1240,N_1055,N_1137);
nand U1241 (N_1241,N_1082,N_1188);
xnor U1242 (N_1242,N_967,In_1244);
xnor U1243 (N_1243,In_808,N_1023);
nor U1244 (N_1244,N_881,N_754);
and U1245 (N_1245,N_1070,N_1170);
xnor U1246 (N_1246,N_1197,In_1111);
xor U1247 (N_1247,N_1152,N_682);
and U1248 (N_1248,N_1104,N_936);
or U1249 (N_1249,In_583,N_69);
nand U1250 (N_1250,In_1094,N_1147);
and U1251 (N_1251,N_1115,N_1116);
nand U1252 (N_1252,N_1005,N_934);
nor U1253 (N_1253,N_846,N_1058);
nand U1254 (N_1254,N_1006,N_943);
xor U1255 (N_1255,N_509,N_718);
nor U1256 (N_1256,N_1192,N_1083);
and U1257 (N_1257,N_1045,N_938);
nand U1258 (N_1258,In_421,N_1140);
nor U1259 (N_1259,N_1026,N_1185);
xor U1260 (N_1260,N_1072,N_1071);
and U1261 (N_1261,In_752,N_1014);
nor U1262 (N_1262,N_36,N_1068);
nand U1263 (N_1263,N_839,N_512);
and U1264 (N_1264,N_1017,N_742);
nand U1265 (N_1265,N_645,N_354);
and U1266 (N_1266,N_1156,N_1069);
nand U1267 (N_1267,N_39,N_281);
or U1268 (N_1268,N_1105,N_1128);
nor U1269 (N_1269,N_1043,In_367);
nand U1270 (N_1270,N_962,N_1113);
xor U1271 (N_1271,N_643,N_1159);
and U1272 (N_1272,N_430,N_1009);
xor U1273 (N_1273,N_1112,N_1167);
or U1274 (N_1274,N_1040,N_1103);
xor U1275 (N_1275,N_1132,In_1290);
xnor U1276 (N_1276,N_984,N_1174);
nand U1277 (N_1277,In_723,N_1096);
nand U1278 (N_1278,N_886,N_1180);
nand U1279 (N_1279,N_1126,N_978);
xnor U1280 (N_1280,N_398,N_1165);
xor U1281 (N_1281,N_532,N_1175);
or U1282 (N_1282,N_1097,N_995);
nand U1283 (N_1283,N_1029,N_1139);
or U1284 (N_1284,N_1038,N_971);
or U1285 (N_1285,N_1182,N_1088);
xor U1286 (N_1286,N_1100,N_930);
xor U1287 (N_1287,N_1052,N_23);
xor U1288 (N_1288,N_549,N_733);
nor U1289 (N_1289,N_1166,N_797);
xnor U1290 (N_1290,N_1130,N_1053);
or U1291 (N_1291,In_176,N_1127);
nor U1292 (N_1292,N_965,N_1030);
xnor U1293 (N_1293,N_998,N_533);
nor U1294 (N_1294,N_1117,In_1341);
nor U1295 (N_1295,In_173,N_1121);
and U1296 (N_1296,N_894,N_383);
nand U1297 (N_1297,N_996,N_1168);
nand U1298 (N_1298,N_1160,N_1093);
nand U1299 (N_1299,N_1157,In_707);
nand U1300 (N_1300,In_595,In_823);
nand U1301 (N_1301,N_316,N_1141);
and U1302 (N_1302,N_1198,N_1179);
nor U1303 (N_1303,N_987,N_997);
xnor U1304 (N_1304,In_1351,N_703);
or U1305 (N_1305,N_961,N_1089);
xnor U1306 (N_1306,N_454,In_874);
xor U1307 (N_1307,N_1146,N_1020);
or U1308 (N_1308,N_97,N_1000);
nand U1309 (N_1309,N_977,N_1019);
or U1310 (N_1310,N_1145,N_1101);
or U1311 (N_1311,N_945,N_807);
or U1312 (N_1312,N_1143,N_1163);
or U1313 (N_1313,N_1066,N_1118);
and U1314 (N_1314,N_734,N_964);
and U1315 (N_1315,N_861,N_1135);
and U1316 (N_1316,N_1037,N_689);
or U1317 (N_1317,In_1289,N_1149);
or U1318 (N_1318,N_766,N_1087);
nor U1319 (N_1319,N_1075,N_1108);
and U1320 (N_1320,N_1031,N_1107);
nand U1321 (N_1321,N_993,N_1110);
xor U1322 (N_1322,N_1003,N_1154);
nor U1323 (N_1323,N_1078,N_1114);
or U1324 (N_1324,N_1054,In_905);
xor U1325 (N_1325,N_1081,N_308);
nand U1326 (N_1326,In_827,N_1099);
and U1327 (N_1327,N_238,N_1153);
nor U1328 (N_1328,N_1122,N_1138);
or U1329 (N_1329,N_1125,N_810);
or U1330 (N_1330,N_1050,N_1120);
xor U1331 (N_1331,N_1091,N_1065);
or U1332 (N_1332,N_1051,N_1042);
or U1333 (N_1333,N_767,N_1036);
xor U1334 (N_1334,N_1191,N_696);
or U1335 (N_1335,N_1183,N_715);
and U1336 (N_1336,N_1061,N_1074);
nand U1337 (N_1337,N_1077,N_1090);
nor U1338 (N_1338,N_950,N_1060);
xor U1339 (N_1339,N_1195,N_1173);
or U1340 (N_1340,N_244,N_1155);
and U1341 (N_1341,N_305,In_591);
nor U1342 (N_1342,N_1057,N_1181);
or U1343 (N_1343,N_1084,In_1495);
nor U1344 (N_1344,N_1133,N_922);
nor U1345 (N_1345,N_1176,N_191);
and U1346 (N_1346,N_1190,N_1119);
xnor U1347 (N_1347,N_1142,N_985);
and U1348 (N_1348,N_1079,In_423);
xor U1349 (N_1349,In_1288,N_1161);
and U1350 (N_1350,N_1328,N_1319);
or U1351 (N_1351,N_1318,N_1220);
xor U1352 (N_1352,N_1298,N_1215);
or U1353 (N_1353,N_1206,N_1279);
xnor U1354 (N_1354,N_1346,N_1272);
or U1355 (N_1355,N_1312,N_1208);
nand U1356 (N_1356,N_1333,N_1256);
or U1357 (N_1357,N_1265,N_1264);
xor U1358 (N_1358,N_1271,N_1300);
or U1359 (N_1359,N_1254,N_1270);
nand U1360 (N_1360,N_1348,N_1224);
nor U1361 (N_1361,N_1291,N_1303);
and U1362 (N_1362,N_1336,N_1221);
xor U1363 (N_1363,N_1246,N_1232);
nand U1364 (N_1364,N_1259,N_1324);
xor U1365 (N_1365,N_1209,N_1268);
and U1366 (N_1366,N_1249,N_1340);
nand U1367 (N_1367,N_1330,N_1280);
and U1368 (N_1368,N_1201,N_1341);
and U1369 (N_1369,N_1299,N_1257);
xor U1370 (N_1370,N_1205,N_1304);
nand U1371 (N_1371,N_1200,N_1229);
nand U1372 (N_1372,N_1210,N_1293);
or U1373 (N_1373,N_1243,N_1316);
and U1374 (N_1374,N_1250,N_1326);
and U1375 (N_1375,N_1202,N_1331);
nor U1376 (N_1376,N_1231,N_1251);
nor U1377 (N_1377,N_1325,N_1218);
and U1378 (N_1378,N_1323,N_1222);
nor U1379 (N_1379,N_1238,N_1241);
and U1380 (N_1380,N_1253,N_1327);
nand U1381 (N_1381,N_1267,N_1347);
xor U1382 (N_1382,N_1236,N_1309);
or U1383 (N_1383,N_1235,N_1296);
xor U1384 (N_1384,N_1301,N_1204);
nor U1385 (N_1385,N_1227,N_1311);
nand U1386 (N_1386,N_1349,N_1219);
nor U1387 (N_1387,N_1307,N_1214);
or U1388 (N_1388,N_1230,N_1226);
and U1389 (N_1389,N_1233,N_1313);
nor U1390 (N_1390,N_1290,N_1344);
and U1391 (N_1391,N_1305,N_1239);
xor U1392 (N_1392,N_1322,N_1203);
nor U1393 (N_1393,N_1286,N_1288);
nand U1394 (N_1394,N_1310,N_1275);
nor U1395 (N_1395,N_1321,N_1345);
or U1396 (N_1396,N_1284,N_1225);
xor U1397 (N_1397,N_1237,N_1252);
nand U1398 (N_1398,N_1337,N_1223);
nor U1399 (N_1399,N_1332,N_1248);
or U1400 (N_1400,N_1295,N_1289);
nand U1401 (N_1401,N_1315,N_1283);
or U1402 (N_1402,N_1244,N_1334);
or U1403 (N_1403,N_1329,N_1217);
or U1404 (N_1404,N_1320,N_1263);
xor U1405 (N_1405,N_1292,N_1281);
nand U1406 (N_1406,N_1234,N_1294);
or U1407 (N_1407,N_1262,N_1306);
nor U1408 (N_1408,N_1317,N_1266);
and U1409 (N_1409,N_1245,N_1278);
nor U1410 (N_1410,N_1285,N_1261);
and U1411 (N_1411,N_1258,N_1314);
nand U1412 (N_1412,N_1240,N_1212);
and U1413 (N_1413,N_1342,N_1242);
nand U1414 (N_1414,N_1255,N_1308);
xor U1415 (N_1415,N_1335,N_1213);
nor U1416 (N_1416,N_1247,N_1228);
nand U1417 (N_1417,N_1273,N_1343);
nor U1418 (N_1418,N_1338,N_1260);
nand U1419 (N_1419,N_1274,N_1302);
nand U1420 (N_1420,N_1297,N_1216);
or U1421 (N_1421,N_1282,N_1211);
nand U1422 (N_1422,N_1276,N_1287);
nand U1423 (N_1423,N_1269,N_1277);
nor U1424 (N_1424,N_1207,N_1339);
nand U1425 (N_1425,N_1280,N_1264);
nor U1426 (N_1426,N_1295,N_1239);
xnor U1427 (N_1427,N_1284,N_1255);
nand U1428 (N_1428,N_1270,N_1253);
and U1429 (N_1429,N_1287,N_1298);
nand U1430 (N_1430,N_1208,N_1248);
and U1431 (N_1431,N_1252,N_1216);
and U1432 (N_1432,N_1216,N_1249);
and U1433 (N_1433,N_1208,N_1327);
nand U1434 (N_1434,N_1287,N_1317);
or U1435 (N_1435,N_1292,N_1288);
nor U1436 (N_1436,N_1343,N_1341);
or U1437 (N_1437,N_1292,N_1301);
xor U1438 (N_1438,N_1314,N_1224);
or U1439 (N_1439,N_1265,N_1290);
nor U1440 (N_1440,N_1234,N_1252);
xnor U1441 (N_1441,N_1322,N_1333);
nor U1442 (N_1442,N_1250,N_1322);
or U1443 (N_1443,N_1209,N_1330);
nor U1444 (N_1444,N_1342,N_1280);
or U1445 (N_1445,N_1313,N_1311);
nand U1446 (N_1446,N_1213,N_1219);
nand U1447 (N_1447,N_1324,N_1276);
xnor U1448 (N_1448,N_1229,N_1242);
nor U1449 (N_1449,N_1242,N_1228);
and U1450 (N_1450,N_1307,N_1246);
and U1451 (N_1451,N_1283,N_1231);
and U1452 (N_1452,N_1339,N_1285);
or U1453 (N_1453,N_1206,N_1230);
nor U1454 (N_1454,N_1282,N_1322);
nor U1455 (N_1455,N_1296,N_1216);
nand U1456 (N_1456,N_1293,N_1243);
or U1457 (N_1457,N_1294,N_1322);
xnor U1458 (N_1458,N_1214,N_1266);
nor U1459 (N_1459,N_1201,N_1231);
xnor U1460 (N_1460,N_1269,N_1328);
nor U1461 (N_1461,N_1253,N_1231);
xor U1462 (N_1462,N_1246,N_1302);
or U1463 (N_1463,N_1308,N_1213);
or U1464 (N_1464,N_1273,N_1240);
xnor U1465 (N_1465,N_1240,N_1200);
nand U1466 (N_1466,N_1289,N_1316);
and U1467 (N_1467,N_1293,N_1255);
nand U1468 (N_1468,N_1293,N_1343);
nand U1469 (N_1469,N_1236,N_1237);
nand U1470 (N_1470,N_1333,N_1277);
xnor U1471 (N_1471,N_1301,N_1281);
nand U1472 (N_1472,N_1253,N_1206);
and U1473 (N_1473,N_1315,N_1253);
nor U1474 (N_1474,N_1206,N_1268);
and U1475 (N_1475,N_1339,N_1211);
nor U1476 (N_1476,N_1237,N_1330);
nand U1477 (N_1477,N_1332,N_1338);
nand U1478 (N_1478,N_1226,N_1338);
nand U1479 (N_1479,N_1205,N_1223);
nor U1480 (N_1480,N_1225,N_1200);
xor U1481 (N_1481,N_1240,N_1305);
or U1482 (N_1482,N_1264,N_1217);
nand U1483 (N_1483,N_1299,N_1324);
xnor U1484 (N_1484,N_1284,N_1327);
or U1485 (N_1485,N_1243,N_1283);
nor U1486 (N_1486,N_1319,N_1344);
nor U1487 (N_1487,N_1213,N_1276);
xor U1488 (N_1488,N_1312,N_1345);
xnor U1489 (N_1489,N_1247,N_1218);
nor U1490 (N_1490,N_1330,N_1315);
nor U1491 (N_1491,N_1201,N_1247);
xor U1492 (N_1492,N_1325,N_1270);
and U1493 (N_1493,N_1307,N_1302);
xor U1494 (N_1494,N_1280,N_1338);
and U1495 (N_1495,N_1285,N_1266);
and U1496 (N_1496,N_1218,N_1212);
nor U1497 (N_1497,N_1218,N_1256);
xor U1498 (N_1498,N_1336,N_1309);
xnor U1499 (N_1499,N_1238,N_1347);
nor U1500 (N_1500,N_1406,N_1389);
or U1501 (N_1501,N_1356,N_1451);
or U1502 (N_1502,N_1439,N_1482);
xnor U1503 (N_1503,N_1428,N_1413);
or U1504 (N_1504,N_1391,N_1432);
xor U1505 (N_1505,N_1447,N_1418);
xnor U1506 (N_1506,N_1452,N_1484);
nand U1507 (N_1507,N_1481,N_1483);
nor U1508 (N_1508,N_1459,N_1416);
or U1509 (N_1509,N_1443,N_1417);
nor U1510 (N_1510,N_1419,N_1373);
xnor U1511 (N_1511,N_1376,N_1380);
nand U1512 (N_1512,N_1393,N_1458);
nand U1513 (N_1513,N_1384,N_1433);
xor U1514 (N_1514,N_1405,N_1404);
xor U1515 (N_1515,N_1388,N_1485);
nand U1516 (N_1516,N_1424,N_1457);
nor U1517 (N_1517,N_1480,N_1397);
nand U1518 (N_1518,N_1449,N_1366);
and U1519 (N_1519,N_1411,N_1392);
nor U1520 (N_1520,N_1446,N_1464);
xnor U1521 (N_1521,N_1492,N_1450);
and U1522 (N_1522,N_1491,N_1420);
nand U1523 (N_1523,N_1364,N_1394);
nand U1524 (N_1524,N_1455,N_1468);
nand U1525 (N_1525,N_1499,N_1495);
and U1526 (N_1526,N_1359,N_1487);
or U1527 (N_1527,N_1367,N_1454);
or U1528 (N_1528,N_1475,N_1461);
and U1529 (N_1529,N_1368,N_1444);
xor U1530 (N_1530,N_1350,N_1382);
nor U1531 (N_1531,N_1498,N_1378);
xnor U1532 (N_1532,N_1442,N_1371);
nand U1533 (N_1533,N_1441,N_1479);
or U1534 (N_1534,N_1425,N_1427);
nand U1535 (N_1535,N_1386,N_1357);
or U1536 (N_1536,N_1438,N_1423);
nand U1537 (N_1537,N_1354,N_1466);
nor U1538 (N_1538,N_1407,N_1390);
xor U1539 (N_1539,N_1414,N_1462);
and U1540 (N_1540,N_1381,N_1401);
and U1541 (N_1541,N_1474,N_1489);
and U1542 (N_1542,N_1396,N_1497);
nor U1543 (N_1543,N_1494,N_1472);
and U1544 (N_1544,N_1403,N_1434);
and U1545 (N_1545,N_1467,N_1365);
or U1546 (N_1546,N_1352,N_1412);
xor U1547 (N_1547,N_1385,N_1470);
and U1548 (N_1548,N_1486,N_1429);
or U1549 (N_1549,N_1476,N_1399);
xor U1550 (N_1550,N_1374,N_1362);
nand U1551 (N_1551,N_1351,N_1400);
or U1552 (N_1552,N_1358,N_1355);
and U1553 (N_1553,N_1426,N_1437);
or U1554 (N_1554,N_1493,N_1421);
xnor U1555 (N_1555,N_1496,N_1463);
xor U1556 (N_1556,N_1456,N_1395);
xor U1557 (N_1557,N_1410,N_1488);
nand U1558 (N_1558,N_1353,N_1473);
and U1559 (N_1559,N_1440,N_1415);
nor U1560 (N_1560,N_1478,N_1422);
nand U1561 (N_1561,N_1375,N_1379);
and U1562 (N_1562,N_1383,N_1430);
xor U1563 (N_1563,N_1372,N_1377);
xnor U1564 (N_1564,N_1402,N_1387);
nand U1565 (N_1565,N_1369,N_1408);
and U1566 (N_1566,N_1361,N_1460);
nor U1567 (N_1567,N_1398,N_1445);
xnor U1568 (N_1568,N_1435,N_1465);
and U1569 (N_1569,N_1436,N_1453);
nor U1570 (N_1570,N_1448,N_1360);
and U1571 (N_1571,N_1477,N_1471);
nand U1572 (N_1572,N_1431,N_1409);
nor U1573 (N_1573,N_1469,N_1370);
nor U1574 (N_1574,N_1363,N_1490);
nand U1575 (N_1575,N_1365,N_1421);
or U1576 (N_1576,N_1478,N_1449);
or U1577 (N_1577,N_1413,N_1494);
nand U1578 (N_1578,N_1434,N_1364);
nor U1579 (N_1579,N_1399,N_1416);
or U1580 (N_1580,N_1463,N_1379);
xnor U1581 (N_1581,N_1489,N_1465);
nand U1582 (N_1582,N_1456,N_1359);
and U1583 (N_1583,N_1373,N_1361);
nand U1584 (N_1584,N_1378,N_1463);
or U1585 (N_1585,N_1401,N_1498);
nor U1586 (N_1586,N_1422,N_1450);
or U1587 (N_1587,N_1386,N_1405);
and U1588 (N_1588,N_1490,N_1384);
xnor U1589 (N_1589,N_1496,N_1410);
and U1590 (N_1590,N_1352,N_1360);
or U1591 (N_1591,N_1400,N_1401);
and U1592 (N_1592,N_1424,N_1397);
nor U1593 (N_1593,N_1393,N_1494);
xnor U1594 (N_1594,N_1407,N_1455);
xnor U1595 (N_1595,N_1451,N_1472);
and U1596 (N_1596,N_1498,N_1437);
xor U1597 (N_1597,N_1366,N_1375);
nand U1598 (N_1598,N_1369,N_1383);
nand U1599 (N_1599,N_1441,N_1386);
xnor U1600 (N_1600,N_1403,N_1452);
and U1601 (N_1601,N_1429,N_1373);
and U1602 (N_1602,N_1470,N_1446);
or U1603 (N_1603,N_1416,N_1468);
xnor U1604 (N_1604,N_1482,N_1446);
nor U1605 (N_1605,N_1461,N_1423);
nor U1606 (N_1606,N_1479,N_1389);
nand U1607 (N_1607,N_1404,N_1351);
xnor U1608 (N_1608,N_1393,N_1449);
xor U1609 (N_1609,N_1456,N_1459);
nor U1610 (N_1610,N_1385,N_1414);
xor U1611 (N_1611,N_1380,N_1385);
nand U1612 (N_1612,N_1414,N_1435);
or U1613 (N_1613,N_1406,N_1487);
or U1614 (N_1614,N_1422,N_1429);
nand U1615 (N_1615,N_1478,N_1440);
xnor U1616 (N_1616,N_1425,N_1473);
or U1617 (N_1617,N_1355,N_1403);
nand U1618 (N_1618,N_1368,N_1448);
nand U1619 (N_1619,N_1494,N_1362);
and U1620 (N_1620,N_1392,N_1378);
or U1621 (N_1621,N_1489,N_1393);
and U1622 (N_1622,N_1383,N_1363);
and U1623 (N_1623,N_1367,N_1364);
and U1624 (N_1624,N_1493,N_1471);
or U1625 (N_1625,N_1416,N_1365);
or U1626 (N_1626,N_1480,N_1463);
nor U1627 (N_1627,N_1374,N_1375);
or U1628 (N_1628,N_1492,N_1429);
nand U1629 (N_1629,N_1392,N_1482);
and U1630 (N_1630,N_1445,N_1433);
nor U1631 (N_1631,N_1394,N_1444);
or U1632 (N_1632,N_1382,N_1380);
nor U1633 (N_1633,N_1483,N_1429);
nand U1634 (N_1634,N_1460,N_1355);
nor U1635 (N_1635,N_1470,N_1464);
or U1636 (N_1636,N_1452,N_1453);
xnor U1637 (N_1637,N_1493,N_1384);
or U1638 (N_1638,N_1440,N_1438);
nand U1639 (N_1639,N_1482,N_1413);
or U1640 (N_1640,N_1490,N_1394);
nor U1641 (N_1641,N_1478,N_1400);
nand U1642 (N_1642,N_1410,N_1424);
xor U1643 (N_1643,N_1370,N_1395);
xor U1644 (N_1644,N_1384,N_1425);
nand U1645 (N_1645,N_1417,N_1431);
nand U1646 (N_1646,N_1499,N_1413);
or U1647 (N_1647,N_1428,N_1492);
and U1648 (N_1648,N_1353,N_1450);
nand U1649 (N_1649,N_1388,N_1409);
xnor U1650 (N_1650,N_1517,N_1548);
or U1651 (N_1651,N_1506,N_1509);
nor U1652 (N_1652,N_1527,N_1616);
and U1653 (N_1653,N_1559,N_1594);
or U1654 (N_1654,N_1565,N_1515);
and U1655 (N_1655,N_1572,N_1573);
nand U1656 (N_1656,N_1525,N_1557);
or U1657 (N_1657,N_1523,N_1599);
xor U1658 (N_1658,N_1537,N_1569);
nor U1659 (N_1659,N_1578,N_1546);
xnor U1660 (N_1660,N_1508,N_1647);
nand U1661 (N_1661,N_1612,N_1634);
and U1662 (N_1662,N_1518,N_1591);
xor U1663 (N_1663,N_1640,N_1528);
or U1664 (N_1664,N_1629,N_1630);
nand U1665 (N_1665,N_1638,N_1598);
nand U1666 (N_1666,N_1574,N_1635);
or U1667 (N_1667,N_1522,N_1532);
or U1668 (N_1668,N_1560,N_1583);
xnor U1669 (N_1669,N_1540,N_1639);
xor U1670 (N_1670,N_1547,N_1534);
xnor U1671 (N_1671,N_1637,N_1632);
or U1672 (N_1672,N_1614,N_1607);
nor U1673 (N_1673,N_1646,N_1502);
nand U1674 (N_1674,N_1580,N_1538);
or U1675 (N_1675,N_1551,N_1643);
or U1676 (N_1676,N_1597,N_1601);
and U1677 (N_1677,N_1567,N_1593);
xnor U1678 (N_1678,N_1558,N_1563);
and U1679 (N_1679,N_1625,N_1617);
or U1680 (N_1680,N_1613,N_1587);
xnor U1681 (N_1681,N_1645,N_1550);
and U1682 (N_1682,N_1556,N_1623);
and U1683 (N_1683,N_1626,N_1619);
nor U1684 (N_1684,N_1592,N_1648);
or U1685 (N_1685,N_1514,N_1504);
nand U1686 (N_1686,N_1622,N_1604);
xnor U1687 (N_1687,N_1606,N_1568);
and U1688 (N_1688,N_1602,N_1519);
and U1689 (N_1689,N_1570,N_1552);
nand U1690 (N_1690,N_1561,N_1649);
xor U1691 (N_1691,N_1596,N_1600);
and U1692 (N_1692,N_1524,N_1544);
or U1693 (N_1693,N_1500,N_1533);
nand U1694 (N_1694,N_1536,N_1605);
nor U1695 (N_1695,N_1571,N_1610);
nor U1696 (N_1696,N_1516,N_1586);
or U1697 (N_1697,N_1590,N_1521);
xnor U1698 (N_1698,N_1642,N_1588);
nor U1699 (N_1699,N_1581,N_1627);
nor U1700 (N_1700,N_1503,N_1566);
xnor U1701 (N_1701,N_1631,N_1620);
or U1702 (N_1702,N_1628,N_1535);
xnor U1703 (N_1703,N_1609,N_1618);
nor U1704 (N_1704,N_1577,N_1520);
nor U1705 (N_1705,N_1553,N_1529);
and U1706 (N_1706,N_1530,N_1621);
nand U1707 (N_1707,N_1531,N_1511);
xor U1708 (N_1708,N_1526,N_1513);
or U1709 (N_1709,N_1608,N_1545);
nand U1710 (N_1710,N_1512,N_1641);
or U1711 (N_1711,N_1541,N_1555);
or U1712 (N_1712,N_1501,N_1505);
nand U1713 (N_1713,N_1615,N_1554);
nor U1714 (N_1714,N_1589,N_1585);
or U1715 (N_1715,N_1507,N_1542);
or U1716 (N_1716,N_1562,N_1584);
xnor U1717 (N_1717,N_1575,N_1576);
and U1718 (N_1718,N_1595,N_1644);
nand U1719 (N_1719,N_1582,N_1603);
or U1720 (N_1720,N_1579,N_1633);
nor U1721 (N_1721,N_1549,N_1624);
xnor U1722 (N_1722,N_1564,N_1543);
nor U1723 (N_1723,N_1539,N_1636);
and U1724 (N_1724,N_1611,N_1510);
xor U1725 (N_1725,N_1628,N_1641);
nand U1726 (N_1726,N_1636,N_1627);
and U1727 (N_1727,N_1519,N_1522);
and U1728 (N_1728,N_1646,N_1579);
xor U1729 (N_1729,N_1609,N_1649);
or U1730 (N_1730,N_1618,N_1508);
xnor U1731 (N_1731,N_1625,N_1586);
and U1732 (N_1732,N_1526,N_1560);
nor U1733 (N_1733,N_1542,N_1617);
nand U1734 (N_1734,N_1646,N_1608);
xor U1735 (N_1735,N_1591,N_1536);
nor U1736 (N_1736,N_1617,N_1631);
or U1737 (N_1737,N_1549,N_1544);
nand U1738 (N_1738,N_1544,N_1608);
nor U1739 (N_1739,N_1626,N_1540);
nand U1740 (N_1740,N_1569,N_1573);
or U1741 (N_1741,N_1533,N_1576);
and U1742 (N_1742,N_1541,N_1517);
and U1743 (N_1743,N_1598,N_1600);
xnor U1744 (N_1744,N_1560,N_1637);
nor U1745 (N_1745,N_1643,N_1629);
nand U1746 (N_1746,N_1536,N_1609);
or U1747 (N_1747,N_1578,N_1551);
and U1748 (N_1748,N_1643,N_1612);
or U1749 (N_1749,N_1518,N_1526);
nor U1750 (N_1750,N_1606,N_1648);
or U1751 (N_1751,N_1530,N_1533);
nand U1752 (N_1752,N_1642,N_1567);
or U1753 (N_1753,N_1503,N_1536);
or U1754 (N_1754,N_1574,N_1616);
nor U1755 (N_1755,N_1520,N_1611);
and U1756 (N_1756,N_1627,N_1542);
or U1757 (N_1757,N_1586,N_1538);
xor U1758 (N_1758,N_1566,N_1501);
xnor U1759 (N_1759,N_1578,N_1575);
nor U1760 (N_1760,N_1608,N_1629);
or U1761 (N_1761,N_1645,N_1580);
nor U1762 (N_1762,N_1636,N_1588);
and U1763 (N_1763,N_1504,N_1564);
and U1764 (N_1764,N_1509,N_1603);
or U1765 (N_1765,N_1606,N_1640);
or U1766 (N_1766,N_1626,N_1530);
xor U1767 (N_1767,N_1639,N_1507);
xor U1768 (N_1768,N_1590,N_1620);
and U1769 (N_1769,N_1625,N_1611);
nand U1770 (N_1770,N_1604,N_1568);
xor U1771 (N_1771,N_1598,N_1590);
xor U1772 (N_1772,N_1573,N_1642);
and U1773 (N_1773,N_1518,N_1587);
and U1774 (N_1774,N_1576,N_1583);
nor U1775 (N_1775,N_1637,N_1528);
nor U1776 (N_1776,N_1616,N_1551);
nor U1777 (N_1777,N_1622,N_1526);
xor U1778 (N_1778,N_1639,N_1601);
nand U1779 (N_1779,N_1621,N_1628);
or U1780 (N_1780,N_1617,N_1564);
nor U1781 (N_1781,N_1627,N_1532);
nand U1782 (N_1782,N_1623,N_1621);
or U1783 (N_1783,N_1628,N_1514);
xnor U1784 (N_1784,N_1546,N_1552);
nor U1785 (N_1785,N_1631,N_1530);
and U1786 (N_1786,N_1560,N_1589);
or U1787 (N_1787,N_1609,N_1563);
and U1788 (N_1788,N_1648,N_1523);
or U1789 (N_1789,N_1575,N_1595);
xor U1790 (N_1790,N_1646,N_1525);
and U1791 (N_1791,N_1623,N_1649);
or U1792 (N_1792,N_1566,N_1632);
nor U1793 (N_1793,N_1536,N_1514);
nand U1794 (N_1794,N_1642,N_1545);
nor U1795 (N_1795,N_1551,N_1612);
nand U1796 (N_1796,N_1565,N_1638);
nand U1797 (N_1797,N_1557,N_1628);
or U1798 (N_1798,N_1587,N_1619);
or U1799 (N_1799,N_1584,N_1539);
or U1800 (N_1800,N_1672,N_1713);
nand U1801 (N_1801,N_1667,N_1693);
nand U1802 (N_1802,N_1790,N_1763);
nand U1803 (N_1803,N_1728,N_1707);
nor U1804 (N_1804,N_1660,N_1676);
nand U1805 (N_1805,N_1739,N_1761);
or U1806 (N_1806,N_1762,N_1651);
nor U1807 (N_1807,N_1653,N_1675);
nor U1808 (N_1808,N_1787,N_1782);
or U1809 (N_1809,N_1753,N_1659);
and U1810 (N_1810,N_1781,N_1696);
and U1811 (N_1811,N_1795,N_1785);
and U1812 (N_1812,N_1686,N_1710);
or U1813 (N_1813,N_1694,N_1722);
xnor U1814 (N_1814,N_1732,N_1727);
nand U1815 (N_1815,N_1768,N_1681);
nor U1816 (N_1816,N_1770,N_1765);
nor U1817 (N_1817,N_1772,N_1759);
xor U1818 (N_1818,N_1690,N_1745);
xor U1819 (N_1819,N_1708,N_1695);
xor U1820 (N_1820,N_1744,N_1726);
or U1821 (N_1821,N_1683,N_1718);
nor U1822 (N_1822,N_1792,N_1774);
and U1823 (N_1823,N_1699,N_1716);
nor U1824 (N_1824,N_1704,N_1777);
and U1825 (N_1825,N_1691,N_1778);
xnor U1826 (N_1826,N_1715,N_1711);
xor U1827 (N_1827,N_1784,N_1666);
nand U1828 (N_1828,N_1735,N_1798);
and U1829 (N_1829,N_1791,N_1658);
and U1830 (N_1830,N_1796,N_1689);
and U1831 (N_1831,N_1794,N_1754);
and U1832 (N_1832,N_1799,N_1712);
or U1833 (N_1833,N_1685,N_1786);
nand U1834 (N_1834,N_1684,N_1797);
and U1835 (N_1835,N_1741,N_1769);
and U1836 (N_1836,N_1734,N_1788);
and U1837 (N_1837,N_1717,N_1655);
or U1838 (N_1838,N_1780,N_1767);
nor U1839 (N_1839,N_1650,N_1652);
and U1840 (N_1840,N_1775,N_1680);
and U1841 (N_1841,N_1789,N_1698);
nor U1842 (N_1842,N_1730,N_1665);
nor U1843 (N_1843,N_1793,N_1682);
xor U1844 (N_1844,N_1721,N_1679);
xnor U1845 (N_1845,N_1674,N_1776);
nand U1846 (N_1846,N_1755,N_1709);
and U1847 (N_1847,N_1697,N_1705);
nor U1848 (N_1848,N_1742,N_1756);
nor U1849 (N_1849,N_1692,N_1714);
xor U1850 (N_1850,N_1751,N_1729);
xor U1851 (N_1851,N_1688,N_1773);
nor U1852 (N_1852,N_1720,N_1673);
nand U1853 (N_1853,N_1764,N_1724);
nor U1854 (N_1854,N_1731,N_1736);
nand U1855 (N_1855,N_1737,N_1725);
nor U1856 (N_1856,N_1757,N_1671);
and U1857 (N_1857,N_1719,N_1752);
nor U1858 (N_1858,N_1743,N_1746);
or U1859 (N_1859,N_1738,N_1703);
xor U1860 (N_1860,N_1771,N_1701);
nand U1861 (N_1861,N_1654,N_1723);
or U1862 (N_1862,N_1748,N_1779);
nand U1863 (N_1863,N_1670,N_1760);
nand U1864 (N_1864,N_1783,N_1687);
nand U1865 (N_1865,N_1664,N_1669);
and U1866 (N_1866,N_1657,N_1678);
and U1867 (N_1867,N_1668,N_1740);
or U1868 (N_1868,N_1747,N_1750);
xnor U1869 (N_1869,N_1702,N_1700);
and U1870 (N_1870,N_1758,N_1733);
nand U1871 (N_1871,N_1662,N_1677);
and U1872 (N_1872,N_1656,N_1661);
xor U1873 (N_1873,N_1706,N_1749);
xnor U1874 (N_1874,N_1663,N_1766);
nor U1875 (N_1875,N_1775,N_1671);
nand U1876 (N_1876,N_1765,N_1798);
or U1877 (N_1877,N_1656,N_1781);
nor U1878 (N_1878,N_1767,N_1758);
nor U1879 (N_1879,N_1768,N_1663);
and U1880 (N_1880,N_1651,N_1685);
nand U1881 (N_1881,N_1785,N_1764);
xnor U1882 (N_1882,N_1686,N_1760);
or U1883 (N_1883,N_1781,N_1743);
nor U1884 (N_1884,N_1698,N_1776);
xor U1885 (N_1885,N_1745,N_1692);
xnor U1886 (N_1886,N_1789,N_1794);
or U1887 (N_1887,N_1691,N_1756);
nand U1888 (N_1888,N_1650,N_1679);
xnor U1889 (N_1889,N_1711,N_1728);
or U1890 (N_1890,N_1789,N_1748);
nor U1891 (N_1891,N_1760,N_1693);
and U1892 (N_1892,N_1718,N_1661);
nand U1893 (N_1893,N_1680,N_1737);
xor U1894 (N_1894,N_1732,N_1748);
nand U1895 (N_1895,N_1717,N_1657);
and U1896 (N_1896,N_1786,N_1711);
nand U1897 (N_1897,N_1735,N_1701);
and U1898 (N_1898,N_1797,N_1679);
nand U1899 (N_1899,N_1719,N_1700);
nor U1900 (N_1900,N_1780,N_1725);
and U1901 (N_1901,N_1717,N_1791);
and U1902 (N_1902,N_1789,N_1715);
nand U1903 (N_1903,N_1667,N_1714);
or U1904 (N_1904,N_1780,N_1749);
nor U1905 (N_1905,N_1682,N_1757);
xnor U1906 (N_1906,N_1788,N_1730);
nand U1907 (N_1907,N_1671,N_1724);
nor U1908 (N_1908,N_1798,N_1715);
nor U1909 (N_1909,N_1710,N_1714);
nand U1910 (N_1910,N_1745,N_1696);
nand U1911 (N_1911,N_1729,N_1695);
nand U1912 (N_1912,N_1664,N_1749);
or U1913 (N_1913,N_1694,N_1758);
xor U1914 (N_1914,N_1775,N_1686);
nand U1915 (N_1915,N_1665,N_1798);
xor U1916 (N_1916,N_1755,N_1748);
nand U1917 (N_1917,N_1676,N_1656);
xnor U1918 (N_1918,N_1792,N_1682);
nor U1919 (N_1919,N_1774,N_1798);
xnor U1920 (N_1920,N_1721,N_1723);
nor U1921 (N_1921,N_1661,N_1680);
or U1922 (N_1922,N_1766,N_1682);
nor U1923 (N_1923,N_1747,N_1739);
or U1924 (N_1924,N_1710,N_1755);
or U1925 (N_1925,N_1708,N_1739);
and U1926 (N_1926,N_1772,N_1698);
or U1927 (N_1927,N_1703,N_1777);
and U1928 (N_1928,N_1697,N_1790);
xnor U1929 (N_1929,N_1766,N_1684);
and U1930 (N_1930,N_1773,N_1690);
nand U1931 (N_1931,N_1774,N_1731);
nand U1932 (N_1932,N_1753,N_1682);
or U1933 (N_1933,N_1724,N_1767);
xor U1934 (N_1934,N_1701,N_1769);
and U1935 (N_1935,N_1798,N_1771);
nand U1936 (N_1936,N_1686,N_1770);
nand U1937 (N_1937,N_1699,N_1779);
nor U1938 (N_1938,N_1708,N_1671);
nand U1939 (N_1939,N_1732,N_1792);
nand U1940 (N_1940,N_1754,N_1750);
and U1941 (N_1941,N_1700,N_1731);
nor U1942 (N_1942,N_1788,N_1781);
and U1943 (N_1943,N_1798,N_1752);
and U1944 (N_1944,N_1704,N_1686);
nand U1945 (N_1945,N_1670,N_1767);
nand U1946 (N_1946,N_1774,N_1777);
nor U1947 (N_1947,N_1659,N_1672);
or U1948 (N_1948,N_1664,N_1733);
and U1949 (N_1949,N_1655,N_1788);
and U1950 (N_1950,N_1811,N_1902);
or U1951 (N_1951,N_1846,N_1942);
nor U1952 (N_1952,N_1801,N_1920);
nand U1953 (N_1953,N_1913,N_1893);
nor U1954 (N_1954,N_1848,N_1935);
xor U1955 (N_1955,N_1886,N_1939);
nand U1956 (N_1956,N_1812,N_1926);
xor U1957 (N_1957,N_1824,N_1905);
and U1958 (N_1958,N_1835,N_1908);
nor U1959 (N_1959,N_1898,N_1851);
nand U1960 (N_1960,N_1829,N_1862);
nor U1961 (N_1961,N_1933,N_1805);
or U1962 (N_1962,N_1889,N_1849);
nor U1963 (N_1963,N_1807,N_1897);
nand U1964 (N_1964,N_1844,N_1883);
nor U1965 (N_1965,N_1860,N_1870);
nor U1966 (N_1966,N_1850,N_1946);
and U1967 (N_1967,N_1852,N_1922);
and U1968 (N_1968,N_1923,N_1872);
or U1969 (N_1969,N_1815,N_1899);
or U1970 (N_1970,N_1839,N_1864);
nand U1971 (N_1971,N_1854,N_1841);
nor U1972 (N_1972,N_1857,N_1924);
nor U1973 (N_1973,N_1855,N_1919);
nand U1974 (N_1974,N_1943,N_1853);
and U1975 (N_1975,N_1840,N_1867);
nor U1976 (N_1976,N_1891,N_1803);
and U1977 (N_1977,N_1944,N_1894);
xnor U1978 (N_1978,N_1847,N_1881);
xor U1979 (N_1979,N_1821,N_1907);
and U1980 (N_1980,N_1877,N_1861);
and U1981 (N_1981,N_1910,N_1875);
xnor U1982 (N_1982,N_1866,N_1836);
or U1983 (N_1983,N_1818,N_1887);
and U1984 (N_1984,N_1930,N_1914);
or U1985 (N_1985,N_1921,N_1822);
or U1986 (N_1986,N_1834,N_1865);
and U1987 (N_1987,N_1929,N_1804);
nor U1988 (N_1988,N_1816,N_1931);
or U1989 (N_1989,N_1869,N_1941);
and U1990 (N_1990,N_1813,N_1884);
nand U1991 (N_1991,N_1856,N_1927);
or U1992 (N_1992,N_1917,N_1817);
and U1993 (N_1993,N_1863,N_1885);
or U1994 (N_1994,N_1871,N_1932);
nor U1995 (N_1995,N_1947,N_1940);
nor U1996 (N_1996,N_1810,N_1858);
nand U1997 (N_1997,N_1895,N_1823);
nand U1998 (N_1998,N_1879,N_1901);
xnor U1999 (N_1999,N_1916,N_1842);
or U2000 (N_2000,N_1903,N_1828);
xnor U2001 (N_2001,N_1938,N_1843);
and U2002 (N_2002,N_1892,N_1802);
or U2003 (N_2003,N_1880,N_1809);
and U2004 (N_2004,N_1826,N_1833);
and U2005 (N_2005,N_1906,N_1874);
xnor U2006 (N_2006,N_1945,N_1825);
and U2007 (N_2007,N_1928,N_1937);
nand U2008 (N_2008,N_1873,N_1949);
nand U2009 (N_2009,N_1936,N_1918);
and U2010 (N_2010,N_1800,N_1900);
nor U2011 (N_2011,N_1878,N_1831);
or U2012 (N_2012,N_1808,N_1832);
nand U2013 (N_2013,N_1909,N_1888);
nor U2014 (N_2014,N_1837,N_1934);
or U2015 (N_2015,N_1876,N_1827);
and U2016 (N_2016,N_1915,N_1820);
nand U2017 (N_2017,N_1845,N_1838);
nor U2018 (N_2018,N_1890,N_1814);
xor U2019 (N_2019,N_1882,N_1868);
xnor U2020 (N_2020,N_1904,N_1911);
or U2021 (N_2021,N_1925,N_1896);
nand U2022 (N_2022,N_1806,N_1948);
and U2023 (N_2023,N_1859,N_1830);
nor U2024 (N_2024,N_1819,N_1912);
nand U2025 (N_2025,N_1865,N_1843);
xnor U2026 (N_2026,N_1861,N_1931);
nand U2027 (N_2027,N_1949,N_1929);
and U2028 (N_2028,N_1923,N_1870);
nand U2029 (N_2029,N_1874,N_1869);
xor U2030 (N_2030,N_1913,N_1906);
and U2031 (N_2031,N_1851,N_1874);
nor U2032 (N_2032,N_1857,N_1852);
or U2033 (N_2033,N_1864,N_1859);
nand U2034 (N_2034,N_1906,N_1853);
xnor U2035 (N_2035,N_1826,N_1924);
and U2036 (N_2036,N_1868,N_1828);
and U2037 (N_2037,N_1938,N_1854);
xor U2038 (N_2038,N_1871,N_1909);
or U2039 (N_2039,N_1820,N_1872);
and U2040 (N_2040,N_1811,N_1861);
and U2041 (N_2041,N_1889,N_1824);
and U2042 (N_2042,N_1925,N_1814);
or U2043 (N_2043,N_1925,N_1902);
nand U2044 (N_2044,N_1882,N_1812);
nor U2045 (N_2045,N_1913,N_1810);
and U2046 (N_2046,N_1868,N_1887);
nand U2047 (N_2047,N_1875,N_1812);
or U2048 (N_2048,N_1899,N_1821);
or U2049 (N_2049,N_1937,N_1827);
nor U2050 (N_2050,N_1809,N_1803);
nor U2051 (N_2051,N_1939,N_1893);
and U2052 (N_2052,N_1935,N_1870);
nor U2053 (N_2053,N_1935,N_1905);
or U2054 (N_2054,N_1812,N_1939);
nand U2055 (N_2055,N_1846,N_1892);
nor U2056 (N_2056,N_1870,N_1861);
and U2057 (N_2057,N_1873,N_1924);
xnor U2058 (N_2058,N_1903,N_1869);
nand U2059 (N_2059,N_1817,N_1832);
nand U2060 (N_2060,N_1833,N_1923);
nand U2061 (N_2061,N_1909,N_1918);
or U2062 (N_2062,N_1846,N_1902);
nor U2063 (N_2063,N_1858,N_1818);
nor U2064 (N_2064,N_1865,N_1912);
and U2065 (N_2065,N_1802,N_1933);
xnor U2066 (N_2066,N_1897,N_1867);
and U2067 (N_2067,N_1806,N_1839);
or U2068 (N_2068,N_1932,N_1938);
nand U2069 (N_2069,N_1902,N_1871);
nand U2070 (N_2070,N_1872,N_1916);
nor U2071 (N_2071,N_1946,N_1904);
nand U2072 (N_2072,N_1883,N_1894);
nor U2073 (N_2073,N_1907,N_1866);
and U2074 (N_2074,N_1860,N_1833);
nand U2075 (N_2075,N_1832,N_1861);
nand U2076 (N_2076,N_1806,N_1877);
nand U2077 (N_2077,N_1917,N_1882);
or U2078 (N_2078,N_1896,N_1924);
and U2079 (N_2079,N_1860,N_1859);
nor U2080 (N_2080,N_1921,N_1899);
and U2081 (N_2081,N_1907,N_1900);
xor U2082 (N_2082,N_1926,N_1903);
or U2083 (N_2083,N_1937,N_1945);
and U2084 (N_2084,N_1815,N_1800);
and U2085 (N_2085,N_1868,N_1929);
xnor U2086 (N_2086,N_1858,N_1853);
nand U2087 (N_2087,N_1894,N_1849);
nor U2088 (N_2088,N_1857,N_1927);
or U2089 (N_2089,N_1928,N_1832);
and U2090 (N_2090,N_1800,N_1832);
or U2091 (N_2091,N_1911,N_1888);
nand U2092 (N_2092,N_1838,N_1843);
or U2093 (N_2093,N_1885,N_1819);
xor U2094 (N_2094,N_1868,N_1856);
and U2095 (N_2095,N_1901,N_1856);
or U2096 (N_2096,N_1807,N_1927);
and U2097 (N_2097,N_1850,N_1903);
nor U2098 (N_2098,N_1860,N_1836);
nand U2099 (N_2099,N_1878,N_1874);
xnor U2100 (N_2100,N_2018,N_2032);
or U2101 (N_2101,N_2033,N_1989);
nor U2102 (N_2102,N_1962,N_2093);
nand U2103 (N_2103,N_2061,N_1994);
nand U2104 (N_2104,N_2057,N_2034);
nor U2105 (N_2105,N_2002,N_1976);
xor U2106 (N_2106,N_1964,N_1971);
xnor U2107 (N_2107,N_1984,N_2029);
and U2108 (N_2108,N_2081,N_2026);
nor U2109 (N_2109,N_2038,N_2072);
nor U2110 (N_2110,N_2082,N_1967);
nand U2111 (N_2111,N_2054,N_2006);
nor U2112 (N_2112,N_2078,N_1997);
or U2113 (N_2113,N_2011,N_2022);
nand U2114 (N_2114,N_2080,N_2027);
xor U2115 (N_2115,N_2064,N_2065);
nor U2116 (N_2116,N_1980,N_1968);
nand U2117 (N_2117,N_2096,N_2053);
xnor U2118 (N_2118,N_1970,N_2076);
nor U2119 (N_2119,N_2025,N_1950);
or U2120 (N_2120,N_2049,N_2028);
xnor U2121 (N_2121,N_2015,N_1969);
nand U2122 (N_2122,N_2036,N_2097);
xor U2123 (N_2123,N_1952,N_1983);
and U2124 (N_2124,N_1963,N_2021);
or U2125 (N_2125,N_2045,N_2004);
xnor U2126 (N_2126,N_2003,N_1973);
and U2127 (N_2127,N_2030,N_2086);
nand U2128 (N_2128,N_2084,N_1960);
and U2129 (N_2129,N_1986,N_1956);
nand U2130 (N_2130,N_2019,N_2068);
nor U2131 (N_2131,N_2014,N_1978);
xnor U2132 (N_2132,N_2007,N_1985);
and U2133 (N_2133,N_1954,N_2090);
or U2134 (N_2134,N_1992,N_2066);
xor U2135 (N_2135,N_2056,N_2005);
or U2136 (N_2136,N_2012,N_2047);
and U2137 (N_2137,N_2071,N_1995);
and U2138 (N_2138,N_2016,N_2060);
nor U2139 (N_2139,N_1981,N_2051);
nand U2140 (N_2140,N_1998,N_2039);
nand U2141 (N_2141,N_1993,N_2094);
nor U2142 (N_2142,N_1953,N_1987);
and U2143 (N_2143,N_2091,N_2062);
or U2144 (N_2144,N_1955,N_1972);
xnor U2145 (N_2145,N_2043,N_1961);
xnor U2146 (N_2146,N_1974,N_2040);
or U2147 (N_2147,N_2079,N_2024);
and U2148 (N_2148,N_2095,N_2046);
and U2149 (N_2149,N_2052,N_2050);
or U2150 (N_2150,N_2031,N_2069);
or U2151 (N_2151,N_1965,N_2075);
xnor U2152 (N_2152,N_1951,N_2009);
nor U2153 (N_2153,N_1982,N_2067);
xor U2154 (N_2154,N_2058,N_2099);
and U2155 (N_2155,N_2098,N_2037);
or U2156 (N_2156,N_2088,N_2010);
or U2157 (N_2157,N_2041,N_2042);
nand U2158 (N_2158,N_1991,N_1999);
and U2159 (N_2159,N_1979,N_2087);
nand U2160 (N_2160,N_1977,N_2000);
and U2161 (N_2161,N_2063,N_2092);
nor U2162 (N_2162,N_2008,N_1975);
and U2163 (N_2163,N_2074,N_2023);
or U2164 (N_2164,N_1966,N_2073);
or U2165 (N_2165,N_2077,N_1988);
nand U2166 (N_2166,N_2089,N_1990);
nand U2167 (N_2167,N_2035,N_2001);
or U2168 (N_2168,N_2083,N_1959);
and U2169 (N_2169,N_2020,N_2013);
nand U2170 (N_2170,N_2044,N_2017);
nand U2171 (N_2171,N_2048,N_1996);
nor U2172 (N_2172,N_1958,N_1957);
nor U2173 (N_2173,N_2055,N_2070);
or U2174 (N_2174,N_2085,N_2059);
nor U2175 (N_2175,N_2060,N_2059);
or U2176 (N_2176,N_2074,N_2046);
nor U2177 (N_2177,N_2068,N_2009);
and U2178 (N_2178,N_2002,N_2015);
nand U2179 (N_2179,N_2005,N_2087);
and U2180 (N_2180,N_2006,N_2055);
nand U2181 (N_2181,N_2038,N_1975);
and U2182 (N_2182,N_2047,N_2089);
or U2183 (N_2183,N_2021,N_1950);
and U2184 (N_2184,N_1965,N_1960);
or U2185 (N_2185,N_2026,N_2001);
xnor U2186 (N_2186,N_2000,N_1980);
nor U2187 (N_2187,N_1963,N_2042);
xnor U2188 (N_2188,N_2062,N_1966);
and U2189 (N_2189,N_2093,N_2011);
nor U2190 (N_2190,N_1963,N_2020);
nand U2191 (N_2191,N_2077,N_1993);
or U2192 (N_2192,N_2021,N_2087);
nor U2193 (N_2193,N_2057,N_1973);
nand U2194 (N_2194,N_2041,N_2027);
nor U2195 (N_2195,N_2086,N_1987);
nor U2196 (N_2196,N_1986,N_2031);
xor U2197 (N_2197,N_2024,N_2096);
nand U2198 (N_2198,N_1980,N_2040);
nand U2199 (N_2199,N_1986,N_2062);
or U2200 (N_2200,N_1950,N_1983);
nor U2201 (N_2201,N_1959,N_2010);
xor U2202 (N_2202,N_2087,N_2069);
or U2203 (N_2203,N_1986,N_2077);
nand U2204 (N_2204,N_2039,N_2061);
or U2205 (N_2205,N_2042,N_1989);
and U2206 (N_2206,N_1968,N_2024);
nor U2207 (N_2207,N_2088,N_2084);
or U2208 (N_2208,N_2029,N_2023);
nor U2209 (N_2209,N_2075,N_2094);
and U2210 (N_2210,N_2082,N_2051);
or U2211 (N_2211,N_2051,N_2031);
nor U2212 (N_2212,N_2052,N_2013);
or U2213 (N_2213,N_1955,N_2017);
and U2214 (N_2214,N_2099,N_2003);
nor U2215 (N_2215,N_1973,N_2048);
xnor U2216 (N_2216,N_2066,N_1950);
and U2217 (N_2217,N_1970,N_2073);
nor U2218 (N_2218,N_2035,N_1953);
and U2219 (N_2219,N_1961,N_2000);
nor U2220 (N_2220,N_2079,N_1990);
nand U2221 (N_2221,N_2046,N_2048);
nand U2222 (N_2222,N_2068,N_2034);
xnor U2223 (N_2223,N_2098,N_2096);
xor U2224 (N_2224,N_2039,N_1989);
nor U2225 (N_2225,N_2091,N_1979);
nand U2226 (N_2226,N_1951,N_1979);
xnor U2227 (N_2227,N_1990,N_2019);
xnor U2228 (N_2228,N_2006,N_2027);
nor U2229 (N_2229,N_2068,N_1968);
and U2230 (N_2230,N_2052,N_1986);
xor U2231 (N_2231,N_2033,N_2047);
and U2232 (N_2232,N_2025,N_1957);
and U2233 (N_2233,N_2043,N_2077);
nor U2234 (N_2234,N_2061,N_1956);
xor U2235 (N_2235,N_2081,N_2009);
and U2236 (N_2236,N_2017,N_2057);
or U2237 (N_2237,N_2010,N_2008);
and U2238 (N_2238,N_2036,N_1954);
or U2239 (N_2239,N_2022,N_2091);
nand U2240 (N_2240,N_1960,N_2096);
or U2241 (N_2241,N_2082,N_2065);
nor U2242 (N_2242,N_2002,N_2044);
nor U2243 (N_2243,N_2039,N_2043);
and U2244 (N_2244,N_2078,N_2026);
and U2245 (N_2245,N_1996,N_2070);
nand U2246 (N_2246,N_1994,N_2096);
nand U2247 (N_2247,N_1957,N_1950);
xor U2248 (N_2248,N_2029,N_1999);
xor U2249 (N_2249,N_2046,N_2004);
and U2250 (N_2250,N_2169,N_2204);
nor U2251 (N_2251,N_2171,N_2207);
xor U2252 (N_2252,N_2190,N_2144);
and U2253 (N_2253,N_2244,N_2226);
nor U2254 (N_2254,N_2248,N_2173);
nand U2255 (N_2255,N_2187,N_2222);
or U2256 (N_2256,N_2161,N_2138);
and U2257 (N_2257,N_2184,N_2140);
nor U2258 (N_2258,N_2163,N_2232);
nor U2259 (N_2259,N_2241,N_2119);
nor U2260 (N_2260,N_2202,N_2164);
and U2261 (N_2261,N_2100,N_2181);
or U2262 (N_2262,N_2194,N_2198);
nand U2263 (N_2263,N_2122,N_2166);
nor U2264 (N_2264,N_2127,N_2154);
nand U2265 (N_2265,N_2175,N_2157);
xnor U2266 (N_2266,N_2113,N_2160);
nand U2267 (N_2267,N_2228,N_2172);
and U2268 (N_2268,N_2239,N_2238);
and U2269 (N_2269,N_2225,N_2180);
nand U2270 (N_2270,N_2199,N_2235);
xor U2271 (N_2271,N_2105,N_2179);
xor U2272 (N_2272,N_2143,N_2106);
xnor U2273 (N_2273,N_2195,N_2185);
nor U2274 (N_2274,N_2242,N_2203);
nor U2275 (N_2275,N_2168,N_2102);
nor U2276 (N_2276,N_2178,N_2126);
or U2277 (N_2277,N_2191,N_2147);
and U2278 (N_2278,N_2223,N_2109);
nor U2279 (N_2279,N_2243,N_2112);
nor U2280 (N_2280,N_2183,N_2189);
or U2281 (N_2281,N_2233,N_2165);
nor U2282 (N_2282,N_2247,N_2141);
nor U2283 (N_2283,N_2249,N_2219);
and U2284 (N_2284,N_2114,N_2123);
xnor U2285 (N_2285,N_2131,N_2116);
nand U2286 (N_2286,N_2214,N_2130);
or U2287 (N_2287,N_2135,N_2156);
xnor U2288 (N_2288,N_2240,N_2150);
xnor U2289 (N_2289,N_2110,N_2149);
and U2290 (N_2290,N_2158,N_2118);
or U2291 (N_2291,N_2176,N_2186);
nand U2292 (N_2292,N_2133,N_2217);
xnor U2293 (N_2293,N_2206,N_2209);
nor U2294 (N_2294,N_2136,N_2237);
nand U2295 (N_2295,N_2128,N_2213);
or U2296 (N_2296,N_2210,N_2231);
nor U2297 (N_2297,N_2196,N_2218);
nor U2298 (N_2298,N_2155,N_2137);
and U2299 (N_2299,N_2236,N_2152);
and U2300 (N_2300,N_2153,N_2142);
and U2301 (N_2301,N_2132,N_2245);
or U2302 (N_2302,N_2201,N_2227);
nor U2303 (N_2303,N_2215,N_2230);
nand U2304 (N_2304,N_2159,N_2221);
or U2305 (N_2305,N_2129,N_2139);
xnor U2306 (N_2306,N_2212,N_2125);
nor U2307 (N_2307,N_2104,N_2182);
xnor U2308 (N_2308,N_2101,N_2220);
nor U2309 (N_2309,N_2134,N_2234);
nor U2310 (N_2310,N_2108,N_2121);
nand U2311 (N_2311,N_2193,N_2145);
nand U2312 (N_2312,N_2208,N_2177);
or U2313 (N_2313,N_2197,N_2174);
nand U2314 (N_2314,N_2216,N_2188);
nand U2315 (N_2315,N_2103,N_2120);
nor U2316 (N_2316,N_2224,N_2162);
nor U2317 (N_2317,N_2115,N_2192);
nand U2318 (N_2318,N_2211,N_2170);
xnor U2319 (N_2319,N_2246,N_2111);
and U2320 (N_2320,N_2205,N_2107);
xor U2321 (N_2321,N_2167,N_2148);
nor U2322 (N_2322,N_2229,N_2117);
xnor U2323 (N_2323,N_2146,N_2200);
nor U2324 (N_2324,N_2124,N_2151);
nor U2325 (N_2325,N_2217,N_2222);
and U2326 (N_2326,N_2148,N_2193);
and U2327 (N_2327,N_2203,N_2181);
and U2328 (N_2328,N_2208,N_2111);
nor U2329 (N_2329,N_2125,N_2164);
or U2330 (N_2330,N_2246,N_2183);
nor U2331 (N_2331,N_2184,N_2125);
nand U2332 (N_2332,N_2173,N_2197);
or U2333 (N_2333,N_2226,N_2155);
or U2334 (N_2334,N_2101,N_2156);
and U2335 (N_2335,N_2224,N_2166);
nand U2336 (N_2336,N_2181,N_2244);
xor U2337 (N_2337,N_2178,N_2140);
or U2338 (N_2338,N_2128,N_2122);
xnor U2339 (N_2339,N_2107,N_2246);
or U2340 (N_2340,N_2133,N_2199);
xor U2341 (N_2341,N_2141,N_2236);
nand U2342 (N_2342,N_2184,N_2217);
nor U2343 (N_2343,N_2185,N_2161);
or U2344 (N_2344,N_2105,N_2135);
xor U2345 (N_2345,N_2198,N_2164);
xor U2346 (N_2346,N_2238,N_2125);
nand U2347 (N_2347,N_2162,N_2158);
xor U2348 (N_2348,N_2189,N_2187);
nor U2349 (N_2349,N_2214,N_2135);
xor U2350 (N_2350,N_2151,N_2104);
nand U2351 (N_2351,N_2212,N_2150);
xor U2352 (N_2352,N_2141,N_2143);
nand U2353 (N_2353,N_2192,N_2197);
nor U2354 (N_2354,N_2156,N_2185);
xnor U2355 (N_2355,N_2170,N_2119);
nor U2356 (N_2356,N_2134,N_2108);
xnor U2357 (N_2357,N_2249,N_2240);
nand U2358 (N_2358,N_2100,N_2203);
nor U2359 (N_2359,N_2135,N_2163);
xnor U2360 (N_2360,N_2232,N_2106);
nand U2361 (N_2361,N_2100,N_2119);
xnor U2362 (N_2362,N_2137,N_2105);
nand U2363 (N_2363,N_2228,N_2126);
and U2364 (N_2364,N_2119,N_2237);
nand U2365 (N_2365,N_2178,N_2196);
nand U2366 (N_2366,N_2206,N_2129);
and U2367 (N_2367,N_2154,N_2209);
and U2368 (N_2368,N_2243,N_2127);
or U2369 (N_2369,N_2140,N_2148);
nand U2370 (N_2370,N_2175,N_2235);
or U2371 (N_2371,N_2249,N_2195);
or U2372 (N_2372,N_2181,N_2194);
nor U2373 (N_2373,N_2238,N_2197);
or U2374 (N_2374,N_2218,N_2244);
or U2375 (N_2375,N_2146,N_2152);
nor U2376 (N_2376,N_2190,N_2180);
nand U2377 (N_2377,N_2214,N_2179);
or U2378 (N_2378,N_2218,N_2192);
and U2379 (N_2379,N_2160,N_2150);
or U2380 (N_2380,N_2188,N_2190);
nor U2381 (N_2381,N_2187,N_2166);
nor U2382 (N_2382,N_2144,N_2228);
nand U2383 (N_2383,N_2173,N_2205);
nand U2384 (N_2384,N_2112,N_2241);
or U2385 (N_2385,N_2125,N_2141);
nor U2386 (N_2386,N_2227,N_2120);
xor U2387 (N_2387,N_2198,N_2219);
and U2388 (N_2388,N_2143,N_2176);
nand U2389 (N_2389,N_2248,N_2147);
nand U2390 (N_2390,N_2222,N_2110);
and U2391 (N_2391,N_2145,N_2202);
nand U2392 (N_2392,N_2105,N_2156);
xnor U2393 (N_2393,N_2139,N_2145);
and U2394 (N_2394,N_2221,N_2240);
or U2395 (N_2395,N_2201,N_2170);
and U2396 (N_2396,N_2175,N_2226);
nor U2397 (N_2397,N_2125,N_2120);
and U2398 (N_2398,N_2118,N_2226);
nand U2399 (N_2399,N_2205,N_2160);
nand U2400 (N_2400,N_2324,N_2355);
xor U2401 (N_2401,N_2352,N_2323);
and U2402 (N_2402,N_2290,N_2288);
and U2403 (N_2403,N_2302,N_2368);
and U2404 (N_2404,N_2348,N_2276);
and U2405 (N_2405,N_2253,N_2345);
nor U2406 (N_2406,N_2370,N_2356);
nor U2407 (N_2407,N_2316,N_2262);
nand U2408 (N_2408,N_2297,N_2284);
and U2409 (N_2409,N_2318,N_2353);
nor U2410 (N_2410,N_2326,N_2396);
xor U2411 (N_2411,N_2340,N_2259);
nand U2412 (N_2412,N_2254,N_2362);
nand U2413 (N_2413,N_2255,N_2369);
or U2414 (N_2414,N_2378,N_2315);
nand U2415 (N_2415,N_2296,N_2344);
or U2416 (N_2416,N_2321,N_2251);
nor U2417 (N_2417,N_2372,N_2335);
nand U2418 (N_2418,N_2338,N_2398);
nand U2419 (N_2419,N_2390,N_2363);
nor U2420 (N_2420,N_2282,N_2392);
nor U2421 (N_2421,N_2379,N_2266);
and U2422 (N_2422,N_2342,N_2314);
nor U2423 (N_2423,N_2377,N_2277);
or U2424 (N_2424,N_2399,N_2359);
or U2425 (N_2425,N_2364,N_2311);
nand U2426 (N_2426,N_2325,N_2319);
or U2427 (N_2427,N_2291,N_2270);
and U2428 (N_2428,N_2328,N_2275);
nand U2429 (N_2429,N_2286,N_2349);
nor U2430 (N_2430,N_2322,N_2386);
nor U2431 (N_2431,N_2272,N_2334);
or U2432 (N_2432,N_2312,N_2394);
nor U2433 (N_2433,N_2267,N_2292);
and U2434 (N_2434,N_2273,N_2330);
or U2435 (N_2435,N_2351,N_2268);
nand U2436 (N_2436,N_2274,N_2350);
and U2437 (N_2437,N_2306,N_2307);
nand U2438 (N_2438,N_2301,N_2365);
nand U2439 (N_2439,N_2382,N_2357);
and U2440 (N_2440,N_2337,N_2391);
and U2441 (N_2441,N_2397,N_2298);
xnor U2442 (N_2442,N_2295,N_2250);
nand U2443 (N_2443,N_2327,N_2380);
nor U2444 (N_2444,N_2260,N_2317);
nand U2445 (N_2445,N_2257,N_2381);
nand U2446 (N_2446,N_2289,N_2261);
and U2447 (N_2447,N_2331,N_2336);
or U2448 (N_2448,N_2281,N_2341);
and U2449 (N_2449,N_2333,N_2387);
and U2450 (N_2450,N_2373,N_2285);
nor U2451 (N_2451,N_2320,N_2310);
or U2452 (N_2452,N_2271,N_2280);
nand U2453 (N_2453,N_2300,N_2308);
xnor U2454 (N_2454,N_2313,N_2343);
xor U2455 (N_2455,N_2376,N_2375);
nand U2456 (N_2456,N_2304,N_2366);
nand U2457 (N_2457,N_2305,N_2279);
nor U2458 (N_2458,N_2389,N_2256);
or U2459 (N_2459,N_2385,N_2293);
xnor U2460 (N_2460,N_2329,N_2263);
nor U2461 (N_2461,N_2374,N_2384);
nor U2462 (N_2462,N_2395,N_2252);
nand U2463 (N_2463,N_2264,N_2258);
nand U2464 (N_2464,N_2278,N_2269);
nor U2465 (N_2465,N_2339,N_2358);
or U2466 (N_2466,N_2393,N_2383);
or U2467 (N_2467,N_2294,N_2346);
nor U2468 (N_2468,N_2265,N_2360);
nand U2469 (N_2469,N_2367,N_2361);
nand U2470 (N_2470,N_2332,N_2309);
or U2471 (N_2471,N_2303,N_2287);
or U2472 (N_2472,N_2299,N_2371);
nand U2473 (N_2473,N_2388,N_2354);
and U2474 (N_2474,N_2347,N_2283);
xor U2475 (N_2475,N_2330,N_2383);
nand U2476 (N_2476,N_2269,N_2384);
and U2477 (N_2477,N_2372,N_2320);
xnor U2478 (N_2478,N_2398,N_2302);
nand U2479 (N_2479,N_2346,N_2371);
and U2480 (N_2480,N_2256,N_2299);
xnor U2481 (N_2481,N_2253,N_2386);
nor U2482 (N_2482,N_2325,N_2322);
or U2483 (N_2483,N_2370,N_2377);
nor U2484 (N_2484,N_2360,N_2336);
xnor U2485 (N_2485,N_2331,N_2270);
nand U2486 (N_2486,N_2294,N_2267);
and U2487 (N_2487,N_2262,N_2335);
xor U2488 (N_2488,N_2397,N_2378);
nor U2489 (N_2489,N_2295,N_2299);
nand U2490 (N_2490,N_2369,N_2374);
nand U2491 (N_2491,N_2281,N_2299);
and U2492 (N_2492,N_2288,N_2368);
and U2493 (N_2493,N_2368,N_2378);
nand U2494 (N_2494,N_2265,N_2258);
xnor U2495 (N_2495,N_2301,N_2397);
xnor U2496 (N_2496,N_2319,N_2324);
or U2497 (N_2497,N_2371,N_2325);
xor U2498 (N_2498,N_2311,N_2277);
or U2499 (N_2499,N_2286,N_2268);
xor U2500 (N_2500,N_2320,N_2265);
nand U2501 (N_2501,N_2312,N_2341);
xor U2502 (N_2502,N_2289,N_2270);
or U2503 (N_2503,N_2351,N_2326);
or U2504 (N_2504,N_2395,N_2290);
nor U2505 (N_2505,N_2289,N_2383);
xor U2506 (N_2506,N_2366,N_2341);
and U2507 (N_2507,N_2313,N_2362);
and U2508 (N_2508,N_2360,N_2308);
xor U2509 (N_2509,N_2300,N_2253);
and U2510 (N_2510,N_2385,N_2265);
nor U2511 (N_2511,N_2333,N_2307);
xor U2512 (N_2512,N_2365,N_2300);
or U2513 (N_2513,N_2341,N_2325);
nand U2514 (N_2514,N_2350,N_2288);
nor U2515 (N_2515,N_2358,N_2291);
nor U2516 (N_2516,N_2342,N_2393);
xnor U2517 (N_2517,N_2285,N_2386);
nor U2518 (N_2518,N_2318,N_2385);
nor U2519 (N_2519,N_2359,N_2295);
nand U2520 (N_2520,N_2290,N_2330);
or U2521 (N_2521,N_2372,N_2284);
and U2522 (N_2522,N_2378,N_2289);
and U2523 (N_2523,N_2370,N_2250);
xnor U2524 (N_2524,N_2347,N_2293);
nand U2525 (N_2525,N_2271,N_2277);
xnor U2526 (N_2526,N_2344,N_2329);
and U2527 (N_2527,N_2335,N_2261);
nand U2528 (N_2528,N_2321,N_2380);
nand U2529 (N_2529,N_2342,N_2286);
nand U2530 (N_2530,N_2274,N_2330);
xnor U2531 (N_2531,N_2340,N_2323);
or U2532 (N_2532,N_2251,N_2382);
and U2533 (N_2533,N_2283,N_2301);
and U2534 (N_2534,N_2387,N_2251);
or U2535 (N_2535,N_2319,N_2326);
xnor U2536 (N_2536,N_2250,N_2347);
and U2537 (N_2537,N_2308,N_2313);
nor U2538 (N_2538,N_2377,N_2357);
xor U2539 (N_2539,N_2328,N_2363);
nand U2540 (N_2540,N_2312,N_2350);
xor U2541 (N_2541,N_2387,N_2316);
nand U2542 (N_2542,N_2287,N_2361);
xnor U2543 (N_2543,N_2260,N_2312);
or U2544 (N_2544,N_2375,N_2315);
nor U2545 (N_2545,N_2315,N_2278);
nand U2546 (N_2546,N_2259,N_2318);
xor U2547 (N_2547,N_2278,N_2317);
and U2548 (N_2548,N_2255,N_2361);
nand U2549 (N_2549,N_2278,N_2321);
xnor U2550 (N_2550,N_2411,N_2430);
xor U2551 (N_2551,N_2510,N_2487);
or U2552 (N_2552,N_2465,N_2436);
nand U2553 (N_2553,N_2531,N_2456);
or U2554 (N_2554,N_2404,N_2418);
nand U2555 (N_2555,N_2495,N_2543);
xnor U2556 (N_2556,N_2403,N_2461);
nor U2557 (N_2557,N_2522,N_2485);
nand U2558 (N_2558,N_2450,N_2410);
nor U2559 (N_2559,N_2412,N_2513);
xnor U2560 (N_2560,N_2529,N_2521);
xnor U2561 (N_2561,N_2439,N_2499);
xnor U2562 (N_2562,N_2435,N_2518);
nor U2563 (N_2563,N_2401,N_2400);
nor U2564 (N_2564,N_2477,N_2471);
or U2565 (N_2565,N_2462,N_2544);
nor U2566 (N_2566,N_2519,N_2492);
nand U2567 (N_2567,N_2420,N_2451);
and U2568 (N_2568,N_2423,N_2445);
xnor U2569 (N_2569,N_2498,N_2490);
nand U2570 (N_2570,N_2429,N_2523);
and U2571 (N_2571,N_2475,N_2511);
and U2572 (N_2572,N_2447,N_2483);
or U2573 (N_2573,N_2524,N_2546);
nor U2574 (N_2574,N_2507,N_2532);
xnor U2575 (N_2575,N_2419,N_2549);
or U2576 (N_2576,N_2496,N_2443);
nand U2577 (N_2577,N_2458,N_2488);
or U2578 (N_2578,N_2448,N_2449);
xor U2579 (N_2579,N_2484,N_2512);
nor U2580 (N_2580,N_2506,N_2446);
and U2581 (N_2581,N_2497,N_2452);
or U2582 (N_2582,N_2427,N_2489);
nor U2583 (N_2583,N_2402,N_2474);
and U2584 (N_2584,N_2520,N_2486);
and U2585 (N_2585,N_2538,N_2541);
nor U2586 (N_2586,N_2501,N_2407);
nor U2587 (N_2587,N_2476,N_2480);
xnor U2588 (N_2588,N_2432,N_2464);
or U2589 (N_2589,N_2516,N_2409);
or U2590 (N_2590,N_2417,N_2455);
xor U2591 (N_2591,N_2548,N_2530);
xor U2592 (N_2592,N_2536,N_2503);
nor U2593 (N_2593,N_2504,N_2508);
nor U2594 (N_2594,N_2437,N_2406);
and U2595 (N_2595,N_2428,N_2424);
nand U2596 (N_2596,N_2470,N_2535);
nand U2597 (N_2597,N_2500,N_2493);
nand U2598 (N_2598,N_2442,N_2468);
nand U2599 (N_2599,N_2405,N_2482);
xnor U2600 (N_2600,N_2509,N_2415);
nand U2601 (N_2601,N_2505,N_2425);
and U2602 (N_2602,N_2413,N_2444);
and U2603 (N_2603,N_2547,N_2416);
and U2604 (N_2604,N_2517,N_2479);
and U2605 (N_2605,N_2526,N_2453);
nor U2606 (N_2606,N_2467,N_2460);
nand U2607 (N_2607,N_2528,N_2481);
nor U2608 (N_2608,N_2441,N_2440);
nor U2609 (N_2609,N_2539,N_2527);
xor U2610 (N_2610,N_2473,N_2472);
nor U2611 (N_2611,N_2459,N_2545);
xnor U2612 (N_2612,N_2494,N_2540);
nor U2613 (N_2613,N_2457,N_2421);
nand U2614 (N_2614,N_2502,N_2463);
nor U2615 (N_2615,N_2426,N_2466);
nand U2616 (N_2616,N_2534,N_2514);
nor U2617 (N_2617,N_2533,N_2431);
or U2618 (N_2618,N_2478,N_2433);
nor U2619 (N_2619,N_2434,N_2454);
nor U2620 (N_2620,N_2542,N_2525);
and U2621 (N_2621,N_2438,N_2408);
xnor U2622 (N_2622,N_2414,N_2537);
nand U2623 (N_2623,N_2422,N_2515);
nor U2624 (N_2624,N_2469,N_2491);
or U2625 (N_2625,N_2527,N_2449);
or U2626 (N_2626,N_2494,N_2504);
nor U2627 (N_2627,N_2522,N_2429);
or U2628 (N_2628,N_2467,N_2535);
nand U2629 (N_2629,N_2508,N_2422);
nand U2630 (N_2630,N_2413,N_2500);
nor U2631 (N_2631,N_2410,N_2534);
nor U2632 (N_2632,N_2465,N_2526);
xnor U2633 (N_2633,N_2424,N_2482);
nor U2634 (N_2634,N_2437,N_2473);
and U2635 (N_2635,N_2429,N_2486);
nand U2636 (N_2636,N_2488,N_2481);
and U2637 (N_2637,N_2509,N_2503);
nand U2638 (N_2638,N_2452,N_2400);
xnor U2639 (N_2639,N_2520,N_2492);
nand U2640 (N_2640,N_2499,N_2403);
nand U2641 (N_2641,N_2489,N_2443);
or U2642 (N_2642,N_2534,N_2432);
nor U2643 (N_2643,N_2441,N_2429);
or U2644 (N_2644,N_2410,N_2419);
nand U2645 (N_2645,N_2456,N_2501);
xnor U2646 (N_2646,N_2415,N_2522);
xnor U2647 (N_2647,N_2424,N_2408);
or U2648 (N_2648,N_2500,N_2528);
or U2649 (N_2649,N_2467,N_2442);
nor U2650 (N_2650,N_2410,N_2470);
nand U2651 (N_2651,N_2425,N_2532);
nor U2652 (N_2652,N_2455,N_2456);
or U2653 (N_2653,N_2459,N_2522);
or U2654 (N_2654,N_2487,N_2548);
or U2655 (N_2655,N_2470,N_2530);
or U2656 (N_2656,N_2518,N_2530);
nor U2657 (N_2657,N_2415,N_2505);
nand U2658 (N_2658,N_2445,N_2420);
or U2659 (N_2659,N_2411,N_2485);
xor U2660 (N_2660,N_2484,N_2533);
xor U2661 (N_2661,N_2408,N_2523);
and U2662 (N_2662,N_2502,N_2454);
xor U2663 (N_2663,N_2448,N_2444);
and U2664 (N_2664,N_2468,N_2439);
and U2665 (N_2665,N_2402,N_2461);
and U2666 (N_2666,N_2433,N_2483);
nand U2667 (N_2667,N_2444,N_2478);
or U2668 (N_2668,N_2541,N_2521);
nor U2669 (N_2669,N_2466,N_2486);
xnor U2670 (N_2670,N_2450,N_2448);
nor U2671 (N_2671,N_2512,N_2516);
nand U2672 (N_2672,N_2491,N_2421);
xnor U2673 (N_2673,N_2518,N_2466);
xor U2674 (N_2674,N_2532,N_2429);
nor U2675 (N_2675,N_2486,N_2499);
or U2676 (N_2676,N_2413,N_2454);
nand U2677 (N_2677,N_2437,N_2413);
and U2678 (N_2678,N_2549,N_2446);
or U2679 (N_2679,N_2455,N_2452);
xor U2680 (N_2680,N_2495,N_2435);
nor U2681 (N_2681,N_2445,N_2548);
nand U2682 (N_2682,N_2526,N_2469);
or U2683 (N_2683,N_2513,N_2436);
and U2684 (N_2684,N_2543,N_2511);
or U2685 (N_2685,N_2475,N_2421);
and U2686 (N_2686,N_2491,N_2525);
nor U2687 (N_2687,N_2445,N_2429);
nor U2688 (N_2688,N_2520,N_2467);
nor U2689 (N_2689,N_2441,N_2508);
xnor U2690 (N_2690,N_2437,N_2537);
xor U2691 (N_2691,N_2474,N_2527);
xnor U2692 (N_2692,N_2531,N_2425);
and U2693 (N_2693,N_2523,N_2431);
and U2694 (N_2694,N_2520,N_2460);
and U2695 (N_2695,N_2511,N_2471);
and U2696 (N_2696,N_2511,N_2460);
nand U2697 (N_2697,N_2537,N_2526);
or U2698 (N_2698,N_2454,N_2458);
or U2699 (N_2699,N_2433,N_2403);
or U2700 (N_2700,N_2620,N_2574);
nor U2701 (N_2701,N_2587,N_2693);
nor U2702 (N_2702,N_2573,N_2662);
and U2703 (N_2703,N_2595,N_2576);
xnor U2704 (N_2704,N_2568,N_2653);
nor U2705 (N_2705,N_2650,N_2624);
nor U2706 (N_2706,N_2691,N_2649);
and U2707 (N_2707,N_2556,N_2641);
and U2708 (N_2708,N_2580,N_2593);
nand U2709 (N_2709,N_2611,N_2644);
or U2710 (N_2710,N_2630,N_2564);
or U2711 (N_2711,N_2670,N_2577);
or U2712 (N_2712,N_2591,N_2553);
xnor U2713 (N_2713,N_2689,N_2654);
or U2714 (N_2714,N_2609,N_2686);
nor U2715 (N_2715,N_2677,N_2652);
xnor U2716 (N_2716,N_2601,N_2661);
nand U2717 (N_2717,N_2598,N_2643);
nand U2718 (N_2718,N_2578,N_2692);
nand U2719 (N_2719,N_2694,N_2665);
xor U2720 (N_2720,N_2600,N_2636);
and U2721 (N_2721,N_2583,N_2680);
and U2722 (N_2722,N_2633,N_2698);
or U2723 (N_2723,N_2596,N_2603);
and U2724 (N_2724,N_2561,N_2687);
nor U2725 (N_2725,N_2555,N_2579);
nor U2726 (N_2726,N_2637,N_2666);
nand U2727 (N_2727,N_2559,N_2554);
or U2728 (N_2728,N_2629,N_2567);
and U2729 (N_2729,N_2639,N_2614);
or U2730 (N_2730,N_2599,N_2594);
or U2731 (N_2731,N_2638,N_2628);
xor U2732 (N_2732,N_2659,N_2563);
or U2733 (N_2733,N_2655,N_2634);
nor U2734 (N_2734,N_2565,N_2642);
or U2735 (N_2735,N_2627,N_2695);
or U2736 (N_2736,N_2612,N_2632);
or U2737 (N_2737,N_2605,N_2604);
nor U2738 (N_2738,N_2571,N_2635);
xor U2739 (N_2739,N_2672,N_2651);
nand U2740 (N_2740,N_2625,N_2613);
and U2741 (N_2741,N_2657,N_2592);
xor U2742 (N_2742,N_2621,N_2688);
or U2743 (N_2743,N_2645,N_2674);
or U2744 (N_2744,N_2615,N_2558);
nor U2745 (N_2745,N_2551,N_2618);
nor U2746 (N_2746,N_2616,N_2572);
nand U2747 (N_2747,N_2685,N_2570);
nand U2748 (N_2748,N_2582,N_2646);
or U2749 (N_2749,N_2682,N_2671);
nand U2750 (N_2750,N_2602,N_2566);
and U2751 (N_2751,N_2562,N_2658);
nand U2752 (N_2752,N_2697,N_2607);
and U2753 (N_2753,N_2699,N_2569);
nor U2754 (N_2754,N_2676,N_2584);
nor U2755 (N_2755,N_2585,N_2631);
or U2756 (N_2756,N_2590,N_2684);
or U2757 (N_2757,N_2656,N_2552);
nor U2758 (N_2758,N_2560,N_2588);
nand U2759 (N_2759,N_2664,N_2660);
and U2760 (N_2760,N_2679,N_2669);
nor U2761 (N_2761,N_2617,N_2608);
nand U2762 (N_2762,N_2581,N_2597);
xor U2763 (N_2763,N_2619,N_2589);
and U2764 (N_2764,N_2626,N_2668);
and U2765 (N_2765,N_2550,N_2696);
and U2766 (N_2766,N_2623,N_2586);
or U2767 (N_2767,N_2683,N_2663);
xor U2768 (N_2768,N_2673,N_2667);
nor U2769 (N_2769,N_2678,N_2610);
xnor U2770 (N_2770,N_2557,N_2647);
nor U2771 (N_2771,N_2648,N_2575);
nand U2772 (N_2772,N_2681,N_2675);
nand U2773 (N_2773,N_2622,N_2690);
or U2774 (N_2774,N_2640,N_2606);
and U2775 (N_2775,N_2625,N_2642);
nand U2776 (N_2776,N_2681,N_2577);
nand U2777 (N_2777,N_2619,N_2591);
nor U2778 (N_2778,N_2556,N_2669);
nand U2779 (N_2779,N_2609,N_2623);
nor U2780 (N_2780,N_2564,N_2619);
nand U2781 (N_2781,N_2558,N_2698);
xnor U2782 (N_2782,N_2632,N_2677);
or U2783 (N_2783,N_2594,N_2603);
xnor U2784 (N_2784,N_2571,N_2593);
xor U2785 (N_2785,N_2691,N_2551);
nand U2786 (N_2786,N_2608,N_2572);
nor U2787 (N_2787,N_2696,N_2615);
nand U2788 (N_2788,N_2653,N_2640);
nand U2789 (N_2789,N_2620,N_2621);
xnor U2790 (N_2790,N_2622,N_2675);
and U2791 (N_2791,N_2620,N_2556);
xnor U2792 (N_2792,N_2558,N_2641);
xnor U2793 (N_2793,N_2693,N_2563);
nor U2794 (N_2794,N_2591,N_2589);
and U2795 (N_2795,N_2697,N_2562);
nand U2796 (N_2796,N_2657,N_2654);
xor U2797 (N_2797,N_2619,N_2562);
and U2798 (N_2798,N_2687,N_2623);
or U2799 (N_2799,N_2562,N_2593);
xor U2800 (N_2800,N_2638,N_2612);
or U2801 (N_2801,N_2558,N_2594);
nand U2802 (N_2802,N_2574,N_2631);
and U2803 (N_2803,N_2639,N_2644);
nand U2804 (N_2804,N_2606,N_2622);
nor U2805 (N_2805,N_2679,N_2568);
nand U2806 (N_2806,N_2636,N_2582);
nand U2807 (N_2807,N_2693,N_2682);
xor U2808 (N_2808,N_2580,N_2639);
nand U2809 (N_2809,N_2677,N_2619);
nand U2810 (N_2810,N_2604,N_2627);
and U2811 (N_2811,N_2579,N_2645);
or U2812 (N_2812,N_2690,N_2670);
or U2813 (N_2813,N_2643,N_2594);
nor U2814 (N_2814,N_2581,N_2646);
or U2815 (N_2815,N_2694,N_2633);
or U2816 (N_2816,N_2658,N_2551);
nor U2817 (N_2817,N_2604,N_2551);
and U2818 (N_2818,N_2620,N_2666);
nor U2819 (N_2819,N_2607,N_2684);
nand U2820 (N_2820,N_2691,N_2591);
or U2821 (N_2821,N_2623,N_2655);
nand U2822 (N_2822,N_2631,N_2591);
nand U2823 (N_2823,N_2595,N_2565);
xnor U2824 (N_2824,N_2625,N_2604);
xor U2825 (N_2825,N_2674,N_2571);
or U2826 (N_2826,N_2609,N_2667);
or U2827 (N_2827,N_2550,N_2609);
nor U2828 (N_2828,N_2618,N_2627);
and U2829 (N_2829,N_2575,N_2662);
nand U2830 (N_2830,N_2664,N_2622);
or U2831 (N_2831,N_2628,N_2606);
xor U2832 (N_2832,N_2642,N_2606);
and U2833 (N_2833,N_2694,N_2654);
nand U2834 (N_2834,N_2648,N_2668);
or U2835 (N_2835,N_2648,N_2593);
and U2836 (N_2836,N_2588,N_2585);
nand U2837 (N_2837,N_2551,N_2608);
nor U2838 (N_2838,N_2690,N_2661);
nand U2839 (N_2839,N_2644,N_2676);
nand U2840 (N_2840,N_2698,N_2695);
xnor U2841 (N_2841,N_2648,N_2622);
and U2842 (N_2842,N_2597,N_2685);
or U2843 (N_2843,N_2603,N_2672);
nand U2844 (N_2844,N_2645,N_2649);
xnor U2845 (N_2845,N_2557,N_2676);
nand U2846 (N_2846,N_2626,N_2606);
or U2847 (N_2847,N_2650,N_2615);
nor U2848 (N_2848,N_2565,N_2588);
nor U2849 (N_2849,N_2586,N_2612);
xor U2850 (N_2850,N_2728,N_2781);
and U2851 (N_2851,N_2755,N_2825);
and U2852 (N_2852,N_2718,N_2784);
nand U2853 (N_2853,N_2743,N_2737);
or U2854 (N_2854,N_2790,N_2747);
nand U2855 (N_2855,N_2705,N_2845);
xor U2856 (N_2856,N_2838,N_2736);
xor U2857 (N_2857,N_2770,N_2836);
nand U2858 (N_2858,N_2815,N_2708);
nand U2859 (N_2859,N_2774,N_2767);
or U2860 (N_2860,N_2734,N_2773);
or U2861 (N_2861,N_2744,N_2745);
nor U2862 (N_2862,N_2811,N_2722);
nand U2863 (N_2863,N_2751,N_2709);
or U2864 (N_2864,N_2814,N_2733);
nand U2865 (N_2865,N_2776,N_2823);
or U2866 (N_2866,N_2843,N_2740);
xor U2867 (N_2867,N_2818,N_2830);
nor U2868 (N_2868,N_2837,N_2804);
or U2869 (N_2869,N_2723,N_2731);
nor U2870 (N_2870,N_2729,N_2765);
xor U2871 (N_2871,N_2735,N_2715);
and U2872 (N_2872,N_2732,N_2748);
or U2873 (N_2873,N_2749,N_2730);
nand U2874 (N_2874,N_2788,N_2824);
nor U2875 (N_2875,N_2721,N_2707);
or U2876 (N_2876,N_2766,N_2758);
or U2877 (N_2877,N_2792,N_2754);
or U2878 (N_2878,N_2704,N_2787);
nor U2879 (N_2879,N_2716,N_2741);
nor U2880 (N_2880,N_2726,N_2817);
nor U2881 (N_2881,N_2701,N_2808);
and U2882 (N_2882,N_2777,N_2757);
or U2883 (N_2883,N_2785,N_2752);
or U2884 (N_2884,N_2848,N_2826);
and U2885 (N_2885,N_2778,N_2783);
nand U2886 (N_2886,N_2812,N_2719);
and U2887 (N_2887,N_2849,N_2798);
nand U2888 (N_2888,N_2759,N_2762);
xor U2889 (N_2889,N_2789,N_2786);
nor U2890 (N_2890,N_2714,N_2793);
and U2891 (N_2891,N_2844,N_2750);
xor U2892 (N_2892,N_2700,N_2780);
nor U2893 (N_2893,N_2713,N_2724);
xor U2894 (N_2894,N_2764,N_2833);
nand U2895 (N_2895,N_2847,N_2829);
xor U2896 (N_2896,N_2822,N_2703);
nor U2897 (N_2897,N_2782,N_2711);
or U2898 (N_2898,N_2720,N_2797);
nor U2899 (N_2899,N_2803,N_2820);
nor U2900 (N_2900,N_2809,N_2763);
nand U2901 (N_2901,N_2839,N_2702);
xor U2902 (N_2902,N_2768,N_2794);
and U2903 (N_2903,N_2710,N_2760);
nand U2904 (N_2904,N_2828,N_2727);
nand U2905 (N_2905,N_2842,N_2835);
nand U2906 (N_2906,N_2746,N_2775);
and U2907 (N_2907,N_2807,N_2706);
and U2908 (N_2908,N_2712,N_2827);
xnor U2909 (N_2909,N_2739,N_2791);
nor U2910 (N_2910,N_2834,N_2772);
or U2911 (N_2911,N_2840,N_2795);
nor U2912 (N_2912,N_2832,N_2846);
nand U2913 (N_2913,N_2753,N_2800);
and U2914 (N_2914,N_2802,N_2779);
and U2915 (N_2915,N_2771,N_2769);
nor U2916 (N_2916,N_2717,N_2725);
and U2917 (N_2917,N_2796,N_2821);
and U2918 (N_2918,N_2816,N_2799);
and U2919 (N_2919,N_2738,N_2813);
nor U2920 (N_2920,N_2742,N_2841);
xnor U2921 (N_2921,N_2756,N_2761);
or U2922 (N_2922,N_2819,N_2831);
nor U2923 (N_2923,N_2806,N_2805);
or U2924 (N_2924,N_2810,N_2801);
nand U2925 (N_2925,N_2814,N_2757);
or U2926 (N_2926,N_2740,N_2847);
nor U2927 (N_2927,N_2829,N_2742);
nor U2928 (N_2928,N_2803,N_2842);
nor U2929 (N_2929,N_2846,N_2728);
xor U2930 (N_2930,N_2743,N_2725);
or U2931 (N_2931,N_2731,N_2704);
xnor U2932 (N_2932,N_2704,N_2806);
nor U2933 (N_2933,N_2811,N_2760);
nor U2934 (N_2934,N_2802,N_2788);
nand U2935 (N_2935,N_2751,N_2824);
nor U2936 (N_2936,N_2777,N_2745);
xor U2937 (N_2937,N_2729,N_2810);
nand U2938 (N_2938,N_2718,N_2768);
or U2939 (N_2939,N_2821,N_2725);
nand U2940 (N_2940,N_2828,N_2811);
or U2941 (N_2941,N_2731,N_2782);
nor U2942 (N_2942,N_2753,N_2812);
nor U2943 (N_2943,N_2819,N_2754);
nor U2944 (N_2944,N_2738,N_2812);
and U2945 (N_2945,N_2830,N_2729);
or U2946 (N_2946,N_2768,N_2715);
nand U2947 (N_2947,N_2811,N_2837);
and U2948 (N_2948,N_2829,N_2719);
nor U2949 (N_2949,N_2803,N_2705);
or U2950 (N_2950,N_2710,N_2746);
nor U2951 (N_2951,N_2715,N_2777);
nand U2952 (N_2952,N_2818,N_2731);
nor U2953 (N_2953,N_2835,N_2769);
nand U2954 (N_2954,N_2740,N_2822);
nor U2955 (N_2955,N_2830,N_2761);
or U2956 (N_2956,N_2804,N_2796);
nand U2957 (N_2957,N_2713,N_2764);
nand U2958 (N_2958,N_2839,N_2786);
and U2959 (N_2959,N_2720,N_2750);
xor U2960 (N_2960,N_2744,N_2830);
or U2961 (N_2961,N_2735,N_2775);
nand U2962 (N_2962,N_2813,N_2700);
xnor U2963 (N_2963,N_2799,N_2798);
nor U2964 (N_2964,N_2727,N_2745);
or U2965 (N_2965,N_2818,N_2771);
xor U2966 (N_2966,N_2783,N_2813);
nand U2967 (N_2967,N_2811,N_2748);
or U2968 (N_2968,N_2715,N_2757);
and U2969 (N_2969,N_2811,N_2790);
nand U2970 (N_2970,N_2740,N_2778);
xnor U2971 (N_2971,N_2751,N_2795);
nand U2972 (N_2972,N_2716,N_2757);
xnor U2973 (N_2973,N_2772,N_2722);
xnor U2974 (N_2974,N_2748,N_2802);
and U2975 (N_2975,N_2729,N_2767);
nor U2976 (N_2976,N_2780,N_2834);
xnor U2977 (N_2977,N_2832,N_2700);
and U2978 (N_2978,N_2760,N_2717);
nand U2979 (N_2979,N_2798,N_2813);
and U2980 (N_2980,N_2811,N_2702);
and U2981 (N_2981,N_2828,N_2758);
or U2982 (N_2982,N_2810,N_2756);
or U2983 (N_2983,N_2759,N_2738);
or U2984 (N_2984,N_2849,N_2755);
xnor U2985 (N_2985,N_2751,N_2842);
and U2986 (N_2986,N_2704,N_2751);
or U2987 (N_2987,N_2711,N_2746);
nor U2988 (N_2988,N_2707,N_2820);
xnor U2989 (N_2989,N_2781,N_2826);
nor U2990 (N_2990,N_2757,N_2843);
nor U2991 (N_2991,N_2716,N_2801);
nor U2992 (N_2992,N_2708,N_2843);
nor U2993 (N_2993,N_2737,N_2803);
or U2994 (N_2994,N_2758,N_2786);
nor U2995 (N_2995,N_2725,N_2728);
nand U2996 (N_2996,N_2731,N_2831);
nand U2997 (N_2997,N_2768,N_2807);
or U2998 (N_2998,N_2801,N_2753);
nor U2999 (N_2999,N_2835,N_2808);
xor U3000 (N_3000,N_2959,N_2958);
xor U3001 (N_3001,N_2895,N_2901);
nor U3002 (N_3002,N_2893,N_2899);
nand U3003 (N_3003,N_2978,N_2871);
and U3004 (N_3004,N_2855,N_2986);
or U3005 (N_3005,N_2993,N_2890);
xnor U3006 (N_3006,N_2902,N_2955);
xnor U3007 (N_3007,N_2939,N_2949);
nand U3008 (N_3008,N_2960,N_2953);
nor U3009 (N_3009,N_2860,N_2966);
nand U3010 (N_3010,N_2905,N_2879);
nor U3011 (N_3011,N_2979,N_2873);
and U3012 (N_3012,N_2883,N_2963);
nand U3013 (N_3013,N_2909,N_2850);
or U3014 (N_3014,N_2919,N_2970);
nor U3015 (N_3015,N_2930,N_2859);
and U3016 (N_3016,N_2863,N_2867);
nor U3017 (N_3017,N_2882,N_2858);
or U3018 (N_3018,N_2932,N_2985);
nor U3019 (N_3019,N_2911,N_2976);
and U3020 (N_3020,N_2968,N_2929);
and U3021 (N_3021,N_2941,N_2887);
and U3022 (N_3022,N_2916,N_2940);
xnor U3023 (N_3023,N_2857,N_2875);
xnor U3024 (N_3024,N_2881,N_2974);
nor U3025 (N_3025,N_2994,N_2935);
or U3026 (N_3026,N_2878,N_2892);
nand U3027 (N_3027,N_2922,N_2945);
and U3028 (N_3028,N_2885,N_2880);
or U3029 (N_3029,N_2972,N_2999);
xor U3030 (N_3030,N_2889,N_2980);
xor U3031 (N_3031,N_2952,N_2977);
or U3032 (N_3032,N_2898,N_2983);
xnor U3033 (N_3033,N_2888,N_2896);
or U3034 (N_3034,N_2884,N_2923);
or U3035 (N_3035,N_2852,N_2915);
xnor U3036 (N_3036,N_2967,N_2965);
and U3037 (N_3037,N_2918,N_2920);
xnor U3038 (N_3038,N_2903,N_2862);
xnor U3039 (N_3039,N_2851,N_2997);
or U3040 (N_3040,N_2856,N_2931);
xnor U3041 (N_3041,N_2897,N_2928);
and U3042 (N_3042,N_2947,N_2942);
nand U3043 (N_3043,N_2962,N_2969);
nor U3044 (N_3044,N_2964,N_2973);
nor U3045 (N_3045,N_2865,N_2908);
and U3046 (N_3046,N_2951,N_2995);
and U3047 (N_3047,N_2938,N_2917);
or U3048 (N_3048,N_2961,N_2944);
or U3049 (N_3049,N_2934,N_2954);
xnor U3050 (N_3050,N_2996,N_2866);
nand U3051 (N_3051,N_2927,N_2872);
or U3052 (N_3052,N_2989,N_2992);
nand U3053 (N_3053,N_2921,N_2988);
nand U3054 (N_3054,N_2891,N_2950);
or U3055 (N_3055,N_2868,N_2990);
xnor U3056 (N_3056,N_2936,N_2913);
or U3057 (N_3057,N_2876,N_2982);
nor U3058 (N_3058,N_2948,N_2877);
or U3059 (N_3059,N_2933,N_2924);
nor U3060 (N_3060,N_2869,N_2925);
nor U3061 (N_3061,N_2907,N_2957);
xor U3062 (N_3062,N_2984,N_2906);
and U3063 (N_3063,N_2854,N_2900);
or U3064 (N_3064,N_2853,N_2937);
nand U3065 (N_3065,N_2946,N_2991);
nand U3066 (N_3066,N_2886,N_2926);
nand U3067 (N_3067,N_2914,N_2912);
nor U3068 (N_3068,N_2956,N_2987);
and U3069 (N_3069,N_2943,N_2861);
nand U3070 (N_3070,N_2998,N_2910);
nand U3071 (N_3071,N_2904,N_2870);
xnor U3072 (N_3072,N_2975,N_2874);
nor U3073 (N_3073,N_2971,N_2981);
and U3074 (N_3074,N_2894,N_2864);
nand U3075 (N_3075,N_2991,N_2930);
nand U3076 (N_3076,N_2974,N_2972);
xor U3077 (N_3077,N_2947,N_2995);
nor U3078 (N_3078,N_2868,N_2925);
xor U3079 (N_3079,N_2875,N_2899);
or U3080 (N_3080,N_2883,N_2980);
nor U3081 (N_3081,N_2946,N_2973);
nor U3082 (N_3082,N_2967,N_2857);
xnor U3083 (N_3083,N_2964,N_2982);
or U3084 (N_3084,N_2878,N_2924);
xnor U3085 (N_3085,N_2905,N_2987);
and U3086 (N_3086,N_2893,N_2953);
nand U3087 (N_3087,N_2857,N_2954);
or U3088 (N_3088,N_2953,N_2972);
nor U3089 (N_3089,N_2876,N_2908);
nor U3090 (N_3090,N_2929,N_2882);
and U3091 (N_3091,N_2941,N_2990);
xor U3092 (N_3092,N_2950,N_2888);
and U3093 (N_3093,N_2963,N_2925);
and U3094 (N_3094,N_2923,N_2915);
nor U3095 (N_3095,N_2921,N_2997);
and U3096 (N_3096,N_2893,N_2947);
or U3097 (N_3097,N_2882,N_2874);
and U3098 (N_3098,N_2872,N_2903);
xnor U3099 (N_3099,N_2857,N_2982);
or U3100 (N_3100,N_2925,N_2883);
or U3101 (N_3101,N_2942,N_2932);
or U3102 (N_3102,N_2979,N_2952);
or U3103 (N_3103,N_2929,N_2877);
or U3104 (N_3104,N_2921,N_2965);
xnor U3105 (N_3105,N_2980,N_2999);
nor U3106 (N_3106,N_2903,N_2973);
nor U3107 (N_3107,N_2956,N_2897);
xor U3108 (N_3108,N_2998,N_2948);
or U3109 (N_3109,N_2998,N_2930);
and U3110 (N_3110,N_2890,N_2960);
and U3111 (N_3111,N_2857,N_2997);
and U3112 (N_3112,N_2900,N_2871);
or U3113 (N_3113,N_2863,N_2971);
nor U3114 (N_3114,N_2927,N_2969);
and U3115 (N_3115,N_2876,N_2857);
nand U3116 (N_3116,N_2912,N_2898);
xnor U3117 (N_3117,N_2875,N_2894);
nand U3118 (N_3118,N_2938,N_2982);
nand U3119 (N_3119,N_2890,N_2952);
or U3120 (N_3120,N_2892,N_2905);
and U3121 (N_3121,N_2864,N_2981);
nand U3122 (N_3122,N_2857,N_2873);
nor U3123 (N_3123,N_2866,N_2959);
nand U3124 (N_3124,N_2933,N_2863);
and U3125 (N_3125,N_2932,N_2988);
or U3126 (N_3126,N_2974,N_2873);
xnor U3127 (N_3127,N_2977,N_2910);
nor U3128 (N_3128,N_2997,N_2928);
and U3129 (N_3129,N_2865,N_2958);
nand U3130 (N_3130,N_2918,N_2987);
nor U3131 (N_3131,N_2887,N_2880);
xor U3132 (N_3132,N_2929,N_2978);
or U3133 (N_3133,N_2998,N_2867);
nor U3134 (N_3134,N_2910,N_2943);
nand U3135 (N_3135,N_2928,N_2947);
nand U3136 (N_3136,N_2875,N_2983);
and U3137 (N_3137,N_2865,N_2872);
nor U3138 (N_3138,N_2934,N_2913);
xor U3139 (N_3139,N_2995,N_2926);
xnor U3140 (N_3140,N_2938,N_2972);
nand U3141 (N_3141,N_2893,N_2866);
xnor U3142 (N_3142,N_2965,N_2982);
or U3143 (N_3143,N_2878,N_2966);
and U3144 (N_3144,N_2878,N_2921);
nand U3145 (N_3145,N_2962,N_2964);
nor U3146 (N_3146,N_2879,N_2888);
nor U3147 (N_3147,N_2991,N_2958);
or U3148 (N_3148,N_2869,N_2897);
nor U3149 (N_3149,N_2952,N_2855);
and U3150 (N_3150,N_3133,N_3015);
or U3151 (N_3151,N_3034,N_3116);
xnor U3152 (N_3152,N_3102,N_3077);
or U3153 (N_3153,N_3089,N_3018);
xor U3154 (N_3154,N_3031,N_3057);
or U3155 (N_3155,N_3060,N_3117);
nor U3156 (N_3156,N_3019,N_3052);
xor U3157 (N_3157,N_3041,N_3097);
or U3158 (N_3158,N_3098,N_3070);
and U3159 (N_3159,N_3064,N_3010);
and U3160 (N_3160,N_3071,N_3056);
xor U3161 (N_3161,N_3037,N_3091);
nand U3162 (N_3162,N_3028,N_3130);
or U3163 (N_3163,N_3027,N_3144);
nor U3164 (N_3164,N_3022,N_3029);
xnor U3165 (N_3165,N_3124,N_3069);
nand U3166 (N_3166,N_3120,N_3007);
nand U3167 (N_3167,N_3093,N_3083);
nand U3168 (N_3168,N_3009,N_3039);
nand U3169 (N_3169,N_3001,N_3136);
xor U3170 (N_3170,N_3067,N_3101);
nor U3171 (N_3171,N_3012,N_3134);
xnor U3172 (N_3172,N_3072,N_3047);
xor U3173 (N_3173,N_3114,N_3055);
or U3174 (N_3174,N_3092,N_3053);
nand U3175 (N_3175,N_3073,N_3075);
xor U3176 (N_3176,N_3129,N_3105);
nand U3177 (N_3177,N_3142,N_3024);
xor U3178 (N_3178,N_3111,N_3032);
xnor U3179 (N_3179,N_3074,N_3004);
xnor U3180 (N_3180,N_3025,N_3100);
xnor U3181 (N_3181,N_3141,N_3016);
and U3182 (N_3182,N_3112,N_3062);
nor U3183 (N_3183,N_3006,N_3148);
and U3184 (N_3184,N_3108,N_3043);
xnor U3185 (N_3185,N_3068,N_3103);
and U3186 (N_3186,N_3138,N_3084);
nand U3187 (N_3187,N_3106,N_3017);
or U3188 (N_3188,N_3125,N_3118);
nor U3189 (N_3189,N_3104,N_3051);
nor U3190 (N_3190,N_3082,N_3132);
or U3191 (N_3191,N_3085,N_3013);
nand U3192 (N_3192,N_3109,N_3059);
nand U3193 (N_3193,N_3128,N_3000);
or U3194 (N_3194,N_3076,N_3137);
or U3195 (N_3195,N_3003,N_3066);
and U3196 (N_3196,N_3095,N_3033);
and U3197 (N_3197,N_3127,N_3040);
nand U3198 (N_3198,N_3061,N_3122);
and U3199 (N_3199,N_3005,N_3119);
and U3200 (N_3200,N_3099,N_3140);
nor U3201 (N_3201,N_3090,N_3081);
nand U3202 (N_3202,N_3079,N_3146);
and U3203 (N_3203,N_3145,N_3065);
nor U3204 (N_3204,N_3054,N_3126);
nand U3205 (N_3205,N_3021,N_3038);
nand U3206 (N_3206,N_3030,N_3049);
nand U3207 (N_3207,N_3045,N_3088);
or U3208 (N_3208,N_3147,N_3149);
xor U3209 (N_3209,N_3096,N_3042);
nand U3210 (N_3210,N_3113,N_3002);
or U3211 (N_3211,N_3086,N_3115);
or U3212 (N_3212,N_3078,N_3046);
or U3213 (N_3213,N_3123,N_3063);
and U3214 (N_3214,N_3026,N_3011);
nand U3215 (N_3215,N_3044,N_3143);
xnor U3216 (N_3216,N_3121,N_3036);
nor U3217 (N_3217,N_3094,N_3080);
nor U3218 (N_3218,N_3050,N_3035);
xor U3219 (N_3219,N_3020,N_3139);
and U3220 (N_3220,N_3131,N_3107);
nand U3221 (N_3221,N_3135,N_3058);
and U3222 (N_3222,N_3048,N_3110);
nand U3223 (N_3223,N_3023,N_3087);
and U3224 (N_3224,N_3014,N_3008);
xnor U3225 (N_3225,N_3030,N_3000);
and U3226 (N_3226,N_3084,N_3093);
xnor U3227 (N_3227,N_3066,N_3136);
nand U3228 (N_3228,N_3003,N_3123);
nand U3229 (N_3229,N_3081,N_3093);
or U3230 (N_3230,N_3088,N_3012);
xnor U3231 (N_3231,N_3026,N_3056);
nor U3232 (N_3232,N_3014,N_3129);
nor U3233 (N_3233,N_3103,N_3073);
xnor U3234 (N_3234,N_3134,N_3097);
nor U3235 (N_3235,N_3023,N_3038);
nor U3236 (N_3236,N_3086,N_3082);
or U3237 (N_3237,N_3030,N_3062);
and U3238 (N_3238,N_3077,N_3047);
nand U3239 (N_3239,N_3040,N_3081);
nor U3240 (N_3240,N_3125,N_3093);
nor U3241 (N_3241,N_3096,N_3043);
or U3242 (N_3242,N_3104,N_3044);
xnor U3243 (N_3243,N_3105,N_3033);
nor U3244 (N_3244,N_3002,N_3054);
or U3245 (N_3245,N_3114,N_3099);
xnor U3246 (N_3246,N_3061,N_3000);
nor U3247 (N_3247,N_3013,N_3020);
xnor U3248 (N_3248,N_3128,N_3031);
or U3249 (N_3249,N_3002,N_3130);
nor U3250 (N_3250,N_3124,N_3131);
xnor U3251 (N_3251,N_3117,N_3020);
xnor U3252 (N_3252,N_3139,N_3080);
xor U3253 (N_3253,N_3133,N_3066);
and U3254 (N_3254,N_3099,N_3145);
or U3255 (N_3255,N_3072,N_3011);
and U3256 (N_3256,N_3026,N_3100);
nand U3257 (N_3257,N_3112,N_3109);
and U3258 (N_3258,N_3067,N_3129);
xor U3259 (N_3259,N_3035,N_3026);
nand U3260 (N_3260,N_3103,N_3115);
nor U3261 (N_3261,N_3121,N_3142);
nor U3262 (N_3262,N_3096,N_3021);
or U3263 (N_3263,N_3119,N_3093);
nor U3264 (N_3264,N_3105,N_3006);
nand U3265 (N_3265,N_3032,N_3057);
xnor U3266 (N_3266,N_3062,N_3045);
and U3267 (N_3267,N_3086,N_3027);
nand U3268 (N_3268,N_3016,N_3012);
and U3269 (N_3269,N_3006,N_3080);
nor U3270 (N_3270,N_3000,N_3063);
xor U3271 (N_3271,N_3072,N_3121);
xor U3272 (N_3272,N_3025,N_3072);
or U3273 (N_3273,N_3117,N_3005);
or U3274 (N_3274,N_3096,N_3102);
or U3275 (N_3275,N_3048,N_3059);
or U3276 (N_3276,N_3149,N_3120);
nand U3277 (N_3277,N_3073,N_3049);
or U3278 (N_3278,N_3075,N_3144);
nand U3279 (N_3279,N_3143,N_3123);
nor U3280 (N_3280,N_3135,N_3136);
xnor U3281 (N_3281,N_3037,N_3016);
xnor U3282 (N_3282,N_3079,N_3125);
nor U3283 (N_3283,N_3051,N_3082);
xnor U3284 (N_3284,N_3105,N_3076);
nand U3285 (N_3285,N_3132,N_3079);
or U3286 (N_3286,N_3037,N_3142);
nand U3287 (N_3287,N_3047,N_3073);
or U3288 (N_3288,N_3045,N_3013);
or U3289 (N_3289,N_3018,N_3122);
nor U3290 (N_3290,N_3133,N_3028);
xnor U3291 (N_3291,N_3116,N_3108);
nor U3292 (N_3292,N_3105,N_3059);
and U3293 (N_3293,N_3090,N_3023);
nor U3294 (N_3294,N_3116,N_3027);
xnor U3295 (N_3295,N_3084,N_3035);
nand U3296 (N_3296,N_3069,N_3040);
nand U3297 (N_3297,N_3100,N_3139);
or U3298 (N_3298,N_3109,N_3061);
nand U3299 (N_3299,N_3119,N_3114);
nand U3300 (N_3300,N_3295,N_3273);
nand U3301 (N_3301,N_3160,N_3233);
and U3302 (N_3302,N_3249,N_3262);
xor U3303 (N_3303,N_3226,N_3252);
nand U3304 (N_3304,N_3247,N_3168);
nand U3305 (N_3305,N_3250,N_3162);
xor U3306 (N_3306,N_3155,N_3152);
nand U3307 (N_3307,N_3203,N_3170);
nor U3308 (N_3308,N_3253,N_3171);
nor U3309 (N_3309,N_3241,N_3198);
nand U3310 (N_3310,N_3150,N_3298);
or U3311 (N_3311,N_3165,N_3275);
nand U3312 (N_3312,N_3191,N_3270);
nand U3313 (N_3313,N_3258,N_3176);
and U3314 (N_3314,N_3267,N_3281);
nand U3315 (N_3315,N_3246,N_3158);
nor U3316 (N_3316,N_3180,N_3172);
and U3317 (N_3317,N_3210,N_3166);
xor U3318 (N_3318,N_3290,N_3257);
or U3319 (N_3319,N_3208,N_3167);
nor U3320 (N_3320,N_3214,N_3201);
or U3321 (N_3321,N_3260,N_3263);
nand U3322 (N_3322,N_3286,N_3211);
and U3323 (N_3323,N_3224,N_3195);
or U3324 (N_3324,N_3175,N_3159);
nand U3325 (N_3325,N_3245,N_3264);
nor U3326 (N_3326,N_3268,N_3261);
xnor U3327 (N_3327,N_3242,N_3219);
xor U3328 (N_3328,N_3157,N_3153);
nand U3329 (N_3329,N_3197,N_3154);
nor U3330 (N_3330,N_3280,N_3234);
xor U3331 (N_3331,N_3240,N_3255);
and U3332 (N_3332,N_3182,N_3248);
or U3333 (N_3333,N_3244,N_3187);
nor U3334 (N_3334,N_3277,N_3215);
xor U3335 (N_3335,N_3254,N_3266);
xor U3336 (N_3336,N_3185,N_3186);
nor U3337 (N_3337,N_3194,N_3289);
xnor U3338 (N_3338,N_3222,N_3299);
or U3339 (N_3339,N_3256,N_3189);
or U3340 (N_3340,N_3223,N_3232);
nand U3341 (N_3341,N_3265,N_3284);
nand U3342 (N_3342,N_3274,N_3251);
xnor U3343 (N_3343,N_3200,N_3163);
or U3344 (N_3344,N_3243,N_3237);
nand U3345 (N_3345,N_3183,N_3178);
xnor U3346 (N_3346,N_3156,N_3294);
xor U3347 (N_3347,N_3221,N_3213);
xor U3348 (N_3348,N_3207,N_3282);
or U3349 (N_3349,N_3283,N_3225);
nor U3350 (N_3350,N_3174,N_3239);
or U3351 (N_3351,N_3271,N_3164);
nor U3352 (N_3352,N_3230,N_3204);
xnor U3353 (N_3353,N_3196,N_3292);
xnor U3354 (N_3354,N_3217,N_3276);
xor U3355 (N_3355,N_3269,N_3288);
and U3356 (N_3356,N_3272,N_3199);
nor U3357 (N_3357,N_3216,N_3179);
nor U3358 (N_3358,N_3293,N_3188);
nand U3359 (N_3359,N_3190,N_3231);
and U3360 (N_3360,N_3184,N_3259);
or U3361 (N_3361,N_3151,N_3218);
xor U3362 (N_3362,N_3181,N_3287);
xnor U3363 (N_3363,N_3202,N_3209);
and U3364 (N_3364,N_3235,N_3161);
nand U3365 (N_3365,N_3220,N_3205);
nand U3366 (N_3366,N_3229,N_3192);
and U3367 (N_3367,N_3238,N_3296);
nand U3368 (N_3368,N_3291,N_3193);
or U3369 (N_3369,N_3285,N_3278);
nand U3370 (N_3370,N_3297,N_3228);
or U3371 (N_3371,N_3279,N_3206);
nor U3372 (N_3372,N_3227,N_3212);
or U3373 (N_3373,N_3177,N_3169);
and U3374 (N_3374,N_3173,N_3236);
xor U3375 (N_3375,N_3167,N_3292);
nor U3376 (N_3376,N_3230,N_3167);
xnor U3377 (N_3377,N_3153,N_3284);
nor U3378 (N_3378,N_3224,N_3285);
nor U3379 (N_3379,N_3158,N_3279);
nor U3380 (N_3380,N_3193,N_3239);
or U3381 (N_3381,N_3220,N_3181);
nand U3382 (N_3382,N_3207,N_3276);
and U3383 (N_3383,N_3214,N_3184);
xor U3384 (N_3384,N_3283,N_3255);
nand U3385 (N_3385,N_3288,N_3159);
and U3386 (N_3386,N_3231,N_3258);
xnor U3387 (N_3387,N_3232,N_3247);
xnor U3388 (N_3388,N_3228,N_3247);
and U3389 (N_3389,N_3297,N_3251);
nor U3390 (N_3390,N_3291,N_3204);
or U3391 (N_3391,N_3165,N_3244);
nand U3392 (N_3392,N_3182,N_3225);
xnor U3393 (N_3393,N_3151,N_3295);
or U3394 (N_3394,N_3220,N_3226);
or U3395 (N_3395,N_3275,N_3152);
nor U3396 (N_3396,N_3163,N_3256);
nor U3397 (N_3397,N_3251,N_3188);
nand U3398 (N_3398,N_3187,N_3295);
and U3399 (N_3399,N_3265,N_3199);
nand U3400 (N_3400,N_3186,N_3275);
xor U3401 (N_3401,N_3236,N_3256);
nor U3402 (N_3402,N_3223,N_3278);
xor U3403 (N_3403,N_3200,N_3204);
and U3404 (N_3404,N_3230,N_3181);
xor U3405 (N_3405,N_3268,N_3154);
nand U3406 (N_3406,N_3201,N_3283);
nand U3407 (N_3407,N_3199,N_3158);
xnor U3408 (N_3408,N_3194,N_3222);
nand U3409 (N_3409,N_3252,N_3233);
and U3410 (N_3410,N_3168,N_3283);
nor U3411 (N_3411,N_3174,N_3203);
xnor U3412 (N_3412,N_3287,N_3256);
nand U3413 (N_3413,N_3295,N_3158);
nand U3414 (N_3414,N_3168,N_3286);
or U3415 (N_3415,N_3196,N_3260);
nand U3416 (N_3416,N_3197,N_3183);
xor U3417 (N_3417,N_3208,N_3239);
or U3418 (N_3418,N_3173,N_3294);
nor U3419 (N_3419,N_3257,N_3177);
nor U3420 (N_3420,N_3150,N_3274);
xor U3421 (N_3421,N_3277,N_3200);
nor U3422 (N_3422,N_3205,N_3288);
nor U3423 (N_3423,N_3211,N_3279);
or U3424 (N_3424,N_3150,N_3188);
or U3425 (N_3425,N_3258,N_3171);
xnor U3426 (N_3426,N_3193,N_3168);
nor U3427 (N_3427,N_3291,N_3277);
nor U3428 (N_3428,N_3224,N_3172);
nor U3429 (N_3429,N_3210,N_3245);
or U3430 (N_3430,N_3239,N_3287);
nand U3431 (N_3431,N_3222,N_3294);
or U3432 (N_3432,N_3243,N_3194);
or U3433 (N_3433,N_3265,N_3299);
or U3434 (N_3434,N_3174,N_3295);
nor U3435 (N_3435,N_3194,N_3156);
or U3436 (N_3436,N_3296,N_3170);
and U3437 (N_3437,N_3251,N_3182);
nor U3438 (N_3438,N_3246,N_3190);
and U3439 (N_3439,N_3270,N_3238);
nand U3440 (N_3440,N_3174,N_3171);
and U3441 (N_3441,N_3262,N_3155);
or U3442 (N_3442,N_3292,N_3176);
nand U3443 (N_3443,N_3217,N_3298);
and U3444 (N_3444,N_3203,N_3181);
xnor U3445 (N_3445,N_3161,N_3176);
nor U3446 (N_3446,N_3291,N_3207);
or U3447 (N_3447,N_3278,N_3156);
and U3448 (N_3448,N_3249,N_3227);
nand U3449 (N_3449,N_3274,N_3237);
nand U3450 (N_3450,N_3373,N_3363);
nand U3451 (N_3451,N_3431,N_3394);
nor U3452 (N_3452,N_3371,N_3445);
nand U3453 (N_3453,N_3393,N_3398);
nand U3454 (N_3454,N_3374,N_3379);
and U3455 (N_3455,N_3355,N_3421);
nor U3456 (N_3456,N_3378,N_3308);
or U3457 (N_3457,N_3361,N_3301);
and U3458 (N_3458,N_3396,N_3399);
or U3459 (N_3459,N_3337,N_3389);
nor U3460 (N_3460,N_3334,N_3365);
xnor U3461 (N_3461,N_3343,N_3325);
or U3462 (N_3462,N_3318,N_3341);
xnor U3463 (N_3463,N_3391,N_3350);
and U3464 (N_3464,N_3364,N_3417);
or U3465 (N_3465,N_3372,N_3369);
or U3466 (N_3466,N_3347,N_3340);
or U3467 (N_3467,N_3446,N_3432);
nor U3468 (N_3468,N_3424,N_3306);
and U3469 (N_3469,N_3412,N_3388);
xnor U3470 (N_3470,N_3336,N_3413);
or U3471 (N_3471,N_3386,N_3332);
and U3472 (N_3472,N_3400,N_3397);
or U3473 (N_3473,N_3305,N_3429);
xor U3474 (N_3474,N_3315,N_3329);
xor U3475 (N_3475,N_3346,N_3444);
or U3476 (N_3476,N_3319,N_3356);
or U3477 (N_3477,N_3426,N_3407);
xnor U3478 (N_3478,N_3404,N_3423);
nand U3479 (N_3479,N_3309,N_3324);
nand U3480 (N_3480,N_3415,N_3302);
and U3481 (N_3481,N_3327,N_3433);
nand U3482 (N_3482,N_3357,N_3442);
nand U3483 (N_3483,N_3408,N_3300);
nor U3484 (N_3484,N_3345,N_3333);
or U3485 (N_3485,N_3360,N_3354);
xor U3486 (N_3486,N_3304,N_3320);
nand U3487 (N_3487,N_3420,N_3339);
nand U3488 (N_3488,N_3367,N_3328);
xnor U3489 (N_3489,N_3335,N_3411);
nand U3490 (N_3490,N_3395,N_3321);
xnor U3491 (N_3491,N_3348,N_3448);
nand U3492 (N_3492,N_3353,N_3358);
nor U3493 (N_3493,N_3414,N_3323);
xnor U3494 (N_3494,N_3359,N_3385);
nand U3495 (N_3495,N_3436,N_3425);
nand U3496 (N_3496,N_3330,N_3387);
xnor U3497 (N_3497,N_3310,N_3438);
xor U3498 (N_3498,N_3307,N_3349);
and U3499 (N_3499,N_3437,N_3322);
xor U3500 (N_3500,N_3439,N_3427);
xor U3501 (N_3501,N_3410,N_3430);
nor U3502 (N_3502,N_3402,N_3326);
nand U3503 (N_3503,N_3383,N_3342);
nand U3504 (N_3504,N_3401,N_3405);
nor U3505 (N_3505,N_3435,N_3380);
nor U3506 (N_3506,N_3312,N_3344);
xor U3507 (N_3507,N_3366,N_3419);
nor U3508 (N_3508,N_3390,N_3418);
nor U3509 (N_3509,N_3409,N_3376);
and U3510 (N_3510,N_3362,N_3311);
or U3511 (N_3511,N_3375,N_3406);
and U3512 (N_3512,N_3441,N_3313);
xor U3513 (N_3513,N_3352,N_3331);
or U3514 (N_3514,N_3370,N_3384);
or U3515 (N_3515,N_3317,N_3447);
nand U3516 (N_3516,N_3449,N_3416);
or U3517 (N_3517,N_3316,N_3303);
and U3518 (N_3518,N_3434,N_3368);
and U3519 (N_3519,N_3314,N_3377);
xnor U3520 (N_3520,N_3392,N_3381);
xor U3521 (N_3521,N_3403,N_3382);
nand U3522 (N_3522,N_3440,N_3351);
and U3523 (N_3523,N_3443,N_3428);
nand U3524 (N_3524,N_3422,N_3338);
xnor U3525 (N_3525,N_3322,N_3343);
xor U3526 (N_3526,N_3340,N_3380);
or U3527 (N_3527,N_3399,N_3344);
xnor U3528 (N_3528,N_3363,N_3369);
nor U3529 (N_3529,N_3407,N_3361);
xnor U3530 (N_3530,N_3379,N_3355);
xor U3531 (N_3531,N_3433,N_3376);
or U3532 (N_3532,N_3381,N_3441);
and U3533 (N_3533,N_3364,N_3437);
or U3534 (N_3534,N_3426,N_3303);
or U3535 (N_3535,N_3352,N_3441);
and U3536 (N_3536,N_3434,N_3396);
nor U3537 (N_3537,N_3374,N_3352);
or U3538 (N_3538,N_3393,N_3356);
nand U3539 (N_3539,N_3360,N_3383);
nor U3540 (N_3540,N_3346,N_3302);
nor U3541 (N_3541,N_3407,N_3317);
nor U3542 (N_3542,N_3384,N_3381);
and U3543 (N_3543,N_3339,N_3390);
nand U3544 (N_3544,N_3409,N_3336);
and U3545 (N_3545,N_3311,N_3337);
xnor U3546 (N_3546,N_3314,N_3368);
nand U3547 (N_3547,N_3431,N_3314);
and U3548 (N_3548,N_3307,N_3447);
nor U3549 (N_3549,N_3304,N_3433);
and U3550 (N_3550,N_3364,N_3337);
xor U3551 (N_3551,N_3367,N_3440);
nor U3552 (N_3552,N_3304,N_3442);
nand U3553 (N_3553,N_3356,N_3376);
nand U3554 (N_3554,N_3401,N_3381);
nor U3555 (N_3555,N_3445,N_3323);
nor U3556 (N_3556,N_3432,N_3404);
or U3557 (N_3557,N_3300,N_3421);
nor U3558 (N_3558,N_3381,N_3410);
or U3559 (N_3559,N_3444,N_3343);
and U3560 (N_3560,N_3389,N_3342);
xor U3561 (N_3561,N_3316,N_3372);
and U3562 (N_3562,N_3322,N_3384);
and U3563 (N_3563,N_3421,N_3315);
and U3564 (N_3564,N_3319,N_3404);
and U3565 (N_3565,N_3414,N_3337);
or U3566 (N_3566,N_3444,N_3389);
nor U3567 (N_3567,N_3327,N_3356);
nor U3568 (N_3568,N_3359,N_3434);
nor U3569 (N_3569,N_3441,N_3347);
and U3570 (N_3570,N_3442,N_3387);
or U3571 (N_3571,N_3415,N_3368);
nand U3572 (N_3572,N_3349,N_3323);
xnor U3573 (N_3573,N_3369,N_3375);
xnor U3574 (N_3574,N_3332,N_3323);
nor U3575 (N_3575,N_3336,N_3374);
or U3576 (N_3576,N_3337,N_3416);
nand U3577 (N_3577,N_3424,N_3440);
xor U3578 (N_3578,N_3354,N_3375);
and U3579 (N_3579,N_3440,N_3427);
or U3580 (N_3580,N_3405,N_3319);
nand U3581 (N_3581,N_3334,N_3345);
and U3582 (N_3582,N_3308,N_3437);
nor U3583 (N_3583,N_3365,N_3423);
nor U3584 (N_3584,N_3315,N_3426);
nor U3585 (N_3585,N_3396,N_3409);
nor U3586 (N_3586,N_3345,N_3428);
nand U3587 (N_3587,N_3321,N_3407);
nor U3588 (N_3588,N_3320,N_3376);
nand U3589 (N_3589,N_3312,N_3410);
nor U3590 (N_3590,N_3391,N_3405);
nor U3591 (N_3591,N_3389,N_3307);
xnor U3592 (N_3592,N_3358,N_3431);
nor U3593 (N_3593,N_3410,N_3440);
nor U3594 (N_3594,N_3315,N_3364);
and U3595 (N_3595,N_3440,N_3392);
nor U3596 (N_3596,N_3331,N_3385);
nor U3597 (N_3597,N_3393,N_3384);
nor U3598 (N_3598,N_3432,N_3319);
nand U3599 (N_3599,N_3361,N_3437);
nor U3600 (N_3600,N_3513,N_3523);
and U3601 (N_3601,N_3508,N_3507);
or U3602 (N_3602,N_3510,N_3572);
or U3603 (N_3603,N_3517,N_3514);
xnor U3604 (N_3604,N_3470,N_3596);
nand U3605 (N_3605,N_3540,N_3575);
xnor U3606 (N_3606,N_3492,N_3546);
or U3607 (N_3607,N_3539,N_3532);
xor U3608 (N_3608,N_3594,N_3469);
and U3609 (N_3609,N_3500,N_3599);
and U3610 (N_3610,N_3473,N_3597);
and U3611 (N_3611,N_3580,N_3561);
xor U3612 (N_3612,N_3495,N_3525);
nor U3613 (N_3613,N_3590,N_3522);
and U3614 (N_3614,N_3544,N_3558);
nor U3615 (N_3615,N_3463,N_3453);
nand U3616 (N_3616,N_3585,N_3550);
xnor U3617 (N_3617,N_3587,N_3545);
xnor U3618 (N_3618,N_3460,N_3511);
and U3619 (N_3619,N_3574,N_3452);
and U3620 (N_3620,N_3551,N_3588);
xnor U3621 (N_3621,N_3466,N_3584);
xnor U3622 (N_3622,N_3455,N_3494);
nand U3623 (N_3623,N_3538,N_3555);
and U3624 (N_3624,N_3484,N_3589);
nor U3625 (N_3625,N_3478,N_3533);
and U3626 (N_3626,N_3553,N_3577);
nand U3627 (N_3627,N_3475,N_3472);
nor U3628 (N_3628,N_3536,N_3465);
or U3629 (N_3629,N_3489,N_3515);
and U3630 (N_3630,N_3526,N_3562);
xor U3631 (N_3631,N_3480,N_3457);
nor U3632 (N_3632,N_3498,N_3481);
xor U3633 (N_3633,N_3506,N_3582);
nand U3634 (N_3634,N_3451,N_3530);
nor U3635 (N_3635,N_3542,N_3598);
and U3636 (N_3636,N_3502,N_3579);
or U3637 (N_3637,N_3456,N_3501);
or U3638 (N_3638,N_3503,N_3578);
nor U3639 (N_3639,N_3459,N_3488);
nor U3640 (N_3640,N_3591,N_3524);
nand U3641 (N_3641,N_3505,N_3583);
xnor U3642 (N_3642,N_3567,N_3581);
xor U3643 (N_3643,N_3563,N_3534);
nand U3644 (N_3644,N_3493,N_3569);
xor U3645 (N_3645,N_3483,N_3593);
nor U3646 (N_3646,N_3471,N_3468);
or U3647 (N_3647,N_3474,N_3477);
xnor U3648 (N_3648,N_3529,N_3499);
xnor U3649 (N_3649,N_3450,N_3541);
nand U3650 (N_3650,N_3566,N_3560);
nand U3651 (N_3651,N_3554,N_3573);
and U3652 (N_3652,N_3504,N_3454);
nand U3653 (N_3653,N_3547,N_3486);
or U3654 (N_3654,N_3535,N_3537);
xor U3655 (N_3655,N_3570,N_3461);
nand U3656 (N_3656,N_3485,N_3592);
and U3657 (N_3657,N_3527,N_3528);
or U3658 (N_3658,N_3496,N_3520);
nand U3659 (N_3659,N_3571,N_3564);
xor U3660 (N_3660,N_3548,N_3519);
and U3661 (N_3661,N_3497,N_3516);
and U3662 (N_3662,N_3462,N_3549);
xor U3663 (N_3663,N_3552,N_3557);
or U3664 (N_3664,N_3482,N_3543);
or U3665 (N_3665,N_3467,N_3595);
or U3666 (N_3666,N_3458,N_3476);
xnor U3667 (N_3667,N_3531,N_3521);
nand U3668 (N_3668,N_3568,N_3479);
or U3669 (N_3669,N_3512,N_3559);
and U3670 (N_3670,N_3491,N_3576);
nor U3671 (N_3671,N_3518,N_3487);
nor U3672 (N_3672,N_3490,N_3565);
xor U3673 (N_3673,N_3586,N_3464);
xnor U3674 (N_3674,N_3556,N_3509);
nand U3675 (N_3675,N_3563,N_3570);
and U3676 (N_3676,N_3461,N_3511);
xor U3677 (N_3677,N_3477,N_3534);
or U3678 (N_3678,N_3455,N_3579);
nor U3679 (N_3679,N_3523,N_3462);
xnor U3680 (N_3680,N_3541,N_3559);
or U3681 (N_3681,N_3569,N_3473);
nand U3682 (N_3682,N_3576,N_3564);
or U3683 (N_3683,N_3467,N_3523);
nor U3684 (N_3684,N_3587,N_3474);
and U3685 (N_3685,N_3473,N_3454);
or U3686 (N_3686,N_3580,N_3539);
xnor U3687 (N_3687,N_3549,N_3574);
or U3688 (N_3688,N_3476,N_3515);
nand U3689 (N_3689,N_3572,N_3539);
nand U3690 (N_3690,N_3542,N_3519);
or U3691 (N_3691,N_3527,N_3465);
nand U3692 (N_3692,N_3526,N_3520);
nor U3693 (N_3693,N_3467,N_3530);
nor U3694 (N_3694,N_3596,N_3487);
and U3695 (N_3695,N_3540,N_3588);
or U3696 (N_3696,N_3480,N_3589);
and U3697 (N_3697,N_3558,N_3559);
nand U3698 (N_3698,N_3561,N_3461);
xor U3699 (N_3699,N_3489,N_3467);
nor U3700 (N_3700,N_3456,N_3580);
xor U3701 (N_3701,N_3520,N_3555);
nor U3702 (N_3702,N_3565,N_3572);
nor U3703 (N_3703,N_3598,N_3505);
nand U3704 (N_3704,N_3555,N_3484);
xnor U3705 (N_3705,N_3465,N_3486);
xnor U3706 (N_3706,N_3538,N_3462);
nor U3707 (N_3707,N_3597,N_3499);
xnor U3708 (N_3708,N_3518,N_3496);
or U3709 (N_3709,N_3561,N_3473);
nand U3710 (N_3710,N_3466,N_3478);
xor U3711 (N_3711,N_3469,N_3569);
nand U3712 (N_3712,N_3565,N_3485);
nand U3713 (N_3713,N_3533,N_3569);
xor U3714 (N_3714,N_3578,N_3536);
nand U3715 (N_3715,N_3470,N_3523);
and U3716 (N_3716,N_3461,N_3574);
xnor U3717 (N_3717,N_3572,N_3462);
xnor U3718 (N_3718,N_3470,N_3457);
and U3719 (N_3719,N_3454,N_3544);
xor U3720 (N_3720,N_3478,N_3551);
nand U3721 (N_3721,N_3535,N_3479);
or U3722 (N_3722,N_3568,N_3538);
xnor U3723 (N_3723,N_3551,N_3523);
nand U3724 (N_3724,N_3485,N_3558);
nor U3725 (N_3725,N_3595,N_3535);
nor U3726 (N_3726,N_3559,N_3587);
nor U3727 (N_3727,N_3494,N_3579);
nor U3728 (N_3728,N_3578,N_3479);
or U3729 (N_3729,N_3452,N_3497);
xnor U3730 (N_3730,N_3480,N_3508);
nand U3731 (N_3731,N_3492,N_3481);
nand U3732 (N_3732,N_3526,N_3560);
nor U3733 (N_3733,N_3506,N_3532);
nor U3734 (N_3734,N_3530,N_3539);
nand U3735 (N_3735,N_3588,N_3563);
nand U3736 (N_3736,N_3546,N_3468);
nor U3737 (N_3737,N_3519,N_3562);
nor U3738 (N_3738,N_3488,N_3512);
and U3739 (N_3739,N_3505,N_3531);
and U3740 (N_3740,N_3500,N_3527);
xnor U3741 (N_3741,N_3509,N_3462);
and U3742 (N_3742,N_3530,N_3498);
nor U3743 (N_3743,N_3547,N_3497);
and U3744 (N_3744,N_3520,N_3530);
nand U3745 (N_3745,N_3476,N_3595);
nand U3746 (N_3746,N_3529,N_3521);
xnor U3747 (N_3747,N_3496,N_3559);
xor U3748 (N_3748,N_3523,N_3538);
nand U3749 (N_3749,N_3553,N_3462);
nor U3750 (N_3750,N_3611,N_3610);
and U3751 (N_3751,N_3604,N_3626);
or U3752 (N_3752,N_3662,N_3699);
nor U3753 (N_3753,N_3726,N_3645);
nor U3754 (N_3754,N_3700,N_3653);
nor U3755 (N_3755,N_3628,N_3693);
or U3756 (N_3756,N_3609,N_3632);
nor U3757 (N_3757,N_3635,N_3740);
nor U3758 (N_3758,N_3607,N_3684);
and U3759 (N_3759,N_3702,N_3728);
nor U3760 (N_3760,N_3741,N_3683);
and U3761 (N_3761,N_3670,N_3660);
and U3762 (N_3762,N_3673,N_3664);
nor U3763 (N_3763,N_3703,N_3633);
nor U3764 (N_3764,N_3727,N_3679);
or U3765 (N_3765,N_3691,N_3682);
nand U3766 (N_3766,N_3712,N_3705);
xor U3767 (N_3767,N_3680,N_3648);
nand U3768 (N_3768,N_3606,N_3644);
nor U3769 (N_3769,N_3643,N_3713);
and U3770 (N_3770,N_3624,N_3636);
or U3771 (N_3771,N_3736,N_3743);
xnor U3772 (N_3772,N_3739,N_3675);
nor U3773 (N_3773,N_3718,N_3689);
nand U3774 (N_3774,N_3646,N_3637);
xnor U3775 (N_3775,N_3711,N_3737);
xnor U3776 (N_3776,N_3733,N_3747);
or U3777 (N_3777,N_3723,N_3735);
xnor U3778 (N_3778,N_3672,N_3627);
and U3779 (N_3779,N_3621,N_3608);
and U3780 (N_3780,N_3663,N_3688);
nor U3781 (N_3781,N_3676,N_3642);
nor U3782 (N_3782,N_3616,N_3707);
and U3783 (N_3783,N_3631,N_3698);
nand U3784 (N_3784,N_3658,N_3701);
nand U3785 (N_3785,N_3744,N_3694);
or U3786 (N_3786,N_3715,N_3629);
xnor U3787 (N_3787,N_3605,N_3685);
nor U3788 (N_3788,N_3746,N_3613);
or U3789 (N_3789,N_3674,N_3710);
xnor U3790 (N_3790,N_3612,N_3615);
nand U3791 (N_3791,N_3742,N_3671);
nor U3792 (N_3792,N_3708,N_3730);
xor U3793 (N_3793,N_3677,N_3668);
or U3794 (N_3794,N_3729,N_3667);
nor U3795 (N_3795,N_3619,N_3652);
xor U3796 (N_3796,N_3654,N_3617);
or U3797 (N_3797,N_3618,N_3602);
xor U3798 (N_3798,N_3650,N_3639);
nor U3799 (N_3799,N_3725,N_3732);
or U3800 (N_3800,N_3620,N_3704);
or U3801 (N_3801,N_3681,N_3669);
nor U3802 (N_3802,N_3656,N_3706);
nor U3803 (N_3803,N_3717,N_3731);
or U3804 (N_3804,N_3745,N_3720);
or U3805 (N_3805,N_3651,N_3666);
xnor U3806 (N_3806,N_3634,N_3665);
xor U3807 (N_3807,N_3600,N_3738);
or U3808 (N_3808,N_3734,N_3709);
nand U3809 (N_3809,N_3696,N_3641);
xor U3810 (N_3810,N_3601,N_3622);
xnor U3811 (N_3811,N_3659,N_3655);
xor U3812 (N_3812,N_3638,N_3647);
xnor U3813 (N_3813,N_3748,N_3603);
nand U3814 (N_3814,N_3687,N_3695);
xnor U3815 (N_3815,N_3678,N_3721);
nand U3816 (N_3816,N_3657,N_3661);
and U3817 (N_3817,N_3716,N_3623);
nor U3818 (N_3818,N_3697,N_3690);
nand U3819 (N_3819,N_3640,N_3724);
nand U3820 (N_3820,N_3692,N_3614);
xor U3821 (N_3821,N_3649,N_3749);
nand U3822 (N_3822,N_3630,N_3719);
or U3823 (N_3823,N_3722,N_3686);
xnor U3824 (N_3824,N_3714,N_3625);
nand U3825 (N_3825,N_3732,N_3645);
nor U3826 (N_3826,N_3710,N_3730);
nor U3827 (N_3827,N_3730,N_3689);
xor U3828 (N_3828,N_3669,N_3718);
or U3829 (N_3829,N_3711,N_3729);
nor U3830 (N_3830,N_3654,N_3703);
or U3831 (N_3831,N_3699,N_3625);
or U3832 (N_3832,N_3733,N_3736);
xor U3833 (N_3833,N_3605,N_3708);
xnor U3834 (N_3834,N_3747,N_3694);
and U3835 (N_3835,N_3729,N_3668);
xnor U3836 (N_3836,N_3668,N_3678);
or U3837 (N_3837,N_3609,N_3641);
and U3838 (N_3838,N_3745,N_3651);
and U3839 (N_3839,N_3608,N_3734);
or U3840 (N_3840,N_3728,N_3705);
or U3841 (N_3841,N_3603,N_3645);
and U3842 (N_3842,N_3738,N_3709);
and U3843 (N_3843,N_3721,N_3694);
nand U3844 (N_3844,N_3609,N_3746);
nor U3845 (N_3845,N_3664,N_3607);
and U3846 (N_3846,N_3655,N_3725);
xor U3847 (N_3847,N_3739,N_3708);
nand U3848 (N_3848,N_3724,N_3721);
nand U3849 (N_3849,N_3688,N_3614);
or U3850 (N_3850,N_3635,N_3620);
nor U3851 (N_3851,N_3648,N_3641);
nand U3852 (N_3852,N_3646,N_3694);
xnor U3853 (N_3853,N_3743,N_3737);
xnor U3854 (N_3854,N_3618,N_3740);
nand U3855 (N_3855,N_3622,N_3658);
nor U3856 (N_3856,N_3746,N_3677);
nor U3857 (N_3857,N_3646,N_3715);
nor U3858 (N_3858,N_3648,N_3677);
or U3859 (N_3859,N_3636,N_3606);
nor U3860 (N_3860,N_3610,N_3704);
nand U3861 (N_3861,N_3640,N_3658);
nand U3862 (N_3862,N_3615,N_3676);
nand U3863 (N_3863,N_3661,N_3665);
or U3864 (N_3864,N_3690,N_3686);
nor U3865 (N_3865,N_3669,N_3691);
or U3866 (N_3866,N_3668,N_3658);
nand U3867 (N_3867,N_3699,N_3664);
nor U3868 (N_3868,N_3716,N_3608);
nand U3869 (N_3869,N_3624,N_3613);
xor U3870 (N_3870,N_3671,N_3632);
nand U3871 (N_3871,N_3747,N_3651);
or U3872 (N_3872,N_3611,N_3700);
nand U3873 (N_3873,N_3647,N_3614);
nor U3874 (N_3874,N_3648,N_3624);
nor U3875 (N_3875,N_3721,N_3720);
xnor U3876 (N_3876,N_3710,N_3680);
nor U3877 (N_3877,N_3661,N_3725);
nand U3878 (N_3878,N_3728,N_3689);
and U3879 (N_3879,N_3634,N_3675);
or U3880 (N_3880,N_3684,N_3737);
nor U3881 (N_3881,N_3609,N_3731);
and U3882 (N_3882,N_3624,N_3638);
nand U3883 (N_3883,N_3689,N_3680);
and U3884 (N_3884,N_3686,N_3701);
xnor U3885 (N_3885,N_3712,N_3612);
nand U3886 (N_3886,N_3643,N_3619);
and U3887 (N_3887,N_3601,N_3704);
and U3888 (N_3888,N_3616,N_3656);
nor U3889 (N_3889,N_3696,N_3620);
or U3890 (N_3890,N_3685,N_3735);
nor U3891 (N_3891,N_3665,N_3671);
and U3892 (N_3892,N_3694,N_3677);
or U3893 (N_3893,N_3705,N_3684);
nor U3894 (N_3894,N_3687,N_3698);
nand U3895 (N_3895,N_3671,N_3682);
and U3896 (N_3896,N_3621,N_3692);
nor U3897 (N_3897,N_3649,N_3639);
nand U3898 (N_3898,N_3727,N_3685);
or U3899 (N_3899,N_3626,N_3720);
nand U3900 (N_3900,N_3826,N_3894);
nor U3901 (N_3901,N_3807,N_3800);
and U3902 (N_3902,N_3750,N_3886);
nor U3903 (N_3903,N_3898,N_3790);
or U3904 (N_3904,N_3844,N_3855);
nor U3905 (N_3905,N_3821,N_3783);
nor U3906 (N_3906,N_3779,N_3815);
nand U3907 (N_3907,N_3824,N_3873);
nor U3908 (N_3908,N_3848,N_3840);
nand U3909 (N_3909,N_3843,N_3789);
nand U3910 (N_3910,N_3769,N_3860);
nand U3911 (N_3911,N_3835,N_3857);
xnor U3912 (N_3912,N_3775,N_3865);
nor U3913 (N_3913,N_3817,N_3761);
nor U3914 (N_3914,N_3890,N_3877);
and U3915 (N_3915,N_3868,N_3820);
xor U3916 (N_3916,N_3842,N_3794);
nor U3917 (N_3917,N_3893,N_3866);
nand U3918 (N_3918,N_3803,N_3767);
nand U3919 (N_3919,N_3787,N_3812);
xnor U3920 (N_3920,N_3780,N_3762);
nand U3921 (N_3921,N_3793,N_3853);
and U3922 (N_3922,N_3784,N_3798);
and U3923 (N_3923,N_3771,N_3796);
and U3924 (N_3924,N_3872,N_3758);
nand U3925 (N_3925,N_3791,N_3804);
or U3926 (N_3926,N_3862,N_3823);
and U3927 (N_3927,N_3773,N_3786);
nor U3928 (N_3928,N_3753,N_3879);
and U3929 (N_3929,N_3871,N_3788);
xnor U3930 (N_3930,N_3852,N_3792);
nor U3931 (N_3931,N_3795,N_3834);
xor U3932 (N_3932,N_3772,N_3829);
or U3933 (N_3933,N_3822,N_3765);
xor U3934 (N_3934,N_3764,N_3858);
nor U3935 (N_3935,N_3899,N_3774);
xnor U3936 (N_3936,N_3751,N_3869);
nor U3937 (N_3937,N_3854,N_3885);
xnor U3938 (N_3938,N_3799,N_3887);
nand U3939 (N_3939,N_3841,N_3828);
or U3940 (N_3940,N_3859,N_3839);
xnor U3941 (N_3941,N_3838,N_3851);
and U3942 (N_3942,N_3831,N_3837);
and U3943 (N_3943,N_3830,N_3802);
nand U3944 (N_3944,N_3864,N_3760);
xnor U3945 (N_3945,N_3881,N_3832);
nor U3946 (N_3946,N_3870,N_3889);
nand U3947 (N_3947,N_3770,N_3861);
and U3948 (N_3948,N_3827,N_3896);
xor U3949 (N_3949,N_3818,N_3875);
or U3950 (N_3950,N_3846,N_3768);
and U3951 (N_3951,N_3884,N_3797);
xor U3952 (N_3952,N_3776,N_3814);
nand U3953 (N_3953,N_3892,N_3782);
nand U3954 (N_3954,N_3806,N_3809);
xor U3955 (N_3955,N_3863,N_3849);
or U3956 (N_3956,N_3888,N_3867);
or U3957 (N_3957,N_3808,N_3876);
and U3958 (N_3958,N_3757,N_3883);
or U3959 (N_3959,N_3777,N_3816);
xor U3960 (N_3960,N_3759,N_3895);
xnor U3961 (N_3961,N_3874,N_3847);
and U3962 (N_3962,N_3778,N_3891);
or U3963 (N_3963,N_3882,N_3880);
or U3964 (N_3964,N_3825,N_3755);
and U3965 (N_3965,N_3781,N_3819);
nand U3966 (N_3966,N_3752,N_3766);
and U3967 (N_3967,N_3805,N_3833);
and U3968 (N_3968,N_3785,N_3763);
nor U3969 (N_3969,N_3850,N_3897);
nor U3970 (N_3970,N_3754,N_3813);
or U3971 (N_3971,N_3810,N_3836);
and U3972 (N_3972,N_3811,N_3756);
or U3973 (N_3973,N_3845,N_3878);
nand U3974 (N_3974,N_3856,N_3801);
xor U3975 (N_3975,N_3802,N_3838);
nand U3976 (N_3976,N_3794,N_3852);
nand U3977 (N_3977,N_3836,N_3772);
nor U3978 (N_3978,N_3831,N_3795);
and U3979 (N_3979,N_3801,N_3839);
nand U3980 (N_3980,N_3887,N_3853);
nor U3981 (N_3981,N_3769,N_3893);
xor U3982 (N_3982,N_3799,N_3894);
nand U3983 (N_3983,N_3759,N_3757);
nor U3984 (N_3984,N_3850,N_3846);
and U3985 (N_3985,N_3807,N_3757);
nand U3986 (N_3986,N_3819,N_3751);
and U3987 (N_3987,N_3798,N_3777);
or U3988 (N_3988,N_3812,N_3803);
nor U3989 (N_3989,N_3776,N_3791);
nand U3990 (N_3990,N_3822,N_3760);
nor U3991 (N_3991,N_3757,N_3787);
and U3992 (N_3992,N_3801,N_3798);
xnor U3993 (N_3993,N_3812,N_3773);
xnor U3994 (N_3994,N_3762,N_3865);
and U3995 (N_3995,N_3845,N_3871);
and U3996 (N_3996,N_3885,N_3893);
nor U3997 (N_3997,N_3851,N_3773);
xnor U3998 (N_3998,N_3758,N_3888);
and U3999 (N_3999,N_3885,N_3768);
and U4000 (N_4000,N_3858,N_3769);
or U4001 (N_4001,N_3876,N_3769);
and U4002 (N_4002,N_3751,N_3784);
nand U4003 (N_4003,N_3763,N_3879);
xnor U4004 (N_4004,N_3890,N_3855);
nand U4005 (N_4005,N_3848,N_3839);
and U4006 (N_4006,N_3789,N_3792);
xnor U4007 (N_4007,N_3809,N_3885);
and U4008 (N_4008,N_3754,N_3824);
and U4009 (N_4009,N_3802,N_3839);
and U4010 (N_4010,N_3854,N_3824);
nor U4011 (N_4011,N_3894,N_3807);
xor U4012 (N_4012,N_3899,N_3877);
xor U4013 (N_4013,N_3875,N_3846);
and U4014 (N_4014,N_3884,N_3808);
nor U4015 (N_4015,N_3870,N_3768);
and U4016 (N_4016,N_3770,N_3788);
nor U4017 (N_4017,N_3796,N_3844);
and U4018 (N_4018,N_3893,N_3873);
or U4019 (N_4019,N_3769,N_3821);
and U4020 (N_4020,N_3896,N_3856);
nor U4021 (N_4021,N_3873,N_3774);
nor U4022 (N_4022,N_3773,N_3839);
xor U4023 (N_4023,N_3786,N_3885);
nand U4024 (N_4024,N_3754,N_3868);
and U4025 (N_4025,N_3896,N_3789);
and U4026 (N_4026,N_3796,N_3787);
or U4027 (N_4027,N_3894,N_3781);
nand U4028 (N_4028,N_3875,N_3866);
xor U4029 (N_4029,N_3893,N_3855);
xnor U4030 (N_4030,N_3835,N_3763);
nor U4031 (N_4031,N_3796,N_3850);
xnor U4032 (N_4032,N_3780,N_3819);
or U4033 (N_4033,N_3816,N_3757);
xnor U4034 (N_4034,N_3806,N_3857);
nor U4035 (N_4035,N_3853,N_3768);
and U4036 (N_4036,N_3891,N_3838);
nor U4037 (N_4037,N_3815,N_3836);
or U4038 (N_4038,N_3842,N_3895);
nor U4039 (N_4039,N_3759,N_3756);
xor U4040 (N_4040,N_3862,N_3877);
nor U4041 (N_4041,N_3856,N_3805);
xor U4042 (N_4042,N_3825,N_3859);
and U4043 (N_4043,N_3761,N_3865);
nor U4044 (N_4044,N_3784,N_3838);
nand U4045 (N_4045,N_3750,N_3821);
nand U4046 (N_4046,N_3889,N_3886);
or U4047 (N_4047,N_3875,N_3826);
and U4048 (N_4048,N_3885,N_3819);
and U4049 (N_4049,N_3830,N_3899);
nand U4050 (N_4050,N_4038,N_3978);
xnor U4051 (N_4051,N_3944,N_4008);
xor U4052 (N_4052,N_3901,N_4010);
and U4053 (N_4053,N_3951,N_3927);
or U4054 (N_4054,N_4042,N_3926);
and U4055 (N_4055,N_4029,N_4030);
or U4056 (N_4056,N_3914,N_3957);
and U4057 (N_4057,N_3938,N_3904);
nand U4058 (N_4058,N_4016,N_3939);
or U4059 (N_4059,N_3965,N_4046);
nand U4060 (N_4060,N_3994,N_3913);
or U4061 (N_4061,N_3910,N_4031);
or U4062 (N_4062,N_3915,N_4025);
nor U4063 (N_4063,N_4026,N_3993);
nor U4064 (N_4064,N_3931,N_4036);
nor U4065 (N_4065,N_3967,N_3902);
and U4066 (N_4066,N_3980,N_3934);
xor U4067 (N_4067,N_3937,N_3973);
xnor U4068 (N_4068,N_4034,N_3961);
xor U4069 (N_4069,N_4019,N_4028);
and U4070 (N_4070,N_3903,N_4023);
nand U4071 (N_4071,N_3974,N_3943);
nand U4072 (N_4072,N_3921,N_3985);
nor U4073 (N_4073,N_4006,N_3955);
nor U4074 (N_4074,N_3996,N_3930);
or U4075 (N_4075,N_4040,N_3979);
or U4076 (N_4076,N_3960,N_3975);
and U4077 (N_4077,N_4000,N_4011);
nor U4078 (N_4078,N_4001,N_3919);
nand U4079 (N_4079,N_3909,N_4027);
or U4080 (N_4080,N_3918,N_3940);
and U4081 (N_4081,N_3995,N_4039);
or U4082 (N_4082,N_3959,N_3947);
nand U4083 (N_4083,N_3968,N_3917);
nand U4084 (N_4084,N_4024,N_3999);
or U4085 (N_4085,N_4022,N_3923);
or U4086 (N_4086,N_3932,N_3977);
or U4087 (N_4087,N_3956,N_3964);
xnor U4088 (N_4088,N_4045,N_3976);
nand U4089 (N_4089,N_3916,N_3941);
nand U4090 (N_4090,N_4033,N_3986);
or U4091 (N_4091,N_3952,N_3922);
nor U4092 (N_4092,N_3990,N_3998);
or U4093 (N_4093,N_4048,N_4004);
nand U4094 (N_4094,N_3935,N_3971);
or U4095 (N_4095,N_4032,N_3950);
and U4096 (N_4096,N_3911,N_3963);
or U4097 (N_4097,N_3908,N_4005);
xnor U4098 (N_4098,N_3946,N_4014);
or U4099 (N_4099,N_3970,N_4003);
nor U4100 (N_4100,N_4015,N_3953);
or U4101 (N_4101,N_3962,N_3987);
nor U4102 (N_4102,N_4020,N_3988);
nor U4103 (N_4103,N_3905,N_3958);
xnor U4104 (N_4104,N_4049,N_3949);
or U4105 (N_4105,N_4021,N_3912);
nand U4106 (N_4106,N_3969,N_3991);
and U4107 (N_4107,N_3906,N_4018);
xnor U4108 (N_4108,N_4035,N_4013);
nand U4109 (N_4109,N_3983,N_3925);
nand U4110 (N_4110,N_3945,N_3982);
nand U4111 (N_4111,N_3954,N_3948);
xor U4112 (N_4112,N_4012,N_3972);
xnor U4113 (N_4113,N_3992,N_3966);
xnor U4114 (N_4114,N_4037,N_3981);
xnor U4115 (N_4115,N_4017,N_3924);
or U4116 (N_4116,N_3936,N_4044);
and U4117 (N_4117,N_3920,N_3942);
nand U4118 (N_4118,N_4002,N_3907);
xor U4119 (N_4119,N_4007,N_4009);
nor U4120 (N_4120,N_3933,N_3900);
nand U4121 (N_4121,N_3984,N_3928);
nand U4122 (N_4122,N_3929,N_4043);
xor U4123 (N_4123,N_3989,N_3997);
or U4124 (N_4124,N_4041,N_4047);
or U4125 (N_4125,N_4030,N_3928);
and U4126 (N_4126,N_4049,N_3935);
or U4127 (N_4127,N_4023,N_4025);
nand U4128 (N_4128,N_3902,N_3917);
nand U4129 (N_4129,N_4009,N_3908);
or U4130 (N_4130,N_3932,N_3987);
xnor U4131 (N_4131,N_3933,N_3948);
and U4132 (N_4132,N_3937,N_3907);
nand U4133 (N_4133,N_3908,N_3936);
and U4134 (N_4134,N_3951,N_3911);
nand U4135 (N_4135,N_3955,N_3972);
or U4136 (N_4136,N_3986,N_4022);
nor U4137 (N_4137,N_3929,N_3940);
nand U4138 (N_4138,N_4026,N_4018);
nor U4139 (N_4139,N_4022,N_3971);
xnor U4140 (N_4140,N_3997,N_4036);
nor U4141 (N_4141,N_3917,N_4004);
nand U4142 (N_4142,N_3995,N_3941);
nand U4143 (N_4143,N_3943,N_3978);
and U4144 (N_4144,N_3944,N_3913);
nand U4145 (N_4145,N_3974,N_3973);
nor U4146 (N_4146,N_4021,N_4035);
xnor U4147 (N_4147,N_4011,N_3988);
nand U4148 (N_4148,N_3970,N_3971);
nand U4149 (N_4149,N_3953,N_3966);
or U4150 (N_4150,N_4006,N_3940);
or U4151 (N_4151,N_3973,N_4024);
nand U4152 (N_4152,N_3901,N_3916);
and U4153 (N_4153,N_3969,N_4038);
and U4154 (N_4154,N_3984,N_4036);
or U4155 (N_4155,N_4049,N_3994);
nor U4156 (N_4156,N_3946,N_3906);
and U4157 (N_4157,N_3964,N_3993);
nand U4158 (N_4158,N_3929,N_4002);
nand U4159 (N_4159,N_3948,N_3965);
and U4160 (N_4160,N_3912,N_3994);
nor U4161 (N_4161,N_3960,N_3900);
or U4162 (N_4162,N_3965,N_3973);
xor U4163 (N_4163,N_3945,N_3987);
nand U4164 (N_4164,N_3938,N_3928);
xor U4165 (N_4165,N_4022,N_4008);
or U4166 (N_4166,N_3913,N_3917);
nor U4167 (N_4167,N_3938,N_3970);
nand U4168 (N_4168,N_3902,N_3903);
or U4169 (N_4169,N_3909,N_4006);
and U4170 (N_4170,N_3963,N_4040);
and U4171 (N_4171,N_4041,N_3948);
nand U4172 (N_4172,N_3981,N_4031);
xor U4173 (N_4173,N_3972,N_3940);
xnor U4174 (N_4174,N_3949,N_4045);
and U4175 (N_4175,N_4011,N_3968);
nor U4176 (N_4176,N_3927,N_4017);
xor U4177 (N_4177,N_3918,N_3923);
nor U4178 (N_4178,N_4020,N_3951);
and U4179 (N_4179,N_3920,N_3962);
nand U4180 (N_4180,N_3970,N_3912);
nand U4181 (N_4181,N_3986,N_4005);
or U4182 (N_4182,N_3967,N_4027);
and U4183 (N_4183,N_3915,N_3943);
xnor U4184 (N_4184,N_3925,N_3936);
xor U4185 (N_4185,N_3948,N_3972);
and U4186 (N_4186,N_3999,N_3987);
nand U4187 (N_4187,N_3950,N_3942);
and U4188 (N_4188,N_4021,N_3934);
or U4189 (N_4189,N_4046,N_4017);
nand U4190 (N_4190,N_3904,N_3942);
nor U4191 (N_4191,N_3910,N_3913);
or U4192 (N_4192,N_3962,N_3937);
or U4193 (N_4193,N_4025,N_3946);
nor U4194 (N_4194,N_3941,N_3988);
and U4195 (N_4195,N_3969,N_3999);
xnor U4196 (N_4196,N_4025,N_3975);
or U4197 (N_4197,N_3988,N_3927);
and U4198 (N_4198,N_4030,N_4036);
nand U4199 (N_4199,N_3980,N_3936);
nor U4200 (N_4200,N_4085,N_4181);
and U4201 (N_4201,N_4099,N_4132);
and U4202 (N_4202,N_4101,N_4195);
nand U4203 (N_4203,N_4112,N_4164);
or U4204 (N_4204,N_4148,N_4091);
and U4205 (N_4205,N_4069,N_4051);
nand U4206 (N_4206,N_4157,N_4086);
and U4207 (N_4207,N_4113,N_4060);
or U4208 (N_4208,N_4054,N_4131);
and U4209 (N_4209,N_4065,N_4122);
nor U4210 (N_4210,N_4196,N_4116);
or U4211 (N_4211,N_4104,N_4100);
nand U4212 (N_4212,N_4120,N_4180);
nor U4213 (N_4213,N_4178,N_4079);
or U4214 (N_4214,N_4059,N_4152);
and U4215 (N_4215,N_4076,N_4078);
nand U4216 (N_4216,N_4055,N_4185);
nor U4217 (N_4217,N_4139,N_4172);
nand U4218 (N_4218,N_4124,N_4056);
nor U4219 (N_4219,N_4128,N_4066);
or U4220 (N_4220,N_4143,N_4098);
or U4221 (N_4221,N_4198,N_4192);
or U4222 (N_4222,N_4077,N_4161);
nor U4223 (N_4223,N_4105,N_4096);
or U4224 (N_4224,N_4163,N_4074);
and U4225 (N_4225,N_4133,N_4063);
or U4226 (N_4226,N_4165,N_4150);
nand U4227 (N_4227,N_4186,N_4193);
and U4228 (N_4228,N_4169,N_4071);
nor U4229 (N_4229,N_4188,N_4061);
nand U4230 (N_4230,N_4121,N_4092);
or U4231 (N_4231,N_4068,N_4166);
nor U4232 (N_4232,N_4126,N_4097);
and U4233 (N_4233,N_4087,N_4108);
nor U4234 (N_4234,N_4050,N_4134);
xnor U4235 (N_4235,N_4135,N_4095);
xor U4236 (N_4236,N_4072,N_4111);
or U4237 (N_4237,N_4197,N_4147);
and U4238 (N_4238,N_4138,N_4117);
nand U4239 (N_4239,N_4094,N_4146);
nand U4240 (N_4240,N_4189,N_4083);
xnor U4241 (N_4241,N_4142,N_4158);
and U4242 (N_4242,N_4114,N_4168);
xor U4243 (N_4243,N_4154,N_4140);
xor U4244 (N_4244,N_4123,N_4171);
nand U4245 (N_4245,N_4102,N_4129);
or U4246 (N_4246,N_4137,N_4183);
xnor U4247 (N_4247,N_4106,N_4151);
nor U4248 (N_4248,N_4075,N_4194);
xor U4249 (N_4249,N_4073,N_4080);
nand U4250 (N_4250,N_4190,N_4081);
and U4251 (N_4251,N_4082,N_4176);
nor U4252 (N_4252,N_4107,N_4052);
or U4253 (N_4253,N_4115,N_4103);
nand U4254 (N_4254,N_4199,N_4093);
or U4255 (N_4255,N_4118,N_4182);
xnor U4256 (N_4256,N_4173,N_4184);
nand U4257 (N_4257,N_4090,N_4175);
xnor U4258 (N_4258,N_4159,N_4067);
xor U4259 (N_4259,N_4153,N_4089);
nand U4260 (N_4260,N_4155,N_4084);
nor U4261 (N_4261,N_4170,N_4191);
or U4262 (N_4262,N_4070,N_4064);
nor U4263 (N_4263,N_4088,N_4058);
xnor U4264 (N_4264,N_4177,N_4062);
or U4265 (N_4265,N_4149,N_4145);
xnor U4266 (N_4266,N_4130,N_4174);
nand U4267 (N_4267,N_4109,N_4110);
xor U4268 (N_4268,N_4167,N_4162);
xor U4269 (N_4269,N_4053,N_4119);
and U4270 (N_4270,N_4127,N_4160);
nand U4271 (N_4271,N_4179,N_4141);
nor U4272 (N_4272,N_4144,N_4156);
nand U4273 (N_4273,N_4187,N_4057);
and U4274 (N_4274,N_4136,N_4125);
xor U4275 (N_4275,N_4064,N_4156);
nor U4276 (N_4276,N_4068,N_4194);
xnor U4277 (N_4277,N_4158,N_4133);
xor U4278 (N_4278,N_4161,N_4131);
nor U4279 (N_4279,N_4155,N_4090);
and U4280 (N_4280,N_4056,N_4135);
nand U4281 (N_4281,N_4065,N_4103);
xor U4282 (N_4282,N_4122,N_4194);
and U4283 (N_4283,N_4119,N_4166);
nor U4284 (N_4284,N_4105,N_4153);
xor U4285 (N_4285,N_4168,N_4071);
and U4286 (N_4286,N_4138,N_4070);
nor U4287 (N_4287,N_4178,N_4194);
nand U4288 (N_4288,N_4173,N_4118);
nand U4289 (N_4289,N_4116,N_4056);
nand U4290 (N_4290,N_4108,N_4130);
nand U4291 (N_4291,N_4127,N_4076);
or U4292 (N_4292,N_4063,N_4139);
xnor U4293 (N_4293,N_4164,N_4087);
nand U4294 (N_4294,N_4158,N_4170);
xor U4295 (N_4295,N_4083,N_4057);
xor U4296 (N_4296,N_4194,N_4088);
nor U4297 (N_4297,N_4189,N_4106);
xnor U4298 (N_4298,N_4106,N_4054);
nor U4299 (N_4299,N_4142,N_4098);
nor U4300 (N_4300,N_4066,N_4093);
or U4301 (N_4301,N_4055,N_4097);
nor U4302 (N_4302,N_4177,N_4050);
and U4303 (N_4303,N_4155,N_4167);
and U4304 (N_4304,N_4141,N_4166);
or U4305 (N_4305,N_4175,N_4104);
nor U4306 (N_4306,N_4073,N_4195);
xor U4307 (N_4307,N_4102,N_4101);
or U4308 (N_4308,N_4076,N_4110);
nand U4309 (N_4309,N_4195,N_4187);
and U4310 (N_4310,N_4087,N_4083);
nor U4311 (N_4311,N_4104,N_4053);
nor U4312 (N_4312,N_4134,N_4092);
nand U4313 (N_4313,N_4197,N_4066);
nand U4314 (N_4314,N_4199,N_4164);
or U4315 (N_4315,N_4189,N_4102);
nor U4316 (N_4316,N_4163,N_4054);
xor U4317 (N_4317,N_4164,N_4151);
nand U4318 (N_4318,N_4145,N_4184);
or U4319 (N_4319,N_4093,N_4172);
nor U4320 (N_4320,N_4106,N_4141);
and U4321 (N_4321,N_4068,N_4111);
nand U4322 (N_4322,N_4072,N_4196);
nand U4323 (N_4323,N_4090,N_4058);
nand U4324 (N_4324,N_4064,N_4114);
nor U4325 (N_4325,N_4070,N_4082);
and U4326 (N_4326,N_4136,N_4146);
xnor U4327 (N_4327,N_4113,N_4120);
nand U4328 (N_4328,N_4156,N_4157);
and U4329 (N_4329,N_4105,N_4173);
and U4330 (N_4330,N_4088,N_4121);
xnor U4331 (N_4331,N_4054,N_4076);
nand U4332 (N_4332,N_4050,N_4152);
xor U4333 (N_4333,N_4064,N_4066);
nor U4334 (N_4334,N_4058,N_4057);
or U4335 (N_4335,N_4116,N_4180);
nand U4336 (N_4336,N_4157,N_4063);
nor U4337 (N_4337,N_4170,N_4052);
and U4338 (N_4338,N_4184,N_4085);
or U4339 (N_4339,N_4175,N_4096);
nor U4340 (N_4340,N_4122,N_4172);
nor U4341 (N_4341,N_4126,N_4054);
nor U4342 (N_4342,N_4178,N_4124);
or U4343 (N_4343,N_4102,N_4169);
nand U4344 (N_4344,N_4150,N_4072);
nand U4345 (N_4345,N_4162,N_4073);
xnor U4346 (N_4346,N_4169,N_4131);
nor U4347 (N_4347,N_4112,N_4160);
xnor U4348 (N_4348,N_4053,N_4146);
nor U4349 (N_4349,N_4078,N_4194);
xor U4350 (N_4350,N_4222,N_4344);
nor U4351 (N_4351,N_4237,N_4308);
or U4352 (N_4352,N_4283,N_4260);
and U4353 (N_4353,N_4349,N_4227);
nand U4354 (N_4354,N_4256,N_4317);
xnor U4355 (N_4355,N_4205,N_4300);
xor U4356 (N_4356,N_4266,N_4303);
xnor U4357 (N_4357,N_4299,N_4270);
nor U4358 (N_4358,N_4312,N_4215);
xor U4359 (N_4359,N_4249,N_4319);
or U4360 (N_4360,N_4209,N_4275);
or U4361 (N_4361,N_4278,N_4327);
nor U4362 (N_4362,N_4238,N_4296);
xnor U4363 (N_4363,N_4293,N_4292);
and U4364 (N_4364,N_4304,N_4217);
or U4365 (N_4365,N_4253,N_4247);
and U4366 (N_4366,N_4264,N_4279);
and U4367 (N_4367,N_4347,N_4298);
nor U4368 (N_4368,N_4269,N_4268);
nor U4369 (N_4369,N_4306,N_4335);
xnor U4370 (N_4370,N_4348,N_4332);
or U4371 (N_4371,N_4294,N_4346);
nor U4372 (N_4372,N_4200,N_4250);
nor U4373 (N_4373,N_4305,N_4324);
nand U4374 (N_4374,N_4336,N_4243);
or U4375 (N_4375,N_4328,N_4244);
nor U4376 (N_4376,N_4239,N_4289);
or U4377 (N_4377,N_4221,N_4320);
xor U4378 (N_4378,N_4333,N_4258);
nor U4379 (N_4379,N_4236,N_4257);
nor U4380 (N_4380,N_4214,N_4220);
nor U4381 (N_4381,N_4255,N_4231);
xor U4382 (N_4382,N_4248,N_4267);
nor U4383 (N_4383,N_4234,N_4224);
xnor U4384 (N_4384,N_4254,N_4232);
nor U4385 (N_4385,N_4242,N_4211);
nand U4386 (N_4386,N_4261,N_4233);
xnor U4387 (N_4387,N_4263,N_4338);
or U4388 (N_4388,N_4216,N_4331);
nor U4389 (N_4389,N_4318,N_4301);
or U4390 (N_4390,N_4281,N_4203);
nand U4391 (N_4391,N_4265,N_4210);
xor U4392 (N_4392,N_4310,N_4201);
xnor U4393 (N_4393,N_4235,N_4316);
or U4394 (N_4394,N_4259,N_4213);
xnor U4395 (N_4395,N_4307,N_4291);
nand U4396 (N_4396,N_4315,N_4342);
nor U4397 (N_4397,N_4271,N_4204);
and U4398 (N_4398,N_4326,N_4273);
or U4399 (N_4399,N_4323,N_4219);
nor U4400 (N_4400,N_4309,N_4339);
xor U4401 (N_4401,N_4208,N_4245);
and U4402 (N_4402,N_4314,N_4313);
or U4403 (N_4403,N_4277,N_4311);
and U4404 (N_4404,N_4345,N_4287);
and U4405 (N_4405,N_4262,N_4282);
or U4406 (N_4406,N_4321,N_4290);
xnor U4407 (N_4407,N_4212,N_4202);
nand U4408 (N_4408,N_4274,N_4341);
nor U4409 (N_4409,N_4329,N_4272);
nor U4410 (N_4410,N_4302,N_4285);
and U4411 (N_4411,N_4206,N_4340);
or U4412 (N_4412,N_4228,N_4337);
or U4413 (N_4413,N_4207,N_4330);
and U4414 (N_4414,N_4218,N_4252);
xnor U4415 (N_4415,N_4322,N_4334);
nand U4416 (N_4416,N_4286,N_4223);
nor U4417 (N_4417,N_4225,N_4276);
nor U4418 (N_4418,N_4251,N_4240);
nor U4419 (N_4419,N_4343,N_4226);
nand U4420 (N_4420,N_4229,N_4284);
nand U4421 (N_4421,N_4280,N_4241);
xnor U4422 (N_4422,N_4246,N_4230);
or U4423 (N_4423,N_4288,N_4295);
nor U4424 (N_4424,N_4297,N_4325);
xor U4425 (N_4425,N_4256,N_4284);
xnor U4426 (N_4426,N_4208,N_4252);
or U4427 (N_4427,N_4239,N_4230);
or U4428 (N_4428,N_4304,N_4263);
and U4429 (N_4429,N_4252,N_4249);
xor U4430 (N_4430,N_4300,N_4341);
xor U4431 (N_4431,N_4348,N_4335);
xnor U4432 (N_4432,N_4204,N_4314);
xor U4433 (N_4433,N_4342,N_4318);
xor U4434 (N_4434,N_4307,N_4286);
nor U4435 (N_4435,N_4282,N_4272);
xor U4436 (N_4436,N_4276,N_4269);
and U4437 (N_4437,N_4258,N_4253);
xor U4438 (N_4438,N_4295,N_4274);
nor U4439 (N_4439,N_4338,N_4238);
xnor U4440 (N_4440,N_4225,N_4294);
or U4441 (N_4441,N_4297,N_4333);
nor U4442 (N_4442,N_4214,N_4227);
and U4443 (N_4443,N_4213,N_4301);
and U4444 (N_4444,N_4298,N_4303);
nand U4445 (N_4445,N_4334,N_4286);
and U4446 (N_4446,N_4289,N_4301);
or U4447 (N_4447,N_4310,N_4273);
nor U4448 (N_4448,N_4306,N_4243);
nor U4449 (N_4449,N_4304,N_4265);
nor U4450 (N_4450,N_4314,N_4238);
nand U4451 (N_4451,N_4317,N_4285);
nand U4452 (N_4452,N_4209,N_4241);
nor U4453 (N_4453,N_4223,N_4338);
or U4454 (N_4454,N_4301,N_4315);
or U4455 (N_4455,N_4223,N_4235);
nand U4456 (N_4456,N_4334,N_4342);
nand U4457 (N_4457,N_4302,N_4283);
xnor U4458 (N_4458,N_4230,N_4243);
nand U4459 (N_4459,N_4278,N_4273);
nand U4460 (N_4460,N_4266,N_4269);
xor U4461 (N_4461,N_4200,N_4262);
nand U4462 (N_4462,N_4253,N_4311);
and U4463 (N_4463,N_4310,N_4247);
nand U4464 (N_4464,N_4248,N_4285);
xnor U4465 (N_4465,N_4232,N_4258);
or U4466 (N_4466,N_4306,N_4329);
nor U4467 (N_4467,N_4208,N_4249);
and U4468 (N_4468,N_4265,N_4248);
and U4469 (N_4469,N_4261,N_4223);
or U4470 (N_4470,N_4302,N_4281);
nor U4471 (N_4471,N_4330,N_4280);
and U4472 (N_4472,N_4255,N_4292);
xnor U4473 (N_4473,N_4221,N_4260);
and U4474 (N_4474,N_4333,N_4345);
xnor U4475 (N_4475,N_4328,N_4236);
nand U4476 (N_4476,N_4232,N_4286);
or U4477 (N_4477,N_4274,N_4302);
nor U4478 (N_4478,N_4205,N_4228);
nor U4479 (N_4479,N_4278,N_4330);
or U4480 (N_4480,N_4291,N_4298);
xnor U4481 (N_4481,N_4326,N_4311);
nand U4482 (N_4482,N_4261,N_4285);
nand U4483 (N_4483,N_4224,N_4340);
xor U4484 (N_4484,N_4266,N_4203);
and U4485 (N_4485,N_4298,N_4228);
or U4486 (N_4486,N_4256,N_4282);
nand U4487 (N_4487,N_4312,N_4297);
and U4488 (N_4488,N_4264,N_4221);
and U4489 (N_4489,N_4347,N_4313);
xor U4490 (N_4490,N_4267,N_4256);
and U4491 (N_4491,N_4314,N_4268);
nor U4492 (N_4492,N_4246,N_4293);
or U4493 (N_4493,N_4277,N_4301);
or U4494 (N_4494,N_4337,N_4290);
and U4495 (N_4495,N_4331,N_4234);
nor U4496 (N_4496,N_4221,N_4250);
nor U4497 (N_4497,N_4230,N_4328);
and U4498 (N_4498,N_4272,N_4266);
or U4499 (N_4499,N_4246,N_4224);
nor U4500 (N_4500,N_4442,N_4433);
nor U4501 (N_4501,N_4369,N_4428);
or U4502 (N_4502,N_4461,N_4435);
or U4503 (N_4503,N_4365,N_4464);
or U4504 (N_4504,N_4403,N_4491);
and U4505 (N_4505,N_4391,N_4423);
xnor U4506 (N_4506,N_4380,N_4355);
or U4507 (N_4507,N_4482,N_4456);
and U4508 (N_4508,N_4432,N_4375);
nand U4509 (N_4509,N_4441,N_4420);
nor U4510 (N_4510,N_4379,N_4489);
or U4511 (N_4511,N_4351,N_4473);
and U4512 (N_4512,N_4478,N_4438);
and U4513 (N_4513,N_4469,N_4465);
xor U4514 (N_4514,N_4429,N_4499);
or U4515 (N_4515,N_4356,N_4483);
xnor U4516 (N_4516,N_4400,N_4404);
nor U4517 (N_4517,N_4446,N_4384);
nor U4518 (N_4518,N_4490,N_4470);
xnor U4519 (N_4519,N_4495,N_4454);
and U4520 (N_4520,N_4437,N_4390);
or U4521 (N_4521,N_4460,N_4484);
nor U4522 (N_4522,N_4416,N_4389);
or U4523 (N_4523,N_4417,N_4422);
and U4524 (N_4524,N_4439,N_4350);
xnor U4525 (N_4525,N_4457,N_4409);
and U4526 (N_4526,N_4430,N_4377);
nor U4527 (N_4527,N_4448,N_4436);
nor U4528 (N_4528,N_4421,N_4393);
nand U4529 (N_4529,N_4359,N_4486);
xnor U4530 (N_4530,N_4397,N_4385);
nand U4531 (N_4531,N_4370,N_4405);
nor U4532 (N_4532,N_4362,N_4498);
nor U4533 (N_4533,N_4467,N_4399);
nor U4534 (N_4534,N_4396,N_4364);
nand U4535 (N_4535,N_4466,N_4458);
or U4536 (N_4536,N_4398,N_4361);
and U4537 (N_4537,N_4407,N_4410);
nor U4538 (N_4538,N_4387,N_4418);
xor U4539 (N_4539,N_4443,N_4431);
and U4540 (N_4540,N_4415,N_4367);
or U4541 (N_4541,N_4382,N_4440);
and U4542 (N_4542,N_4494,N_4371);
or U4543 (N_4543,N_4471,N_4474);
or U4544 (N_4544,N_4477,N_4475);
nand U4545 (N_4545,N_4357,N_4434);
nor U4546 (N_4546,N_4449,N_4411);
nor U4547 (N_4547,N_4360,N_4394);
and U4548 (N_4548,N_4488,N_4383);
xnor U4549 (N_4549,N_4386,N_4493);
and U4550 (N_4550,N_4424,N_4374);
nand U4551 (N_4551,N_4485,N_4392);
and U4552 (N_4552,N_4481,N_4492);
and U4553 (N_4553,N_4408,N_4455);
and U4554 (N_4554,N_4354,N_4363);
nand U4555 (N_4555,N_4358,N_4479);
and U4556 (N_4556,N_4487,N_4402);
xnor U4557 (N_4557,N_4453,N_4406);
nor U4558 (N_4558,N_4445,N_4444);
nor U4559 (N_4559,N_4468,N_4395);
or U4560 (N_4560,N_4425,N_4401);
or U4561 (N_4561,N_4497,N_4476);
or U4562 (N_4562,N_4451,N_4426);
or U4563 (N_4563,N_4447,N_4414);
and U4564 (N_4564,N_4472,N_4376);
xor U4565 (N_4565,N_4373,N_4353);
xor U4566 (N_4566,N_4372,N_4419);
xnor U4567 (N_4567,N_4459,N_4450);
xnor U4568 (N_4568,N_4413,N_4388);
nand U4569 (N_4569,N_4463,N_4378);
and U4570 (N_4570,N_4462,N_4427);
nand U4571 (N_4571,N_4366,N_4368);
xnor U4572 (N_4572,N_4452,N_4496);
nand U4573 (N_4573,N_4480,N_4412);
nand U4574 (N_4574,N_4352,N_4381);
nand U4575 (N_4575,N_4458,N_4355);
nand U4576 (N_4576,N_4491,N_4368);
and U4577 (N_4577,N_4473,N_4427);
and U4578 (N_4578,N_4408,N_4463);
and U4579 (N_4579,N_4410,N_4384);
xnor U4580 (N_4580,N_4383,N_4442);
xor U4581 (N_4581,N_4453,N_4462);
and U4582 (N_4582,N_4454,N_4434);
xnor U4583 (N_4583,N_4496,N_4398);
nand U4584 (N_4584,N_4400,N_4420);
and U4585 (N_4585,N_4478,N_4375);
xor U4586 (N_4586,N_4482,N_4433);
nand U4587 (N_4587,N_4474,N_4424);
nand U4588 (N_4588,N_4451,N_4477);
xor U4589 (N_4589,N_4372,N_4407);
nand U4590 (N_4590,N_4391,N_4410);
nand U4591 (N_4591,N_4363,N_4404);
xor U4592 (N_4592,N_4493,N_4434);
xnor U4593 (N_4593,N_4448,N_4403);
nand U4594 (N_4594,N_4395,N_4463);
and U4595 (N_4595,N_4352,N_4466);
nor U4596 (N_4596,N_4445,N_4494);
nand U4597 (N_4597,N_4359,N_4426);
nor U4598 (N_4598,N_4365,N_4388);
or U4599 (N_4599,N_4379,N_4430);
xnor U4600 (N_4600,N_4418,N_4455);
nor U4601 (N_4601,N_4388,N_4447);
and U4602 (N_4602,N_4451,N_4386);
or U4603 (N_4603,N_4476,N_4459);
or U4604 (N_4604,N_4438,N_4499);
and U4605 (N_4605,N_4387,N_4433);
xor U4606 (N_4606,N_4355,N_4382);
or U4607 (N_4607,N_4460,N_4368);
xnor U4608 (N_4608,N_4420,N_4486);
or U4609 (N_4609,N_4412,N_4422);
or U4610 (N_4610,N_4439,N_4444);
or U4611 (N_4611,N_4382,N_4404);
or U4612 (N_4612,N_4371,N_4433);
nand U4613 (N_4613,N_4384,N_4459);
nand U4614 (N_4614,N_4356,N_4495);
and U4615 (N_4615,N_4434,N_4400);
xnor U4616 (N_4616,N_4413,N_4371);
xor U4617 (N_4617,N_4499,N_4396);
nand U4618 (N_4618,N_4448,N_4480);
xnor U4619 (N_4619,N_4386,N_4362);
nor U4620 (N_4620,N_4454,N_4478);
nand U4621 (N_4621,N_4466,N_4491);
nand U4622 (N_4622,N_4377,N_4436);
nor U4623 (N_4623,N_4368,N_4481);
nand U4624 (N_4624,N_4451,N_4488);
nand U4625 (N_4625,N_4478,N_4435);
nor U4626 (N_4626,N_4446,N_4427);
and U4627 (N_4627,N_4422,N_4493);
nor U4628 (N_4628,N_4439,N_4360);
and U4629 (N_4629,N_4411,N_4366);
nand U4630 (N_4630,N_4458,N_4428);
nand U4631 (N_4631,N_4369,N_4395);
nand U4632 (N_4632,N_4433,N_4352);
xor U4633 (N_4633,N_4476,N_4470);
nand U4634 (N_4634,N_4482,N_4353);
and U4635 (N_4635,N_4408,N_4392);
or U4636 (N_4636,N_4380,N_4407);
nand U4637 (N_4637,N_4496,N_4406);
and U4638 (N_4638,N_4491,N_4376);
xor U4639 (N_4639,N_4381,N_4350);
or U4640 (N_4640,N_4477,N_4412);
xnor U4641 (N_4641,N_4444,N_4487);
or U4642 (N_4642,N_4487,N_4471);
nand U4643 (N_4643,N_4483,N_4446);
nand U4644 (N_4644,N_4481,N_4477);
xnor U4645 (N_4645,N_4437,N_4497);
or U4646 (N_4646,N_4356,N_4418);
and U4647 (N_4647,N_4473,N_4434);
nor U4648 (N_4648,N_4475,N_4462);
and U4649 (N_4649,N_4406,N_4423);
xor U4650 (N_4650,N_4630,N_4531);
and U4651 (N_4651,N_4540,N_4587);
nand U4652 (N_4652,N_4552,N_4574);
or U4653 (N_4653,N_4565,N_4567);
xor U4654 (N_4654,N_4614,N_4588);
xor U4655 (N_4655,N_4523,N_4564);
nor U4656 (N_4656,N_4607,N_4563);
nand U4657 (N_4657,N_4584,N_4507);
and U4658 (N_4658,N_4591,N_4511);
nor U4659 (N_4659,N_4643,N_4649);
or U4660 (N_4660,N_4506,N_4516);
and U4661 (N_4661,N_4503,N_4606);
xnor U4662 (N_4662,N_4637,N_4553);
xor U4663 (N_4663,N_4510,N_4605);
nor U4664 (N_4664,N_4534,N_4515);
nor U4665 (N_4665,N_4586,N_4538);
nand U4666 (N_4666,N_4526,N_4561);
and U4667 (N_4667,N_4570,N_4556);
or U4668 (N_4668,N_4529,N_4522);
xnor U4669 (N_4669,N_4544,N_4647);
nor U4670 (N_4670,N_4550,N_4558);
or U4671 (N_4671,N_4504,N_4543);
and U4672 (N_4672,N_4596,N_4512);
or U4673 (N_4673,N_4648,N_4572);
and U4674 (N_4674,N_4594,N_4546);
nand U4675 (N_4675,N_4537,N_4545);
nand U4676 (N_4676,N_4639,N_4547);
nand U4677 (N_4677,N_4617,N_4542);
nor U4678 (N_4678,N_4592,N_4579);
and U4679 (N_4679,N_4622,N_4536);
nand U4680 (N_4680,N_4636,N_4530);
nor U4681 (N_4681,N_4548,N_4518);
and U4682 (N_4682,N_4627,N_4533);
nand U4683 (N_4683,N_4585,N_4551);
and U4684 (N_4684,N_4597,N_4632);
nor U4685 (N_4685,N_4608,N_4620);
xor U4686 (N_4686,N_4535,N_4619);
nand U4687 (N_4687,N_4615,N_4559);
and U4688 (N_4688,N_4527,N_4610);
and U4689 (N_4689,N_4593,N_4578);
nand U4690 (N_4690,N_4568,N_4566);
or U4691 (N_4691,N_4638,N_4613);
nor U4692 (N_4692,N_4539,N_4560);
nor U4693 (N_4693,N_4573,N_4595);
and U4694 (N_4694,N_4508,N_4618);
nand U4695 (N_4695,N_4582,N_4521);
nor U4696 (N_4696,N_4590,N_4517);
nand U4697 (N_4697,N_4635,N_4621);
nor U4698 (N_4698,N_4623,N_4532);
nor U4699 (N_4699,N_4645,N_4604);
and U4700 (N_4700,N_4589,N_4525);
and U4701 (N_4701,N_4626,N_4611);
xor U4702 (N_4702,N_4612,N_4520);
nand U4703 (N_4703,N_4513,N_4519);
or U4704 (N_4704,N_4646,N_4599);
nor U4705 (N_4705,N_4602,N_4577);
or U4706 (N_4706,N_4501,N_4600);
or U4707 (N_4707,N_4580,N_4631);
and U4708 (N_4708,N_4575,N_4500);
nor U4709 (N_4709,N_4562,N_4541);
nor U4710 (N_4710,N_4571,N_4616);
xor U4711 (N_4711,N_4601,N_4514);
nand U4712 (N_4712,N_4505,N_4502);
or U4713 (N_4713,N_4557,N_4640);
nor U4714 (N_4714,N_4528,N_4634);
and U4715 (N_4715,N_4624,N_4598);
nand U4716 (N_4716,N_4603,N_4581);
or U4717 (N_4717,N_4509,N_4524);
nand U4718 (N_4718,N_4549,N_4555);
or U4719 (N_4719,N_4554,N_4644);
or U4720 (N_4720,N_4629,N_4576);
nand U4721 (N_4721,N_4569,N_4642);
or U4722 (N_4722,N_4641,N_4628);
nor U4723 (N_4723,N_4583,N_4609);
nor U4724 (N_4724,N_4625,N_4633);
or U4725 (N_4725,N_4601,N_4645);
and U4726 (N_4726,N_4548,N_4556);
nand U4727 (N_4727,N_4511,N_4500);
nor U4728 (N_4728,N_4592,N_4580);
xor U4729 (N_4729,N_4540,N_4598);
and U4730 (N_4730,N_4641,N_4571);
nand U4731 (N_4731,N_4622,N_4615);
or U4732 (N_4732,N_4601,N_4578);
nand U4733 (N_4733,N_4595,N_4569);
xnor U4734 (N_4734,N_4615,N_4586);
xnor U4735 (N_4735,N_4558,N_4534);
nor U4736 (N_4736,N_4529,N_4535);
xor U4737 (N_4737,N_4604,N_4596);
xnor U4738 (N_4738,N_4501,N_4577);
or U4739 (N_4739,N_4576,N_4596);
or U4740 (N_4740,N_4553,N_4629);
nor U4741 (N_4741,N_4596,N_4504);
or U4742 (N_4742,N_4575,N_4562);
xnor U4743 (N_4743,N_4567,N_4615);
or U4744 (N_4744,N_4516,N_4628);
and U4745 (N_4745,N_4610,N_4548);
or U4746 (N_4746,N_4591,N_4552);
and U4747 (N_4747,N_4519,N_4539);
or U4748 (N_4748,N_4546,N_4611);
nand U4749 (N_4749,N_4629,N_4523);
and U4750 (N_4750,N_4544,N_4594);
nor U4751 (N_4751,N_4647,N_4511);
nor U4752 (N_4752,N_4623,N_4619);
or U4753 (N_4753,N_4539,N_4583);
nor U4754 (N_4754,N_4617,N_4521);
or U4755 (N_4755,N_4509,N_4634);
nor U4756 (N_4756,N_4526,N_4643);
xor U4757 (N_4757,N_4645,N_4605);
nor U4758 (N_4758,N_4634,N_4595);
nand U4759 (N_4759,N_4520,N_4643);
and U4760 (N_4760,N_4514,N_4645);
or U4761 (N_4761,N_4518,N_4583);
nor U4762 (N_4762,N_4521,N_4577);
and U4763 (N_4763,N_4569,N_4579);
nand U4764 (N_4764,N_4569,N_4563);
or U4765 (N_4765,N_4563,N_4596);
and U4766 (N_4766,N_4520,N_4564);
nor U4767 (N_4767,N_4510,N_4609);
nor U4768 (N_4768,N_4617,N_4569);
xnor U4769 (N_4769,N_4562,N_4530);
nor U4770 (N_4770,N_4555,N_4573);
nand U4771 (N_4771,N_4599,N_4633);
or U4772 (N_4772,N_4561,N_4587);
nor U4773 (N_4773,N_4548,N_4568);
or U4774 (N_4774,N_4584,N_4610);
nor U4775 (N_4775,N_4573,N_4600);
xnor U4776 (N_4776,N_4632,N_4634);
xnor U4777 (N_4777,N_4565,N_4519);
or U4778 (N_4778,N_4538,N_4567);
nor U4779 (N_4779,N_4528,N_4562);
and U4780 (N_4780,N_4580,N_4622);
and U4781 (N_4781,N_4513,N_4557);
nor U4782 (N_4782,N_4531,N_4555);
xor U4783 (N_4783,N_4540,N_4531);
xor U4784 (N_4784,N_4607,N_4545);
or U4785 (N_4785,N_4636,N_4608);
and U4786 (N_4786,N_4614,N_4594);
and U4787 (N_4787,N_4547,N_4509);
xnor U4788 (N_4788,N_4621,N_4543);
and U4789 (N_4789,N_4526,N_4504);
and U4790 (N_4790,N_4576,N_4604);
nand U4791 (N_4791,N_4608,N_4625);
nand U4792 (N_4792,N_4532,N_4546);
xor U4793 (N_4793,N_4607,N_4511);
nor U4794 (N_4794,N_4510,N_4566);
nand U4795 (N_4795,N_4615,N_4509);
nor U4796 (N_4796,N_4630,N_4626);
nand U4797 (N_4797,N_4590,N_4632);
xnor U4798 (N_4798,N_4637,N_4608);
nand U4799 (N_4799,N_4565,N_4586);
xnor U4800 (N_4800,N_4791,N_4738);
xor U4801 (N_4801,N_4735,N_4776);
xnor U4802 (N_4802,N_4726,N_4699);
or U4803 (N_4803,N_4799,N_4660);
and U4804 (N_4804,N_4667,N_4692);
xor U4805 (N_4805,N_4666,N_4793);
nand U4806 (N_4806,N_4688,N_4741);
nand U4807 (N_4807,N_4707,N_4782);
nor U4808 (N_4808,N_4676,N_4654);
nand U4809 (N_4809,N_4796,N_4760);
or U4810 (N_4810,N_4655,N_4729);
xnor U4811 (N_4811,N_4790,N_4718);
or U4812 (N_4812,N_4708,N_4710);
or U4813 (N_4813,N_4664,N_4734);
nand U4814 (N_4814,N_4771,N_4720);
xnor U4815 (N_4815,N_4716,N_4768);
nor U4816 (N_4816,N_4744,N_4794);
nand U4817 (N_4817,N_4671,N_4766);
xor U4818 (N_4818,N_4731,N_4789);
and U4819 (N_4819,N_4657,N_4795);
xnor U4820 (N_4820,N_4714,N_4728);
xnor U4821 (N_4821,N_4769,N_4770);
or U4822 (N_4822,N_4725,N_4775);
or U4823 (N_4823,N_4787,N_4695);
and U4824 (N_4824,N_4717,N_4745);
xor U4825 (N_4825,N_4797,N_4669);
nand U4826 (N_4826,N_4673,N_4747);
and U4827 (N_4827,N_4751,N_4665);
nor U4828 (N_4828,N_4722,N_4719);
xor U4829 (N_4829,N_4706,N_4761);
nor U4830 (N_4830,N_4704,N_4778);
nor U4831 (N_4831,N_4650,N_4685);
xor U4832 (N_4832,N_4689,N_4697);
nand U4833 (N_4833,N_4663,N_4672);
or U4834 (N_4834,N_4691,N_4723);
nand U4835 (N_4835,N_4736,N_4755);
nand U4836 (N_4836,N_4727,N_4756);
nand U4837 (N_4837,N_4653,N_4792);
or U4838 (N_4838,N_4694,N_4737);
and U4839 (N_4839,N_4740,N_4730);
nand U4840 (N_4840,N_4788,N_4652);
and U4841 (N_4841,N_4674,N_4743);
or U4842 (N_4842,N_4656,N_4679);
xnor U4843 (N_4843,N_4703,N_4773);
or U4844 (N_4844,N_4668,N_4739);
xor U4845 (N_4845,N_4701,N_4780);
or U4846 (N_4846,N_4754,N_4758);
xor U4847 (N_4847,N_4732,N_4750);
or U4848 (N_4848,N_4680,N_4784);
nor U4849 (N_4849,N_4715,N_4693);
nand U4850 (N_4850,N_4724,N_4774);
nor U4851 (N_4851,N_4690,N_4687);
or U4852 (N_4852,N_4705,N_4702);
or U4853 (N_4853,N_4711,N_4662);
nand U4854 (N_4854,N_4681,N_4762);
nand U4855 (N_4855,N_4742,N_4748);
and U4856 (N_4856,N_4698,N_4783);
or U4857 (N_4857,N_4651,N_4767);
and U4858 (N_4858,N_4753,N_4659);
nand U4859 (N_4859,N_4779,N_4686);
nor U4860 (N_4860,N_4721,N_4765);
or U4861 (N_4861,N_4733,N_4709);
or U4862 (N_4862,N_4764,N_4786);
nor U4863 (N_4863,N_4684,N_4670);
xnor U4864 (N_4864,N_4700,N_4661);
nor U4865 (N_4865,N_4696,N_4763);
nand U4866 (N_4866,N_4713,N_4757);
or U4867 (N_4867,N_4682,N_4658);
xnor U4868 (N_4868,N_4772,N_4683);
and U4869 (N_4869,N_4746,N_4677);
nand U4870 (N_4870,N_4785,N_4752);
xor U4871 (N_4871,N_4678,N_4759);
nand U4872 (N_4872,N_4777,N_4798);
or U4873 (N_4873,N_4712,N_4749);
and U4874 (N_4874,N_4781,N_4675);
xnor U4875 (N_4875,N_4758,N_4717);
nand U4876 (N_4876,N_4707,N_4721);
xnor U4877 (N_4877,N_4760,N_4733);
or U4878 (N_4878,N_4715,N_4699);
xor U4879 (N_4879,N_4670,N_4675);
nand U4880 (N_4880,N_4780,N_4708);
nand U4881 (N_4881,N_4709,N_4665);
nand U4882 (N_4882,N_4744,N_4717);
and U4883 (N_4883,N_4656,N_4789);
xor U4884 (N_4884,N_4736,N_4722);
nand U4885 (N_4885,N_4772,N_4733);
nor U4886 (N_4886,N_4676,N_4671);
nor U4887 (N_4887,N_4652,N_4674);
nand U4888 (N_4888,N_4669,N_4766);
or U4889 (N_4889,N_4753,N_4768);
or U4890 (N_4890,N_4715,N_4787);
and U4891 (N_4891,N_4658,N_4782);
and U4892 (N_4892,N_4796,N_4758);
nor U4893 (N_4893,N_4678,N_4789);
nor U4894 (N_4894,N_4662,N_4670);
xor U4895 (N_4895,N_4664,N_4773);
and U4896 (N_4896,N_4742,N_4660);
xnor U4897 (N_4897,N_4703,N_4784);
xnor U4898 (N_4898,N_4752,N_4691);
nand U4899 (N_4899,N_4718,N_4672);
or U4900 (N_4900,N_4779,N_4681);
or U4901 (N_4901,N_4777,N_4766);
xor U4902 (N_4902,N_4670,N_4781);
nor U4903 (N_4903,N_4754,N_4798);
or U4904 (N_4904,N_4758,N_4677);
and U4905 (N_4905,N_4685,N_4680);
nand U4906 (N_4906,N_4793,N_4743);
nand U4907 (N_4907,N_4735,N_4685);
xnor U4908 (N_4908,N_4773,N_4764);
or U4909 (N_4909,N_4678,N_4695);
or U4910 (N_4910,N_4705,N_4681);
and U4911 (N_4911,N_4761,N_4735);
or U4912 (N_4912,N_4787,N_4710);
or U4913 (N_4913,N_4789,N_4795);
and U4914 (N_4914,N_4708,N_4744);
xnor U4915 (N_4915,N_4798,N_4716);
or U4916 (N_4916,N_4650,N_4797);
nand U4917 (N_4917,N_4652,N_4689);
nor U4918 (N_4918,N_4697,N_4678);
xor U4919 (N_4919,N_4758,N_4766);
nor U4920 (N_4920,N_4793,N_4752);
nand U4921 (N_4921,N_4752,N_4799);
xor U4922 (N_4922,N_4683,N_4728);
nand U4923 (N_4923,N_4674,N_4693);
xnor U4924 (N_4924,N_4697,N_4707);
or U4925 (N_4925,N_4773,N_4738);
and U4926 (N_4926,N_4671,N_4683);
and U4927 (N_4927,N_4675,N_4699);
and U4928 (N_4928,N_4692,N_4713);
nand U4929 (N_4929,N_4779,N_4652);
nand U4930 (N_4930,N_4777,N_4702);
or U4931 (N_4931,N_4766,N_4789);
nor U4932 (N_4932,N_4659,N_4781);
nor U4933 (N_4933,N_4789,N_4702);
nand U4934 (N_4934,N_4777,N_4738);
or U4935 (N_4935,N_4734,N_4758);
xor U4936 (N_4936,N_4673,N_4713);
nor U4937 (N_4937,N_4659,N_4748);
nand U4938 (N_4938,N_4714,N_4696);
nand U4939 (N_4939,N_4690,N_4701);
and U4940 (N_4940,N_4730,N_4667);
and U4941 (N_4941,N_4714,N_4695);
nand U4942 (N_4942,N_4737,N_4788);
and U4943 (N_4943,N_4665,N_4702);
xnor U4944 (N_4944,N_4767,N_4689);
or U4945 (N_4945,N_4788,N_4668);
or U4946 (N_4946,N_4659,N_4796);
nand U4947 (N_4947,N_4762,N_4707);
and U4948 (N_4948,N_4726,N_4753);
xor U4949 (N_4949,N_4744,N_4700);
xor U4950 (N_4950,N_4902,N_4858);
xnor U4951 (N_4951,N_4914,N_4900);
or U4952 (N_4952,N_4854,N_4882);
or U4953 (N_4953,N_4844,N_4946);
xnor U4954 (N_4954,N_4945,N_4865);
and U4955 (N_4955,N_4892,N_4846);
nand U4956 (N_4956,N_4856,N_4903);
or U4957 (N_4957,N_4904,N_4826);
nand U4958 (N_4958,N_4804,N_4916);
xor U4959 (N_4959,N_4811,N_4843);
and U4960 (N_4960,N_4889,N_4823);
nand U4961 (N_4961,N_4940,N_4937);
nand U4962 (N_4962,N_4939,N_4813);
or U4963 (N_4963,N_4947,N_4942);
xnor U4964 (N_4964,N_4887,N_4810);
xnor U4965 (N_4965,N_4881,N_4899);
xnor U4966 (N_4966,N_4905,N_4840);
and U4967 (N_4967,N_4873,N_4819);
xor U4968 (N_4968,N_4895,N_4825);
xor U4969 (N_4969,N_4809,N_4851);
xnor U4970 (N_4970,N_4883,N_4886);
nand U4971 (N_4971,N_4816,N_4925);
xnor U4972 (N_4972,N_4867,N_4839);
xnor U4973 (N_4973,N_4808,N_4872);
or U4974 (N_4974,N_4885,N_4864);
xnor U4975 (N_4975,N_4820,N_4803);
nor U4976 (N_4976,N_4822,N_4802);
and U4977 (N_4977,N_4909,N_4836);
nor U4978 (N_4978,N_4814,N_4866);
or U4979 (N_4979,N_4801,N_4868);
nor U4980 (N_4980,N_4841,N_4936);
nand U4981 (N_4981,N_4862,N_4850);
xor U4982 (N_4982,N_4926,N_4806);
xnor U4983 (N_4983,N_4842,N_4857);
nand U4984 (N_4984,N_4929,N_4941);
xor U4985 (N_4985,N_4919,N_4934);
and U4986 (N_4986,N_4908,N_4894);
or U4987 (N_4987,N_4915,N_4875);
nand U4988 (N_4988,N_4906,N_4920);
or U4989 (N_4989,N_4827,N_4834);
nand U4990 (N_4990,N_4821,N_4817);
or U4991 (N_4991,N_4924,N_4800);
nand U4992 (N_4992,N_4884,N_4829);
nand U4993 (N_4993,N_4910,N_4860);
and U4994 (N_4994,N_4832,N_4879);
xnor U4995 (N_4995,N_4838,N_4880);
or U4996 (N_4996,N_4930,N_4876);
or U4997 (N_4997,N_4943,N_4847);
or U4998 (N_4998,N_4853,N_4888);
and U4999 (N_4999,N_4912,N_4831);
nand U5000 (N_5000,N_4877,N_4849);
and U5001 (N_5001,N_4935,N_4855);
or U5002 (N_5002,N_4835,N_4944);
xor U5003 (N_5003,N_4896,N_4852);
nor U5004 (N_5004,N_4893,N_4891);
or U5005 (N_5005,N_4830,N_4932);
and U5006 (N_5006,N_4907,N_4848);
xor U5007 (N_5007,N_4861,N_4913);
nand U5008 (N_5008,N_4807,N_4923);
nand U5009 (N_5009,N_4859,N_4911);
nor U5010 (N_5010,N_4833,N_4878);
nand U5011 (N_5011,N_4869,N_4874);
xnor U5012 (N_5012,N_4948,N_4949);
nor U5013 (N_5013,N_4818,N_4921);
and U5014 (N_5014,N_4918,N_4805);
nor U5015 (N_5015,N_4812,N_4828);
nor U5016 (N_5016,N_4922,N_4815);
and U5017 (N_5017,N_4901,N_4931);
and U5018 (N_5018,N_4890,N_4928);
nor U5019 (N_5019,N_4938,N_4933);
and U5020 (N_5020,N_4897,N_4863);
and U5021 (N_5021,N_4824,N_4917);
nor U5022 (N_5022,N_4845,N_4870);
nand U5023 (N_5023,N_4898,N_4837);
or U5024 (N_5024,N_4871,N_4927);
xnor U5025 (N_5025,N_4945,N_4911);
or U5026 (N_5026,N_4948,N_4847);
nor U5027 (N_5027,N_4939,N_4929);
and U5028 (N_5028,N_4852,N_4923);
nand U5029 (N_5029,N_4919,N_4850);
and U5030 (N_5030,N_4933,N_4879);
nand U5031 (N_5031,N_4883,N_4812);
and U5032 (N_5032,N_4818,N_4944);
xnor U5033 (N_5033,N_4824,N_4834);
nor U5034 (N_5034,N_4841,N_4940);
xor U5035 (N_5035,N_4850,N_4904);
and U5036 (N_5036,N_4862,N_4860);
nand U5037 (N_5037,N_4810,N_4831);
nand U5038 (N_5038,N_4947,N_4890);
nor U5039 (N_5039,N_4926,N_4949);
nand U5040 (N_5040,N_4832,N_4897);
xnor U5041 (N_5041,N_4847,N_4877);
or U5042 (N_5042,N_4933,N_4815);
nor U5043 (N_5043,N_4889,N_4809);
nand U5044 (N_5044,N_4826,N_4902);
and U5045 (N_5045,N_4900,N_4851);
xnor U5046 (N_5046,N_4838,N_4829);
or U5047 (N_5047,N_4848,N_4807);
or U5048 (N_5048,N_4901,N_4934);
or U5049 (N_5049,N_4812,N_4805);
nand U5050 (N_5050,N_4886,N_4942);
nand U5051 (N_5051,N_4814,N_4899);
nor U5052 (N_5052,N_4913,N_4906);
nand U5053 (N_5053,N_4906,N_4855);
and U5054 (N_5054,N_4875,N_4855);
or U5055 (N_5055,N_4901,N_4844);
xor U5056 (N_5056,N_4805,N_4860);
nand U5057 (N_5057,N_4914,N_4874);
xnor U5058 (N_5058,N_4854,N_4883);
and U5059 (N_5059,N_4851,N_4874);
nand U5060 (N_5060,N_4886,N_4828);
nand U5061 (N_5061,N_4845,N_4853);
nand U5062 (N_5062,N_4849,N_4833);
nor U5063 (N_5063,N_4878,N_4938);
and U5064 (N_5064,N_4855,N_4834);
nor U5065 (N_5065,N_4904,N_4845);
and U5066 (N_5066,N_4897,N_4940);
and U5067 (N_5067,N_4949,N_4815);
nand U5068 (N_5068,N_4840,N_4895);
nand U5069 (N_5069,N_4813,N_4947);
or U5070 (N_5070,N_4919,N_4825);
and U5071 (N_5071,N_4923,N_4937);
nor U5072 (N_5072,N_4816,N_4914);
nand U5073 (N_5073,N_4886,N_4896);
or U5074 (N_5074,N_4925,N_4917);
nand U5075 (N_5075,N_4897,N_4877);
nand U5076 (N_5076,N_4939,N_4902);
nor U5077 (N_5077,N_4927,N_4884);
nor U5078 (N_5078,N_4922,N_4854);
xor U5079 (N_5079,N_4856,N_4941);
xor U5080 (N_5080,N_4947,N_4800);
nor U5081 (N_5081,N_4862,N_4834);
and U5082 (N_5082,N_4845,N_4889);
or U5083 (N_5083,N_4871,N_4840);
or U5084 (N_5084,N_4929,N_4949);
and U5085 (N_5085,N_4944,N_4842);
nor U5086 (N_5086,N_4920,N_4837);
or U5087 (N_5087,N_4929,N_4839);
nor U5088 (N_5088,N_4848,N_4935);
or U5089 (N_5089,N_4925,N_4871);
or U5090 (N_5090,N_4822,N_4840);
nand U5091 (N_5091,N_4902,N_4868);
nand U5092 (N_5092,N_4815,N_4927);
or U5093 (N_5093,N_4939,N_4932);
xnor U5094 (N_5094,N_4857,N_4912);
xor U5095 (N_5095,N_4831,N_4818);
and U5096 (N_5096,N_4881,N_4872);
nand U5097 (N_5097,N_4823,N_4896);
or U5098 (N_5098,N_4849,N_4886);
xnor U5099 (N_5099,N_4852,N_4808);
nand U5100 (N_5100,N_4981,N_5080);
xnor U5101 (N_5101,N_5048,N_5088);
and U5102 (N_5102,N_5050,N_4963);
xor U5103 (N_5103,N_5057,N_5095);
or U5104 (N_5104,N_5068,N_4962);
nor U5105 (N_5105,N_4955,N_5028);
nor U5106 (N_5106,N_5055,N_5045);
nand U5107 (N_5107,N_5069,N_5024);
xor U5108 (N_5108,N_4959,N_5004);
nor U5109 (N_5109,N_5007,N_5011);
xor U5110 (N_5110,N_5083,N_4980);
xor U5111 (N_5111,N_5060,N_4971);
xnor U5112 (N_5112,N_5000,N_5089);
xnor U5113 (N_5113,N_4997,N_5046);
nor U5114 (N_5114,N_5031,N_4983);
or U5115 (N_5115,N_5023,N_5064);
or U5116 (N_5116,N_5033,N_5078);
and U5117 (N_5117,N_5085,N_5072);
xor U5118 (N_5118,N_5098,N_4982);
nand U5119 (N_5119,N_4992,N_5010);
or U5120 (N_5120,N_4999,N_5021);
and U5121 (N_5121,N_5030,N_4979);
or U5122 (N_5122,N_5073,N_5036);
nor U5123 (N_5123,N_5096,N_4977);
or U5124 (N_5124,N_5099,N_4964);
xor U5125 (N_5125,N_5092,N_5086);
and U5126 (N_5126,N_4985,N_5090);
xor U5127 (N_5127,N_5067,N_4958);
nand U5128 (N_5128,N_5018,N_4988);
nand U5129 (N_5129,N_5084,N_4950);
nand U5130 (N_5130,N_5029,N_4973);
nor U5131 (N_5131,N_5094,N_5074);
nor U5132 (N_5132,N_5001,N_5075);
xnor U5133 (N_5133,N_4960,N_5081);
and U5134 (N_5134,N_4990,N_4967);
or U5135 (N_5135,N_5016,N_4975);
nand U5136 (N_5136,N_5040,N_4998);
nor U5137 (N_5137,N_5022,N_5049);
nand U5138 (N_5138,N_5054,N_5027);
and U5139 (N_5139,N_5008,N_5061);
xor U5140 (N_5140,N_5043,N_5053);
nand U5141 (N_5141,N_5003,N_5062);
or U5142 (N_5142,N_4995,N_4952);
nor U5143 (N_5143,N_5052,N_5093);
and U5144 (N_5144,N_4965,N_4951);
xor U5145 (N_5145,N_5009,N_5097);
nand U5146 (N_5146,N_5005,N_5058);
and U5147 (N_5147,N_4978,N_5038);
and U5148 (N_5148,N_5047,N_5070);
nor U5149 (N_5149,N_4954,N_4986);
nand U5150 (N_5150,N_5056,N_5013);
nand U5151 (N_5151,N_5019,N_5012);
nand U5152 (N_5152,N_5026,N_5079);
xnor U5153 (N_5153,N_4957,N_4972);
or U5154 (N_5154,N_5077,N_5063);
xnor U5155 (N_5155,N_5044,N_4989);
nand U5156 (N_5156,N_4991,N_4956);
and U5157 (N_5157,N_4976,N_4974);
and U5158 (N_5158,N_5032,N_5041);
xnor U5159 (N_5159,N_5087,N_4987);
and U5160 (N_5160,N_4968,N_4966);
xnor U5161 (N_5161,N_5020,N_5059);
xor U5162 (N_5162,N_5034,N_4969);
or U5163 (N_5163,N_5014,N_5076);
and U5164 (N_5164,N_5082,N_5025);
nand U5165 (N_5165,N_4970,N_5002);
nand U5166 (N_5166,N_4994,N_5035);
or U5167 (N_5167,N_5015,N_5091);
xnor U5168 (N_5168,N_5037,N_5066);
nor U5169 (N_5169,N_5065,N_5006);
nand U5170 (N_5170,N_5071,N_4993);
xnor U5171 (N_5171,N_5039,N_4961);
nand U5172 (N_5172,N_5051,N_5017);
or U5173 (N_5173,N_4953,N_4984);
nand U5174 (N_5174,N_4996,N_5042);
or U5175 (N_5175,N_5001,N_4990);
nor U5176 (N_5176,N_4974,N_5094);
xnor U5177 (N_5177,N_5086,N_4974);
or U5178 (N_5178,N_5037,N_5087);
and U5179 (N_5179,N_4959,N_4993);
nor U5180 (N_5180,N_5057,N_5066);
nor U5181 (N_5181,N_4956,N_5076);
or U5182 (N_5182,N_5043,N_5096);
xor U5183 (N_5183,N_5020,N_4989);
nand U5184 (N_5184,N_5090,N_4953);
nand U5185 (N_5185,N_4954,N_4976);
xor U5186 (N_5186,N_4993,N_5016);
and U5187 (N_5187,N_5042,N_5011);
or U5188 (N_5188,N_5091,N_5050);
or U5189 (N_5189,N_5036,N_5084);
and U5190 (N_5190,N_4972,N_5095);
and U5191 (N_5191,N_4953,N_5035);
nand U5192 (N_5192,N_5099,N_5041);
nand U5193 (N_5193,N_4989,N_5058);
nor U5194 (N_5194,N_5066,N_4982);
or U5195 (N_5195,N_4994,N_5076);
or U5196 (N_5196,N_5050,N_5087);
nand U5197 (N_5197,N_4965,N_5056);
xor U5198 (N_5198,N_5073,N_5029);
and U5199 (N_5199,N_4980,N_5096);
and U5200 (N_5200,N_5057,N_4970);
and U5201 (N_5201,N_4953,N_5010);
and U5202 (N_5202,N_5034,N_5088);
or U5203 (N_5203,N_5048,N_4989);
nand U5204 (N_5204,N_4970,N_4958);
or U5205 (N_5205,N_5001,N_5002);
and U5206 (N_5206,N_5028,N_5053);
and U5207 (N_5207,N_4978,N_5064);
or U5208 (N_5208,N_5072,N_5070);
nand U5209 (N_5209,N_5057,N_4952);
or U5210 (N_5210,N_4952,N_4958);
xnor U5211 (N_5211,N_4968,N_4994);
xor U5212 (N_5212,N_4986,N_5091);
and U5213 (N_5213,N_4977,N_5073);
or U5214 (N_5214,N_4960,N_5057);
nand U5215 (N_5215,N_5021,N_4970);
xor U5216 (N_5216,N_5049,N_5014);
nor U5217 (N_5217,N_4992,N_5086);
and U5218 (N_5218,N_4976,N_4980);
xor U5219 (N_5219,N_5095,N_5087);
nor U5220 (N_5220,N_4952,N_5043);
nand U5221 (N_5221,N_5021,N_4994);
nor U5222 (N_5222,N_5076,N_5018);
or U5223 (N_5223,N_5032,N_5005);
and U5224 (N_5224,N_5072,N_4998);
nor U5225 (N_5225,N_4992,N_5041);
nand U5226 (N_5226,N_5083,N_5039);
or U5227 (N_5227,N_5071,N_5075);
nand U5228 (N_5228,N_4983,N_5036);
xnor U5229 (N_5229,N_5097,N_4987);
and U5230 (N_5230,N_5077,N_4961);
nor U5231 (N_5231,N_4988,N_5084);
and U5232 (N_5232,N_4999,N_5085);
nand U5233 (N_5233,N_5087,N_5058);
nor U5234 (N_5234,N_5086,N_5008);
nand U5235 (N_5235,N_5081,N_4975);
nor U5236 (N_5236,N_5041,N_4954);
nor U5237 (N_5237,N_5046,N_5077);
and U5238 (N_5238,N_4985,N_5036);
xor U5239 (N_5239,N_4975,N_5012);
nand U5240 (N_5240,N_4969,N_5025);
xnor U5241 (N_5241,N_5091,N_5090);
nor U5242 (N_5242,N_4987,N_5029);
or U5243 (N_5243,N_5030,N_4962);
or U5244 (N_5244,N_4964,N_5062);
xnor U5245 (N_5245,N_5027,N_4992);
and U5246 (N_5246,N_4981,N_5056);
and U5247 (N_5247,N_5033,N_5051);
or U5248 (N_5248,N_4969,N_4957);
and U5249 (N_5249,N_4985,N_5093);
nand U5250 (N_5250,N_5138,N_5127);
xnor U5251 (N_5251,N_5173,N_5179);
nand U5252 (N_5252,N_5186,N_5215);
nand U5253 (N_5253,N_5151,N_5180);
or U5254 (N_5254,N_5107,N_5199);
and U5255 (N_5255,N_5115,N_5174);
nor U5256 (N_5256,N_5229,N_5102);
or U5257 (N_5257,N_5206,N_5228);
or U5258 (N_5258,N_5247,N_5128);
xor U5259 (N_5259,N_5101,N_5100);
nor U5260 (N_5260,N_5243,N_5142);
or U5261 (N_5261,N_5133,N_5210);
or U5262 (N_5262,N_5230,N_5197);
nor U5263 (N_5263,N_5181,N_5246);
and U5264 (N_5264,N_5217,N_5124);
and U5265 (N_5265,N_5166,N_5112);
nand U5266 (N_5266,N_5191,N_5139);
nand U5267 (N_5267,N_5204,N_5244);
and U5268 (N_5268,N_5104,N_5103);
nor U5269 (N_5269,N_5198,N_5220);
nand U5270 (N_5270,N_5120,N_5123);
and U5271 (N_5271,N_5235,N_5249);
nand U5272 (N_5272,N_5185,N_5209);
and U5273 (N_5273,N_5126,N_5130);
nand U5274 (N_5274,N_5109,N_5105);
and U5275 (N_5275,N_5207,N_5145);
and U5276 (N_5276,N_5158,N_5194);
or U5277 (N_5277,N_5135,N_5169);
xor U5278 (N_5278,N_5141,N_5156);
and U5279 (N_5279,N_5171,N_5154);
nand U5280 (N_5280,N_5153,N_5231);
nor U5281 (N_5281,N_5195,N_5225);
and U5282 (N_5282,N_5222,N_5203);
xnor U5283 (N_5283,N_5237,N_5146);
nand U5284 (N_5284,N_5177,N_5182);
and U5285 (N_5285,N_5147,N_5116);
xor U5286 (N_5286,N_5205,N_5200);
or U5287 (N_5287,N_5183,N_5233);
nor U5288 (N_5288,N_5121,N_5172);
nor U5289 (N_5289,N_5211,N_5152);
and U5290 (N_5290,N_5106,N_5201);
nor U5291 (N_5291,N_5214,N_5188);
or U5292 (N_5292,N_5196,N_5162);
nor U5293 (N_5293,N_5132,N_5122);
and U5294 (N_5294,N_5178,N_5125);
xnor U5295 (N_5295,N_5149,N_5176);
nor U5296 (N_5296,N_5187,N_5248);
nor U5297 (N_5297,N_5190,N_5165);
xnor U5298 (N_5298,N_5212,N_5114);
nor U5299 (N_5299,N_5161,N_5108);
or U5300 (N_5300,N_5208,N_5164);
or U5301 (N_5301,N_5245,N_5226);
and U5302 (N_5302,N_5155,N_5219);
nor U5303 (N_5303,N_5232,N_5144);
or U5304 (N_5304,N_5227,N_5216);
and U5305 (N_5305,N_5148,N_5113);
nand U5306 (N_5306,N_5134,N_5111);
nand U5307 (N_5307,N_5159,N_5170);
nand U5308 (N_5308,N_5241,N_5119);
nor U5309 (N_5309,N_5137,N_5129);
and U5310 (N_5310,N_5239,N_5157);
xnor U5311 (N_5311,N_5242,N_5175);
and U5312 (N_5312,N_5238,N_5189);
nor U5313 (N_5313,N_5168,N_5234);
nor U5314 (N_5314,N_5240,N_5218);
nand U5315 (N_5315,N_5131,N_5163);
or U5316 (N_5316,N_5224,N_5160);
nor U5317 (N_5317,N_5150,N_5221);
and U5318 (N_5318,N_5184,N_5236);
nor U5319 (N_5319,N_5193,N_5143);
nand U5320 (N_5320,N_5136,N_5202);
nor U5321 (N_5321,N_5167,N_5110);
and U5322 (N_5322,N_5118,N_5117);
and U5323 (N_5323,N_5192,N_5223);
nor U5324 (N_5324,N_5213,N_5140);
xor U5325 (N_5325,N_5200,N_5177);
nand U5326 (N_5326,N_5126,N_5224);
or U5327 (N_5327,N_5164,N_5177);
and U5328 (N_5328,N_5163,N_5193);
xnor U5329 (N_5329,N_5124,N_5108);
nor U5330 (N_5330,N_5240,N_5178);
and U5331 (N_5331,N_5118,N_5142);
and U5332 (N_5332,N_5215,N_5103);
nor U5333 (N_5333,N_5135,N_5233);
and U5334 (N_5334,N_5135,N_5216);
nand U5335 (N_5335,N_5207,N_5177);
and U5336 (N_5336,N_5173,N_5217);
or U5337 (N_5337,N_5110,N_5112);
and U5338 (N_5338,N_5231,N_5234);
nand U5339 (N_5339,N_5135,N_5105);
or U5340 (N_5340,N_5156,N_5180);
xnor U5341 (N_5341,N_5132,N_5116);
nor U5342 (N_5342,N_5122,N_5110);
nor U5343 (N_5343,N_5174,N_5150);
nand U5344 (N_5344,N_5148,N_5235);
nor U5345 (N_5345,N_5162,N_5205);
nor U5346 (N_5346,N_5154,N_5117);
or U5347 (N_5347,N_5153,N_5141);
nand U5348 (N_5348,N_5193,N_5196);
nand U5349 (N_5349,N_5205,N_5176);
xor U5350 (N_5350,N_5198,N_5234);
nor U5351 (N_5351,N_5153,N_5235);
and U5352 (N_5352,N_5146,N_5125);
nand U5353 (N_5353,N_5175,N_5205);
or U5354 (N_5354,N_5174,N_5176);
nor U5355 (N_5355,N_5180,N_5193);
xnor U5356 (N_5356,N_5196,N_5121);
or U5357 (N_5357,N_5164,N_5116);
nand U5358 (N_5358,N_5179,N_5125);
xor U5359 (N_5359,N_5206,N_5233);
and U5360 (N_5360,N_5242,N_5150);
xnor U5361 (N_5361,N_5219,N_5127);
xor U5362 (N_5362,N_5243,N_5236);
xor U5363 (N_5363,N_5208,N_5212);
or U5364 (N_5364,N_5242,N_5219);
nand U5365 (N_5365,N_5103,N_5185);
xnor U5366 (N_5366,N_5200,N_5171);
and U5367 (N_5367,N_5219,N_5118);
xor U5368 (N_5368,N_5236,N_5207);
and U5369 (N_5369,N_5125,N_5242);
xor U5370 (N_5370,N_5233,N_5113);
and U5371 (N_5371,N_5174,N_5113);
and U5372 (N_5372,N_5190,N_5193);
or U5373 (N_5373,N_5212,N_5185);
or U5374 (N_5374,N_5117,N_5159);
or U5375 (N_5375,N_5143,N_5117);
and U5376 (N_5376,N_5213,N_5184);
or U5377 (N_5377,N_5110,N_5215);
nor U5378 (N_5378,N_5168,N_5235);
or U5379 (N_5379,N_5181,N_5204);
or U5380 (N_5380,N_5107,N_5244);
or U5381 (N_5381,N_5183,N_5176);
or U5382 (N_5382,N_5130,N_5218);
nor U5383 (N_5383,N_5118,N_5145);
and U5384 (N_5384,N_5169,N_5167);
and U5385 (N_5385,N_5141,N_5202);
or U5386 (N_5386,N_5208,N_5176);
and U5387 (N_5387,N_5213,N_5155);
nor U5388 (N_5388,N_5138,N_5223);
nor U5389 (N_5389,N_5220,N_5128);
or U5390 (N_5390,N_5126,N_5102);
nor U5391 (N_5391,N_5211,N_5123);
and U5392 (N_5392,N_5223,N_5119);
nor U5393 (N_5393,N_5100,N_5234);
nor U5394 (N_5394,N_5131,N_5232);
nand U5395 (N_5395,N_5192,N_5218);
and U5396 (N_5396,N_5155,N_5153);
xnor U5397 (N_5397,N_5116,N_5228);
nor U5398 (N_5398,N_5216,N_5126);
nor U5399 (N_5399,N_5123,N_5232);
or U5400 (N_5400,N_5389,N_5287);
xor U5401 (N_5401,N_5291,N_5350);
nand U5402 (N_5402,N_5385,N_5295);
and U5403 (N_5403,N_5357,N_5352);
nor U5404 (N_5404,N_5361,N_5337);
xnor U5405 (N_5405,N_5344,N_5383);
xor U5406 (N_5406,N_5293,N_5380);
and U5407 (N_5407,N_5390,N_5369);
nor U5408 (N_5408,N_5281,N_5331);
and U5409 (N_5409,N_5274,N_5360);
xnor U5410 (N_5410,N_5256,N_5268);
nand U5411 (N_5411,N_5300,N_5263);
nor U5412 (N_5412,N_5366,N_5261);
nand U5413 (N_5413,N_5325,N_5269);
xor U5414 (N_5414,N_5393,N_5250);
or U5415 (N_5415,N_5345,N_5388);
or U5416 (N_5416,N_5272,N_5286);
or U5417 (N_5417,N_5399,N_5260);
nor U5418 (N_5418,N_5373,N_5283);
nor U5419 (N_5419,N_5306,N_5301);
and U5420 (N_5420,N_5333,N_5296);
nor U5421 (N_5421,N_5270,N_5336);
nand U5422 (N_5422,N_5315,N_5328);
or U5423 (N_5423,N_5258,N_5313);
and U5424 (N_5424,N_5298,N_5288);
nand U5425 (N_5425,N_5307,N_5358);
or U5426 (N_5426,N_5367,N_5303);
nor U5427 (N_5427,N_5353,N_5365);
xor U5428 (N_5428,N_5392,N_5304);
and U5429 (N_5429,N_5310,N_5339);
xor U5430 (N_5430,N_5319,N_5271);
xnor U5431 (N_5431,N_5276,N_5252);
nand U5432 (N_5432,N_5267,N_5302);
or U5433 (N_5433,N_5318,N_5334);
nor U5434 (N_5434,N_5395,N_5356);
and U5435 (N_5435,N_5259,N_5320);
xor U5436 (N_5436,N_5265,N_5262);
xnor U5437 (N_5437,N_5362,N_5381);
nand U5438 (N_5438,N_5377,N_5305);
nand U5439 (N_5439,N_5290,N_5343);
nand U5440 (N_5440,N_5351,N_5285);
xnor U5441 (N_5441,N_5257,N_5321);
xnor U5442 (N_5442,N_5317,N_5363);
or U5443 (N_5443,N_5278,N_5289);
or U5444 (N_5444,N_5264,N_5398);
xnor U5445 (N_5445,N_5338,N_5299);
or U5446 (N_5446,N_5348,N_5326);
or U5447 (N_5447,N_5375,N_5311);
xnor U5448 (N_5448,N_5266,N_5359);
xnor U5449 (N_5449,N_5371,N_5275);
xor U5450 (N_5450,N_5335,N_5308);
nand U5451 (N_5451,N_5394,N_5284);
or U5452 (N_5452,N_5378,N_5327);
or U5453 (N_5453,N_5316,N_5294);
xor U5454 (N_5454,N_5391,N_5251);
nor U5455 (N_5455,N_5355,N_5372);
and U5456 (N_5456,N_5370,N_5322);
and U5457 (N_5457,N_5349,N_5292);
or U5458 (N_5458,N_5323,N_5282);
and U5459 (N_5459,N_5364,N_5346);
or U5460 (N_5460,N_5332,N_5329);
or U5461 (N_5461,N_5314,N_5280);
and U5462 (N_5462,N_5279,N_5386);
or U5463 (N_5463,N_5382,N_5297);
and U5464 (N_5464,N_5255,N_5379);
or U5465 (N_5465,N_5374,N_5254);
nand U5466 (N_5466,N_5396,N_5368);
nor U5467 (N_5467,N_5340,N_5387);
or U5468 (N_5468,N_5273,N_5330);
nor U5469 (N_5469,N_5309,N_5277);
and U5470 (N_5470,N_5376,N_5354);
nand U5471 (N_5471,N_5384,N_5253);
nor U5472 (N_5472,N_5312,N_5341);
or U5473 (N_5473,N_5397,N_5342);
xnor U5474 (N_5474,N_5347,N_5324);
or U5475 (N_5475,N_5380,N_5347);
nor U5476 (N_5476,N_5258,N_5290);
xnor U5477 (N_5477,N_5333,N_5267);
xnor U5478 (N_5478,N_5394,N_5348);
nand U5479 (N_5479,N_5321,N_5311);
nand U5480 (N_5480,N_5321,N_5324);
and U5481 (N_5481,N_5283,N_5260);
and U5482 (N_5482,N_5271,N_5345);
or U5483 (N_5483,N_5364,N_5361);
xor U5484 (N_5484,N_5320,N_5276);
xor U5485 (N_5485,N_5380,N_5264);
nand U5486 (N_5486,N_5395,N_5367);
or U5487 (N_5487,N_5340,N_5326);
nand U5488 (N_5488,N_5375,N_5285);
nor U5489 (N_5489,N_5374,N_5337);
nand U5490 (N_5490,N_5359,N_5368);
nor U5491 (N_5491,N_5311,N_5340);
xor U5492 (N_5492,N_5266,N_5375);
or U5493 (N_5493,N_5287,N_5349);
nor U5494 (N_5494,N_5380,N_5333);
or U5495 (N_5495,N_5352,N_5370);
xor U5496 (N_5496,N_5386,N_5306);
or U5497 (N_5497,N_5368,N_5341);
xor U5498 (N_5498,N_5278,N_5286);
or U5499 (N_5499,N_5356,N_5353);
nand U5500 (N_5500,N_5300,N_5311);
nor U5501 (N_5501,N_5264,N_5262);
nor U5502 (N_5502,N_5303,N_5348);
and U5503 (N_5503,N_5368,N_5312);
xor U5504 (N_5504,N_5353,N_5318);
xor U5505 (N_5505,N_5312,N_5316);
nor U5506 (N_5506,N_5344,N_5253);
or U5507 (N_5507,N_5280,N_5392);
nand U5508 (N_5508,N_5254,N_5356);
nand U5509 (N_5509,N_5280,N_5302);
xnor U5510 (N_5510,N_5265,N_5370);
nand U5511 (N_5511,N_5295,N_5378);
nand U5512 (N_5512,N_5314,N_5251);
nor U5513 (N_5513,N_5381,N_5382);
or U5514 (N_5514,N_5332,N_5372);
nor U5515 (N_5515,N_5313,N_5364);
nand U5516 (N_5516,N_5329,N_5328);
or U5517 (N_5517,N_5358,N_5352);
nand U5518 (N_5518,N_5362,N_5298);
and U5519 (N_5519,N_5325,N_5275);
nor U5520 (N_5520,N_5260,N_5372);
xor U5521 (N_5521,N_5314,N_5270);
nor U5522 (N_5522,N_5374,N_5334);
xnor U5523 (N_5523,N_5384,N_5335);
xor U5524 (N_5524,N_5253,N_5378);
and U5525 (N_5525,N_5365,N_5328);
or U5526 (N_5526,N_5351,N_5256);
nor U5527 (N_5527,N_5307,N_5285);
and U5528 (N_5528,N_5326,N_5309);
nor U5529 (N_5529,N_5334,N_5280);
xnor U5530 (N_5530,N_5344,N_5365);
or U5531 (N_5531,N_5329,N_5373);
or U5532 (N_5532,N_5366,N_5255);
nand U5533 (N_5533,N_5316,N_5372);
and U5534 (N_5534,N_5283,N_5384);
or U5535 (N_5535,N_5326,N_5287);
and U5536 (N_5536,N_5262,N_5260);
nand U5537 (N_5537,N_5397,N_5350);
nor U5538 (N_5538,N_5363,N_5337);
or U5539 (N_5539,N_5365,N_5340);
and U5540 (N_5540,N_5274,N_5332);
nor U5541 (N_5541,N_5317,N_5297);
xor U5542 (N_5542,N_5350,N_5297);
nand U5543 (N_5543,N_5343,N_5377);
xor U5544 (N_5544,N_5273,N_5333);
xnor U5545 (N_5545,N_5265,N_5324);
nand U5546 (N_5546,N_5391,N_5298);
nor U5547 (N_5547,N_5256,N_5363);
and U5548 (N_5548,N_5291,N_5290);
nor U5549 (N_5549,N_5291,N_5284);
nand U5550 (N_5550,N_5541,N_5506);
and U5551 (N_5551,N_5429,N_5520);
and U5552 (N_5552,N_5544,N_5440);
nor U5553 (N_5553,N_5519,N_5532);
and U5554 (N_5554,N_5524,N_5513);
nand U5555 (N_5555,N_5542,N_5503);
and U5556 (N_5556,N_5401,N_5465);
and U5557 (N_5557,N_5430,N_5482);
xnor U5558 (N_5558,N_5433,N_5468);
and U5559 (N_5559,N_5435,N_5421);
nor U5560 (N_5560,N_5529,N_5515);
xnor U5561 (N_5561,N_5490,N_5470);
or U5562 (N_5562,N_5415,N_5497);
or U5563 (N_5563,N_5459,N_5498);
nand U5564 (N_5564,N_5548,N_5514);
nor U5565 (N_5565,N_5450,N_5537);
nand U5566 (N_5566,N_5422,N_5405);
xor U5567 (N_5567,N_5424,N_5500);
xnor U5568 (N_5568,N_5456,N_5413);
and U5569 (N_5569,N_5525,N_5484);
and U5570 (N_5570,N_5501,N_5475);
nand U5571 (N_5571,N_5521,N_5425);
or U5572 (N_5572,N_5442,N_5463);
or U5573 (N_5573,N_5485,N_5474);
xor U5574 (N_5574,N_5464,N_5439);
xor U5575 (N_5575,N_5434,N_5473);
nand U5576 (N_5576,N_5476,N_5438);
or U5577 (N_5577,N_5527,N_5437);
and U5578 (N_5578,N_5409,N_5414);
nand U5579 (N_5579,N_5528,N_5451);
or U5580 (N_5580,N_5426,N_5436);
nand U5581 (N_5581,N_5518,N_5545);
xor U5582 (N_5582,N_5423,N_5417);
nor U5583 (N_5583,N_5479,N_5471);
nand U5584 (N_5584,N_5457,N_5510);
xor U5585 (N_5585,N_5408,N_5496);
nand U5586 (N_5586,N_5508,N_5522);
or U5587 (N_5587,N_5488,N_5432);
nor U5588 (N_5588,N_5411,N_5507);
and U5589 (N_5589,N_5540,N_5509);
xor U5590 (N_5590,N_5543,N_5511);
nand U5591 (N_5591,N_5418,N_5517);
nand U5592 (N_5592,N_5505,N_5491);
nand U5593 (N_5593,N_5523,N_5416);
nor U5594 (N_5594,N_5480,N_5494);
nor U5595 (N_5595,N_5486,N_5404);
xor U5596 (N_5596,N_5460,N_5536);
or U5597 (N_5597,N_5504,N_5431);
nor U5598 (N_5598,N_5402,N_5462);
xnor U5599 (N_5599,N_5478,N_5526);
nand U5600 (N_5600,N_5495,N_5492);
nand U5601 (N_5601,N_5441,N_5487);
and U5602 (N_5602,N_5502,N_5535);
nor U5603 (N_5603,N_5533,N_5469);
and U5604 (N_5604,N_5512,N_5400);
nor U5605 (N_5605,N_5403,N_5534);
nand U5606 (N_5606,N_5427,N_5458);
and U5607 (N_5607,N_5531,N_5547);
or U5608 (N_5608,N_5449,N_5452);
xor U5609 (N_5609,N_5467,N_5493);
and U5610 (N_5610,N_5481,N_5466);
nor U5611 (N_5611,N_5407,N_5419);
nand U5612 (N_5612,N_5539,N_5455);
xnor U5613 (N_5613,N_5412,N_5428);
or U5614 (N_5614,N_5443,N_5448);
and U5615 (N_5615,N_5453,N_5445);
nand U5616 (N_5616,N_5406,N_5444);
nand U5617 (N_5617,N_5446,N_5516);
nand U5618 (N_5618,N_5410,N_5472);
nand U5619 (N_5619,N_5420,N_5530);
nor U5620 (N_5620,N_5499,N_5483);
nor U5621 (N_5621,N_5546,N_5549);
xnor U5622 (N_5622,N_5454,N_5538);
nand U5623 (N_5623,N_5489,N_5477);
nor U5624 (N_5624,N_5447,N_5461);
xor U5625 (N_5625,N_5423,N_5406);
or U5626 (N_5626,N_5453,N_5432);
xor U5627 (N_5627,N_5445,N_5450);
and U5628 (N_5628,N_5531,N_5537);
nand U5629 (N_5629,N_5409,N_5513);
or U5630 (N_5630,N_5424,N_5538);
or U5631 (N_5631,N_5481,N_5429);
nand U5632 (N_5632,N_5463,N_5426);
nand U5633 (N_5633,N_5514,N_5505);
and U5634 (N_5634,N_5505,N_5420);
or U5635 (N_5635,N_5499,N_5497);
nor U5636 (N_5636,N_5492,N_5536);
nand U5637 (N_5637,N_5474,N_5491);
nor U5638 (N_5638,N_5473,N_5460);
or U5639 (N_5639,N_5500,N_5466);
and U5640 (N_5640,N_5499,N_5447);
or U5641 (N_5641,N_5491,N_5439);
and U5642 (N_5642,N_5455,N_5419);
xor U5643 (N_5643,N_5478,N_5443);
or U5644 (N_5644,N_5403,N_5528);
xor U5645 (N_5645,N_5463,N_5465);
nand U5646 (N_5646,N_5459,N_5432);
or U5647 (N_5647,N_5535,N_5441);
xnor U5648 (N_5648,N_5533,N_5535);
and U5649 (N_5649,N_5482,N_5547);
and U5650 (N_5650,N_5493,N_5513);
nor U5651 (N_5651,N_5411,N_5436);
xor U5652 (N_5652,N_5499,N_5545);
nor U5653 (N_5653,N_5464,N_5475);
or U5654 (N_5654,N_5475,N_5507);
nor U5655 (N_5655,N_5489,N_5548);
nor U5656 (N_5656,N_5443,N_5496);
and U5657 (N_5657,N_5424,N_5401);
or U5658 (N_5658,N_5460,N_5521);
nand U5659 (N_5659,N_5443,N_5400);
nor U5660 (N_5660,N_5443,N_5450);
and U5661 (N_5661,N_5496,N_5511);
or U5662 (N_5662,N_5409,N_5464);
xor U5663 (N_5663,N_5426,N_5487);
xnor U5664 (N_5664,N_5450,N_5473);
nand U5665 (N_5665,N_5412,N_5485);
or U5666 (N_5666,N_5537,N_5500);
xnor U5667 (N_5667,N_5490,N_5425);
and U5668 (N_5668,N_5494,N_5490);
or U5669 (N_5669,N_5481,N_5492);
and U5670 (N_5670,N_5406,N_5493);
or U5671 (N_5671,N_5539,N_5525);
nor U5672 (N_5672,N_5427,N_5457);
or U5673 (N_5673,N_5513,N_5494);
nand U5674 (N_5674,N_5458,N_5428);
nand U5675 (N_5675,N_5427,N_5484);
nand U5676 (N_5676,N_5526,N_5427);
xnor U5677 (N_5677,N_5528,N_5492);
or U5678 (N_5678,N_5428,N_5481);
nand U5679 (N_5679,N_5444,N_5520);
and U5680 (N_5680,N_5416,N_5455);
nor U5681 (N_5681,N_5456,N_5466);
nor U5682 (N_5682,N_5503,N_5416);
xor U5683 (N_5683,N_5449,N_5483);
nor U5684 (N_5684,N_5434,N_5412);
nand U5685 (N_5685,N_5435,N_5410);
and U5686 (N_5686,N_5492,N_5546);
xor U5687 (N_5687,N_5481,N_5412);
xnor U5688 (N_5688,N_5453,N_5424);
nand U5689 (N_5689,N_5516,N_5457);
or U5690 (N_5690,N_5432,N_5526);
xnor U5691 (N_5691,N_5490,N_5478);
nor U5692 (N_5692,N_5410,N_5492);
nor U5693 (N_5693,N_5457,N_5444);
nand U5694 (N_5694,N_5429,N_5546);
xnor U5695 (N_5695,N_5543,N_5496);
xor U5696 (N_5696,N_5528,N_5525);
nor U5697 (N_5697,N_5526,N_5474);
nor U5698 (N_5698,N_5440,N_5409);
or U5699 (N_5699,N_5507,N_5546);
nand U5700 (N_5700,N_5692,N_5695);
or U5701 (N_5701,N_5566,N_5567);
or U5702 (N_5702,N_5680,N_5641);
xnor U5703 (N_5703,N_5614,N_5634);
nand U5704 (N_5704,N_5611,N_5665);
nand U5705 (N_5705,N_5554,N_5594);
nor U5706 (N_5706,N_5593,N_5645);
or U5707 (N_5707,N_5698,N_5596);
xnor U5708 (N_5708,N_5666,N_5619);
and U5709 (N_5709,N_5561,N_5588);
and U5710 (N_5710,N_5616,N_5575);
nand U5711 (N_5711,N_5660,N_5696);
and U5712 (N_5712,N_5558,N_5550);
xnor U5713 (N_5713,N_5656,N_5565);
nor U5714 (N_5714,N_5639,N_5652);
and U5715 (N_5715,N_5642,N_5636);
and U5716 (N_5716,N_5590,N_5581);
xnor U5717 (N_5717,N_5605,N_5600);
xnor U5718 (N_5718,N_5556,N_5640);
xnor U5719 (N_5719,N_5675,N_5607);
nor U5720 (N_5720,N_5626,N_5623);
and U5721 (N_5721,N_5670,N_5551);
nor U5722 (N_5722,N_5583,N_5635);
xor U5723 (N_5723,N_5685,N_5598);
xor U5724 (N_5724,N_5679,N_5563);
and U5725 (N_5725,N_5622,N_5689);
nand U5726 (N_5726,N_5668,N_5699);
or U5727 (N_5727,N_5691,N_5597);
nand U5728 (N_5728,N_5643,N_5632);
xor U5729 (N_5729,N_5667,N_5673);
and U5730 (N_5730,N_5559,N_5627);
and U5731 (N_5731,N_5585,N_5592);
or U5732 (N_5732,N_5638,N_5648);
and U5733 (N_5733,N_5604,N_5571);
nor U5734 (N_5734,N_5628,N_5587);
xor U5735 (N_5735,N_5662,N_5621);
or U5736 (N_5736,N_5663,N_5618);
xor U5737 (N_5737,N_5672,N_5580);
nand U5738 (N_5738,N_5577,N_5657);
and U5739 (N_5739,N_5630,N_5674);
nand U5740 (N_5740,N_5620,N_5644);
or U5741 (N_5741,N_5671,N_5637);
nand U5742 (N_5742,N_5684,N_5568);
xor U5743 (N_5743,N_5601,N_5669);
nand U5744 (N_5744,N_5564,N_5570);
nor U5745 (N_5745,N_5678,N_5687);
or U5746 (N_5746,N_5629,N_5688);
xnor U5747 (N_5747,N_5589,N_5661);
nand U5748 (N_5748,N_5574,N_5625);
or U5749 (N_5749,N_5608,N_5681);
nor U5750 (N_5750,N_5610,N_5690);
xor U5751 (N_5751,N_5555,N_5693);
xor U5752 (N_5752,N_5578,N_5557);
nand U5753 (N_5753,N_5603,N_5647);
and U5754 (N_5754,N_5682,N_5631);
and U5755 (N_5755,N_5633,N_5697);
nand U5756 (N_5756,N_5651,N_5586);
nor U5757 (N_5757,N_5599,N_5584);
or U5758 (N_5758,N_5653,N_5617);
xor U5759 (N_5759,N_5572,N_5573);
nor U5760 (N_5760,N_5553,N_5552);
and U5761 (N_5761,N_5664,N_5677);
nand U5762 (N_5762,N_5560,N_5650);
nor U5763 (N_5763,N_5591,N_5613);
and U5764 (N_5764,N_5649,N_5602);
xor U5765 (N_5765,N_5582,N_5659);
and U5766 (N_5766,N_5562,N_5658);
xor U5767 (N_5767,N_5569,N_5612);
nor U5768 (N_5768,N_5615,N_5576);
and U5769 (N_5769,N_5676,N_5579);
nor U5770 (N_5770,N_5654,N_5646);
xor U5771 (N_5771,N_5609,N_5595);
nand U5772 (N_5772,N_5683,N_5686);
and U5773 (N_5773,N_5606,N_5655);
or U5774 (N_5774,N_5624,N_5694);
xnor U5775 (N_5775,N_5586,N_5668);
xnor U5776 (N_5776,N_5647,N_5599);
or U5777 (N_5777,N_5600,N_5657);
nor U5778 (N_5778,N_5668,N_5654);
nor U5779 (N_5779,N_5650,N_5672);
and U5780 (N_5780,N_5598,N_5664);
and U5781 (N_5781,N_5645,N_5660);
xnor U5782 (N_5782,N_5688,N_5613);
and U5783 (N_5783,N_5699,N_5676);
or U5784 (N_5784,N_5636,N_5569);
and U5785 (N_5785,N_5671,N_5655);
nand U5786 (N_5786,N_5579,N_5660);
nand U5787 (N_5787,N_5695,N_5625);
and U5788 (N_5788,N_5654,N_5566);
nor U5789 (N_5789,N_5684,N_5566);
nor U5790 (N_5790,N_5643,N_5626);
nand U5791 (N_5791,N_5628,N_5697);
nand U5792 (N_5792,N_5666,N_5699);
or U5793 (N_5793,N_5628,N_5684);
nand U5794 (N_5794,N_5572,N_5579);
and U5795 (N_5795,N_5623,N_5550);
xnor U5796 (N_5796,N_5636,N_5584);
nor U5797 (N_5797,N_5633,N_5568);
nor U5798 (N_5798,N_5642,N_5652);
nor U5799 (N_5799,N_5588,N_5646);
or U5800 (N_5800,N_5665,N_5690);
nand U5801 (N_5801,N_5608,N_5602);
and U5802 (N_5802,N_5640,N_5597);
or U5803 (N_5803,N_5580,N_5608);
and U5804 (N_5804,N_5594,N_5645);
and U5805 (N_5805,N_5594,N_5567);
and U5806 (N_5806,N_5667,N_5698);
xnor U5807 (N_5807,N_5660,N_5598);
nor U5808 (N_5808,N_5666,N_5590);
and U5809 (N_5809,N_5570,N_5562);
and U5810 (N_5810,N_5693,N_5649);
and U5811 (N_5811,N_5615,N_5657);
nand U5812 (N_5812,N_5554,N_5693);
xor U5813 (N_5813,N_5672,N_5559);
or U5814 (N_5814,N_5626,N_5550);
nor U5815 (N_5815,N_5612,N_5663);
or U5816 (N_5816,N_5585,N_5645);
and U5817 (N_5817,N_5645,N_5625);
or U5818 (N_5818,N_5616,N_5654);
nor U5819 (N_5819,N_5585,N_5551);
and U5820 (N_5820,N_5556,N_5623);
xnor U5821 (N_5821,N_5582,N_5588);
nor U5822 (N_5822,N_5694,N_5685);
or U5823 (N_5823,N_5564,N_5554);
and U5824 (N_5824,N_5672,N_5667);
nor U5825 (N_5825,N_5617,N_5606);
nor U5826 (N_5826,N_5676,N_5636);
nand U5827 (N_5827,N_5691,N_5652);
and U5828 (N_5828,N_5653,N_5553);
xor U5829 (N_5829,N_5582,N_5612);
and U5830 (N_5830,N_5551,N_5558);
nand U5831 (N_5831,N_5665,N_5632);
xor U5832 (N_5832,N_5573,N_5644);
xor U5833 (N_5833,N_5635,N_5577);
xnor U5834 (N_5834,N_5605,N_5620);
nand U5835 (N_5835,N_5623,N_5577);
or U5836 (N_5836,N_5635,N_5579);
nand U5837 (N_5837,N_5550,N_5681);
or U5838 (N_5838,N_5627,N_5691);
or U5839 (N_5839,N_5643,N_5675);
xnor U5840 (N_5840,N_5611,N_5637);
or U5841 (N_5841,N_5582,N_5561);
or U5842 (N_5842,N_5581,N_5655);
and U5843 (N_5843,N_5576,N_5577);
xor U5844 (N_5844,N_5666,N_5643);
xor U5845 (N_5845,N_5550,N_5629);
nand U5846 (N_5846,N_5650,N_5576);
nand U5847 (N_5847,N_5619,N_5680);
and U5848 (N_5848,N_5552,N_5699);
or U5849 (N_5849,N_5590,N_5584);
xor U5850 (N_5850,N_5724,N_5820);
or U5851 (N_5851,N_5754,N_5792);
xor U5852 (N_5852,N_5725,N_5824);
xnor U5853 (N_5853,N_5746,N_5778);
or U5854 (N_5854,N_5809,N_5702);
nor U5855 (N_5855,N_5729,N_5831);
nand U5856 (N_5856,N_5737,N_5722);
nor U5857 (N_5857,N_5848,N_5711);
and U5858 (N_5858,N_5753,N_5757);
xnor U5859 (N_5859,N_5841,N_5706);
and U5860 (N_5860,N_5822,N_5721);
xor U5861 (N_5861,N_5821,N_5832);
xor U5862 (N_5862,N_5780,N_5811);
or U5863 (N_5863,N_5783,N_5715);
and U5864 (N_5864,N_5731,N_5834);
and U5865 (N_5865,N_5723,N_5843);
and U5866 (N_5866,N_5726,N_5703);
and U5867 (N_5867,N_5713,N_5798);
xor U5868 (N_5868,N_5768,N_5714);
nor U5869 (N_5869,N_5829,N_5733);
or U5870 (N_5870,N_5741,N_5847);
nor U5871 (N_5871,N_5838,N_5787);
or U5872 (N_5872,N_5727,N_5817);
or U5873 (N_5873,N_5794,N_5769);
and U5874 (N_5874,N_5779,N_5846);
xnor U5875 (N_5875,N_5774,N_5804);
xor U5876 (N_5876,N_5710,N_5799);
and U5877 (N_5877,N_5776,N_5717);
or U5878 (N_5878,N_5803,N_5755);
and U5879 (N_5879,N_5819,N_5839);
nand U5880 (N_5880,N_5815,N_5795);
and U5881 (N_5881,N_5771,N_5782);
xor U5882 (N_5882,N_5813,N_5718);
or U5883 (N_5883,N_5784,N_5766);
nand U5884 (N_5884,N_5770,N_5788);
xor U5885 (N_5885,N_5700,N_5767);
or U5886 (N_5886,N_5738,N_5775);
xnor U5887 (N_5887,N_5801,N_5818);
or U5888 (N_5888,N_5742,N_5734);
and U5889 (N_5889,N_5840,N_5772);
xnor U5890 (N_5890,N_5719,N_5827);
xor U5891 (N_5891,N_5751,N_5762);
nor U5892 (N_5892,N_5773,N_5743);
xnor U5893 (N_5893,N_5793,N_5777);
and U5894 (N_5894,N_5705,N_5740);
nor U5895 (N_5895,N_5752,N_5806);
nor U5896 (N_5896,N_5761,N_5844);
xor U5897 (N_5897,N_5786,N_5797);
xor U5898 (N_5898,N_5790,N_5730);
nor U5899 (N_5899,N_5744,N_5732);
nor U5900 (N_5900,N_5802,N_5745);
or U5901 (N_5901,N_5759,N_5764);
and U5902 (N_5902,N_5739,N_5736);
xor U5903 (N_5903,N_5835,N_5748);
and U5904 (N_5904,N_5785,N_5765);
or U5905 (N_5905,N_5750,N_5707);
and U5906 (N_5906,N_5716,N_5720);
or U5907 (N_5907,N_5781,N_5796);
nor U5908 (N_5908,N_5747,N_5816);
and U5909 (N_5909,N_5763,N_5760);
or U5910 (N_5910,N_5708,N_5758);
and U5911 (N_5911,N_5842,N_5704);
nor U5912 (N_5912,N_5837,N_5826);
nand U5913 (N_5913,N_5709,N_5825);
or U5914 (N_5914,N_5800,N_5810);
xnor U5915 (N_5915,N_5808,N_5791);
xor U5916 (N_5916,N_5712,N_5845);
xor U5917 (N_5917,N_5728,N_5735);
or U5918 (N_5918,N_5830,N_5812);
nor U5919 (N_5919,N_5756,N_5833);
nand U5920 (N_5920,N_5807,N_5701);
or U5921 (N_5921,N_5828,N_5814);
xnor U5922 (N_5922,N_5805,N_5749);
xor U5923 (N_5923,N_5823,N_5789);
xnor U5924 (N_5924,N_5836,N_5849);
nor U5925 (N_5925,N_5713,N_5766);
and U5926 (N_5926,N_5738,N_5763);
xor U5927 (N_5927,N_5817,N_5736);
nand U5928 (N_5928,N_5816,N_5717);
and U5929 (N_5929,N_5708,N_5719);
and U5930 (N_5930,N_5746,N_5825);
and U5931 (N_5931,N_5739,N_5700);
nand U5932 (N_5932,N_5779,N_5826);
and U5933 (N_5933,N_5799,N_5844);
xnor U5934 (N_5934,N_5765,N_5773);
or U5935 (N_5935,N_5716,N_5738);
nand U5936 (N_5936,N_5728,N_5749);
and U5937 (N_5937,N_5704,N_5799);
xnor U5938 (N_5938,N_5795,N_5844);
nor U5939 (N_5939,N_5734,N_5733);
nand U5940 (N_5940,N_5733,N_5799);
nand U5941 (N_5941,N_5729,N_5828);
nand U5942 (N_5942,N_5808,N_5835);
or U5943 (N_5943,N_5733,N_5714);
nor U5944 (N_5944,N_5703,N_5757);
nand U5945 (N_5945,N_5719,N_5747);
and U5946 (N_5946,N_5811,N_5738);
nor U5947 (N_5947,N_5767,N_5717);
nand U5948 (N_5948,N_5840,N_5820);
and U5949 (N_5949,N_5777,N_5841);
nor U5950 (N_5950,N_5717,N_5812);
nor U5951 (N_5951,N_5784,N_5702);
xor U5952 (N_5952,N_5846,N_5732);
nor U5953 (N_5953,N_5754,N_5730);
and U5954 (N_5954,N_5803,N_5763);
xor U5955 (N_5955,N_5712,N_5759);
and U5956 (N_5956,N_5760,N_5786);
and U5957 (N_5957,N_5716,N_5768);
nand U5958 (N_5958,N_5815,N_5753);
or U5959 (N_5959,N_5792,N_5781);
nand U5960 (N_5960,N_5786,N_5785);
and U5961 (N_5961,N_5836,N_5714);
xor U5962 (N_5962,N_5831,N_5750);
and U5963 (N_5963,N_5807,N_5735);
nor U5964 (N_5964,N_5832,N_5717);
nand U5965 (N_5965,N_5779,N_5759);
and U5966 (N_5966,N_5766,N_5767);
nand U5967 (N_5967,N_5745,N_5782);
xnor U5968 (N_5968,N_5829,N_5794);
nor U5969 (N_5969,N_5819,N_5762);
and U5970 (N_5970,N_5840,N_5752);
or U5971 (N_5971,N_5761,N_5769);
xnor U5972 (N_5972,N_5739,N_5772);
xnor U5973 (N_5973,N_5734,N_5745);
nand U5974 (N_5974,N_5707,N_5768);
xnor U5975 (N_5975,N_5807,N_5740);
or U5976 (N_5976,N_5727,N_5820);
xnor U5977 (N_5977,N_5769,N_5749);
nand U5978 (N_5978,N_5745,N_5791);
xnor U5979 (N_5979,N_5802,N_5730);
nand U5980 (N_5980,N_5802,N_5807);
and U5981 (N_5981,N_5724,N_5824);
nand U5982 (N_5982,N_5778,N_5783);
or U5983 (N_5983,N_5776,N_5752);
and U5984 (N_5984,N_5832,N_5707);
nand U5985 (N_5985,N_5730,N_5847);
xnor U5986 (N_5986,N_5784,N_5764);
xor U5987 (N_5987,N_5753,N_5711);
nand U5988 (N_5988,N_5723,N_5834);
nand U5989 (N_5989,N_5720,N_5774);
nand U5990 (N_5990,N_5739,N_5759);
nor U5991 (N_5991,N_5820,N_5815);
or U5992 (N_5992,N_5755,N_5727);
and U5993 (N_5993,N_5831,N_5808);
and U5994 (N_5994,N_5839,N_5738);
or U5995 (N_5995,N_5711,N_5728);
nand U5996 (N_5996,N_5749,N_5778);
and U5997 (N_5997,N_5747,N_5790);
xnor U5998 (N_5998,N_5721,N_5849);
nor U5999 (N_5999,N_5708,N_5759);
nor U6000 (N_6000,N_5967,N_5916);
nand U6001 (N_6001,N_5866,N_5982);
xor U6002 (N_6002,N_5968,N_5922);
or U6003 (N_6003,N_5964,N_5981);
nand U6004 (N_6004,N_5954,N_5986);
nor U6005 (N_6005,N_5972,N_5929);
and U6006 (N_6006,N_5991,N_5868);
xor U6007 (N_6007,N_5927,N_5897);
nand U6008 (N_6008,N_5860,N_5978);
xnor U6009 (N_6009,N_5975,N_5898);
and U6010 (N_6010,N_5990,N_5886);
or U6011 (N_6011,N_5891,N_5935);
nand U6012 (N_6012,N_5977,N_5883);
nand U6013 (N_6013,N_5948,N_5874);
and U6014 (N_6014,N_5920,N_5885);
and U6015 (N_6015,N_5933,N_5973);
xnor U6016 (N_6016,N_5934,N_5942);
nand U6017 (N_6017,N_5931,N_5987);
nor U6018 (N_6018,N_5884,N_5945);
nand U6019 (N_6019,N_5992,N_5899);
and U6020 (N_6020,N_5867,N_5900);
nor U6021 (N_6021,N_5993,N_5914);
and U6022 (N_6022,N_5923,N_5877);
xnor U6023 (N_6023,N_5869,N_5911);
nand U6024 (N_6024,N_5984,N_5994);
or U6025 (N_6025,N_5949,N_5937);
xnor U6026 (N_6026,N_5976,N_5940);
or U6027 (N_6027,N_5960,N_5952);
xor U6028 (N_6028,N_5851,N_5974);
and U6029 (N_6029,N_5999,N_5958);
and U6030 (N_6030,N_5928,N_5996);
or U6031 (N_6031,N_5910,N_5896);
nand U6032 (N_6032,N_5893,N_5907);
xor U6033 (N_6033,N_5962,N_5998);
and U6034 (N_6034,N_5957,N_5895);
nor U6035 (N_6035,N_5915,N_5947);
or U6036 (N_6036,N_5950,N_5863);
or U6037 (N_6037,N_5901,N_5862);
xor U6038 (N_6038,N_5989,N_5983);
or U6039 (N_6039,N_5985,N_5970);
nor U6040 (N_6040,N_5938,N_5889);
or U6041 (N_6041,N_5906,N_5941);
xor U6042 (N_6042,N_5879,N_5882);
and U6043 (N_6043,N_5857,N_5888);
nand U6044 (N_6044,N_5953,N_5850);
xor U6045 (N_6045,N_5925,N_5959);
and U6046 (N_6046,N_5939,N_5873);
nand U6047 (N_6047,N_5890,N_5870);
and U6048 (N_6048,N_5909,N_5887);
nand U6049 (N_6049,N_5965,N_5852);
or U6050 (N_6050,N_5944,N_5971);
and U6051 (N_6051,N_5858,N_5904);
nand U6052 (N_6052,N_5912,N_5913);
nand U6053 (N_6053,N_5865,N_5936);
or U6054 (N_6054,N_5864,N_5963);
nor U6055 (N_6055,N_5854,N_5997);
nand U6056 (N_6056,N_5903,N_5892);
xor U6057 (N_6057,N_5871,N_5979);
and U6058 (N_6058,N_5861,N_5988);
nand U6059 (N_6059,N_5951,N_5946);
nor U6060 (N_6060,N_5917,N_5955);
or U6061 (N_6061,N_5995,N_5853);
nand U6062 (N_6062,N_5918,N_5878);
or U6063 (N_6063,N_5905,N_5926);
nand U6064 (N_6064,N_5980,N_5856);
nand U6065 (N_6065,N_5969,N_5966);
xnor U6066 (N_6066,N_5876,N_5956);
nand U6067 (N_6067,N_5881,N_5902);
or U6068 (N_6068,N_5943,N_5855);
xnor U6069 (N_6069,N_5919,N_5872);
xnor U6070 (N_6070,N_5880,N_5961);
or U6071 (N_6071,N_5921,N_5930);
or U6072 (N_6072,N_5932,N_5875);
nand U6073 (N_6073,N_5908,N_5859);
and U6074 (N_6074,N_5924,N_5894);
nor U6075 (N_6075,N_5936,N_5899);
or U6076 (N_6076,N_5962,N_5913);
nand U6077 (N_6077,N_5872,N_5959);
and U6078 (N_6078,N_5921,N_5977);
and U6079 (N_6079,N_5936,N_5941);
nand U6080 (N_6080,N_5947,N_5946);
nor U6081 (N_6081,N_5986,N_5908);
nor U6082 (N_6082,N_5911,N_5948);
xor U6083 (N_6083,N_5858,N_5943);
or U6084 (N_6084,N_5940,N_5921);
nor U6085 (N_6085,N_5968,N_5884);
nand U6086 (N_6086,N_5908,N_5985);
xnor U6087 (N_6087,N_5933,N_5978);
nor U6088 (N_6088,N_5891,N_5968);
and U6089 (N_6089,N_5860,N_5987);
xnor U6090 (N_6090,N_5893,N_5946);
and U6091 (N_6091,N_5973,N_5904);
and U6092 (N_6092,N_5924,N_5883);
or U6093 (N_6093,N_5920,N_5871);
or U6094 (N_6094,N_5869,N_5885);
and U6095 (N_6095,N_5899,N_5931);
xor U6096 (N_6096,N_5955,N_5918);
xor U6097 (N_6097,N_5883,N_5855);
nand U6098 (N_6098,N_5962,N_5894);
nand U6099 (N_6099,N_5980,N_5926);
or U6100 (N_6100,N_5971,N_5909);
or U6101 (N_6101,N_5948,N_5962);
nand U6102 (N_6102,N_5963,N_5940);
nor U6103 (N_6103,N_5951,N_5880);
nor U6104 (N_6104,N_5991,N_5947);
xor U6105 (N_6105,N_5883,N_5885);
nor U6106 (N_6106,N_5888,N_5990);
xnor U6107 (N_6107,N_5921,N_5953);
xnor U6108 (N_6108,N_5911,N_5910);
nor U6109 (N_6109,N_5992,N_5860);
nand U6110 (N_6110,N_5908,N_5923);
or U6111 (N_6111,N_5944,N_5976);
xnor U6112 (N_6112,N_5920,N_5911);
and U6113 (N_6113,N_5896,N_5999);
or U6114 (N_6114,N_5919,N_5924);
or U6115 (N_6115,N_5940,N_5917);
nor U6116 (N_6116,N_5970,N_5962);
nor U6117 (N_6117,N_5866,N_5874);
or U6118 (N_6118,N_5890,N_5925);
xor U6119 (N_6119,N_5887,N_5968);
or U6120 (N_6120,N_5999,N_5991);
or U6121 (N_6121,N_5969,N_5942);
nand U6122 (N_6122,N_5969,N_5950);
or U6123 (N_6123,N_5867,N_5986);
and U6124 (N_6124,N_5921,N_5945);
or U6125 (N_6125,N_5911,N_5956);
or U6126 (N_6126,N_5918,N_5915);
nor U6127 (N_6127,N_5936,N_5870);
nor U6128 (N_6128,N_5957,N_5922);
and U6129 (N_6129,N_5852,N_5983);
xor U6130 (N_6130,N_5873,N_5979);
or U6131 (N_6131,N_5952,N_5956);
nand U6132 (N_6132,N_5944,N_5967);
or U6133 (N_6133,N_5997,N_5945);
and U6134 (N_6134,N_5909,N_5852);
nor U6135 (N_6135,N_5855,N_5940);
nand U6136 (N_6136,N_5927,N_5922);
or U6137 (N_6137,N_5955,N_5957);
nor U6138 (N_6138,N_5976,N_5860);
nor U6139 (N_6139,N_5898,N_5927);
nor U6140 (N_6140,N_5867,N_5933);
nor U6141 (N_6141,N_5972,N_5903);
nor U6142 (N_6142,N_5850,N_5933);
and U6143 (N_6143,N_5858,N_5886);
or U6144 (N_6144,N_5902,N_5927);
or U6145 (N_6145,N_5977,N_5919);
nand U6146 (N_6146,N_5892,N_5928);
and U6147 (N_6147,N_5864,N_5980);
and U6148 (N_6148,N_5978,N_5903);
xnor U6149 (N_6149,N_5938,N_5910);
and U6150 (N_6150,N_6070,N_6025);
nand U6151 (N_6151,N_6126,N_6086);
nor U6152 (N_6152,N_6013,N_6038);
xnor U6153 (N_6153,N_6137,N_6135);
or U6154 (N_6154,N_6067,N_6011);
nand U6155 (N_6155,N_6015,N_6007);
or U6156 (N_6156,N_6010,N_6099);
and U6157 (N_6157,N_6064,N_6050);
or U6158 (N_6158,N_6029,N_6016);
xnor U6159 (N_6159,N_6018,N_6049);
nor U6160 (N_6160,N_6066,N_6083);
xnor U6161 (N_6161,N_6035,N_6096);
nand U6162 (N_6162,N_6109,N_6047);
and U6163 (N_6163,N_6146,N_6044);
nor U6164 (N_6164,N_6001,N_6118);
and U6165 (N_6165,N_6002,N_6115);
or U6166 (N_6166,N_6054,N_6012);
nand U6167 (N_6167,N_6143,N_6131);
nand U6168 (N_6168,N_6021,N_6114);
nor U6169 (N_6169,N_6072,N_6142);
and U6170 (N_6170,N_6125,N_6145);
and U6171 (N_6171,N_6149,N_6017);
nand U6172 (N_6172,N_6073,N_6004);
or U6173 (N_6173,N_6101,N_6034);
or U6174 (N_6174,N_6023,N_6055);
nand U6175 (N_6175,N_6046,N_6030);
and U6176 (N_6176,N_6090,N_6121);
and U6177 (N_6177,N_6059,N_6130);
nor U6178 (N_6178,N_6092,N_6129);
and U6179 (N_6179,N_6048,N_6019);
or U6180 (N_6180,N_6144,N_6009);
or U6181 (N_6181,N_6033,N_6141);
nand U6182 (N_6182,N_6040,N_6106);
and U6183 (N_6183,N_6043,N_6133);
or U6184 (N_6184,N_6039,N_6108);
or U6185 (N_6185,N_6102,N_6031);
nor U6186 (N_6186,N_6136,N_6078);
or U6187 (N_6187,N_6091,N_6095);
xnor U6188 (N_6188,N_6085,N_6022);
and U6189 (N_6189,N_6127,N_6062);
nand U6190 (N_6190,N_6024,N_6051);
and U6191 (N_6191,N_6061,N_6113);
nor U6192 (N_6192,N_6110,N_6116);
and U6193 (N_6193,N_6005,N_6063);
or U6194 (N_6194,N_6105,N_6076);
nor U6195 (N_6195,N_6088,N_6100);
xnor U6196 (N_6196,N_6053,N_6000);
nand U6197 (N_6197,N_6148,N_6068);
or U6198 (N_6198,N_6094,N_6060);
or U6199 (N_6199,N_6120,N_6074);
xnor U6200 (N_6200,N_6071,N_6057);
nand U6201 (N_6201,N_6107,N_6028);
and U6202 (N_6202,N_6077,N_6003);
nand U6203 (N_6203,N_6140,N_6014);
nand U6204 (N_6204,N_6032,N_6079);
nor U6205 (N_6205,N_6134,N_6139);
and U6206 (N_6206,N_6080,N_6097);
and U6207 (N_6207,N_6036,N_6132);
and U6208 (N_6208,N_6041,N_6065);
nand U6209 (N_6209,N_6104,N_6112);
or U6210 (N_6210,N_6084,N_6069);
or U6211 (N_6211,N_6026,N_6058);
xnor U6212 (N_6212,N_6081,N_6056);
xor U6213 (N_6213,N_6042,N_6119);
xnor U6214 (N_6214,N_6087,N_6020);
and U6215 (N_6215,N_6093,N_6006);
or U6216 (N_6216,N_6075,N_6117);
nor U6217 (N_6217,N_6037,N_6138);
or U6218 (N_6218,N_6027,N_6111);
and U6219 (N_6219,N_6052,N_6045);
nand U6220 (N_6220,N_6122,N_6008);
nor U6221 (N_6221,N_6123,N_6124);
nand U6222 (N_6222,N_6128,N_6098);
and U6223 (N_6223,N_6103,N_6147);
nand U6224 (N_6224,N_6089,N_6082);
xnor U6225 (N_6225,N_6103,N_6063);
or U6226 (N_6226,N_6081,N_6064);
nor U6227 (N_6227,N_6006,N_6019);
xnor U6228 (N_6228,N_6015,N_6126);
or U6229 (N_6229,N_6037,N_6062);
nor U6230 (N_6230,N_6048,N_6100);
nor U6231 (N_6231,N_6070,N_6036);
nor U6232 (N_6232,N_6144,N_6038);
xor U6233 (N_6233,N_6063,N_6059);
nor U6234 (N_6234,N_6013,N_6005);
or U6235 (N_6235,N_6068,N_6006);
nor U6236 (N_6236,N_6034,N_6144);
nor U6237 (N_6237,N_6043,N_6021);
or U6238 (N_6238,N_6099,N_6054);
nor U6239 (N_6239,N_6081,N_6011);
xor U6240 (N_6240,N_6073,N_6104);
nand U6241 (N_6241,N_6009,N_6033);
nor U6242 (N_6242,N_6049,N_6034);
xnor U6243 (N_6243,N_6117,N_6120);
or U6244 (N_6244,N_6025,N_6127);
nor U6245 (N_6245,N_6116,N_6134);
xor U6246 (N_6246,N_6108,N_6010);
xnor U6247 (N_6247,N_6044,N_6121);
nor U6248 (N_6248,N_6031,N_6081);
xor U6249 (N_6249,N_6046,N_6073);
or U6250 (N_6250,N_6147,N_6149);
or U6251 (N_6251,N_6055,N_6102);
nor U6252 (N_6252,N_6001,N_6060);
nand U6253 (N_6253,N_6051,N_6014);
nand U6254 (N_6254,N_6030,N_6144);
nand U6255 (N_6255,N_6127,N_6058);
nor U6256 (N_6256,N_6086,N_6098);
nand U6257 (N_6257,N_6114,N_6077);
and U6258 (N_6258,N_6101,N_6130);
or U6259 (N_6259,N_6060,N_6076);
or U6260 (N_6260,N_6114,N_6136);
and U6261 (N_6261,N_6038,N_6047);
nand U6262 (N_6262,N_6016,N_6110);
or U6263 (N_6263,N_6074,N_6105);
xnor U6264 (N_6264,N_6072,N_6120);
and U6265 (N_6265,N_6047,N_6067);
nor U6266 (N_6266,N_6109,N_6057);
nand U6267 (N_6267,N_6016,N_6113);
or U6268 (N_6268,N_6063,N_6060);
and U6269 (N_6269,N_6016,N_6013);
nand U6270 (N_6270,N_6070,N_6128);
xnor U6271 (N_6271,N_6043,N_6052);
nor U6272 (N_6272,N_6145,N_6065);
xor U6273 (N_6273,N_6100,N_6083);
nor U6274 (N_6274,N_6104,N_6059);
xnor U6275 (N_6275,N_6064,N_6120);
nand U6276 (N_6276,N_6068,N_6127);
or U6277 (N_6277,N_6117,N_6014);
nand U6278 (N_6278,N_6015,N_6117);
nand U6279 (N_6279,N_6117,N_6083);
xor U6280 (N_6280,N_6000,N_6086);
nor U6281 (N_6281,N_6141,N_6007);
or U6282 (N_6282,N_6089,N_6076);
and U6283 (N_6283,N_6140,N_6139);
nand U6284 (N_6284,N_6011,N_6128);
nor U6285 (N_6285,N_6120,N_6012);
nand U6286 (N_6286,N_6043,N_6068);
nor U6287 (N_6287,N_6131,N_6093);
and U6288 (N_6288,N_6000,N_6074);
xnor U6289 (N_6289,N_6111,N_6055);
and U6290 (N_6290,N_6109,N_6105);
nand U6291 (N_6291,N_6020,N_6000);
or U6292 (N_6292,N_6088,N_6046);
xnor U6293 (N_6293,N_6117,N_6105);
and U6294 (N_6294,N_6074,N_6102);
or U6295 (N_6295,N_6141,N_6100);
nor U6296 (N_6296,N_6137,N_6091);
and U6297 (N_6297,N_6142,N_6087);
nand U6298 (N_6298,N_6127,N_6099);
nor U6299 (N_6299,N_6080,N_6115);
nand U6300 (N_6300,N_6283,N_6295);
or U6301 (N_6301,N_6236,N_6221);
and U6302 (N_6302,N_6237,N_6177);
xnor U6303 (N_6303,N_6269,N_6279);
nor U6304 (N_6304,N_6262,N_6153);
or U6305 (N_6305,N_6179,N_6292);
nor U6306 (N_6306,N_6233,N_6247);
nand U6307 (N_6307,N_6263,N_6214);
or U6308 (N_6308,N_6175,N_6248);
and U6309 (N_6309,N_6165,N_6245);
nand U6310 (N_6310,N_6171,N_6272);
nor U6311 (N_6311,N_6257,N_6297);
and U6312 (N_6312,N_6244,N_6216);
nor U6313 (N_6313,N_6170,N_6241);
xor U6314 (N_6314,N_6189,N_6169);
xnor U6315 (N_6315,N_6256,N_6196);
or U6316 (N_6316,N_6222,N_6178);
nand U6317 (N_6317,N_6265,N_6215);
and U6318 (N_6318,N_6194,N_6249);
xnor U6319 (N_6319,N_6151,N_6229);
or U6320 (N_6320,N_6186,N_6208);
or U6321 (N_6321,N_6240,N_6299);
or U6322 (N_6322,N_6288,N_6250);
nand U6323 (N_6323,N_6187,N_6289);
and U6324 (N_6324,N_6156,N_6238);
and U6325 (N_6325,N_6202,N_6173);
or U6326 (N_6326,N_6176,N_6264);
nand U6327 (N_6327,N_6282,N_6252);
or U6328 (N_6328,N_6191,N_6158);
xor U6329 (N_6329,N_6218,N_6205);
xnor U6330 (N_6330,N_6183,N_6155);
nand U6331 (N_6331,N_6152,N_6164);
nor U6332 (N_6332,N_6226,N_6168);
nand U6333 (N_6333,N_6174,N_6296);
and U6334 (N_6334,N_6200,N_6231);
xnor U6335 (N_6335,N_6217,N_6284);
and U6336 (N_6336,N_6286,N_6150);
and U6337 (N_6337,N_6277,N_6246);
or U6338 (N_6338,N_6162,N_6172);
and U6339 (N_6339,N_6223,N_6157);
xor U6340 (N_6340,N_6207,N_6239);
nand U6341 (N_6341,N_6224,N_6180);
and U6342 (N_6342,N_6161,N_6273);
xor U6343 (N_6343,N_6227,N_6213);
or U6344 (N_6344,N_6259,N_6235);
or U6345 (N_6345,N_6285,N_6181);
and U6346 (N_6346,N_6210,N_6290);
nor U6347 (N_6347,N_6192,N_6188);
nand U6348 (N_6348,N_6209,N_6298);
xnor U6349 (N_6349,N_6254,N_6190);
or U6350 (N_6350,N_6159,N_6291);
nor U6351 (N_6351,N_6182,N_6267);
nor U6352 (N_6352,N_6278,N_6225);
nand U6353 (N_6353,N_6275,N_6185);
nand U6354 (N_6354,N_6204,N_6266);
nand U6355 (N_6355,N_6228,N_6163);
or U6356 (N_6356,N_6234,N_6203);
or U6357 (N_6357,N_6167,N_6206);
and U6358 (N_6358,N_6287,N_6197);
and U6359 (N_6359,N_6255,N_6198);
nand U6360 (N_6360,N_6258,N_6160);
nor U6361 (N_6361,N_6251,N_6260);
and U6362 (N_6362,N_6211,N_6154);
nand U6363 (N_6363,N_6199,N_6230);
xor U6364 (N_6364,N_6212,N_6184);
nor U6365 (N_6365,N_6293,N_6195);
and U6366 (N_6366,N_6253,N_6274);
xor U6367 (N_6367,N_6261,N_6281);
nand U6368 (N_6368,N_6276,N_6271);
xor U6369 (N_6369,N_6270,N_6219);
or U6370 (N_6370,N_6232,N_6243);
or U6371 (N_6371,N_6294,N_6242);
nor U6372 (N_6372,N_6201,N_6166);
and U6373 (N_6373,N_6268,N_6280);
nor U6374 (N_6374,N_6220,N_6193);
nand U6375 (N_6375,N_6201,N_6232);
and U6376 (N_6376,N_6232,N_6200);
and U6377 (N_6377,N_6192,N_6213);
nand U6378 (N_6378,N_6273,N_6152);
nor U6379 (N_6379,N_6269,N_6280);
nor U6380 (N_6380,N_6288,N_6223);
or U6381 (N_6381,N_6275,N_6257);
xor U6382 (N_6382,N_6241,N_6260);
nor U6383 (N_6383,N_6262,N_6266);
and U6384 (N_6384,N_6189,N_6183);
nor U6385 (N_6385,N_6283,N_6278);
nor U6386 (N_6386,N_6255,N_6268);
xnor U6387 (N_6387,N_6264,N_6297);
nand U6388 (N_6388,N_6219,N_6207);
nand U6389 (N_6389,N_6250,N_6193);
and U6390 (N_6390,N_6261,N_6191);
nand U6391 (N_6391,N_6176,N_6299);
xnor U6392 (N_6392,N_6253,N_6213);
and U6393 (N_6393,N_6192,N_6214);
or U6394 (N_6394,N_6197,N_6185);
xor U6395 (N_6395,N_6251,N_6220);
nand U6396 (N_6396,N_6296,N_6230);
xnor U6397 (N_6397,N_6284,N_6280);
nand U6398 (N_6398,N_6229,N_6271);
nor U6399 (N_6399,N_6260,N_6291);
or U6400 (N_6400,N_6191,N_6228);
nor U6401 (N_6401,N_6262,N_6226);
and U6402 (N_6402,N_6205,N_6179);
nor U6403 (N_6403,N_6296,N_6165);
nor U6404 (N_6404,N_6156,N_6288);
nor U6405 (N_6405,N_6222,N_6169);
xor U6406 (N_6406,N_6203,N_6291);
xnor U6407 (N_6407,N_6226,N_6298);
xor U6408 (N_6408,N_6250,N_6261);
xor U6409 (N_6409,N_6223,N_6272);
or U6410 (N_6410,N_6297,N_6286);
xor U6411 (N_6411,N_6253,N_6259);
and U6412 (N_6412,N_6196,N_6179);
nor U6413 (N_6413,N_6243,N_6299);
xor U6414 (N_6414,N_6181,N_6150);
and U6415 (N_6415,N_6167,N_6276);
and U6416 (N_6416,N_6171,N_6238);
xor U6417 (N_6417,N_6281,N_6232);
nand U6418 (N_6418,N_6208,N_6241);
xnor U6419 (N_6419,N_6204,N_6182);
or U6420 (N_6420,N_6242,N_6197);
xnor U6421 (N_6421,N_6211,N_6162);
xnor U6422 (N_6422,N_6242,N_6198);
nand U6423 (N_6423,N_6207,N_6253);
or U6424 (N_6424,N_6255,N_6295);
or U6425 (N_6425,N_6212,N_6200);
or U6426 (N_6426,N_6264,N_6170);
and U6427 (N_6427,N_6254,N_6221);
and U6428 (N_6428,N_6196,N_6284);
nand U6429 (N_6429,N_6154,N_6165);
nand U6430 (N_6430,N_6272,N_6167);
nor U6431 (N_6431,N_6261,N_6214);
xnor U6432 (N_6432,N_6229,N_6177);
nand U6433 (N_6433,N_6236,N_6162);
nand U6434 (N_6434,N_6202,N_6179);
and U6435 (N_6435,N_6292,N_6157);
nor U6436 (N_6436,N_6250,N_6251);
xor U6437 (N_6437,N_6176,N_6189);
and U6438 (N_6438,N_6167,N_6287);
and U6439 (N_6439,N_6223,N_6262);
nor U6440 (N_6440,N_6249,N_6290);
and U6441 (N_6441,N_6227,N_6196);
or U6442 (N_6442,N_6260,N_6228);
nand U6443 (N_6443,N_6235,N_6192);
or U6444 (N_6444,N_6160,N_6157);
and U6445 (N_6445,N_6211,N_6202);
nor U6446 (N_6446,N_6188,N_6232);
and U6447 (N_6447,N_6162,N_6246);
xor U6448 (N_6448,N_6299,N_6241);
or U6449 (N_6449,N_6169,N_6291);
nor U6450 (N_6450,N_6423,N_6303);
nand U6451 (N_6451,N_6430,N_6422);
nor U6452 (N_6452,N_6406,N_6304);
and U6453 (N_6453,N_6443,N_6447);
and U6454 (N_6454,N_6433,N_6344);
nand U6455 (N_6455,N_6311,N_6431);
nor U6456 (N_6456,N_6347,N_6320);
nor U6457 (N_6457,N_6338,N_6398);
xnor U6458 (N_6458,N_6389,N_6315);
xor U6459 (N_6459,N_6381,N_6400);
nand U6460 (N_6460,N_6333,N_6355);
nor U6461 (N_6461,N_6441,N_6301);
nand U6462 (N_6462,N_6378,N_6349);
nor U6463 (N_6463,N_6409,N_6343);
and U6464 (N_6464,N_6421,N_6382);
or U6465 (N_6465,N_6438,N_6385);
nor U6466 (N_6466,N_6387,N_6354);
nand U6467 (N_6467,N_6312,N_6351);
or U6468 (N_6468,N_6346,N_6405);
or U6469 (N_6469,N_6370,N_6436);
nand U6470 (N_6470,N_6363,N_6313);
or U6471 (N_6471,N_6439,N_6377);
xor U6472 (N_6472,N_6413,N_6371);
xnor U6473 (N_6473,N_6364,N_6330);
nand U6474 (N_6474,N_6305,N_6309);
or U6475 (N_6475,N_6306,N_6420);
xnor U6476 (N_6476,N_6345,N_6324);
nor U6477 (N_6477,N_6412,N_6392);
xnor U6478 (N_6478,N_6322,N_6310);
nor U6479 (N_6479,N_6339,N_6327);
or U6480 (N_6480,N_6359,N_6360);
nor U6481 (N_6481,N_6326,N_6318);
and U6482 (N_6482,N_6362,N_6367);
and U6483 (N_6483,N_6337,N_6300);
xor U6484 (N_6484,N_6384,N_6323);
nand U6485 (N_6485,N_6428,N_6314);
and U6486 (N_6486,N_6435,N_6341);
xnor U6487 (N_6487,N_6444,N_6336);
nor U6488 (N_6488,N_6434,N_6308);
nand U6489 (N_6489,N_6365,N_6368);
or U6490 (N_6490,N_6342,N_6448);
xor U6491 (N_6491,N_6325,N_6358);
xor U6492 (N_6492,N_6316,N_6429);
and U6493 (N_6493,N_6375,N_6395);
xnor U6494 (N_6494,N_6426,N_6376);
or U6495 (N_6495,N_6366,N_6383);
nand U6496 (N_6496,N_6414,N_6356);
xor U6497 (N_6497,N_6357,N_6393);
or U6498 (N_6498,N_6348,N_6374);
and U6499 (N_6499,N_6307,N_6399);
nor U6500 (N_6500,N_6379,N_6416);
nor U6501 (N_6501,N_6396,N_6334);
or U6502 (N_6502,N_6449,N_6390);
or U6503 (N_6503,N_6440,N_6361);
nor U6504 (N_6504,N_6302,N_6332);
xnor U6505 (N_6505,N_6394,N_6445);
nor U6506 (N_6506,N_6408,N_6419);
or U6507 (N_6507,N_6415,N_6319);
or U6508 (N_6508,N_6340,N_6391);
or U6509 (N_6509,N_6403,N_6424);
nor U6510 (N_6510,N_6352,N_6410);
or U6511 (N_6511,N_6386,N_6437);
and U6512 (N_6512,N_6417,N_6432);
nand U6513 (N_6513,N_6418,N_6401);
nand U6514 (N_6514,N_6411,N_6321);
or U6515 (N_6515,N_6397,N_6335);
nor U6516 (N_6516,N_6380,N_6373);
xor U6517 (N_6517,N_6402,N_6442);
xor U6518 (N_6518,N_6353,N_6369);
and U6519 (N_6519,N_6388,N_6407);
and U6520 (N_6520,N_6350,N_6331);
or U6521 (N_6521,N_6372,N_6329);
nor U6522 (N_6522,N_6404,N_6446);
and U6523 (N_6523,N_6425,N_6427);
nor U6524 (N_6524,N_6317,N_6328);
xor U6525 (N_6525,N_6442,N_6376);
and U6526 (N_6526,N_6366,N_6416);
nor U6527 (N_6527,N_6375,N_6437);
or U6528 (N_6528,N_6433,N_6436);
nor U6529 (N_6529,N_6424,N_6300);
or U6530 (N_6530,N_6328,N_6334);
xnor U6531 (N_6531,N_6339,N_6439);
and U6532 (N_6532,N_6416,N_6391);
and U6533 (N_6533,N_6331,N_6359);
and U6534 (N_6534,N_6325,N_6343);
xor U6535 (N_6535,N_6384,N_6391);
nor U6536 (N_6536,N_6391,N_6362);
nor U6537 (N_6537,N_6341,N_6420);
xnor U6538 (N_6538,N_6348,N_6339);
nor U6539 (N_6539,N_6436,N_6445);
nor U6540 (N_6540,N_6360,N_6383);
nor U6541 (N_6541,N_6335,N_6389);
nand U6542 (N_6542,N_6374,N_6340);
and U6543 (N_6543,N_6393,N_6300);
or U6544 (N_6544,N_6336,N_6367);
xnor U6545 (N_6545,N_6444,N_6357);
nand U6546 (N_6546,N_6304,N_6390);
or U6547 (N_6547,N_6300,N_6440);
and U6548 (N_6548,N_6357,N_6441);
and U6549 (N_6549,N_6424,N_6416);
nand U6550 (N_6550,N_6447,N_6420);
nor U6551 (N_6551,N_6306,N_6387);
nand U6552 (N_6552,N_6377,N_6337);
nor U6553 (N_6553,N_6331,N_6349);
or U6554 (N_6554,N_6342,N_6326);
nand U6555 (N_6555,N_6314,N_6396);
xor U6556 (N_6556,N_6425,N_6433);
nor U6557 (N_6557,N_6348,N_6417);
and U6558 (N_6558,N_6351,N_6424);
nand U6559 (N_6559,N_6421,N_6302);
xor U6560 (N_6560,N_6396,N_6356);
nand U6561 (N_6561,N_6395,N_6304);
nor U6562 (N_6562,N_6321,N_6425);
and U6563 (N_6563,N_6422,N_6361);
xor U6564 (N_6564,N_6447,N_6395);
xnor U6565 (N_6565,N_6365,N_6401);
nor U6566 (N_6566,N_6340,N_6439);
nand U6567 (N_6567,N_6404,N_6417);
nand U6568 (N_6568,N_6422,N_6353);
nor U6569 (N_6569,N_6320,N_6406);
nor U6570 (N_6570,N_6350,N_6408);
nor U6571 (N_6571,N_6316,N_6326);
nor U6572 (N_6572,N_6403,N_6356);
nand U6573 (N_6573,N_6330,N_6344);
nor U6574 (N_6574,N_6371,N_6385);
or U6575 (N_6575,N_6300,N_6426);
nor U6576 (N_6576,N_6360,N_6388);
xnor U6577 (N_6577,N_6348,N_6308);
or U6578 (N_6578,N_6418,N_6373);
nand U6579 (N_6579,N_6389,N_6371);
and U6580 (N_6580,N_6353,N_6366);
and U6581 (N_6581,N_6411,N_6337);
xnor U6582 (N_6582,N_6427,N_6440);
and U6583 (N_6583,N_6355,N_6424);
xnor U6584 (N_6584,N_6369,N_6364);
and U6585 (N_6585,N_6443,N_6406);
nor U6586 (N_6586,N_6373,N_6302);
xnor U6587 (N_6587,N_6363,N_6393);
nor U6588 (N_6588,N_6320,N_6307);
nand U6589 (N_6589,N_6372,N_6439);
nand U6590 (N_6590,N_6444,N_6330);
or U6591 (N_6591,N_6394,N_6343);
nor U6592 (N_6592,N_6314,N_6349);
or U6593 (N_6593,N_6398,N_6361);
nor U6594 (N_6594,N_6372,N_6397);
nor U6595 (N_6595,N_6421,N_6414);
or U6596 (N_6596,N_6418,N_6422);
xor U6597 (N_6597,N_6391,N_6369);
nand U6598 (N_6598,N_6366,N_6328);
and U6599 (N_6599,N_6337,N_6342);
nor U6600 (N_6600,N_6571,N_6562);
nand U6601 (N_6601,N_6503,N_6526);
nor U6602 (N_6602,N_6501,N_6461);
and U6603 (N_6603,N_6468,N_6467);
and U6604 (N_6604,N_6482,N_6545);
or U6605 (N_6605,N_6560,N_6491);
nand U6606 (N_6606,N_6579,N_6575);
nand U6607 (N_6607,N_6546,N_6540);
nand U6608 (N_6608,N_6553,N_6493);
nor U6609 (N_6609,N_6475,N_6597);
and U6610 (N_6610,N_6511,N_6578);
xnor U6611 (N_6611,N_6543,N_6478);
xor U6612 (N_6612,N_6515,N_6507);
nor U6613 (N_6613,N_6529,N_6498);
and U6614 (N_6614,N_6520,N_6470);
or U6615 (N_6615,N_6544,N_6476);
nand U6616 (N_6616,N_6554,N_6508);
nand U6617 (N_6617,N_6559,N_6487);
or U6618 (N_6618,N_6580,N_6466);
nand U6619 (N_6619,N_6492,N_6594);
nor U6620 (N_6620,N_6464,N_6458);
and U6621 (N_6621,N_6576,N_6518);
nor U6622 (N_6622,N_6586,N_6537);
and U6623 (N_6623,N_6506,N_6539);
nor U6624 (N_6624,N_6532,N_6598);
nand U6625 (N_6625,N_6552,N_6499);
or U6626 (N_6626,N_6463,N_6460);
nand U6627 (N_6627,N_6523,N_6457);
or U6628 (N_6628,N_6516,N_6484);
nand U6629 (N_6629,N_6572,N_6531);
xnor U6630 (N_6630,N_6533,N_6509);
and U6631 (N_6631,N_6477,N_6556);
or U6632 (N_6632,N_6459,N_6517);
and U6633 (N_6633,N_6500,N_6558);
xnor U6634 (N_6634,N_6455,N_6521);
xor U6635 (N_6635,N_6599,N_6592);
xnor U6636 (N_6636,N_6569,N_6583);
xnor U6637 (N_6637,N_6547,N_6590);
xnor U6638 (N_6638,N_6538,N_6452);
nor U6639 (N_6639,N_6469,N_6564);
nor U6640 (N_6640,N_6595,N_6502);
xor U6641 (N_6641,N_6584,N_6534);
and U6642 (N_6642,N_6550,N_6485);
or U6643 (N_6643,N_6587,N_6591);
xnor U6644 (N_6644,N_6574,N_6541);
and U6645 (N_6645,N_6483,N_6514);
or U6646 (N_6646,N_6549,N_6593);
nor U6647 (N_6647,N_6462,N_6504);
or U6648 (N_6648,N_6596,N_6454);
nand U6649 (N_6649,N_6474,N_6530);
and U6650 (N_6650,N_6585,N_6570);
nand U6651 (N_6651,N_6565,N_6573);
nor U6652 (N_6652,N_6519,N_6465);
nand U6653 (N_6653,N_6490,N_6488);
or U6654 (N_6654,N_6557,N_6528);
nor U6655 (N_6655,N_6536,N_6456);
and U6656 (N_6656,N_6567,N_6563);
and U6657 (N_6657,N_6561,N_6566);
and U6658 (N_6658,N_6480,N_6486);
nand U6659 (N_6659,N_6588,N_6568);
nand U6660 (N_6660,N_6473,N_6471);
xnor U6661 (N_6661,N_6555,N_6522);
nand U6662 (N_6662,N_6510,N_6551);
nor U6663 (N_6663,N_6451,N_6527);
nand U6664 (N_6664,N_6496,N_6548);
xor U6665 (N_6665,N_6472,N_6497);
nand U6666 (N_6666,N_6582,N_6535);
and U6667 (N_6667,N_6495,N_6542);
nand U6668 (N_6668,N_6494,N_6512);
and U6669 (N_6669,N_6513,N_6505);
nor U6670 (N_6670,N_6453,N_6581);
nand U6671 (N_6671,N_6525,N_6577);
and U6672 (N_6672,N_6589,N_6524);
nor U6673 (N_6673,N_6479,N_6481);
nand U6674 (N_6674,N_6489,N_6450);
nand U6675 (N_6675,N_6482,N_6522);
and U6676 (N_6676,N_6566,N_6460);
and U6677 (N_6677,N_6584,N_6545);
nand U6678 (N_6678,N_6569,N_6579);
nand U6679 (N_6679,N_6496,N_6499);
and U6680 (N_6680,N_6460,N_6556);
xor U6681 (N_6681,N_6571,N_6588);
and U6682 (N_6682,N_6487,N_6555);
xor U6683 (N_6683,N_6519,N_6521);
and U6684 (N_6684,N_6567,N_6514);
or U6685 (N_6685,N_6551,N_6486);
xnor U6686 (N_6686,N_6538,N_6489);
nand U6687 (N_6687,N_6532,N_6531);
and U6688 (N_6688,N_6463,N_6550);
and U6689 (N_6689,N_6462,N_6545);
and U6690 (N_6690,N_6586,N_6459);
nor U6691 (N_6691,N_6463,N_6506);
nor U6692 (N_6692,N_6510,N_6464);
and U6693 (N_6693,N_6563,N_6508);
nand U6694 (N_6694,N_6450,N_6546);
nor U6695 (N_6695,N_6594,N_6466);
nand U6696 (N_6696,N_6462,N_6585);
xnor U6697 (N_6697,N_6503,N_6591);
and U6698 (N_6698,N_6451,N_6471);
or U6699 (N_6699,N_6488,N_6528);
and U6700 (N_6700,N_6546,N_6550);
nand U6701 (N_6701,N_6471,N_6561);
and U6702 (N_6702,N_6547,N_6584);
xnor U6703 (N_6703,N_6535,N_6563);
xnor U6704 (N_6704,N_6472,N_6552);
or U6705 (N_6705,N_6452,N_6518);
nand U6706 (N_6706,N_6538,N_6567);
nor U6707 (N_6707,N_6481,N_6525);
nor U6708 (N_6708,N_6506,N_6579);
and U6709 (N_6709,N_6573,N_6464);
and U6710 (N_6710,N_6545,N_6563);
nor U6711 (N_6711,N_6457,N_6598);
xnor U6712 (N_6712,N_6595,N_6531);
nor U6713 (N_6713,N_6494,N_6468);
xnor U6714 (N_6714,N_6536,N_6573);
xor U6715 (N_6715,N_6480,N_6509);
nand U6716 (N_6716,N_6571,N_6516);
nor U6717 (N_6717,N_6506,N_6488);
nor U6718 (N_6718,N_6483,N_6591);
nand U6719 (N_6719,N_6545,N_6529);
or U6720 (N_6720,N_6501,N_6519);
nand U6721 (N_6721,N_6464,N_6587);
nand U6722 (N_6722,N_6456,N_6575);
nor U6723 (N_6723,N_6504,N_6540);
and U6724 (N_6724,N_6538,N_6553);
xnor U6725 (N_6725,N_6583,N_6475);
or U6726 (N_6726,N_6552,N_6498);
nand U6727 (N_6727,N_6488,N_6501);
and U6728 (N_6728,N_6471,N_6486);
and U6729 (N_6729,N_6577,N_6497);
or U6730 (N_6730,N_6502,N_6522);
nand U6731 (N_6731,N_6496,N_6535);
or U6732 (N_6732,N_6469,N_6535);
and U6733 (N_6733,N_6500,N_6571);
nand U6734 (N_6734,N_6579,N_6521);
nor U6735 (N_6735,N_6491,N_6498);
nor U6736 (N_6736,N_6519,N_6516);
and U6737 (N_6737,N_6585,N_6542);
and U6738 (N_6738,N_6514,N_6532);
and U6739 (N_6739,N_6529,N_6586);
nor U6740 (N_6740,N_6509,N_6498);
and U6741 (N_6741,N_6476,N_6466);
or U6742 (N_6742,N_6508,N_6507);
or U6743 (N_6743,N_6502,N_6494);
and U6744 (N_6744,N_6470,N_6519);
nand U6745 (N_6745,N_6515,N_6534);
xor U6746 (N_6746,N_6588,N_6491);
nand U6747 (N_6747,N_6569,N_6577);
or U6748 (N_6748,N_6480,N_6523);
nor U6749 (N_6749,N_6548,N_6491);
nor U6750 (N_6750,N_6610,N_6640);
or U6751 (N_6751,N_6708,N_6709);
nand U6752 (N_6752,N_6749,N_6647);
nand U6753 (N_6753,N_6734,N_6643);
nand U6754 (N_6754,N_6644,N_6724);
and U6755 (N_6755,N_6726,N_6690);
nand U6756 (N_6756,N_6639,N_6665);
nand U6757 (N_6757,N_6674,N_6682);
nand U6758 (N_6758,N_6613,N_6636);
and U6759 (N_6759,N_6646,N_6730);
nor U6760 (N_6760,N_6736,N_6687);
xor U6761 (N_6761,N_6660,N_6729);
or U6762 (N_6762,N_6655,N_6680);
xor U6763 (N_6763,N_6686,N_6629);
nand U6764 (N_6764,N_6676,N_6648);
nand U6765 (N_6765,N_6616,N_6635);
nand U6766 (N_6766,N_6735,N_6620);
nor U6767 (N_6767,N_6714,N_6723);
or U6768 (N_6768,N_6611,N_6684);
nand U6769 (N_6769,N_6657,N_6731);
xnor U6770 (N_6770,N_6642,N_6738);
xnor U6771 (N_6771,N_6626,N_6614);
nand U6772 (N_6772,N_6733,N_6727);
and U6773 (N_6773,N_6663,N_6630);
xor U6774 (N_6774,N_6710,N_6720);
or U6775 (N_6775,N_6671,N_6719);
xnor U6776 (N_6776,N_6740,N_6633);
and U6777 (N_6777,N_6741,N_6677);
or U6778 (N_6778,N_6668,N_6745);
nor U6779 (N_6779,N_6669,N_6716);
xor U6780 (N_6780,N_6624,N_6732);
and U6781 (N_6781,N_6623,N_6693);
and U6782 (N_6782,N_6600,N_6702);
nand U6783 (N_6783,N_6698,N_6696);
or U6784 (N_6784,N_6689,N_6707);
nor U6785 (N_6785,N_6743,N_6654);
nor U6786 (N_6786,N_6706,N_6737);
nor U6787 (N_6787,N_6603,N_6704);
or U6788 (N_6788,N_6747,N_6744);
or U6789 (N_6789,N_6746,N_6649);
nand U6790 (N_6790,N_6681,N_6670);
nor U6791 (N_6791,N_6748,N_6703);
and U6792 (N_6792,N_6664,N_6632);
nor U6793 (N_6793,N_6661,N_6675);
xnor U6794 (N_6794,N_6625,N_6617);
nor U6795 (N_6795,N_6673,N_6615);
nor U6796 (N_6796,N_6608,N_6695);
xnor U6797 (N_6797,N_6631,N_6725);
xnor U6798 (N_6798,N_6638,N_6622);
and U6799 (N_6799,N_6679,N_6658);
and U6800 (N_6800,N_6672,N_6742);
xor U6801 (N_6801,N_6666,N_6662);
nor U6802 (N_6802,N_6634,N_6712);
nor U6803 (N_6803,N_6605,N_6637);
xnor U6804 (N_6804,N_6721,N_6728);
xor U6805 (N_6805,N_6602,N_6645);
nand U6806 (N_6806,N_6717,N_6641);
xnor U6807 (N_6807,N_6678,N_6628);
and U6808 (N_6808,N_6601,N_6692);
or U6809 (N_6809,N_6694,N_6685);
xnor U6810 (N_6810,N_6722,N_6713);
or U6811 (N_6811,N_6604,N_6699);
nand U6812 (N_6812,N_6683,N_6656);
or U6813 (N_6813,N_6650,N_6651);
nor U6814 (N_6814,N_6607,N_6688);
nor U6815 (N_6815,N_6653,N_6705);
and U6816 (N_6816,N_6691,N_6718);
or U6817 (N_6817,N_6715,N_6697);
nand U6818 (N_6818,N_6667,N_6619);
nand U6819 (N_6819,N_6700,N_6612);
nand U6820 (N_6820,N_6711,N_6652);
nor U6821 (N_6821,N_6739,N_6621);
xnor U6822 (N_6822,N_6618,N_6701);
nand U6823 (N_6823,N_6609,N_6606);
nand U6824 (N_6824,N_6659,N_6627);
nor U6825 (N_6825,N_6663,N_6618);
xnor U6826 (N_6826,N_6647,N_6622);
and U6827 (N_6827,N_6744,N_6635);
or U6828 (N_6828,N_6689,N_6600);
or U6829 (N_6829,N_6666,N_6625);
and U6830 (N_6830,N_6632,N_6667);
nor U6831 (N_6831,N_6610,N_6688);
xor U6832 (N_6832,N_6719,N_6711);
or U6833 (N_6833,N_6666,N_6715);
nand U6834 (N_6834,N_6634,N_6607);
xnor U6835 (N_6835,N_6723,N_6718);
nand U6836 (N_6836,N_6745,N_6613);
xor U6837 (N_6837,N_6739,N_6724);
and U6838 (N_6838,N_6650,N_6744);
or U6839 (N_6839,N_6740,N_6641);
and U6840 (N_6840,N_6735,N_6689);
xnor U6841 (N_6841,N_6704,N_6692);
nand U6842 (N_6842,N_6681,N_6715);
or U6843 (N_6843,N_6713,N_6693);
nand U6844 (N_6844,N_6689,N_6725);
xnor U6845 (N_6845,N_6693,N_6688);
xnor U6846 (N_6846,N_6665,N_6605);
xnor U6847 (N_6847,N_6605,N_6612);
nor U6848 (N_6848,N_6645,N_6673);
and U6849 (N_6849,N_6725,N_6697);
and U6850 (N_6850,N_6735,N_6665);
xnor U6851 (N_6851,N_6699,N_6696);
nand U6852 (N_6852,N_6682,N_6720);
xnor U6853 (N_6853,N_6659,N_6731);
nand U6854 (N_6854,N_6609,N_6678);
or U6855 (N_6855,N_6601,N_6615);
nor U6856 (N_6856,N_6642,N_6746);
nand U6857 (N_6857,N_6655,N_6719);
nand U6858 (N_6858,N_6608,N_6659);
nor U6859 (N_6859,N_6705,N_6642);
nand U6860 (N_6860,N_6707,N_6654);
xor U6861 (N_6861,N_6642,N_6605);
and U6862 (N_6862,N_6742,N_6671);
and U6863 (N_6863,N_6748,N_6606);
or U6864 (N_6864,N_6640,N_6742);
or U6865 (N_6865,N_6624,N_6600);
or U6866 (N_6866,N_6632,N_6622);
nand U6867 (N_6867,N_6692,N_6730);
nor U6868 (N_6868,N_6644,N_6746);
nand U6869 (N_6869,N_6639,N_6632);
and U6870 (N_6870,N_6693,N_6606);
or U6871 (N_6871,N_6687,N_6749);
xnor U6872 (N_6872,N_6646,N_6721);
nor U6873 (N_6873,N_6694,N_6706);
or U6874 (N_6874,N_6726,N_6694);
nor U6875 (N_6875,N_6691,N_6703);
nor U6876 (N_6876,N_6671,N_6604);
nor U6877 (N_6877,N_6654,N_6727);
nand U6878 (N_6878,N_6733,N_6654);
nand U6879 (N_6879,N_6724,N_6617);
and U6880 (N_6880,N_6622,N_6726);
nand U6881 (N_6881,N_6694,N_6658);
and U6882 (N_6882,N_6653,N_6706);
nand U6883 (N_6883,N_6682,N_6723);
nand U6884 (N_6884,N_6639,N_6737);
or U6885 (N_6885,N_6615,N_6690);
xor U6886 (N_6886,N_6625,N_6681);
nand U6887 (N_6887,N_6702,N_6603);
or U6888 (N_6888,N_6717,N_6653);
or U6889 (N_6889,N_6683,N_6711);
and U6890 (N_6890,N_6736,N_6688);
and U6891 (N_6891,N_6678,N_6696);
nand U6892 (N_6892,N_6687,N_6677);
or U6893 (N_6893,N_6657,N_6709);
xor U6894 (N_6894,N_6659,N_6723);
or U6895 (N_6895,N_6632,N_6658);
and U6896 (N_6896,N_6690,N_6723);
and U6897 (N_6897,N_6654,N_6741);
xor U6898 (N_6898,N_6614,N_6618);
xor U6899 (N_6899,N_6709,N_6723);
nand U6900 (N_6900,N_6760,N_6784);
or U6901 (N_6901,N_6827,N_6837);
nor U6902 (N_6902,N_6890,N_6835);
xnor U6903 (N_6903,N_6805,N_6814);
or U6904 (N_6904,N_6782,N_6775);
or U6905 (N_6905,N_6802,N_6886);
or U6906 (N_6906,N_6860,N_6830);
nand U6907 (N_6907,N_6893,N_6799);
or U6908 (N_6908,N_6845,N_6843);
nand U6909 (N_6909,N_6808,N_6778);
and U6910 (N_6910,N_6761,N_6881);
nor U6911 (N_6911,N_6822,N_6882);
nand U6912 (N_6912,N_6826,N_6764);
nand U6913 (N_6913,N_6896,N_6884);
or U6914 (N_6914,N_6820,N_6792);
nor U6915 (N_6915,N_6870,N_6769);
nand U6916 (N_6916,N_6880,N_6758);
xor U6917 (N_6917,N_6829,N_6768);
xor U6918 (N_6918,N_6865,N_6848);
and U6919 (N_6919,N_6877,N_6800);
or U6920 (N_6920,N_6867,N_6872);
or U6921 (N_6921,N_6895,N_6810);
nor U6922 (N_6922,N_6840,N_6853);
and U6923 (N_6923,N_6846,N_6888);
xnor U6924 (N_6924,N_6780,N_6815);
nor U6925 (N_6925,N_6875,N_6757);
or U6926 (N_6926,N_6817,N_6879);
xnor U6927 (N_6927,N_6813,N_6816);
xor U6928 (N_6928,N_6833,N_6771);
xnor U6929 (N_6929,N_6798,N_6862);
nand U6930 (N_6930,N_6839,N_6750);
xor U6931 (N_6931,N_6852,N_6844);
xnor U6932 (N_6932,N_6795,N_6801);
or U6933 (N_6933,N_6765,N_6766);
nand U6934 (N_6934,N_6783,N_6767);
nor U6935 (N_6935,N_6831,N_6756);
or U6936 (N_6936,N_6791,N_6803);
and U6937 (N_6937,N_6894,N_6762);
and U6938 (N_6938,N_6823,N_6832);
and U6939 (N_6939,N_6873,N_6856);
or U6940 (N_6940,N_6824,N_6786);
and U6941 (N_6941,N_6889,N_6869);
and U6942 (N_6942,N_6776,N_6759);
nand U6943 (N_6943,N_6863,N_6770);
xor U6944 (N_6944,N_6796,N_6849);
nor U6945 (N_6945,N_6797,N_6781);
xor U6946 (N_6946,N_6804,N_6885);
xnor U6947 (N_6947,N_6772,N_6811);
or U6948 (N_6948,N_6858,N_6854);
or U6949 (N_6949,N_6898,N_6874);
xor U6950 (N_6950,N_6892,N_6807);
or U6951 (N_6951,N_6754,N_6752);
xor U6952 (N_6952,N_6779,N_6773);
nor U6953 (N_6953,N_6794,N_6883);
xor U6954 (N_6954,N_6855,N_6790);
and U6955 (N_6955,N_6812,N_6847);
nor U6956 (N_6956,N_6842,N_6763);
nor U6957 (N_6957,N_6806,N_6818);
nand U6958 (N_6958,N_6785,N_6871);
and U6959 (N_6959,N_6866,N_6777);
nand U6960 (N_6960,N_6899,N_6868);
nor U6961 (N_6961,N_6793,N_6841);
or U6962 (N_6962,N_6751,N_6850);
or U6963 (N_6963,N_6891,N_6861);
xor U6964 (N_6964,N_6864,N_6821);
xnor U6965 (N_6965,N_6878,N_6819);
nor U6966 (N_6966,N_6828,N_6857);
or U6967 (N_6967,N_6876,N_6838);
xnor U6968 (N_6968,N_6809,N_6851);
nand U6969 (N_6969,N_6887,N_6788);
xor U6970 (N_6970,N_6859,N_6834);
xor U6971 (N_6971,N_6787,N_6774);
and U6972 (N_6972,N_6755,N_6753);
nand U6973 (N_6973,N_6825,N_6897);
xor U6974 (N_6974,N_6789,N_6836);
nor U6975 (N_6975,N_6800,N_6868);
xor U6976 (N_6976,N_6831,N_6887);
nand U6977 (N_6977,N_6761,N_6788);
nand U6978 (N_6978,N_6822,N_6791);
nand U6979 (N_6979,N_6881,N_6782);
or U6980 (N_6980,N_6816,N_6772);
xor U6981 (N_6981,N_6774,N_6823);
nand U6982 (N_6982,N_6814,N_6761);
xor U6983 (N_6983,N_6750,N_6822);
and U6984 (N_6984,N_6873,N_6849);
nand U6985 (N_6985,N_6849,N_6792);
or U6986 (N_6986,N_6824,N_6882);
xnor U6987 (N_6987,N_6788,N_6826);
xor U6988 (N_6988,N_6867,N_6760);
or U6989 (N_6989,N_6818,N_6899);
or U6990 (N_6990,N_6843,N_6897);
nand U6991 (N_6991,N_6771,N_6772);
or U6992 (N_6992,N_6821,N_6855);
or U6993 (N_6993,N_6890,N_6833);
or U6994 (N_6994,N_6875,N_6874);
nor U6995 (N_6995,N_6821,N_6840);
nand U6996 (N_6996,N_6862,N_6892);
and U6997 (N_6997,N_6772,N_6854);
nor U6998 (N_6998,N_6853,N_6823);
nor U6999 (N_6999,N_6842,N_6856);
or U7000 (N_7000,N_6793,N_6858);
nand U7001 (N_7001,N_6758,N_6792);
or U7002 (N_7002,N_6858,N_6784);
nand U7003 (N_7003,N_6792,N_6876);
xor U7004 (N_7004,N_6860,N_6871);
nor U7005 (N_7005,N_6896,N_6872);
or U7006 (N_7006,N_6767,N_6802);
and U7007 (N_7007,N_6751,N_6851);
or U7008 (N_7008,N_6785,N_6891);
nand U7009 (N_7009,N_6777,N_6874);
and U7010 (N_7010,N_6887,N_6888);
nor U7011 (N_7011,N_6837,N_6785);
xor U7012 (N_7012,N_6787,N_6845);
and U7013 (N_7013,N_6872,N_6844);
nand U7014 (N_7014,N_6860,N_6765);
nand U7015 (N_7015,N_6783,N_6848);
xnor U7016 (N_7016,N_6829,N_6826);
or U7017 (N_7017,N_6847,N_6772);
nand U7018 (N_7018,N_6782,N_6784);
nand U7019 (N_7019,N_6821,N_6843);
or U7020 (N_7020,N_6877,N_6861);
xnor U7021 (N_7021,N_6758,N_6777);
xnor U7022 (N_7022,N_6876,N_6770);
xnor U7023 (N_7023,N_6886,N_6885);
and U7024 (N_7024,N_6780,N_6783);
and U7025 (N_7025,N_6883,N_6889);
nand U7026 (N_7026,N_6851,N_6857);
and U7027 (N_7027,N_6802,N_6798);
or U7028 (N_7028,N_6780,N_6879);
nor U7029 (N_7029,N_6788,N_6806);
or U7030 (N_7030,N_6793,N_6855);
nand U7031 (N_7031,N_6775,N_6814);
and U7032 (N_7032,N_6871,N_6890);
and U7033 (N_7033,N_6886,N_6767);
xnor U7034 (N_7034,N_6862,N_6790);
nor U7035 (N_7035,N_6849,N_6835);
xor U7036 (N_7036,N_6760,N_6824);
xor U7037 (N_7037,N_6825,N_6771);
xor U7038 (N_7038,N_6873,N_6766);
nor U7039 (N_7039,N_6854,N_6830);
nor U7040 (N_7040,N_6831,N_6761);
nand U7041 (N_7041,N_6754,N_6785);
or U7042 (N_7042,N_6823,N_6811);
xnor U7043 (N_7043,N_6839,N_6760);
and U7044 (N_7044,N_6829,N_6766);
nor U7045 (N_7045,N_6843,N_6860);
or U7046 (N_7046,N_6851,N_6838);
xor U7047 (N_7047,N_6836,N_6809);
and U7048 (N_7048,N_6867,N_6853);
xnor U7049 (N_7049,N_6830,N_6783);
and U7050 (N_7050,N_6952,N_7049);
xor U7051 (N_7051,N_6925,N_7033);
nor U7052 (N_7052,N_6961,N_7001);
nor U7053 (N_7053,N_6971,N_7002);
nand U7054 (N_7054,N_7020,N_6994);
nor U7055 (N_7055,N_7010,N_6986);
nand U7056 (N_7056,N_6911,N_6956);
nor U7057 (N_7057,N_6988,N_6972);
nand U7058 (N_7058,N_6917,N_6923);
and U7059 (N_7059,N_7027,N_6977);
or U7060 (N_7060,N_6950,N_6936);
and U7061 (N_7061,N_6938,N_6939);
xnor U7062 (N_7062,N_6935,N_6963);
nand U7063 (N_7063,N_7000,N_6906);
xor U7064 (N_7064,N_6933,N_6975);
nor U7065 (N_7065,N_6990,N_6954);
nor U7066 (N_7066,N_7031,N_7038);
nand U7067 (N_7067,N_7030,N_6995);
nand U7068 (N_7068,N_6996,N_6944);
and U7069 (N_7069,N_6930,N_7046);
nor U7070 (N_7070,N_6929,N_6949);
nor U7071 (N_7071,N_6909,N_6968);
nor U7072 (N_7072,N_6965,N_6919);
and U7073 (N_7073,N_6907,N_6970);
nand U7074 (N_7074,N_7014,N_6916);
nor U7075 (N_7075,N_6985,N_6918);
nor U7076 (N_7076,N_7012,N_6964);
nand U7077 (N_7077,N_6959,N_6951);
or U7078 (N_7078,N_6905,N_6931);
xor U7079 (N_7079,N_7044,N_6903);
or U7080 (N_7080,N_6958,N_6943);
nor U7081 (N_7081,N_6924,N_6922);
nand U7082 (N_7082,N_6978,N_6908);
nand U7083 (N_7083,N_6976,N_6955);
xnor U7084 (N_7084,N_6904,N_7021);
or U7085 (N_7085,N_6913,N_7018);
nor U7086 (N_7086,N_6902,N_7042);
nand U7087 (N_7087,N_7013,N_7032);
nand U7088 (N_7088,N_6983,N_6914);
and U7089 (N_7089,N_6934,N_6942);
xnor U7090 (N_7090,N_6960,N_6987);
nor U7091 (N_7091,N_6973,N_6998);
nand U7092 (N_7092,N_7026,N_7011);
nor U7093 (N_7093,N_6948,N_7037);
nor U7094 (N_7094,N_6940,N_7035);
nor U7095 (N_7095,N_6997,N_7025);
nand U7096 (N_7096,N_7039,N_6927);
or U7097 (N_7097,N_7043,N_7036);
xor U7098 (N_7098,N_6969,N_7003);
or U7099 (N_7099,N_6966,N_6992);
nand U7100 (N_7100,N_7006,N_7034);
xor U7101 (N_7101,N_7017,N_6947);
or U7102 (N_7102,N_7007,N_7009);
nor U7103 (N_7103,N_6981,N_7023);
and U7104 (N_7104,N_6915,N_6957);
and U7105 (N_7105,N_6928,N_7040);
or U7106 (N_7106,N_7047,N_6920);
xor U7107 (N_7107,N_6912,N_6999);
or U7108 (N_7108,N_6941,N_6980);
xnor U7109 (N_7109,N_6937,N_6989);
or U7110 (N_7110,N_7015,N_6926);
nor U7111 (N_7111,N_6932,N_6921);
nor U7112 (N_7112,N_7022,N_6900);
xnor U7113 (N_7113,N_7005,N_6910);
nor U7114 (N_7114,N_7041,N_7029);
xnor U7115 (N_7115,N_6962,N_6979);
xor U7116 (N_7116,N_6953,N_6982);
xor U7117 (N_7117,N_6984,N_6991);
or U7118 (N_7118,N_7016,N_7045);
or U7119 (N_7119,N_6945,N_6974);
or U7120 (N_7120,N_7024,N_7048);
or U7121 (N_7121,N_6993,N_6967);
and U7122 (N_7122,N_7004,N_6946);
or U7123 (N_7123,N_7019,N_7028);
and U7124 (N_7124,N_7008,N_6901);
or U7125 (N_7125,N_6945,N_6995);
or U7126 (N_7126,N_6969,N_6968);
xor U7127 (N_7127,N_7026,N_6992);
or U7128 (N_7128,N_6932,N_7021);
nand U7129 (N_7129,N_7044,N_6979);
and U7130 (N_7130,N_6976,N_6945);
nor U7131 (N_7131,N_7019,N_7038);
and U7132 (N_7132,N_6947,N_6988);
xor U7133 (N_7133,N_6983,N_7046);
nand U7134 (N_7134,N_6930,N_6992);
nand U7135 (N_7135,N_6981,N_7022);
and U7136 (N_7136,N_6993,N_7012);
and U7137 (N_7137,N_6992,N_6901);
nand U7138 (N_7138,N_6922,N_7022);
and U7139 (N_7139,N_6982,N_7031);
nand U7140 (N_7140,N_7010,N_6980);
xor U7141 (N_7141,N_7030,N_7014);
or U7142 (N_7142,N_6996,N_6925);
xor U7143 (N_7143,N_7048,N_6972);
or U7144 (N_7144,N_6975,N_6947);
or U7145 (N_7145,N_6933,N_6949);
xnor U7146 (N_7146,N_7018,N_6946);
xor U7147 (N_7147,N_6981,N_6979);
or U7148 (N_7148,N_6999,N_6934);
xnor U7149 (N_7149,N_6975,N_6969);
or U7150 (N_7150,N_6959,N_6953);
nor U7151 (N_7151,N_6944,N_6982);
nor U7152 (N_7152,N_7038,N_6974);
or U7153 (N_7153,N_7041,N_6900);
nor U7154 (N_7154,N_6933,N_6989);
xor U7155 (N_7155,N_7025,N_7048);
or U7156 (N_7156,N_6901,N_6945);
nor U7157 (N_7157,N_7028,N_7000);
nand U7158 (N_7158,N_6982,N_6904);
and U7159 (N_7159,N_6924,N_6987);
xnor U7160 (N_7160,N_6911,N_6947);
and U7161 (N_7161,N_7006,N_7015);
or U7162 (N_7162,N_6974,N_7037);
nor U7163 (N_7163,N_6982,N_6960);
xnor U7164 (N_7164,N_6960,N_7004);
or U7165 (N_7165,N_6968,N_6913);
xor U7166 (N_7166,N_6995,N_7024);
nor U7167 (N_7167,N_6999,N_7038);
nand U7168 (N_7168,N_6925,N_6914);
nand U7169 (N_7169,N_6940,N_6989);
nand U7170 (N_7170,N_7045,N_7046);
xnor U7171 (N_7171,N_7035,N_6978);
and U7172 (N_7172,N_7049,N_6995);
nand U7173 (N_7173,N_6948,N_7029);
nand U7174 (N_7174,N_7029,N_7026);
xnor U7175 (N_7175,N_6976,N_7037);
or U7176 (N_7176,N_6917,N_7018);
xor U7177 (N_7177,N_6948,N_6914);
nor U7178 (N_7178,N_7040,N_6945);
nor U7179 (N_7179,N_6999,N_7039);
xnor U7180 (N_7180,N_6910,N_6986);
or U7181 (N_7181,N_7038,N_6919);
or U7182 (N_7182,N_7027,N_6970);
nor U7183 (N_7183,N_7049,N_6958);
and U7184 (N_7184,N_6950,N_6987);
or U7185 (N_7185,N_6995,N_6973);
or U7186 (N_7186,N_7010,N_6954);
or U7187 (N_7187,N_6991,N_6961);
and U7188 (N_7188,N_6913,N_6906);
or U7189 (N_7189,N_6987,N_6973);
and U7190 (N_7190,N_7007,N_7030);
nand U7191 (N_7191,N_7031,N_6971);
nand U7192 (N_7192,N_7020,N_6996);
nand U7193 (N_7193,N_6969,N_6912);
and U7194 (N_7194,N_6984,N_6928);
nor U7195 (N_7195,N_6957,N_7007);
or U7196 (N_7196,N_6944,N_6936);
nor U7197 (N_7197,N_7006,N_6974);
nand U7198 (N_7198,N_7006,N_7024);
nand U7199 (N_7199,N_6978,N_7041);
nand U7200 (N_7200,N_7156,N_7142);
and U7201 (N_7201,N_7161,N_7127);
nand U7202 (N_7202,N_7162,N_7122);
xor U7203 (N_7203,N_7182,N_7132);
nor U7204 (N_7204,N_7185,N_7195);
and U7205 (N_7205,N_7148,N_7149);
or U7206 (N_7206,N_7056,N_7123);
nor U7207 (N_7207,N_7146,N_7138);
and U7208 (N_7208,N_7104,N_7091);
and U7209 (N_7209,N_7141,N_7112);
nand U7210 (N_7210,N_7083,N_7118);
nand U7211 (N_7211,N_7128,N_7092);
and U7212 (N_7212,N_7119,N_7144);
and U7213 (N_7213,N_7090,N_7114);
or U7214 (N_7214,N_7199,N_7184);
xnor U7215 (N_7215,N_7135,N_7110);
nand U7216 (N_7216,N_7067,N_7097);
xnor U7217 (N_7217,N_7160,N_7168);
xnor U7218 (N_7218,N_7106,N_7134);
nor U7219 (N_7219,N_7145,N_7166);
or U7220 (N_7220,N_7074,N_7191);
or U7221 (N_7221,N_7159,N_7050);
nor U7222 (N_7222,N_7170,N_7163);
xor U7223 (N_7223,N_7054,N_7131);
nor U7224 (N_7224,N_7124,N_7193);
nand U7225 (N_7225,N_7059,N_7070);
and U7226 (N_7226,N_7103,N_7117);
nand U7227 (N_7227,N_7126,N_7096);
xor U7228 (N_7228,N_7081,N_7073);
nor U7229 (N_7229,N_7174,N_7157);
and U7230 (N_7230,N_7194,N_7158);
nand U7231 (N_7231,N_7064,N_7115);
nand U7232 (N_7232,N_7155,N_7075);
and U7233 (N_7233,N_7066,N_7113);
or U7234 (N_7234,N_7078,N_7190);
and U7235 (N_7235,N_7069,N_7084);
nor U7236 (N_7236,N_7068,N_7062);
or U7237 (N_7237,N_7133,N_7150);
and U7238 (N_7238,N_7071,N_7139);
and U7239 (N_7239,N_7105,N_7055);
or U7240 (N_7240,N_7082,N_7178);
or U7241 (N_7241,N_7186,N_7086);
or U7242 (N_7242,N_7094,N_7058);
or U7243 (N_7243,N_7169,N_7088);
xor U7244 (N_7244,N_7188,N_7057);
nand U7245 (N_7245,N_7154,N_7052);
nand U7246 (N_7246,N_7108,N_7181);
nor U7247 (N_7247,N_7063,N_7140);
and U7248 (N_7248,N_7143,N_7171);
nor U7249 (N_7249,N_7093,N_7130);
nor U7250 (N_7250,N_7120,N_7065);
and U7251 (N_7251,N_7085,N_7060);
or U7252 (N_7252,N_7125,N_7192);
and U7253 (N_7253,N_7164,N_7102);
nor U7254 (N_7254,N_7196,N_7072);
or U7255 (N_7255,N_7121,N_7100);
xor U7256 (N_7256,N_7153,N_7099);
xnor U7257 (N_7257,N_7151,N_7079);
and U7258 (N_7258,N_7175,N_7198);
or U7259 (N_7259,N_7172,N_7147);
nand U7260 (N_7260,N_7189,N_7165);
or U7261 (N_7261,N_7076,N_7173);
nor U7262 (N_7262,N_7109,N_7152);
and U7263 (N_7263,N_7176,N_7051);
and U7264 (N_7264,N_7179,N_7080);
nor U7265 (N_7265,N_7095,N_7089);
and U7266 (N_7266,N_7187,N_7053);
and U7267 (N_7267,N_7101,N_7111);
or U7268 (N_7268,N_7137,N_7129);
nand U7269 (N_7269,N_7136,N_7077);
nor U7270 (N_7270,N_7183,N_7107);
or U7271 (N_7271,N_7197,N_7180);
xor U7272 (N_7272,N_7087,N_7167);
or U7273 (N_7273,N_7177,N_7061);
nand U7274 (N_7274,N_7098,N_7116);
nor U7275 (N_7275,N_7147,N_7101);
or U7276 (N_7276,N_7131,N_7080);
xnor U7277 (N_7277,N_7116,N_7066);
or U7278 (N_7278,N_7184,N_7096);
nor U7279 (N_7279,N_7053,N_7163);
nor U7280 (N_7280,N_7170,N_7147);
xor U7281 (N_7281,N_7181,N_7183);
nor U7282 (N_7282,N_7199,N_7125);
or U7283 (N_7283,N_7089,N_7115);
nand U7284 (N_7284,N_7112,N_7053);
nand U7285 (N_7285,N_7059,N_7085);
or U7286 (N_7286,N_7090,N_7080);
or U7287 (N_7287,N_7105,N_7119);
nand U7288 (N_7288,N_7181,N_7173);
or U7289 (N_7289,N_7163,N_7118);
xnor U7290 (N_7290,N_7147,N_7161);
xnor U7291 (N_7291,N_7068,N_7180);
and U7292 (N_7292,N_7125,N_7121);
nor U7293 (N_7293,N_7195,N_7072);
xnor U7294 (N_7294,N_7155,N_7086);
nor U7295 (N_7295,N_7193,N_7199);
or U7296 (N_7296,N_7119,N_7126);
nand U7297 (N_7297,N_7104,N_7192);
nor U7298 (N_7298,N_7146,N_7126);
xor U7299 (N_7299,N_7078,N_7146);
or U7300 (N_7300,N_7150,N_7080);
nor U7301 (N_7301,N_7143,N_7190);
nor U7302 (N_7302,N_7052,N_7198);
xor U7303 (N_7303,N_7168,N_7147);
xnor U7304 (N_7304,N_7153,N_7189);
nand U7305 (N_7305,N_7155,N_7127);
and U7306 (N_7306,N_7111,N_7098);
nor U7307 (N_7307,N_7118,N_7148);
nor U7308 (N_7308,N_7127,N_7083);
nor U7309 (N_7309,N_7074,N_7175);
nor U7310 (N_7310,N_7084,N_7136);
nand U7311 (N_7311,N_7145,N_7135);
and U7312 (N_7312,N_7115,N_7162);
nor U7313 (N_7313,N_7067,N_7162);
nand U7314 (N_7314,N_7140,N_7081);
and U7315 (N_7315,N_7185,N_7178);
nor U7316 (N_7316,N_7188,N_7078);
nand U7317 (N_7317,N_7126,N_7100);
nor U7318 (N_7318,N_7122,N_7102);
nor U7319 (N_7319,N_7125,N_7122);
nand U7320 (N_7320,N_7116,N_7126);
nor U7321 (N_7321,N_7181,N_7086);
or U7322 (N_7322,N_7103,N_7075);
and U7323 (N_7323,N_7123,N_7108);
or U7324 (N_7324,N_7185,N_7065);
nand U7325 (N_7325,N_7105,N_7068);
nand U7326 (N_7326,N_7171,N_7146);
and U7327 (N_7327,N_7103,N_7069);
or U7328 (N_7328,N_7180,N_7058);
xnor U7329 (N_7329,N_7087,N_7198);
nor U7330 (N_7330,N_7090,N_7130);
and U7331 (N_7331,N_7188,N_7094);
and U7332 (N_7332,N_7056,N_7065);
and U7333 (N_7333,N_7071,N_7070);
or U7334 (N_7334,N_7091,N_7093);
or U7335 (N_7335,N_7138,N_7078);
xnor U7336 (N_7336,N_7097,N_7197);
nand U7337 (N_7337,N_7153,N_7193);
nor U7338 (N_7338,N_7189,N_7135);
or U7339 (N_7339,N_7169,N_7194);
xnor U7340 (N_7340,N_7105,N_7092);
or U7341 (N_7341,N_7068,N_7174);
and U7342 (N_7342,N_7074,N_7167);
or U7343 (N_7343,N_7163,N_7153);
or U7344 (N_7344,N_7154,N_7199);
nand U7345 (N_7345,N_7168,N_7170);
xnor U7346 (N_7346,N_7102,N_7099);
and U7347 (N_7347,N_7140,N_7071);
nor U7348 (N_7348,N_7115,N_7057);
and U7349 (N_7349,N_7121,N_7112);
xnor U7350 (N_7350,N_7294,N_7318);
nor U7351 (N_7351,N_7257,N_7330);
xnor U7352 (N_7352,N_7266,N_7272);
or U7353 (N_7353,N_7249,N_7218);
or U7354 (N_7354,N_7329,N_7310);
nor U7355 (N_7355,N_7251,N_7215);
nand U7356 (N_7356,N_7301,N_7282);
nor U7357 (N_7357,N_7327,N_7345);
xor U7358 (N_7358,N_7237,N_7271);
and U7359 (N_7359,N_7295,N_7307);
or U7360 (N_7360,N_7267,N_7228);
xor U7361 (N_7361,N_7244,N_7250);
and U7362 (N_7362,N_7346,N_7313);
or U7363 (N_7363,N_7339,N_7326);
nor U7364 (N_7364,N_7247,N_7320);
xor U7365 (N_7365,N_7241,N_7205);
nand U7366 (N_7366,N_7223,N_7274);
nand U7367 (N_7367,N_7328,N_7283);
or U7368 (N_7368,N_7342,N_7233);
nor U7369 (N_7369,N_7308,N_7319);
nand U7370 (N_7370,N_7254,N_7240);
nor U7371 (N_7371,N_7279,N_7265);
nor U7372 (N_7372,N_7252,N_7211);
nand U7373 (N_7373,N_7332,N_7296);
nor U7374 (N_7374,N_7323,N_7298);
and U7375 (N_7375,N_7206,N_7312);
xnor U7376 (N_7376,N_7226,N_7219);
xnor U7377 (N_7377,N_7341,N_7280);
xor U7378 (N_7378,N_7288,N_7300);
xnor U7379 (N_7379,N_7297,N_7213);
nand U7380 (N_7380,N_7284,N_7204);
or U7381 (N_7381,N_7275,N_7200);
xor U7382 (N_7382,N_7304,N_7315);
and U7383 (N_7383,N_7246,N_7348);
nor U7384 (N_7384,N_7210,N_7347);
xnor U7385 (N_7385,N_7349,N_7278);
and U7386 (N_7386,N_7259,N_7209);
and U7387 (N_7387,N_7314,N_7248);
nor U7388 (N_7388,N_7268,N_7343);
xor U7389 (N_7389,N_7335,N_7291);
and U7390 (N_7390,N_7273,N_7344);
and U7391 (N_7391,N_7292,N_7225);
or U7392 (N_7392,N_7212,N_7258);
and U7393 (N_7393,N_7333,N_7286);
nand U7394 (N_7394,N_7316,N_7340);
or U7395 (N_7395,N_7281,N_7262);
nor U7396 (N_7396,N_7331,N_7317);
or U7397 (N_7397,N_7229,N_7245);
nor U7398 (N_7398,N_7227,N_7299);
or U7399 (N_7399,N_7276,N_7270);
xor U7400 (N_7400,N_7221,N_7201);
or U7401 (N_7401,N_7239,N_7285);
nand U7402 (N_7402,N_7234,N_7287);
and U7403 (N_7403,N_7216,N_7238);
or U7404 (N_7404,N_7235,N_7236);
xnor U7405 (N_7405,N_7214,N_7261);
or U7406 (N_7406,N_7302,N_7321);
or U7407 (N_7407,N_7224,N_7277);
nand U7408 (N_7408,N_7311,N_7269);
nor U7409 (N_7409,N_7325,N_7322);
or U7410 (N_7410,N_7338,N_7202);
xnor U7411 (N_7411,N_7309,N_7232);
nand U7412 (N_7412,N_7305,N_7255);
or U7413 (N_7413,N_7289,N_7222);
or U7414 (N_7414,N_7334,N_7260);
and U7415 (N_7415,N_7290,N_7242);
nand U7416 (N_7416,N_7220,N_7324);
xnor U7417 (N_7417,N_7203,N_7256);
nand U7418 (N_7418,N_7231,N_7303);
and U7419 (N_7419,N_7263,N_7293);
xnor U7420 (N_7420,N_7208,N_7253);
and U7421 (N_7421,N_7336,N_7264);
xnor U7422 (N_7422,N_7207,N_7230);
xnor U7423 (N_7423,N_7243,N_7306);
nor U7424 (N_7424,N_7337,N_7217);
nand U7425 (N_7425,N_7243,N_7234);
xnor U7426 (N_7426,N_7223,N_7201);
nand U7427 (N_7427,N_7284,N_7343);
nand U7428 (N_7428,N_7274,N_7332);
or U7429 (N_7429,N_7208,N_7218);
or U7430 (N_7430,N_7238,N_7329);
nand U7431 (N_7431,N_7265,N_7346);
nand U7432 (N_7432,N_7282,N_7298);
or U7433 (N_7433,N_7316,N_7260);
nand U7434 (N_7434,N_7225,N_7220);
xnor U7435 (N_7435,N_7262,N_7297);
nor U7436 (N_7436,N_7216,N_7305);
nor U7437 (N_7437,N_7322,N_7291);
nand U7438 (N_7438,N_7324,N_7258);
nand U7439 (N_7439,N_7298,N_7297);
or U7440 (N_7440,N_7323,N_7265);
nor U7441 (N_7441,N_7230,N_7314);
and U7442 (N_7442,N_7344,N_7309);
or U7443 (N_7443,N_7272,N_7253);
nor U7444 (N_7444,N_7285,N_7206);
nand U7445 (N_7445,N_7302,N_7323);
and U7446 (N_7446,N_7314,N_7287);
or U7447 (N_7447,N_7207,N_7327);
xnor U7448 (N_7448,N_7291,N_7278);
nor U7449 (N_7449,N_7268,N_7213);
or U7450 (N_7450,N_7274,N_7312);
and U7451 (N_7451,N_7252,N_7244);
xor U7452 (N_7452,N_7282,N_7318);
and U7453 (N_7453,N_7244,N_7308);
nor U7454 (N_7454,N_7236,N_7219);
nor U7455 (N_7455,N_7282,N_7308);
nand U7456 (N_7456,N_7305,N_7294);
and U7457 (N_7457,N_7285,N_7266);
and U7458 (N_7458,N_7256,N_7276);
and U7459 (N_7459,N_7335,N_7206);
nor U7460 (N_7460,N_7202,N_7248);
nor U7461 (N_7461,N_7201,N_7246);
and U7462 (N_7462,N_7218,N_7203);
nand U7463 (N_7463,N_7215,N_7336);
or U7464 (N_7464,N_7207,N_7219);
nor U7465 (N_7465,N_7252,N_7276);
and U7466 (N_7466,N_7343,N_7201);
or U7467 (N_7467,N_7249,N_7200);
and U7468 (N_7468,N_7339,N_7255);
nor U7469 (N_7469,N_7331,N_7242);
and U7470 (N_7470,N_7217,N_7329);
nor U7471 (N_7471,N_7238,N_7343);
and U7472 (N_7472,N_7216,N_7224);
nor U7473 (N_7473,N_7213,N_7326);
or U7474 (N_7474,N_7308,N_7299);
nand U7475 (N_7475,N_7204,N_7305);
or U7476 (N_7476,N_7341,N_7209);
xnor U7477 (N_7477,N_7337,N_7284);
xor U7478 (N_7478,N_7268,N_7347);
nor U7479 (N_7479,N_7265,N_7246);
xnor U7480 (N_7480,N_7239,N_7221);
nor U7481 (N_7481,N_7291,N_7340);
nand U7482 (N_7482,N_7348,N_7334);
or U7483 (N_7483,N_7343,N_7302);
nand U7484 (N_7484,N_7347,N_7221);
xor U7485 (N_7485,N_7245,N_7202);
nor U7486 (N_7486,N_7226,N_7283);
xnor U7487 (N_7487,N_7338,N_7292);
or U7488 (N_7488,N_7317,N_7344);
xnor U7489 (N_7489,N_7206,N_7345);
and U7490 (N_7490,N_7310,N_7211);
and U7491 (N_7491,N_7260,N_7349);
and U7492 (N_7492,N_7339,N_7327);
nor U7493 (N_7493,N_7340,N_7234);
nor U7494 (N_7494,N_7251,N_7219);
nor U7495 (N_7495,N_7250,N_7344);
nand U7496 (N_7496,N_7240,N_7332);
or U7497 (N_7497,N_7311,N_7226);
nor U7498 (N_7498,N_7337,N_7231);
or U7499 (N_7499,N_7276,N_7301);
and U7500 (N_7500,N_7462,N_7478);
or U7501 (N_7501,N_7488,N_7415);
and U7502 (N_7502,N_7464,N_7422);
nand U7503 (N_7503,N_7376,N_7426);
nor U7504 (N_7504,N_7489,N_7452);
nand U7505 (N_7505,N_7466,N_7449);
nor U7506 (N_7506,N_7368,N_7497);
nor U7507 (N_7507,N_7362,N_7438);
nor U7508 (N_7508,N_7386,N_7402);
or U7509 (N_7509,N_7470,N_7428);
nand U7510 (N_7510,N_7433,N_7467);
nor U7511 (N_7511,N_7377,N_7465);
or U7512 (N_7512,N_7354,N_7492);
nor U7513 (N_7513,N_7460,N_7390);
nor U7514 (N_7514,N_7490,N_7397);
or U7515 (N_7515,N_7364,N_7420);
and U7516 (N_7516,N_7425,N_7417);
or U7517 (N_7517,N_7430,N_7398);
xnor U7518 (N_7518,N_7394,N_7392);
nand U7519 (N_7519,N_7382,N_7375);
xnor U7520 (N_7520,N_7483,N_7499);
nor U7521 (N_7521,N_7419,N_7409);
and U7522 (N_7522,N_7444,N_7410);
xor U7523 (N_7523,N_7448,N_7423);
nand U7524 (N_7524,N_7401,N_7472);
nor U7525 (N_7525,N_7477,N_7369);
xor U7526 (N_7526,N_7479,N_7481);
nor U7527 (N_7527,N_7381,N_7475);
and U7528 (N_7528,N_7455,N_7427);
and U7529 (N_7529,N_7447,N_7495);
and U7530 (N_7530,N_7442,N_7491);
or U7531 (N_7531,N_7357,N_7383);
or U7532 (N_7532,N_7469,N_7451);
nor U7533 (N_7533,N_7461,N_7360);
or U7534 (N_7534,N_7391,N_7434);
nand U7535 (N_7535,N_7476,N_7367);
xor U7536 (N_7536,N_7387,N_7421);
nor U7537 (N_7537,N_7453,N_7432);
nand U7538 (N_7538,N_7403,N_7411);
nand U7539 (N_7539,N_7431,N_7471);
and U7540 (N_7540,N_7473,N_7463);
nor U7541 (N_7541,N_7408,N_7440);
nor U7542 (N_7542,N_7358,N_7365);
xor U7543 (N_7543,N_7493,N_7412);
and U7544 (N_7544,N_7446,N_7456);
or U7545 (N_7545,N_7485,N_7443);
nand U7546 (N_7546,N_7379,N_7416);
nor U7547 (N_7547,N_7496,N_7359);
and U7548 (N_7548,N_7424,N_7395);
and U7549 (N_7549,N_7413,N_7389);
or U7550 (N_7550,N_7482,N_7399);
and U7551 (N_7551,N_7457,N_7370);
nand U7552 (N_7552,N_7445,N_7361);
or U7553 (N_7553,N_7436,N_7400);
or U7554 (N_7554,N_7498,N_7484);
xnor U7555 (N_7555,N_7350,N_7486);
nor U7556 (N_7556,N_7352,N_7384);
nand U7557 (N_7557,N_7378,N_7385);
nand U7558 (N_7558,N_7393,N_7407);
xor U7559 (N_7559,N_7355,N_7435);
xor U7560 (N_7560,N_7405,N_7450);
nand U7561 (N_7561,N_7363,N_7474);
nor U7562 (N_7562,N_7351,N_7441);
xor U7563 (N_7563,N_7374,N_7414);
and U7564 (N_7564,N_7480,N_7388);
nor U7565 (N_7565,N_7487,N_7356);
nor U7566 (N_7566,N_7404,N_7458);
xnor U7567 (N_7567,N_7372,N_7437);
nor U7568 (N_7568,N_7406,N_7373);
nand U7569 (N_7569,N_7454,N_7494);
or U7570 (N_7570,N_7371,N_7396);
nor U7571 (N_7571,N_7418,N_7459);
and U7572 (N_7572,N_7429,N_7468);
xor U7573 (N_7573,N_7366,N_7353);
and U7574 (N_7574,N_7380,N_7439);
xor U7575 (N_7575,N_7485,N_7436);
and U7576 (N_7576,N_7496,N_7477);
or U7577 (N_7577,N_7373,N_7409);
nor U7578 (N_7578,N_7434,N_7483);
nand U7579 (N_7579,N_7442,N_7374);
nand U7580 (N_7580,N_7381,N_7498);
nor U7581 (N_7581,N_7482,N_7400);
nand U7582 (N_7582,N_7402,N_7428);
nand U7583 (N_7583,N_7381,N_7417);
xnor U7584 (N_7584,N_7372,N_7470);
or U7585 (N_7585,N_7368,N_7433);
or U7586 (N_7586,N_7494,N_7394);
xor U7587 (N_7587,N_7470,N_7413);
and U7588 (N_7588,N_7350,N_7430);
and U7589 (N_7589,N_7494,N_7391);
xnor U7590 (N_7590,N_7387,N_7439);
nor U7591 (N_7591,N_7412,N_7408);
or U7592 (N_7592,N_7438,N_7366);
and U7593 (N_7593,N_7452,N_7474);
nor U7594 (N_7594,N_7467,N_7453);
xor U7595 (N_7595,N_7423,N_7416);
nand U7596 (N_7596,N_7423,N_7390);
and U7597 (N_7597,N_7432,N_7472);
nor U7598 (N_7598,N_7352,N_7491);
and U7599 (N_7599,N_7401,N_7475);
nor U7600 (N_7600,N_7422,N_7434);
and U7601 (N_7601,N_7364,N_7452);
and U7602 (N_7602,N_7386,N_7422);
or U7603 (N_7603,N_7397,N_7413);
and U7604 (N_7604,N_7470,N_7473);
and U7605 (N_7605,N_7457,N_7386);
nand U7606 (N_7606,N_7381,N_7427);
or U7607 (N_7607,N_7401,N_7476);
xnor U7608 (N_7608,N_7422,N_7456);
nor U7609 (N_7609,N_7450,N_7472);
or U7610 (N_7610,N_7468,N_7401);
xnor U7611 (N_7611,N_7413,N_7465);
xor U7612 (N_7612,N_7414,N_7366);
and U7613 (N_7613,N_7473,N_7462);
nor U7614 (N_7614,N_7398,N_7350);
xnor U7615 (N_7615,N_7452,N_7459);
xor U7616 (N_7616,N_7488,N_7406);
nand U7617 (N_7617,N_7456,N_7477);
xnor U7618 (N_7618,N_7450,N_7376);
nand U7619 (N_7619,N_7439,N_7490);
nor U7620 (N_7620,N_7403,N_7380);
or U7621 (N_7621,N_7411,N_7457);
xor U7622 (N_7622,N_7439,N_7381);
nor U7623 (N_7623,N_7480,N_7460);
and U7624 (N_7624,N_7418,N_7369);
or U7625 (N_7625,N_7390,N_7414);
nand U7626 (N_7626,N_7359,N_7385);
xnor U7627 (N_7627,N_7409,N_7446);
and U7628 (N_7628,N_7446,N_7376);
or U7629 (N_7629,N_7478,N_7375);
xnor U7630 (N_7630,N_7409,N_7499);
and U7631 (N_7631,N_7474,N_7457);
nor U7632 (N_7632,N_7387,N_7492);
xnor U7633 (N_7633,N_7366,N_7470);
or U7634 (N_7634,N_7375,N_7449);
nand U7635 (N_7635,N_7484,N_7495);
nand U7636 (N_7636,N_7475,N_7405);
or U7637 (N_7637,N_7477,N_7432);
xor U7638 (N_7638,N_7456,N_7416);
or U7639 (N_7639,N_7384,N_7391);
or U7640 (N_7640,N_7405,N_7353);
or U7641 (N_7641,N_7408,N_7483);
or U7642 (N_7642,N_7408,N_7404);
and U7643 (N_7643,N_7443,N_7429);
nand U7644 (N_7644,N_7438,N_7399);
or U7645 (N_7645,N_7398,N_7483);
and U7646 (N_7646,N_7455,N_7375);
and U7647 (N_7647,N_7380,N_7480);
and U7648 (N_7648,N_7439,N_7431);
or U7649 (N_7649,N_7427,N_7354);
xor U7650 (N_7650,N_7543,N_7631);
nand U7651 (N_7651,N_7507,N_7635);
and U7652 (N_7652,N_7583,N_7634);
or U7653 (N_7653,N_7597,N_7557);
and U7654 (N_7654,N_7630,N_7622);
xor U7655 (N_7655,N_7590,N_7516);
and U7656 (N_7656,N_7616,N_7528);
or U7657 (N_7657,N_7527,N_7552);
nor U7658 (N_7658,N_7504,N_7524);
or U7659 (N_7659,N_7633,N_7586);
and U7660 (N_7660,N_7601,N_7611);
or U7661 (N_7661,N_7511,N_7648);
nor U7662 (N_7662,N_7535,N_7540);
and U7663 (N_7663,N_7539,N_7637);
nor U7664 (N_7664,N_7506,N_7588);
or U7665 (N_7665,N_7626,N_7649);
or U7666 (N_7666,N_7639,N_7549);
or U7667 (N_7667,N_7580,N_7561);
xor U7668 (N_7668,N_7545,N_7550);
and U7669 (N_7669,N_7546,N_7577);
or U7670 (N_7670,N_7615,N_7595);
nor U7671 (N_7671,N_7646,N_7569);
nand U7672 (N_7672,N_7579,N_7530);
nand U7673 (N_7673,N_7592,N_7536);
or U7674 (N_7674,N_7612,N_7613);
nor U7675 (N_7675,N_7562,N_7610);
xnor U7676 (N_7676,N_7531,N_7570);
or U7677 (N_7677,N_7560,N_7578);
or U7678 (N_7678,N_7605,N_7532);
or U7679 (N_7679,N_7573,N_7591);
xor U7680 (N_7680,N_7525,N_7603);
or U7681 (N_7681,N_7505,N_7521);
nor U7682 (N_7682,N_7641,N_7618);
and U7683 (N_7683,N_7534,N_7510);
nor U7684 (N_7684,N_7519,N_7542);
nand U7685 (N_7685,N_7628,N_7568);
or U7686 (N_7686,N_7643,N_7640);
xor U7687 (N_7687,N_7620,N_7556);
and U7688 (N_7688,N_7515,N_7607);
xnor U7689 (N_7689,N_7567,N_7596);
nand U7690 (N_7690,N_7623,N_7500);
nand U7691 (N_7691,N_7617,N_7582);
and U7692 (N_7692,N_7645,N_7501);
or U7693 (N_7693,N_7564,N_7587);
xor U7694 (N_7694,N_7608,N_7508);
and U7695 (N_7695,N_7513,N_7619);
nor U7696 (N_7696,N_7584,N_7554);
nor U7697 (N_7697,N_7502,N_7538);
or U7698 (N_7698,N_7518,N_7576);
and U7699 (N_7699,N_7537,N_7551);
xor U7700 (N_7700,N_7632,N_7565);
or U7701 (N_7701,N_7572,N_7589);
nor U7702 (N_7702,N_7559,N_7594);
xnor U7703 (N_7703,N_7606,N_7598);
nor U7704 (N_7704,N_7602,N_7614);
nor U7705 (N_7705,N_7644,N_7571);
xnor U7706 (N_7706,N_7593,N_7548);
and U7707 (N_7707,N_7509,N_7636);
nand U7708 (N_7708,N_7574,N_7585);
and U7709 (N_7709,N_7517,N_7638);
nand U7710 (N_7710,N_7522,N_7544);
or U7711 (N_7711,N_7647,N_7621);
or U7712 (N_7712,N_7558,N_7503);
nor U7713 (N_7713,N_7529,N_7599);
and U7714 (N_7714,N_7523,N_7526);
nor U7715 (N_7715,N_7520,N_7563);
nor U7716 (N_7716,N_7581,N_7555);
and U7717 (N_7717,N_7553,N_7541);
nand U7718 (N_7718,N_7514,N_7566);
and U7719 (N_7719,N_7512,N_7642);
and U7720 (N_7720,N_7627,N_7600);
nand U7721 (N_7721,N_7533,N_7604);
xor U7722 (N_7722,N_7609,N_7624);
nand U7723 (N_7723,N_7629,N_7625);
xor U7724 (N_7724,N_7547,N_7575);
xnor U7725 (N_7725,N_7529,N_7629);
or U7726 (N_7726,N_7550,N_7637);
nor U7727 (N_7727,N_7643,N_7520);
nor U7728 (N_7728,N_7649,N_7637);
nor U7729 (N_7729,N_7509,N_7573);
xor U7730 (N_7730,N_7554,N_7512);
xor U7731 (N_7731,N_7563,N_7636);
and U7732 (N_7732,N_7552,N_7627);
nor U7733 (N_7733,N_7635,N_7632);
nor U7734 (N_7734,N_7596,N_7530);
nor U7735 (N_7735,N_7542,N_7545);
xnor U7736 (N_7736,N_7607,N_7551);
and U7737 (N_7737,N_7598,N_7592);
nor U7738 (N_7738,N_7615,N_7521);
nor U7739 (N_7739,N_7519,N_7504);
xor U7740 (N_7740,N_7602,N_7526);
xnor U7741 (N_7741,N_7548,N_7500);
and U7742 (N_7742,N_7559,N_7604);
nand U7743 (N_7743,N_7500,N_7646);
nand U7744 (N_7744,N_7620,N_7630);
nor U7745 (N_7745,N_7519,N_7613);
or U7746 (N_7746,N_7611,N_7618);
and U7747 (N_7747,N_7589,N_7641);
nand U7748 (N_7748,N_7579,N_7551);
nand U7749 (N_7749,N_7589,N_7523);
nand U7750 (N_7750,N_7587,N_7634);
nor U7751 (N_7751,N_7531,N_7648);
and U7752 (N_7752,N_7559,N_7590);
xnor U7753 (N_7753,N_7569,N_7586);
and U7754 (N_7754,N_7535,N_7524);
and U7755 (N_7755,N_7511,N_7527);
xnor U7756 (N_7756,N_7643,N_7566);
xor U7757 (N_7757,N_7526,N_7583);
nand U7758 (N_7758,N_7646,N_7579);
xnor U7759 (N_7759,N_7636,N_7600);
and U7760 (N_7760,N_7587,N_7604);
or U7761 (N_7761,N_7548,N_7585);
nor U7762 (N_7762,N_7646,N_7575);
xnor U7763 (N_7763,N_7531,N_7530);
nor U7764 (N_7764,N_7595,N_7512);
xnor U7765 (N_7765,N_7599,N_7611);
nand U7766 (N_7766,N_7564,N_7601);
nand U7767 (N_7767,N_7615,N_7610);
and U7768 (N_7768,N_7634,N_7532);
and U7769 (N_7769,N_7592,N_7551);
xnor U7770 (N_7770,N_7524,N_7514);
nor U7771 (N_7771,N_7501,N_7625);
xnor U7772 (N_7772,N_7536,N_7505);
nor U7773 (N_7773,N_7583,N_7561);
nand U7774 (N_7774,N_7513,N_7501);
and U7775 (N_7775,N_7577,N_7560);
or U7776 (N_7776,N_7580,N_7512);
or U7777 (N_7777,N_7549,N_7597);
and U7778 (N_7778,N_7617,N_7634);
nor U7779 (N_7779,N_7616,N_7567);
or U7780 (N_7780,N_7525,N_7616);
and U7781 (N_7781,N_7642,N_7601);
nor U7782 (N_7782,N_7507,N_7542);
xnor U7783 (N_7783,N_7561,N_7579);
and U7784 (N_7784,N_7577,N_7598);
and U7785 (N_7785,N_7575,N_7501);
xor U7786 (N_7786,N_7625,N_7637);
or U7787 (N_7787,N_7593,N_7569);
or U7788 (N_7788,N_7522,N_7598);
nor U7789 (N_7789,N_7593,N_7540);
and U7790 (N_7790,N_7562,N_7609);
and U7791 (N_7791,N_7635,N_7518);
nor U7792 (N_7792,N_7645,N_7560);
nor U7793 (N_7793,N_7538,N_7559);
and U7794 (N_7794,N_7625,N_7623);
nor U7795 (N_7795,N_7559,N_7625);
xnor U7796 (N_7796,N_7526,N_7550);
nand U7797 (N_7797,N_7575,N_7523);
or U7798 (N_7798,N_7603,N_7533);
nor U7799 (N_7799,N_7639,N_7505);
nor U7800 (N_7800,N_7764,N_7654);
or U7801 (N_7801,N_7794,N_7787);
nor U7802 (N_7802,N_7774,N_7712);
or U7803 (N_7803,N_7781,N_7742);
nand U7804 (N_7804,N_7782,N_7759);
and U7805 (N_7805,N_7695,N_7678);
xnor U7806 (N_7806,N_7657,N_7660);
and U7807 (N_7807,N_7670,N_7739);
nand U7808 (N_7808,N_7771,N_7734);
xnor U7809 (N_7809,N_7724,N_7681);
and U7810 (N_7810,N_7761,N_7760);
xnor U7811 (N_7811,N_7668,N_7752);
xnor U7812 (N_7812,N_7777,N_7715);
nor U7813 (N_7813,N_7688,N_7758);
nand U7814 (N_7814,N_7686,N_7755);
or U7815 (N_7815,N_7746,N_7676);
nor U7816 (N_7816,N_7780,N_7701);
nor U7817 (N_7817,N_7662,N_7737);
nor U7818 (N_7818,N_7677,N_7756);
nor U7819 (N_7819,N_7692,N_7793);
and U7820 (N_7820,N_7797,N_7791);
xor U7821 (N_7821,N_7773,N_7727);
or U7822 (N_7822,N_7730,N_7738);
xor U7823 (N_7823,N_7725,N_7786);
xnor U7824 (N_7824,N_7747,N_7723);
nand U7825 (N_7825,N_7673,N_7753);
nand U7826 (N_7826,N_7702,N_7748);
nor U7827 (N_7827,N_7699,N_7736);
or U7828 (N_7828,N_7762,N_7792);
or U7829 (N_7829,N_7783,N_7785);
xor U7830 (N_7830,N_7745,N_7731);
nand U7831 (N_7831,N_7703,N_7666);
or U7832 (N_7832,N_7705,N_7659);
nor U7833 (N_7833,N_7722,N_7704);
nand U7834 (N_7834,N_7691,N_7751);
nand U7835 (N_7835,N_7663,N_7711);
nor U7836 (N_7836,N_7721,N_7683);
and U7837 (N_7837,N_7682,N_7652);
or U7838 (N_7838,N_7735,N_7798);
nand U7839 (N_7839,N_7697,N_7726);
nor U7840 (N_7840,N_7744,N_7728);
or U7841 (N_7841,N_7687,N_7720);
nand U7842 (N_7842,N_7719,N_7706);
xor U7843 (N_7843,N_7733,N_7749);
nor U7844 (N_7844,N_7698,N_7768);
and U7845 (N_7845,N_7754,N_7740);
nand U7846 (N_7846,N_7743,N_7675);
nor U7847 (N_7847,N_7779,N_7696);
nand U7848 (N_7848,N_7799,N_7651);
or U7849 (N_7849,N_7784,N_7694);
and U7850 (N_7850,N_7795,N_7655);
and U7851 (N_7851,N_7658,N_7684);
nand U7852 (N_7852,N_7708,N_7685);
or U7853 (N_7853,N_7776,N_7707);
nand U7854 (N_7854,N_7656,N_7772);
and U7855 (N_7855,N_7789,N_7674);
xnor U7856 (N_7856,N_7750,N_7757);
and U7857 (N_7857,N_7718,N_7664);
xor U7858 (N_7858,N_7693,N_7672);
or U7859 (N_7859,N_7680,N_7788);
and U7860 (N_7860,N_7717,N_7775);
and U7861 (N_7861,N_7763,N_7650);
and U7862 (N_7862,N_7766,N_7689);
or U7863 (N_7863,N_7778,N_7769);
nor U7864 (N_7864,N_7653,N_7732);
nor U7865 (N_7865,N_7671,N_7790);
nor U7866 (N_7866,N_7669,N_7713);
and U7867 (N_7867,N_7716,N_7665);
xnor U7868 (N_7868,N_7709,N_7661);
xnor U7869 (N_7869,N_7714,N_7767);
xor U7870 (N_7870,N_7729,N_7667);
or U7871 (N_7871,N_7796,N_7765);
xnor U7872 (N_7872,N_7690,N_7679);
nand U7873 (N_7873,N_7700,N_7741);
nand U7874 (N_7874,N_7710,N_7770);
xor U7875 (N_7875,N_7695,N_7680);
and U7876 (N_7876,N_7796,N_7694);
xnor U7877 (N_7877,N_7687,N_7689);
xor U7878 (N_7878,N_7795,N_7797);
and U7879 (N_7879,N_7681,N_7714);
nor U7880 (N_7880,N_7789,N_7655);
and U7881 (N_7881,N_7730,N_7710);
xnor U7882 (N_7882,N_7776,N_7652);
nor U7883 (N_7883,N_7681,N_7796);
nand U7884 (N_7884,N_7779,N_7798);
nand U7885 (N_7885,N_7760,N_7692);
or U7886 (N_7886,N_7665,N_7708);
and U7887 (N_7887,N_7657,N_7724);
nor U7888 (N_7888,N_7742,N_7787);
xor U7889 (N_7889,N_7679,N_7790);
and U7890 (N_7890,N_7728,N_7738);
or U7891 (N_7891,N_7686,N_7672);
and U7892 (N_7892,N_7699,N_7684);
nor U7893 (N_7893,N_7770,N_7761);
and U7894 (N_7894,N_7660,N_7656);
or U7895 (N_7895,N_7760,N_7763);
or U7896 (N_7896,N_7799,N_7721);
xnor U7897 (N_7897,N_7724,N_7752);
and U7898 (N_7898,N_7710,N_7686);
nor U7899 (N_7899,N_7726,N_7752);
nor U7900 (N_7900,N_7782,N_7691);
nand U7901 (N_7901,N_7779,N_7660);
nor U7902 (N_7902,N_7787,N_7781);
nand U7903 (N_7903,N_7690,N_7741);
xor U7904 (N_7904,N_7754,N_7655);
xor U7905 (N_7905,N_7750,N_7754);
or U7906 (N_7906,N_7755,N_7731);
nand U7907 (N_7907,N_7766,N_7720);
or U7908 (N_7908,N_7758,N_7769);
xor U7909 (N_7909,N_7744,N_7721);
or U7910 (N_7910,N_7774,N_7739);
nor U7911 (N_7911,N_7712,N_7727);
or U7912 (N_7912,N_7688,N_7691);
nor U7913 (N_7913,N_7748,N_7737);
or U7914 (N_7914,N_7668,N_7672);
nor U7915 (N_7915,N_7700,N_7778);
nor U7916 (N_7916,N_7723,N_7655);
nand U7917 (N_7917,N_7721,N_7782);
xor U7918 (N_7918,N_7727,N_7771);
or U7919 (N_7919,N_7659,N_7687);
xor U7920 (N_7920,N_7789,N_7753);
nor U7921 (N_7921,N_7737,N_7681);
nor U7922 (N_7922,N_7755,N_7788);
xor U7923 (N_7923,N_7659,N_7793);
nand U7924 (N_7924,N_7678,N_7709);
and U7925 (N_7925,N_7667,N_7708);
nor U7926 (N_7926,N_7796,N_7672);
or U7927 (N_7927,N_7677,N_7700);
nand U7928 (N_7928,N_7797,N_7662);
nor U7929 (N_7929,N_7656,N_7729);
xor U7930 (N_7930,N_7784,N_7752);
and U7931 (N_7931,N_7798,N_7799);
nand U7932 (N_7932,N_7722,N_7711);
nand U7933 (N_7933,N_7729,N_7699);
nand U7934 (N_7934,N_7724,N_7668);
xnor U7935 (N_7935,N_7781,N_7706);
nand U7936 (N_7936,N_7715,N_7736);
and U7937 (N_7937,N_7707,N_7766);
xor U7938 (N_7938,N_7684,N_7677);
or U7939 (N_7939,N_7798,N_7706);
and U7940 (N_7940,N_7745,N_7736);
xor U7941 (N_7941,N_7687,N_7737);
nand U7942 (N_7942,N_7748,N_7691);
xor U7943 (N_7943,N_7676,N_7661);
or U7944 (N_7944,N_7688,N_7732);
and U7945 (N_7945,N_7734,N_7744);
nor U7946 (N_7946,N_7738,N_7746);
or U7947 (N_7947,N_7662,N_7793);
xor U7948 (N_7948,N_7764,N_7736);
xor U7949 (N_7949,N_7700,N_7699);
xnor U7950 (N_7950,N_7896,N_7815);
or U7951 (N_7951,N_7855,N_7801);
nor U7952 (N_7952,N_7837,N_7907);
nor U7953 (N_7953,N_7880,N_7808);
xnor U7954 (N_7954,N_7913,N_7942);
xnor U7955 (N_7955,N_7824,N_7811);
nor U7956 (N_7956,N_7848,N_7851);
or U7957 (N_7957,N_7829,N_7823);
or U7958 (N_7958,N_7885,N_7862);
xnor U7959 (N_7959,N_7891,N_7927);
nor U7960 (N_7960,N_7912,N_7935);
nor U7961 (N_7961,N_7939,N_7832);
nor U7962 (N_7962,N_7931,N_7943);
or U7963 (N_7963,N_7817,N_7821);
and U7964 (N_7964,N_7904,N_7853);
nand U7965 (N_7965,N_7842,N_7870);
or U7966 (N_7966,N_7889,N_7921);
xor U7967 (N_7967,N_7864,N_7923);
and U7968 (N_7968,N_7892,N_7879);
nor U7969 (N_7969,N_7914,N_7813);
or U7970 (N_7970,N_7905,N_7833);
nand U7971 (N_7971,N_7881,N_7814);
xor U7972 (N_7972,N_7859,N_7852);
nand U7973 (N_7973,N_7838,N_7888);
and U7974 (N_7974,N_7899,N_7920);
xor U7975 (N_7975,N_7841,N_7947);
and U7976 (N_7976,N_7856,N_7906);
nand U7977 (N_7977,N_7877,N_7940);
and U7978 (N_7978,N_7810,N_7925);
and U7979 (N_7979,N_7893,N_7916);
xor U7980 (N_7980,N_7876,N_7825);
and U7981 (N_7981,N_7860,N_7936);
nand U7982 (N_7982,N_7918,N_7886);
xor U7983 (N_7983,N_7865,N_7805);
and U7984 (N_7984,N_7804,N_7868);
and U7985 (N_7985,N_7948,N_7839);
and U7986 (N_7986,N_7874,N_7944);
nand U7987 (N_7987,N_7894,N_7901);
nand U7988 (N_7988,N_7900,N_7867);
and U7989 (N_7989,N_7895,N_7945);
xnor U7990 (N_7990,N_7937,N_7828);
nand U7991 (N_7991,N_7875,N_7926);
nand U7992 (N_7992,N_7869,N_7934);
nand U7993 (N_7993,N_7812,N_7816);
xor U7994 (N_7994,N_7844,N_7917);
and U7995 (N_7995,N_7857,N_7932);
xnor U7996 (N_7996,N_7807,N_7903);
nand U7997 (N_7997,N_7858,N_7846);
nand U7998 (N_7998,N_7882,N_7831);
xor U7999 (N_7999,N_7949,N_7866);
or U8000 (N_8000,N_7806,N_7930);
xor U8001 (N_8001,N_7941,N_7800);
and U8002 (N_8002,N_7861,N_7909);
nor U8003 (N_8003,N_7884,N_7822);
xor U8004 (N_8004,N_7890,N_7834);
and U8005 (N_8005,N_7840,N_7938);
xnor U8006 (N_8006,N_7922,N_7845);
and U8007 (N_8007,N_7902,N_7827);
xor U8008 (N_8008,N_7871,N_7849);
or U8009 (N_8009,N_7802,N_7933);
and U8010 (N_8010,N_7836,N_7820);
and U8011 (N_8011,N_7887,N_7830);
or U8012 (N_8012,N_7898,N_7878);
nor U8013 (N_8013,N_7929,N_7854);
nor U8014 (N_8014,N_7835,N_7826);
nand U8015 (N_8015,N_7850,N_7872);
or U8016 (N_8016,N_7863,N_7915);
nor U8017 (N_8017,N_7928,N_7910);
and U8018 (N_8018,N_7883,N_7911);
or U8019 (N_8019,N_7803,N_7908);
xnor U8020 (N_8020,N_7809,N_7924);
nor U8021 (N_8021,N_7843,N_7818);
or U8022 (N_8022,N_7819,N_7873);
xor U8023 (N_8023,N_7919,N_7847);
nand U8024 (N_8024,N_7897,N_7946);
and U8025 (N_8025,N_7939,N_7821);
xnor U8026 (N_8026,N_7862,N_7802);
and U8027 (N_8027,N_7813,N_7821);
nand U8028 (N_8028,N_7850,N_7828);
xor U8029 (N_8029,N_7928,N_7805);
and U8030 (N_8030,N_7818,N_7891);
and U8031 (N_8031,N_7927,N_7821);
nor U8032 (N_8032,N_7947,N_7913);
or U8033 (N_8033,N_7849,N_7922);
xor U8034 (N_8034,N_7823,N_7857);
nand U8035 (N_8035,N_7913,N_7800);
and U8036 (N_8036,N_7844,N_7837);
and U8037 (N_8037,N_7833,N_7829);
nand U8038 (N_8038,N_7817,N_7849);
nor U8039 (N_8039,N_7868,N_7896);
xnor U8040 (N_8040,N_7947,N_7809);
xnor U8041 (N_8041,N_7887,N_7869);
nor U8042 (N_8042,N_7863,N_7885);
or U8043 (N_8043,N_7933,N_7888);
nor U8044 (N_8044,N_7821,N_7804);
or U8045 (N_8045,N_7812,N_7906);
nor U8046 (N_8046,N_7910,N_7860);
xor U8047 (N_8047,N_7804,N_7934);
nor U8048 (N_8048,N_7840,N_7876);
and U8049 (N_8049,N_7921,N_7867);
or U8050 (N_8050,N_7858,N_7866);
xnor U8051 (N_8051,N_7917,N_7931);
xnor U8052 (N_8052,N_7887,N_7811);
xnor U8053 (N_8053,N_7907,N_7825);
nand U8054 (N_8054,N_7866,N_7819);
nand U8055 (N_8055,N_7924,N_7805);
xor U8056 (N_8056,N_7835,N_7942);
and U8057 (N_8057,N_7854,N_7915);
and U8058 (N_8058,N_7926,N_7932);
or U8059 (N_8059,N_7830,N_7820);
xor U8060 (N_8060,N_7867,N_7807);
nand U8061 (N_8061,N_7804,N_7829);
xnor U8062 (N_8062,N_7900,N_7837);
and U8063 (N_8063,N_7851,N_7844);
xor U8064 (N_8064,N_7823,N_7840);
nor U8065 (N_8065,N_7914,N_7858);
nand U8066 (N_8066,N_7931,N_7838);
xnor U8067 (N_8067,N_7841,N_7938);
nor U8068 (N_8068,N_7850,N_7874);
or U8069 (N_8069,N_7866,N_7803);
nand U8070 (N_8070,N_7878,N_7909);
nor U8071 (N_8071,N_7842,N_7866);
nor U8072 (N_8072,N_7912,N_7871);
xor U8073 (N_8073,N_7833,N_7851);
and U8074 (N_8074,N_7807,N_7846);
or U8075 (N_8075,N_7915,N_7883);
or U8076 (N_8076,N_7807,N_7919);
nand U8077 (N_8077,N_7855,N_7869);
nor U8078 (N_8078,N_7862,N_7841);
nand U8079 (N_8079,N_7852,N_7843);
and U8080 (N_8080,N_7823,N_7826);
or U8081 (N_8081,N_7895,N_7941);
xor U8082 (N_8082,N_7889,N_7899);
or U8083 (N_8083,N_7920,N_7817);
xor U8084 (N_8084,N_7820,N_7881);
xor U8085 (N_8085,N_7848,N_7944);
and U8086 (N_8086,N_7892,N_7855);
nor U8087 (N_8087,N_7831,N_7878);
and U8088 (N_8088,N_7833,N_7902);
xnor U8089 (N_8089,N_7908,N_7853);
and U8090 (N_8090,N_7936,N_7940);
and U8091 (N_8091,N_7833,N_7824);
and U8092 (N_8092,N_7829,N_7861);
nor U8093 (N_8093,N_7815,N_7811);
and U8094 (N_8094,N_7801,N_7891);
nor U8095 (N_8095,N_7900,N_7854);
xor U8096 (N_8096,N_7947,N_7892);
or U8097 (N_8097,N_7839,N_7838);
nor U8098 (N_8098,N_7841,N_7913);
xnor U8099 (N_8099,N_7813,N_7934);
and U8100 (N_8100,N_8025,N_8099);
and U8101 (N_8101,N_8069,N_8036);
nand U8102 (N_8102,N_8072,N_7972);
nand U8103 (N_8103,N_8028,N_8034);
nor U8104 (N_8104,N_8096,N_7988);
xor U8105 (N_8105,N_7969,N_8066);
nand U8106 (N_8106,N_8078,N_8063);
xor U8107 (N_8107,N_8048,N_7998);
or U8108 (N_8108,N_8016,N_7967);
nor U8109 (N_8109,N_7975,N_8038);
or U8110 (N_8110,N_8056,N_8093);
and U8111 (N_8111,N_8027,N_7957);
nand U8112 (N_8112,N_7953,N_8032);
and U8113 (N_8113,N_8089,N_8044);
and U8114 (N_8114,N_8074,N_8065);
or U8115 (N_8115,N_7983,N_8053);
nor U8116 (N_8116,N_8021,N_7996);
nor U8117 (N_8117,N_7984,N_8083);
nor U8118 (N_8118,N_8002,N_8098);
nand U8119 (N_8119,N_7987,N_8046);
and U8120 (N_8120,N_7960,N_8067);
nand U8121 (N_8121,N_7995,N_7959);
xor U8122 (N_8122,N_7961,N_8071);
xor U8123 (N_8123,N_8033,N_7958);
and U8124 (N_8124,N_8085,N_8084);
nor U8125 (N_8125,N_8051,N_8006);
or U8126 (N_8126,N_8076,N_8020);
nor U8127 (N_8127,N_7970,N_8041);
nand U8128 (N_8128,N_8011,N_8091);
nor U8129 (N_8129,N_8068,N_8008);
nand U8130 (N_8130,N_8024,N_7991);
xor U8131 (N_8131,N_7979,N_8014);
or U8132 (N_8132,N_7965,N_7989);
nand U8133 (N_8133,N_8088,N_8019);
nand U8134 (N_8134,N_8055,N_7976);
nor U8135 (N_8135,N_8062,N_8054);
xor U8136 (N_8136,N_7986,N_8061);
and U8137 (N_8137,N_7980,N_7994);
and U8138 (N_8138,N_8050,N_8081);
nand U8139 (N_8139,N_7964,N_7974);
and U8140 (N_8140,N_8092,N_8090);
or U8141 (N_8141,N_8080,N_8023);
and U8142 (N_8142,N_8029,N_8035);
nand U8143 (N_8143,N_8086,N_8043);
xnor U8144 (N_8144,N_8079,N_8039);
nand U8145 (N_8145,N_7951,N_8000);
nand U8146 (N_8146,N_7963,N_7997);
xnor U8147 (N_8147,N_8075,N_7973);
nor U8148 (N_8148,N_8004,N_8070);
nand U8149 (N_8149,N_7954,N_8094);
nand U8150 (N_8150,N_7985,N_8007);
or U8151 (N_8151,N_8087,N_8064);
nor U8152 (N_8152,N_7978,N_8052);
nor U8153 (N_8153,N_7955,N_7968);
nand U8154 (N_8154,N_8042,N_8095);
nor U8155 (N_8155,N_7981,N_8058);
or U8156 (N_8156,N_8057,N_8022);
and U8157 (N_8157,N_8030,N_7990);
or U8158 (N_8158,N_8082,N_8073);
or U8159 (N_8159,N_8017,N_7999);
or U8160 (N_8160,N_7982,N_8037);
xor U8161 (N_8161,N_8005,N_7971);
xnor U8162 (N_8162,N_7977,N_8097);
or U8163 (N_8163,N_8047,N_8026);
xor U8164 (N_8164,N_8060,N_7962);
xnor U8165 (N_8165,N_8013,N_8040);
nand U8166 (N_8166,N_7966,N_8018);
and U8167 (N_8167,N_8031,N_8012);
nand U8168 (N_8168,N_8077,N_7993);
nand U8169 (N_8169,N_7950,N_8059);
nor U8170 (N_8170,N_7956,N_8009);
or U8171 (N_8171,N_8003,N_7952);
or U8172 (N_8172,N_8001,N_8015);
or U8173 (N_8173,N_8049,N_8045);
nor U8174 (N_8174,N_7992,N_8010);
xor U8175 (N_8175,N_8014,N_8090);
and U8176 (N_8176,N_8080,N_7964);
nor U8177 (N_8177,N_8016,N_7974);
or U8178 (N_8178,N_8083,N_7951);
nand U8179 (N_8179,N_7985,N_8049);
or U8180 (N_8180,N_7968,N_8015);
nor U8181 (N_8181,N_8072,N_8047);
nor U8182 (N_8182,N_7978,N_8099);
or U8183 (N_8183,N_8046,N_7954);
and U8184 (N_8184,N_7967,N_8057);
nand U8185 (N_8185,N_8092,N_7975);
or U8186 (N_8186,N_7966,N_8023);
nor U8187 (N_8187,N_7958,N_8023);
or U8188 (N_8188,N_8079,N_8056);
and U8189 (N_8189,N_7967,N_8019);
nand U8190 (N_8190,N_8038,N_8092);
nor U8191 (N_8191,N_7963,N_8083);
and U8192 (N_8192,N_7973,N_8099);
nor U8193 (N_8193,N_8045,N_7976);
xor U8194 (N_8194,N_7998,N_8097);
or U8195 (N_8195,N_8012,N_8059);
nand U8196 (N_8196,N_8066,N_7950);
nor U8197 (N_8197,N_7984,N_7956);
nand U8198 (N_8198,N_8085,N_8028);
nor U8199 (N_8199,N_8049,N_8087);
and U8200 (N_8200,N_7981,N_7976);
nor U8201 (N_8201,N_8025,N_7961);
and U8202 (N_8202,N_7963,N_8061);
nor U8203 (N_8203,N_8020,N_7964);
nor U8204 (N_8204,N_8050,N_8031);
or U8205 (N_8205,N_7988,N_7992);
or U8206 (N_8206,N_7956,N_7999);
and U8207 (N_8207,N_8089,N_7993);
and U8208 (N_8208,N_7995,N_8006);
nor U8209 (N_8209,N_8017,N_7988);
nand U8210 (N_8210,N_7990,N_8013);
or U8211 (N_8211,N_7987,N_8059);
and U8212 (N_8212,N_8043,N_8033);
xnor U8213 (N_8213,N_8051,N_8026);
nand U8214 (N_8214,N_8064,N_8078);
nor U8215 (N_8215,N_8050,N_8095);
nand U8216 (N_8216,N_8059,N_8066);
nor U8217 (N_8217,N_7971,N_8045);
xnor U8218 (N_8218,N_8063,N_8064);
nor U8219 (N_8219,N_7968,N_7976);
or U8220 (N_8220,N_8035,N_7999);
or U8221 (N_8221,N_7987,N_8065);
nor U8222 (N_8222,N_8084,N_8075);
and U8223 (N_8223,N_8048,N_8075);
and U8224 (N_8224,N_7952,N_7969);
nand U8225 (N_8225,N_7968,N_8086);
and U8226 (N_8226,N_7988,N_8098);
and U8227 (N_8227,N_8003,N_8021);
or U8228 (N_8228,N_7973,N_8084);
or U8229 (N_8229,N_8037,N_8025);
nor U8230 (N_8230,N_7981,N_8011);
and U8231 (N_8231,N_7964,N_7951);
and U8232 (N_8232,N_7989,N_8049);
nand U8233 (N_8233,N_8099,N_7960);
nand U8234 (N_8234,N_8011,N_7998);
and U8235 (N_8235,N_7980,N_8067);
or U8236 (N_8236,N_7963,N_8033);
nand U8237 (N_8237,N_7971,N_7980);
xnor U8238 (N_8238,N_8023,N_8090);
xnor U8239 (N_8239,N_8050,N_8072);
or U8240 (N_8240,N_8010,N_7951);
nor U8241 (N_8241,N_8004,N_7963);
nand U8242 (N_8242,N_7953,N_8020);
nand U8243 (N_8243,N_7987,N_8096);
nor U8244 (N_8244,N_7978,N_8032);
nor U8245 (N_8245,N_7951,N_7988);
nor U8246 (N_8246,N_8049,N_7992);
and U8247 (N_8247,N_8047,N_7976);
nand U8248 (N_8248,N_8083,N_7992);
and U8249 (N_8249,N_8089,N_8023);
and U8250 (N_8250,N_8192,N_8159);
nor U8251 (N_8251,N_8249,N_8138);
and U8252 (N_8252,N_8220,N_8225);
nand U8253 (N_8253,N_8127,N_8204);
and U8254 (N_8254,N_8196,N_8155);
xnor U8255 (N_8255,N_8247,N_8200);
or U8256 (N_8256,N_8132,N_8181);
xnor U8257 (N_8257,N_8115,N_8121);
xnor U8258 (N_8258,N_8153,N_8116);
and U8259 (N_8259,N_8122,N_8112);
or U8260 (N_8260,N_8142,N_8169);
and U8261 (N_8261,N_8154,N_8179);
nor U8262 (N_8262,N_8139,N_8193);
and U8263 (N_8263,N_8214,N_8203);
or U8264 (N_8264,N_8108,N_8207);
xor U8265 (N_8265,N_8237,N_8157);
and U8266 (N_8266,N_8114,N_8136);
and U8267 (N_8267,N_8131,N_8143);
nand U8268 (N_8268,N_8189,N_8218);
xnor U8269 (N_8269,N_8182,N_8240);
nand U8270 (N_8270,N_8156,N_8152);
nor U8271 (N_8271,N_8219,N_8197);
and U8272 (N_8272,N_8160,N_8184);
nand U8273 (N_8273,N_8126,N_8227);
nand U8274 (N_8274,N_8113,N_8205);
or U8275 (N_8275,N_8177,N_8109);
nor U8276 (N_8276,N_8150,N_8148);
and U8277 (N_8277,N_8103,N_8133);
xnor U8278 (N_8278,N_8232,N_8228);
xor U8279 (N_8279,N_8168,N_8244);
nand U8280 (N_8280,N_8101,N_8238);
or U8281 (N_8281,N_8165,N_8129);
or U8282 (N_8282,N_8164,N_8167);
or U8283 (N_8283,N_8202,N_8212);
nand U8284 (N_8284,N_8120,N_8147);
and U8285 (N_8285,N_8183,N_8178);
nor U8286 (N_8286,N_8248,N_8117);
xor U8287 (N_8287,N_8124,N_8130);
or U8288 (N_8288,N_8198,N_8145);
nor U8289 (N_8289,N_8162,N_8226);
nand U8290 (N_8290,N_8146,N_8208);
nor U8291 (N_8291,N_8123,N_8188);
xnor U8292 (N_8292,N_8137,N_8102);
nand U8293 (N_8293,N_8187,N_8118);
xnor U8294 (N_8294,N_8106,N_8215);
nand U8295 (N_8295,N_8206,N_8230);
nand U8296 (N_8296,N_8144,N_8140);
nor U8297 (N_8297,N_8107,N_8185);
and U8298 (N_8298,N_8158,N_8191);
or U8299 (N_8299,N_8173,N_8229);
nand U8300 (N_8300,N_8100,N_8234);
nand U8301 (N_8301,N_8171,N_8245);
nor U8302 (N_8302,N_8176,N_8210);
nand U8303 (N_8303,N_8190,N_8175);
or U8304 (N_8304,N_8217,N_8161);
or U8305 (N_8305,N_8211,N_8236);
or U8306 (N_8306,N_8105,N_8151);
xor U8307 (N_8307,N_8104,N_8128);
or U8308 (N_8308,N_8216,N_8163);
xnor U8309 (N_8309,N_8235,N_8170);
and U8310 (N_8310,N_8195,N_8119);
nand U8311 (N_8311,N_8166,N_8111);
or U8312 (N_8312,N_8199,N_8149);
and U8313 (N_8313,N_8243,N_8201);
xor U8314 (N_8314,N_8172,N_8209);
nand U8315 (N_8315,N_8180,N_8125);
and U8316 (N_8316,N_8246,N_8186);
and U8317 (N_8317,N_8194,N_8242);
xnor U8318 (N_8318,N_8174,N_8241);
or U8319 (N_8319,N_8110,N_8224);
xnor U8320 (N_8320,N_8221,N_8223);
nor U8321 (N_8321,N_8141,N_8239);
nand U8322 (N_8322,N_8222,N_8213);
nand U8323 (N_8323,N_8134,N_8233);
or U8324 (N_8324,N_8135,N_8231);
xor U8325 (N_8325,N_8223,N_8176);
or U8326 (N_8326,N_8200,N_8160);
xor U8327 (N_8327,N_8148,N_8115);
or U8328 (N_8328,N_8112,N_8233);
nand U8329 (N_8329,N_8109,N_8205);
or U8330 (N_8330,N_8219,N_8173);
nor U8331 (N_8331,N_8141,N_8151);
nand U8332 (N_8332,N_8152,N_8176);
nand U8333 (N_8333,N_8222,N_8231);
or U8334 (N_8334,N_8138,N_8185);
nand U8335 (N_8335,N_8247,N_8123);
and U8336 (N_8336,N_8105,N_8192);
nor U8337 (N_8337,N_8180,N_8184);
and U8338 (N_8338,N_8109,N_8206);
xor U8339 (N_8339,N_8213,N_8170);
or U8340 (N_8340,N_8245,N_8116);
nand U8341 (N_8341,N_8220,N_8175);
and U8342 (N_8342,N_8178,N_8155);
xor U8343 (N_8343,N_8222,N_8200);
xor U8344 (N_8344,N_8243,N_8187);
xnor U8345 (N_8345,N_8127,N_8198);
nor U8346 (N_8346,N_8161,N_8190);
xor U8347 (N_8347,N_8129,N_8146);
or U8348 (N_8348,N_8104,N_8102);
nand U8349 (N_8349,N_8204,N_8156);
xor U8350 (N_8350,N_8233,N_8130);
nand U8351 (N_8351,N_8134,N_8176);
nand U8352 (N_8352,N_8139,N_8104);
nand U8353 (N_8353,N_8188,N_8218);
and U8354 (N_8354,N_8100,N_8131);
or U8355 (N_8355,N_8158,N_8212);
or U8356 (N_8356,N_8100,N_8246);
xor U8357 (N_8357,N_8159,N_8146);
and U8358 (N_8358,N_8181,N_8203);
nand U8359 (N_8359,N_8217,N_8166);
nor U8360 (N_8360,N_8226,N_8107);
and U8361 (N_8361,N_8136,N_8103);
and U8362 (N_8362,N_8217,N_8108);
nor U8363 (N_8363,N_8134,N_8139);
xnor U8364 (N_8364,N_8241,N_8212);
or U8365 (N_8365,N_8169,N_8126);
xnor U8366 (N_8366,N_8120,N_8216);
or U8367 (N_8367,N_8229,N_8114);
or U8368 (N_8368,N_8137,N_8247);
and U8369 (N_8369,N_8247,N_8129);
xor U8370 (N_8370,N_8104,N_8178);
and U8371 (N_8371,N_8130,N_8173);
nor U8372 (N_8372,N_8190,N_8198);
and U8373 (N_8373,N_8177,N_8139);
xor U8374 (N_8374,N_8104,N_8143);
nand U8375 (N_8375,N_8138,N_8215);
xor U8376 (N_8376,N_8150,N_8130);
and U8377 (N_8377,N_8234,N_8113);
and U8378 (N_8378,N_8171,N_8142);
and U8379 (N_8379,N_8215,N_8235);
and U8380 (N_8380,N_8128,N_8178);
or U8381 (N_8381,N_8223,N_8202);
nor U8382 (N_8382,N_8140,N_8236);
and U8383 (N_8383,N_8147,N_8184);
and U8384 (N_8384,N_8158,N_8161);
and U8385 (N_8385,N_8186,N_8132);
xnor U8386 (N_8386,N_8150,N_8192);
nor U8387 (N_8387,N_8140,N_8113);
nor U8388 (N_8388,N_8139,N_8105);
nor U8389 (N_8389,N_8178,N_8164);
or U8390 (N_8390,N_8244,N_8169);
xnor U8391 (N_8391,N_8134,N_8229);
nand U8392 (N_8392,N_8217,N_8195);
nand U8393 (N_8393,N_8116,N_8119);
xor U8394 (N_8394,N_8225,N_8171);
nor U8395 (N_8395,N_8245,N_8230);
nor U8396 (N_8396,N_8209,N_8197);
nand U8397 (N_8397,N_8237,N_8134);
nand U8398 (N_8398,N_8155,N_8150);
or U8399 (N_8399,N_8204,N_8163);
nor U8400 (N_8400,N_8388,N_8351);
or U8401 (N_8401,N_8383,N_8258);
nor U8402 (N_8402,N_8386,N_8357);
nor U8403 (N_8403,N_8370,N_8347);
or U8404 (N_8404,N_8300,N_8314);
and U8405 (N_8405,N_8255,N_8358);
nor U8406 (N_8406,N_8311,N_8272);
or U8407 (N_8407,N_8296,N_8372);
nor U8408 (N_8408,N_8338,N_8327);
xnor U8409 (N_8409,N_8260,N_8355);
nor U8410 (N_8410,N_8251,N_8374);
xor U8411 (N_8411,N_8324,N_8375);
nor U8412 (N_8412,N_8377,N_8328);
nor U8413 (N_8413,N_8385,N_8331);
nand U8414 (N_8414,N_8335,N_8390);
nand U8415 (N_8415,N_8278,N_8349);
xnor U8416 (N_8416,N_8320,N_8264);
xor U8417 (N_8417,N_8270,N_8330);
nor U8418 (N_8418,N_8392,N_8302);
nand U8419 (N_8419,N_8287,N_8282);
xnor U8420 (N_8420,N_8274,N_8306);
nor U8421 (N_8421,N_8290,N_8268);
and U8422 (N_8422,N_8384,N_8319);
nor U8423 (N_8423,N_8257,N_8360);
xor U8424 (N_8424,N_8309,N_8397);
and U8425 (N_8425,N_8298,N_8277);
nor U8426 (N_8426,N_8362,N_8299);
and U8427 (N_8427,N_8350,N_8295);
and U8428 (N_8428,N_8376,N_8323);
or U8429 (N_8429,N_8253,N_8305);
and U8430 (N_8430,N_8389,N_8281);
nor U8431 (N_8431,N_8326,N_8345);
xnor U8432 (N_8432,N_8337,N_8322);
and U8433 (N_8433,N_8252,N_8286);
nor U8434 (N_8434,N_8380,N_8361);
or U8435 (N_8435,N_8363,N_8315);
nor U8436 (N_8436,N_8303,N_8250);
nor U8437 (N_8437,N_8334,N_8381);
or U8438 (N_8438,N_8364,N_8378);
nor U8439 (N_8439,N_8279,N_8359);
and U8440 (N_8440,N_8373,N_8321);
and U8441 (N_8441,N_8395,N_8371);
nand U8442 (N_8442,N_8280,N_8365);
xnor U8443 (N_8443,N_8316,N_8329);
and U8444 (N_8444,N_8340,N_8353);
or U8445 (N_8445,N_8291,N_8292);
or U8446 (N_8446,N_8399,N_8382);
nor U8447 (N_8447,N_8307,N_8267);
nand U8448 (N_8448,N_8288,N_8368);
nand U8449 (N_8449,N_8343,N_8394);
nor U8450 (N_8450,N_8263,N_8333);
xnor U8451 (N_8451,N_8256,N_8336);
nor U8452 (N_8452,N_8393,N_8332);
and U8453 (N_8453,N_8297,N_8294);
and U8454 (N_8454,N_8275,N_8341);
nor U8455 (N_8455,N_8387,N_8293);
xnor U8456 (N_8456,N_8273,N_8339);
nor U8457 (N_8457,N_8342,N_8352);
or U8458 (N_8458,N_8391,N_8276);
and U8459 (N_8459,N_8344,N_8284);
nand U8460 (N_8460,N_8354,N_8259);
nor U8461 (N_8461,N_8318,N_8254);
nor U8462 (N_8462,N_8367,N_8366);
and U8463 (N_8463,N_8310,N_8266);
xnor U8464 (N_8464,N_8269,N_8325);
and U8465 (N_8465,N_8398,N_8312);
xnor U8466 (N_8466,N_8265,N_8379);
nor U8467 (N_8467,N_8262,N_8369);
and U8468 (N_8468,N_8283,N_8261);
nand U8469 (N_8469,N_8356,N_8313);
or U8470 (N_8470,N_8348,N_8285);
nor U8471 (N_8471,N_8304,N_8317);
and U8472 (N_8472,N_8346,N_8396);
nor U8473 (N_8473,N_8301,N_8271);
and U8474 (N_8474,N_8289,N_8308);
nand U8475 (N_8475,N_8297,N_8263);
xnor U8476 (N_8476,N_8347,N_8348);
and U8477 (N_8477,N_8287,N_8350);
xor U8478 (N_8478,N_8290,N_8326);
and U8479 (N_8479,N_8297,N_8392);
nor U8480 (N_8480,N_8288,N_8394);
nand U8481 (N_8481,N_8251,N_8298);
or U8482 (N_8482,N_8329,N_8323);
xor U8483 (N_8483,N_8255,N_8331);
nand U8484 (N_8484,N_8393,N_8373);
xor U8485 (N_8485,N_8350,N_8271);
nand U8486 (N_8486,N_8391,N_8343);
or U8487 (N_8487,N_8270,N_8298);
and U8488 (N_8488,N_8381,N_8263);
or U8489 (N_8489,N_8270,N_8278);
or U8490 (N_8490,N_8378,N_8273);
and U8491 (N_8491,N_8268,N_8302);
and U8492 (N_8492,N_8304,N_8297);
nand U8493 (N_8493,N_8268,N_8366);
and U8494 (N_8494,N_8259,N_8291);
and U8495 (N_8495,N_8287,N_8370);
and U8496 (N_8496,N_8336,N_8250);
xnor U8497 (N_8497,N_8384,N_8370);
and U8498 (N_8498,N_8339,N_8350);
nor U8499 (N_8499,N_8399,N_8342);
xor U8500 (N_8500,N_8348,N_8376);
or U8501 (N_8501,N_8393,N_8294);
or U8502 (N_8502,N_8392,N_8303);
nor U8503 (N_8503,N_8271,N_8325);
nand U8504 (N_8504,N_8319,N_8365);
nand U8505 (N_8505,N_8390,N_8281);
nand U8506 (N_8506,N_8363,N_8287);
nand U8507 (N_8507,N_8272,N_8369);
and U8508 (N_8508,N_8371,N_8336);
nor U8509 (N_8509,N_8327,N_8342);
xor U8510 (N_8510,N_8284,N_8332);
nand U8511 (N_8511,N_8288,N_8373);
and U8512 (N_8512,N_8293,N_8289);
nor U8513 (N_8513,N_8363,N_8290);
and U8514 (N_8514,N_8335,N_8269);
or U8515 (N_8515,N_8368,N_8311);
nand U8516 (N_8516,N_8388,N_8266);
nand U8517 (N_8517,N_8313,N_8309);
nor U8518 (N_8518,N_8272,N_8251);
and U8519 (N_8519,N_8307,N_8325);
and U8520 (N_8520,N_8375,N_8386);
nand U8521 (N_8521,N_8272,N_8332);
nor U8522 (N_8522,N_8279,N_8339);
and U8523 (N_8523,N_8309,N_8394);
nand U8524 (N_8524,N_8300,N_8301);
xnor U8525 (N_8525,N_8395,N_8269);
nand U8526 (N_8526,N_8369,N_8284);
and U8527 (N_8527,N_8311,N_8302);
or U8528 (N_8528,N_8389,N_8294);
and U8529 (N_8529,N_8346,N_8287);
and U8530 (N_8530,N_8338,N_8288);
nor U8531 (N_8531,N_8323,N_8384);
and U8532 (N_8532,N_8338,N_8295);
and U8533 (N_8533,N_8371,N_8324);
nor U8534 (N_8534,N_8316,N_8352);
or U8535 (N_8535,N_8260,N_8399);
and U8536 (N_8536,N_8375,N_8280);
and U8537 (N_8537,N_8308,N_8319);
and U8538 (N_8538,N_8278,N_8271);
nand U8539 (N_8539,N_8318,N_8366);
nand U8540 (N_8540,N_8255,N_8334);
xor U8541 (N_8541,N_8384,N_8353);
xnor U8542 (N_8542,N_8287,N_8296);
and U8543 (N_8543,N_8378,N_8315);
nand U8544 (N_8544,N_8296,N_8251);
or U8545 (N_8545,N_8316,N_8358);
or U8546 (N_8546,N_8381,N_8252);
nor U8547 (N_8547,N_8269,N_8338);
nor U8548 (N_8548,N_8258,N_8368);
xor U8549 (N_8549,N_8369,N_8295);
nor U8550 (N_8550,N_8479,N_8492);
or U8551 (N_8551,N_8508,N_8516);
and U8552 (N_8552,N_8418,N_8476);
nand U8553 (N_8553,N_8459,N_8420);
nand U8554 (N_8554,N_8434,N_8511);
nor U8555 (N_8555,N_8438,N_8460);
nand U8556 (N_8556,N_8456,N_8437);
xor U8557 (N_8557,N_8472,N_8452);
xnor U8558 (N_8558,N_8501,N_8401);
or U8559 (N_8559,N_8515,N_8417);
xnor U8560 (N_8560,N_8458,N_8538);
nor U8561 (N_8561,N_8523,N_8485);
xnor U8562 (N_8562,N_8474,N_8510);
nor U8563 (N_8563,N_8414,N_8500);
and U8564 (N_8564,N_8528,N_8412);
xnor U8565 (N_8565,N_8426,N_8490);
xnor U8566 (N_8566,N_8537,N_8431);
and U8567 (N_8567,N_8406,N_8536);
and U8568 (N_8568,N_8546,N_8525);
or U8569 (N_8569,N_8497,N_8453);
or U8570 (N_8570,N_8503,N_8483);
nand U8571 (N_8571,N_8475,N_8439);
and U8572 (N_8572,N_8409,N_8512);
and U8573 (N_8573,N_8522,N_8466);
nand U8574 (N_8574,N_8505,N_8498);
and U8575 (N_8575,N_8446,N_8404);
and U8576 (N_8576,N_8496,N_8405);
xor U8577 (N_8577,N_8461,N_8448);
nand U8578 (N_8578,N_8504,N_8436);
nand U8579 (N_8579,N_8402,N_8468);
nand U8580 (N_8580,N_8532,N_8462);
xor U8581 (N_8581,N_8445,N_8425);
xor U8582 (N_8582,N_8544,N_8543);
and U8583 (N_8583,N_8403,N_8545);
nand U8584 (N_8584,N_8509,N_8502);
or U8585 (N_8585,N_8530,N_8484);
and U8586 (N_8586,N_8527,N_8440);
nand U8587 (N_8587,N_8407,N_8526);
xor U8588 (N_8588,N_8514,N_8540);
xor U8589 (N_8589,N_8427,N_8535);
nor U8590 (N_8590,N_8488,N_8531);
nand U8591 (N_8591,N_8493,N_8482);
xor U8592 (N_8592,N_8430,N_8541);
or U8593 (N_8593,N_8506,N_8499);
or U8594 (N_8594,N_8471,N_8521);
nor U8595 (N_8595,N_8518,N_8421);
nand U8596 (N_8596,N_8443,N_8539);
and U8597 (N_8597,N_8428,N_8520);
xor U8598 (N_8598,N_8429,N_8548);
xnor U8599 (N_8599,N_8464,N_8534);
xnor U8600 (N_8600,N_8422,N_8533);
or U8601 (N_8601,N_8416,N_8524);
nand U8602 (N_8602,N_8519,N_8451);
and U8603 (N_8603,N_8467,N_8432);
or U8604 (N_8604,N_8457,N_8450);
nor U8605 (N_8605,N_8495,N_8549);
xnor U8606 (N_8606,N_8473,N_8477);
xor U8607 (N_8607,N_8419,N_8442);
nor U8608 (N_8608,N_8542,N_8494);
and U8609 (N_8609,N_8441,N_8481);
nor U8610 (N_8610,N_8478,N_8411);
xnor U8611 (N_8611,N_8517,N_8486);
and U8612 (N_8612,N_8423,N_8413);
and U8613 (N_8613,N_8480,N_8455);
nor U8614 (N_8614,N_8529,N_8410);
and U8615 (N_8615,N_8424,N_8415);
and U8616 (N_8616,N_8513,N_8400);
and U8617 (N_8617,N_8454,N_8447);
nand U8618 (N_8618,N_8435,N_8547);
xnor U8619 (N_8619,N_8433,N_8463);
and U8620 (N_8620,N_8507,N_8449);
xnor U8621 (N_8621,N_8408,N_8469);
nor U8622 (N_8622,N_8465,N_8489);
nand U8623 (N_8623,N_8444,N_8487);
and U8624 (N_8624,N_8491,N_8470);
and U8625 (N_8625,N_8471,N_8510);
or U8626 (N_8626,N_8420,N_8469);
xnor U8627 (N_8627,N_8430,N_8476);
or U8628 (N_8628,N_8475,N_8505);
nor U8629 (N_8629,N_8539,N_8438);
and U8630 (N_8630,N_8504,N_8495);
xnor U8631 (N_8631,N_8447,N_8518);
nand U8632 (N_8632,N_8434,N_8448);
or U8633 (N_8633,N_8529,N_8515);
and U8634 (N_8634,N_8475,N_8449);
nor U8635 (N_8635,N_8524,N_8400);
nor U8636 (N_8636,N_8437,N_8516);
nor U8637 (N_8637,N_8498,N_8430);
xor U8638 (N_8638,N_8471,N_8522);
or U8639 (N_8639,N_8424,N_8456);
nor U8640 (N_8640,N_8438,N_8455);
xnor U8641 (N_8641,N_8517,N_8519);
nor U8642 (N_8642,N_8495,N_8414);
nand U8643 (N_8643,N_8455,N_8547);
and U8644 (N_8644,N_8500,N_8451);
xor U8645 (N_8645,N_8436,N_8417);
nand U8646 (N_8646,N_8532,N_8480);
xor U8647 (N_8647,N_8480,N_8518);
xnor U8648 (N_8648,N_8510,N_8490);
and U8649 (N_8649,N_8507,N_8438);
and U8650 (N_8650,N_8539,N_8440);
nor U8651 (N_8651,N_8535,N_8490);
or U8652 (N_8652,N_8526,N_8521);
xnor U8653 (N_8653,N_8519,N_8421);
and U8654 (N_8654,N_8480,N_8493);
nor U8655 (N_8655,N_8405,N_8510);
nor U8656 (N_8656,N_8532,N_8498);
nand U8657 (N_8657,N_8511,N_8454);
and U8658 (N_8658,N_8539,N_8489);
and U8659 (N_8659,N_8452,N_8424);
or U8660 (N_8660,N_8457,N_8548);
or U8661 (N_8661,N_8459,N_8428);
and U8662 (N_8662,N_8521,N_8407);
and U8663 (N_8663,N_8518,N_8405);
nand U8664 (N_8664,N_8480,N_8536);
and U8665 (N_8665,N_8490,N_8427);
or U8666 (N_8666,N_8413,N_8405);
nor U8667 (N_8667,N_8424,N_8502);
and U8668 (N_8668,N_8532,N_8423);
nand U8669 (N_8669,N_8432,N_8537);
nor U8670 (N_8670,N_8440,N_8420);
or U8671 (N_8671,N_8543,N_8449);
nor U8672 (N_8672,N_8487,N_8514);
and U8673 (N_8673,N_8467,N_8466);
xnor U8674 (N_8674,N_8510,N_8512);
and U8675 (N_8675,N_8417,N_8530);
nor U8676 (N_8676,N_8412,N_8405);
and U8677 (N_8677,N_8408,N_8401);
or U8678 (N_8678,N_8506,N_8408);
and U8679 (N_8679,N_8533,N_8527);
xor U8680 (N_8680,N_8530,N_8424);
and U8681 (N_8681,N_8471,N_8506);
nand U8682 (N_8682,N_8432,N_8458);
and U8683 (N_8683,N_8548,N_8455);
nor U8684 (N_8684,N_8447,N_8400);
or U8685 (N_8685,N_8476,N_8514);
and U8686 (N_8686,N_8458,N_8406);
nor U8687 (N_8687,N_8525,N_8468);
nor U8688 (N_8688,N_8432,N_8444);
nand U8689 (N_8689,N_8513,N_8524);
nand U8690 (N_8690,N_8444,N_8401);
nor U8691 (N_8691,N_8496,N_8494);
xor U8692 (N_8692,N_8502,N_8479);
xnor U8693 (N_8693,N_8527,N_8506);
or U8694 (N_8694,N_8466,N_8482);
and U8695 (N_8695,N_8434,N_8415);
nor U8696 (N_8696,N_8429,N_8512);
or U8697 (N_8697,N_8433,N_8535);
nand U8698 (N_8698,N_8486,N_8456);
xnor U8699 (N_8699,N_8466,N_8458);
and U8700 (N_8700,N_8572,N_8695);
xor U8701 (N_8701,N_8553,N_8659);
and U8702 (N_8702,N_8573,N_8614);
and U8703 (N_8703,N_8627,N_8582);
xor U8704 (N_8704,N_8691,N_8611);
or U8705 (N_8705,N_8636,N_8690);
nand U8706 (N_8706,N_8588,N_8696);
nand U8707 (N_8707,N_8612,N_8625);
or U8708 (N_8708,N_8666,N_8687);
and U8709 (N_8709,N_8604,N_8568);
or U8710 (N_8710,N_8587,N_8560);
and U8711 (N_8711,N_8603,N_8571);
nand U8712 (N_8712,N_8590,N_8686);
or U8713 (N_8713,N_8610,N_8682);
nand U8714 (N_8714,N_8652,N_8673);
xor U8715 (N_8715,N_8600,N_8576);
nand U8716 (N_8716,N_8606,N_8599);
or U8717 (N_8717,N_8658,N_8685);
nand U8718 (N_8718,N_8583,N_8679);
or U8719 (N_8719,N_8593,N_8563);
nand U8720 (N_8720,N_8675,N_8684);
nor U8721 (N_8721,N_8668,N_8562);
xnor U8722 (N_8722,N_8575,N_8592);
or U8723 (N_8723,N_8649,N_8594);
or U8724 (N_8724,N_8567,N_8683);
nand U8725 (N_8725,N_8569,N_8676);
and U8726 (N_8726,N_8623,N_8608);
or U8727 (N_8727,N_8597,N_8556);
xnor U8728 (N_8728,N_8619,N_8585);
xor U8729 (N_8729,N_8660,N_8579);
nor U8730 (N_8730,N_8626,N_8662);
nand U8731 (N_8731,N_8574,N_8609);
xor U8732 (N_8732,N_8694,N_8570);
xnor U8733 (N_8733,N_8564,N_8596);
nand U8734 (N_8734,N_8656,N_8578);
nand U8735 (N_8735,N_8616,N_8663);
or U8736 (N_8736,N_8601,N_8650);
and U8737 (N_8737,N_8628,N_8622);
xor U8738 (N_8738,N_8671,N_8566);
and U8739 (N_8739,N_8565,N_8584);
or U8740 (N_8740,N_8613,N_8654);
xor U8741 (N_8741,N_8637,N_8618);
nand U8742 (N_8742,N_8629,N_8697);
nand U8743 (N_8743,N_8641,N_8591);
and U8744 (N_8744,N_8624,N_8665);
nand U8745 (N_8745,N_8643,N_8698);
nor U8746 (N_8746,N_8639,N_8620);
and U8747 (N_8747,N_8699,N_8551);
and U8748 (N_8748,N_8552,N_8670);
or U8749 (N_8749,N_8633,N_8580);
nand U8750 (N_8750,N_8648,N_8681);
nand U8751 (N_8751,N_8598,N_8647);
or U8752 (N_8752,N_8595,N_8638);
or U8753 (N_8753,N_8577,N_8631);
xnor U8754 (N_8754,N_8693,N_8634);
or U8755 (N_8755,N_8692,N_8630);
xnor U8756 (N_8756,N_8661,N_8680);
xnor U8757 (N_8757,N_8651,N_8674);
or U8758 (N_8758,N_8586,N_8605);
nand U8759 (N_8759,N_8635,N_8669);
and U8760 (N_8760,N_8664,N_8561);
and U8761 (N_8761,N_8607,N_8688);
xnor U8762 (N_8762,N_8617,N_8646);
or U8763 (N_8763,N_8555,N_8615);
and U8764 (N_8764,N_8558,N_8655);
nor U8765 (N_8765,N_8557,N_8678);
or U8766 (N_8766,N_8621,N_8642);
or U8767 (N_8767,N_8689,N_8657);
nand U8768 (N_8768,N_8589,N_8644);
or U8769 (N_8769,N_8632,N_8653);
nor U8770 (N_8770,N_8672,N_8640);
xnor U8771 (N_8771,N_8550,N_8645);
and U8772 (N_8772,N_8602,N_8559);
nor U8773 (N_8773,N_8667,N_8581);
nand U8774 (N_8774,N_8554,N_8677);
nand U8775 (N_8775,N_8594,N_8672);
nand U8776 (N_8776,N_8644,N_8561);
nand U8777 (N_8777,N_8666,N_8635);
and U8778 (N_8778,N_8597,N_8670);
and U8779 (N_8779,N_8621,N_8560);
and U8780 (N_8780,N_8598,N_8672);
xor U8781 (N_8781,N_8577,N_8596);
and U8782 (N_8782,N_8651,N_8634);
nand U8783 (N_8783,N_8576,N_8631);
nand U8784 (N_8784,N_8687,N_8558);
or U8785 (N_8785,N_8660,N_8650);
nand U8786 (N_8786,N_8698,N_8654);
nand U8787 (N_8787,N_8608,N_8672);
nor U8788 (N_8788,N_8558,N_8570);
nand U8789 (N_8789,N_8625,N_8691);
nand U8790 (N_8790,N_8688,N_8692);
nand U8791 (N_8791,N_8654,N_8683);
or U8792 (N_8792,N_8639,N_8599);
and U8793 (N_8793,N_8696,N_8553);
xor U8794 (N_8794,N_8612,N_8687);
nand U8795 (N_8795,N_8614,N_8570);
and U8796 (N_8796,N_8664,N_8575);
nor U8797 (N_8797,N_8555,N_8660);
nand U8798 (N_8798,N_8551,N_8589);
and U8799 (N_8799,N_8579,N_8689);
nor U8800 (N_8800,N_8687,N_8620);
nand U8801 (N_8801,N_8590,N_8678);
nand U8802 (N_8802,N_8610,N_8600);
nor U8803 (N_8803,N_8670,N_8628);
nand U8804 (N_8804,N_8651,N_8601);
xor U8805 (N_8805,N_8573,N_8649);
and U8806 (N_8806,N_8649,N_8583);
and U8807 (N_8807,N_8690,N_8659);
and U8808 (N_8808,N_8699,N_8659);
xor U8809 (N_8809,N_8675,N_8670);
nor U8810 (N_8810,N_8614,N_8589);
xnor U8811 (N_8811,N_8685,N_8605);
and U8812 (N_8812,N_8604,N_8559);
nor U8813 (N_8813,N_8665,N_8634);
nand U8814 (N_8814,N_8651,N_8662);
and U8815 (N_8815,N_8684,N_8694);
xor U8816 (N_8816,N_8573,N_8673);
or U8817 (N_8817,N_8635,N_8647);
xor U8818 (N_8818,N_8583,N_8603);
nor U8819 (N_8819,N_8654,N_8626);
xor U8820 (N_8820,N_8621,N_8662);
nor U8821 (N_8821,N_8690,N_8650);
nor U8822 (N_8822,N_8696,N_8590);
or U8823 (N_8823,N_8618,N_8660);
nor U8824 (N_8824,N_8581,N_8654);
xor U8825 (N_8825,N_8694,N_8569);
nand U8826 (N_8826,N_8578,N_8668);
nor U8827 (N_8827,N_8580,N_8687);
nand U8828 (N_8828,N_8567,N_8584);
and U8829 (N_8829,N_8635,N_8621);
xnor U8830 (N_8830,N_8563,N_8662);
or U8831 (N_8831,N_8584,N_8693);
or U8832 (N_8832,N_8657,N_8680);
nor U8833 (N_8833,N_8663,N_8606);
or U8834 (N_8834,N_8683,N_8642);
and U8835 (N_8835,N_8575,N_8659);
and U8836 (N_8836,N_8563,N_8608);
xor U8837 (N_8837,N_8587,N_8614);
nor U8838 (N_8838,N_8588,N_8686);
xor U8839 (N_8839,N_8597,N_8593);
and U8840 (N_8840,N_8631,N_8691);
xor U8841 (N_8841,N_8666,N_8699);
nand U8842 (N_8842,N_8673,N_8580);
or U8843 (N_8843,N_8680,N_8662);
or U8844 (N_8844,N_8576,N_8665);
or U8845 (N_8845,N_8655,N_8589);
or U8846 (N_8846,N_8562,N_8614);
nor U8847 (N_8847,N_8687,N_8642);
nand U8848 (N_8848,N_8647,N_8624);
xnor U8849 (N_8849,N_8699,N_8584);
or U8850 (N_8850,N_8798,N_8783);
or U8851 (N_8851,N_8701,N_8714);
nand U8852 (N_8852,N_8777,N_8781);
or U8853 (N_8853,N_8794,N_8722);
nor U8854 (N_8854,N_8825,N_8782);
or U8855 (N_8855,N_8743,N_8841);
nor U8856 (N_8856,N_8809,N_8827);
xnor U8857 (N_8857,N_8778,N_8761);
nor U8858 (N_8858,N_8744,N_8708);
or U8859 (N_8859,N_8765,N_8760);
and U8860 (N_8860,N_8713,N_8715);
and U8861 (N_8861,N_8788,N_8751);
nor U8862 (N_8862,N_8768,N_8797);
and U8863 (N_8863,N_8800,N_8835);
and U8864 (N_8864,N_8824,N_8753);
nand U8865 (N_8865,N_8845,N_8717);
and U8866 (N_8866,N_8740,N_8769);
and U8867 (N_8867,N_8805,N_8821);
nand U8868 (N_8868,N_8804,N_8729);
or U8869 (N_8869,N_8846,N_8774);
xor U8870 (N_8870,N_8739,N_8834);
nor U8871 (N_8871,N_8775,N_8726);
and U8872 (N_8872,N_8773,N_8801);
nor U8873 (N_8873,N_8732,N_8840);
xor U8874 (N_8874,N_8815,N_8741);
xor U8875 (N_8875,N_8810,N_8816);
or U8876 (N_8876,N_8730,N_8847);
and U8877 (N_8877,N_8747,N_8784);
or U8878 (N_8878,N_8745,N_8749);
nor U8879 (N_8879,N_8791,N_8818);
nor U8880 (N_8880,N_8826,N_8704);
and U8881 (N_8881,N_8796,N_8808);
or U8882 (N_8882,N_8787,N_8723);
and U8883 (N_8883,N_8716,N_8721);
nor U8884 (N_8884,N_8819,N_8706);
or U8885 (N_8885,N_8750,N_8737);
or U8886 (N_8886,N_8837,N_8833);
and U8887 (N_8887,N_8817,N_8718);
or U8888 (N_8888,N_8842,N_8820);
and U8889 (N_8889,N_8725,N_8823);
and U8890 (N_8890,N_8812,N_8789);
nand U8891 (N_8891,N_8811,N_8839);
nand U8892 (N_8892,N_8703,N_8830);
and U8893 (N_8893,N_8832,N_8844);
and U8894 (N_8894,N_8720,N_8710);
xor U8895 (N_8895,N_8836,N_8790);
xor U8896 (N_8896,N_8709,N_8727);
or U8897 (N_8897,N_8780,N_8776);
or U8898 (N_8898,N_8712,N_8838);
xor U8899 (N_8899,N_8779,N_8799);
or U8900 (N_8900,N_8806,N_8785);
xnor U8901 (N_8901,N_8772,N_8711);
xor U8902 (N_8902,N_8763,N_8762);
xnor U8903 (N_8903,N_8767,N_8766);
or U8904 (N_8904,N_8829,N_8802);
xnor U8905 (N_8905,N_8754,N_8759);
or U8906 (N_8906,N_8707,N_8728);
xor U8907 (N_8907,N_8724,N_8738);
or U8908 (N_8908,N_8813,N_8734);
or U8909 (N_8909,N_8700,N_8786);
and U8910 (N_8910,N_8770,N_8795);
and U8911 (N_8911,N_8702,N_8849);
nand U8912 (N_8912,N_8756,N_8719);
or U8913 (N_8913,N_8848,N_8828);
and U8914 (N_8914,N_8705,N_8807);
or U8915 (N_8915,N_8735,N_8736);
nor U8916 (N_8916,N_8814,N_8822);
nor U8917 (N_8917,N_8752,N_8748);
nand U8918 (N_8918,N_8803,N_8758);
and U8919 (N_8919,N_8733,N_8731);
and U8920 (N_8920,N_8843,N_8746);
or U8921 (N_8921,N_8755,N_8771);
nand U8922 (N_8922,N_8742,N_8764);
nand U8923 (N_8923,N_8793,N_8757);
or U8924 (N_8924,N_8792,N_8831);
or U8925 (N_8925,N_8793,N_8803);
and U8926 (N_8926,N_8757,N_8700);
and U8927 (N_8927,N_8735,N_8794);
and U8928 (N_8928,N_8764,N_8815);
nand U8929 (N_8929,N_8755,N_8732);
nand U8930 (N_8930,N_8779,N_8782);
nor U8931 (N_8931,N_8786,N_8738);
xor U8932 (N_8932,N_8727,N_8817);
xor U8933 (N_8933,N_8783,N_8738);
or U8934 (N_8934,N_8826,N_8816);
nor U8935 (N_8935,N_8726,N_8703);
nand U8936 (N_8936,N_8772,N_8790);
nand U8937 (N_8937,N_8795,N_8720);
and U8938 (N_8938,N_8715,N_8769);
and U8939 (N_8939,N_8834,N_8787);
and U8940 (N_8940,N_8777,N_8832);
nor U8941 (N_8941,N_8700,N_8717);
and U8942 (N_8942,N_8756,N_8743);
nand U8943 (N_8943,N_8807,N_8735);
xor U8944 (N_8944,N_8771,N_8708);
and U8945 (N_8945,N_8831,N_8755);
nor U8946 (N_8946,N_8797,N_8750);
and U8947 (N_8947,N_8844,N_8831);
xor U8948 (N_8948,N_8829,N_8719);
xnor U8949 (N_8949,N_8788,N_8738);
nor U8950 (N_8950,N_8707,N_8848);
xor U8951 (N_8951,N_8749,N_8816);
nand U8952 (N_8952,N_8795,N_8766);
and U8953 (N_8953,N_8847,N_8781);
nand U8954 (N_8954,N_8836,N_8777);
xor U8955 (N_8955,N_8725,N_8829);
nand U8956 (N_8956,N_8742,N_8723);
nand U8957 (N_8957,N_8746,N_8717);
and U8958 (N_8958,N_8730,N_8796);
or U8959 (N_8959,N_8848,N_8770);
and U8960 (N_8960,N_8845,N_8754);
or U8961 (N_8961,N_8835,N_8806);
or U8962 (N_8962,N_8794,N_8744);
and U8963 (N_8963,N_8752,N_8705);
nor U8964 (N_8964,N_8781,N_8798);
nand U8965 (N_8965,N_8701,N_8765);
and U8966 (N_8966,N_8729,N_8836);
nand U8967 (N_8967,N_8812,N_8781);
xor U8968 (N_8968,N_8839,N_8720);
nand U8969 (N_8969,N_8838,N_8766);
nor U8970 (N_8970,N_8839,N_8700);
xor U8971 (N_8971,N_8744,N_8742);
xnor U8972 (N_8972,N_8805,N_8734);
and U8973 (N_8973,N_8803,N_8721);
xnor U8974 (N_8974,N_8811,N_8832);
and U8975 (N_8975,N_8839,N_8739);
and U8976 (N_8976,N_8821,N_8791);
xnor U8977 (N_8977,N_8736,N_8741);
nand U8978 (N_8978,N_8813,N_8742);
xor U8979 (N_8979,N_8769,N_8818);
or U8980 (N_8980,N_8844,N_8737);
and U8981 (N_8981,N_8771,N_8739);
and U8982 (N_8982,N_8720,N_8841);
nand U8983 (N_8983,N_8717,N_8802);
or U8984 (N_8984,N_8716,N_8737);
nor U8985 (N_8985,N_8762,N_8750);
nand U8986 (N_8986,N_8712,N_8797);
or U8987 (N_8987,N_8729,N_8762);
nor U8988 (N_8988,N_8701,N_8709);
xnor U8989 (N_8989,N_8706,N_8752);
and U8990 (N_8990,N_8758,N_8784);
nand U8991 (N_8991,N_8822,N_8807);
xnor U8992 (N_8992,N_8707,N_8725);
and U8993 (N_8993,N_8746,N_8774);
and U8994 (N_8994,N_8839,N_8796);
or U8995 (N_8995,N_8723,N_8781);
xnor U8996 (N_8996,N_8721,N_8713);
or U8997 (N_8997,N_8843,N_8748);
or U8998 (N_8998,N_8813,N_8740);
xnor U8999 (N_8999,N_8745,N_8816);
nor U9000 (N_9000,N_8954,N_8987);
nor U9001 (N_9001,N_8870,N_8999);
nand U9002 (N_9002,N_8887,N_8906);
xnor U9003 (N_9003,N_8967,N_8941);
and U9004 (N_9004,N_8964,N_8945);
nor U9005 (N_9005,N_8983,N_8867);
and U9006 (N_9006,N_8921,N_8981);
and U9007 (N_9007,N_8884,N_8863);
xnor U9008 (N_9008,N_8955,N_8907);
nor U9009 (N_9009,N_8950,N_8929);
nand U9010 (N_9010,N_8868,N_8880);
nand U9011 (N_9011,N_8854,N_8899);
xor U9012 (N_9012,N_8966,N_8936);
or U9013 (N_9013,N_8869,N_8856);
nand U9014 (N_9014,N_8919,N_8877);
and U9015 (N_9015,N_8930,N_8938);
xor U9016 (N_9016,N_8914,N_8969);
and U9017 (N_9017,N_8944,N_8898);
nor U9018 (N_9018,N_8988,N_8928);
and U9019 (N_9019,N_8927,N_8939);
or U9020 (N_9020,N_8989,N_8952);
xnor U9021 (N_9021,N_8943,N_8960);
nand U9022 (N_9022,N_8962,N_8916);
nand U9023 (N_9023,N_8975,N_8861);
xnor U9024 (N_9024,N_8900,N_8893);
xor U9025 (N_9025,N_8892,N_8897);
xnor U9026 (N_9026,N_8991,N_8917);
xor U9027 (N_9027,N_8881,N_8973);
and U9028 (N_9028,N_8993,N_8926);
or U9029 (N_9029,N_8890,N_8915);
xnor U9030 (N_9030,N_8970,N_8865);
nor U9031 (N_9031,N_8978,N_8949);
and U9032 (N_9032,N_8997,N_8985);
or U9033 (N_9033,N_8982,N_8998);
or U9034 (N_9034,N_8937,N_8908);
and U9035 (N_9035,N_8913,N_8860);
nand U9036 (N_9036,N_8951,N_8851);
xnor U9037 (N_9037,N_8953,N_8855);
xnor U9038 (N_9038,N_8963,N_8891);
nor U9039 (N_9039,N_8931,N_8976);
nand U9040 (N_9040,N_8871,N_8958);
nand U9041 (N_9041,N_8894,N_8852);
and U9042 (N_9042,N_8957,N_8896);
nor U9043 (N_9043,N_8972,N_8918);
or U9044 (N_9044,N_8876,N_8864);
nand U9045 (N_9045,N_8912,N_8911);
or U9046 (N_9046,N_8909,N_8942);
nand U9047 (N_9047,N_8933,N_8886);
nor U9048 (N_9048,N_8986,N_8857);
nand U9049 (N_9049,N_8940,N_8934);
nor U9050 (N_9050,N_8922,N_8935);
nor U9051 (N_9051,N_8878,N_8895);
nor U9052 (N_9052,N_8977,N_8885);
nand U9053 (N_9053,N_8948,N_8959);
nor U9054 (N_9054,N_8853,N_8923);
nand U9055 (N_9055,N_8901,N_8902);
nand U9056 (N_9056,N_8859,N_8910);
or U9057 (N_9057,N_8992,N_8883);
xnor U9058 (N_9058,N_8996,N_8903);
xnor U9059 (N_9059,N_8920,N_8872);
or U9060 (N_9060,N_8961,N_8956);
and U9061 (N_9061,N_8904,N_8874);
and U9062 (N_9062,N_8889,N_8873);
xor U9063 (N_9063,N_8888,N_8850);
nor U9064 (N_9064,N_8971,N_8979);
nand U9065 (N_9065,N_8994,N_8984);
and U9066 (N_9066,N_8968,N_8866);
or U9067 (N_9067,N_8882,N_8905);
and U9068 (N_9068,N_8932,N_8974);
or U9069 (N_9069,N_8980,N_8858);
and U9070 (N_9070,N_8879,N_8924);
and U9071 (N_9071,N_8947,N_8875);
and U9072 (N_9072,N_8862,N_8995);
nor U9073 (N_9073,N_8990,N_8965);
and U9074 (N_9074,N_8946,N_8925);
and U9075 (N_9075,N_8906,N_8966);
or U9076 (N_9076,N_8926,N_8863);
and U9077 (N_9077,N_8938,N_8893);
nand U9078 (N_9078,N_8910,N_8911);
or U9079 (N_9079,N_8965,N_8910);
xor U9080 (N_9080,N_8897,N_8854);
xor U9081 (N_9081,N_8886,N_8924);
nor U9082 (N_9082,N_8973,N_8985);
nand U9083 (N_9083,N_8971,N_8905);
xnor U9084 (N_9084,N_8944,N_8904);
xnor U9085 (N_9085,N_8966,N_8886);
nor U9086 (N_9086,N_8900,N_8865);
nand U9087 (N_9087,N_8943,N_8980);
nand U9088 (N_9088,N_8941,N_8926);
xnor U9089 (N_9089,N_8943,N_8974);
xnor U9090 (N_9090,N_8895,N_8911);
or U9091 (N_9091,N_8875,N_8953);
xnor U9092 (N_9092,N_8990,N_8873);
and U9093 (N_9093,N_8923,N_8940);
xnor U9094 (N_9094,N_8893,N_8955);
nand U9095 (N_9095,N_8853,N_8937);
xor U9096 (N_9096,N_8850,N_8857);
nand U9097 (N_9097,N_8987,N_8903);
nand U9098 (N_9098,N_8885,N_8889);
and U9099 (N_9099,N_8977,N_8860);
xor U9100 (N_9100,N_8862,N_8989);
xor U9101 (N_9101,N_8862,N_8933);
nand U9102 (N_9102,N_8907,N_8928);
nand U9103 (N_9103,N_8990,N_8971);
nor U9104 (N_9104,N_8975,N_8867);
and U9105 (N_9105,N_8968,N_8973);
nor U9106 (N_9106,N_8919,N_8959);
and U9107 (N_9107,N_8880,N_8973);
xnor U9108 (N_9108,N_8935,N_8970);
or U9109 (N_9109,N_8921,N_8869);
nand U9110 (N_9110,N_8865,N_8880);
and U9111 (N_9111,N_8949,N_8892);
nor U9112 (N_9112,N_8864,N_8929);
or U9113 (N_9113,N_8968,N_8932);
nor U9114 (N_9114,N_8944,N_8851);
nor U9115 (N_9115,N_8958,N_8899);
nand U9116 (N_9116,N_8963,N_8941);
nor U9117 (N_9117,N_8936,N_8957);
nand U9118 (N_9118,N_8944,N_8958);
nand U9119 (N_9119,N_8893,N_8921);
or U9120 (N_9120,N_8892,N_8950);
and U9121 (N_9121,N_8871,N_8852);
nand U9122 (N_9122,N_8911,N_8971);
xnor U9123 (N_9123,N_8896,N_8950);
and U9124 (N_9124,N_8984,N_8858);
nor U9125 (N_9125,N_8929,N_8853);
nor U9126 (N_9126,N_8859,N_8960);
xor U9127 (N_9127,N_8949,N_8899);
nand U9128 (N_9128,N_8956,N_8859);
and U9129 (N_9129,N_8987,N_8971);
or U9130 (N_9130,N_8903,N_8868);
and U9131 (N_9131,N_8947,N_8883);
xnor U9132 (N_9132,N_8979,N_8986);
and U9133 (N_9133,N_8906,N_8996);
or U9134 (N_9134,N_8997,N_8929);
nand U9135 (N_9135,N_8917,N_8873);
nand U9136 (N_9136,N_8878,N_8953);
or U9137 (N_9137,N_8958,N_8922);
nand U9138 (N_9138,N_8990,N_8994);
and U9139 (N_9139,N_8951,N_8982);
or U9140 (N_9140,N_8918,N_8999);
or U9141 (N_9141,N_8984,N_8981);
xnor U9142 (N_9142,N_8955,N_8913);
nand U9143 (N_9143,N_8987,N_8917);
xor U9144 (N_9144,N_8953,N_8918);
and U9145 (N_9145,N_8995,N_8949);
xor U9146 (N_9146,N_8975,N_8957);
nor U9147 (N_9147,N_8866,N_8889);
nand U9148 (N_9148,N_8981,N_8919);
nor U9149 (N_9149,N_8960,N_8982);
nand U9150 (N_9150,N_9047,N_9082);
xnor U9151 (N_9151,N_9066,N_9124);
and U9152 (N_9152,N_9000,N_9063);
or U9153 (N_9153,N_9083,N_9113);
nand U9154 (N_9154,N_9035,N_9108);
xnor U9155 (N_9155,N_9045,N_9128);
or U9156 (N_9156,N_9146,N_9107);
nor U9157 (N_9157,N_9010,N_9139);
nand U9158 (N_9158,N_9004,N_9133);
and U9159 (N_9159,N_9149,N_9123);
and U9160 (N_9160,N_9001,N_9041);
and U9161 (N_9161,N_9080,N_9037);
and U9162 (N_9162,N_9094,N_9016);
xnor U9163 (N_9163,N_9119,N_9009);
nor U9164 (N_9164,N_9079,N_9011);
nor U9165 (N_9165,N_9012,N_9057);
and U9166 (N_9166,N_9007,N_9144);
nor U9167 (N_9167,N_9071,N_9086);
xnor U9168 (N_9168,N_9058,N_9088);
or U9169 (N_9169,N_9053,N_9143);
or U9170 (N_9170,N_9131,N_9021);
xnor U9171 (N_9171,N_9019,N_9118);
and U9172 (N_9172,N_9038,N_9085);
nand U9173 (N_9173,N_9008,N_9034);
xor U9174 (N_9174,N_9109,N_9048);
and U9175 (N_9175,N_9121,N_9039);
nor U9176 (N_9176,N_9032,N_9033);
and U9177 (N_9177,N_9100,N_9103);
xor U9178 (N_9178,N_9116,N_9060);
and U9179 (N_9179,N_9022,N_9138);
nand U9180 (N_9180,N_9068,N_9115);
and U9181 (N_9181,N_9028,N_9140);
nand U9182 (N_9182,N_9102,N_9061);
and U9183 (N_9183,N_9117,N_9042);
nor U9184 (N_9184,N_9091,N_9056);
and U9185 (N_9185,N_9130,N_9036);
nand U9186 (N_9186,N_9114,N_9067);
nand U9187 (N_9187,N_9129,N_9135);
xnor U9188 (N_9188,N_9052,N_9147);
nand U9189 (N_9189,N_9134,N_9126);
or U9190 (N_9190,N_9122,N_9142);
nand U9191 (N_9191,N_9106,N_9084);
xnor U9192 (N_9192,N_9062,N_9020);
nor U9193 (N_9193,N_9077,N_9070);
nor U9194 (N_9194,N_9029,N_9025);
xnor U9195 (N_9195,N_9145,N_9093);
xor U9196 (N_9196,N_9148,N_9096);
nand U9197 (N_9197,N_9111,N_9141);
nand U9198 (N_9198,N_9076,N_9030);
xor U9199 (N_9199,N_9026,N_9003);
nor U9200 (N_9200,N_9027,N_9072);
or U9201 (N_9201,N_9137,N_9043);
nand U9202 (N_9202,N_9074,N_9044);
nor U9203 (N_9203,N_9018,N_9006);
nor U9204 (N_9204,N_9046,N_9104);
and U9205 (N_9205,N_9099,N_9023);
nand U9206 (N_9206,N_9120,N_9081);
nor U9207 (N_9207,N_9040,N_9078);
xor U9208 (N_9208,N_9049,N_9002);
nand U9209 (N_9209,N_9073,N_9069);
and U9210 (N_9210,N_9031,N_9051);
and U9211 (N_9211,N_9014,N_9101);
xor U9212 (N_9212,N_9127,N_9054);
or U9213 (N_9213,N_9089,N_9095);
or U9214 (N_9214,N_9098,N_9059);
xor U9215 (N_9215,N_9005,N_9090);
nor U9216 (N_9216,N_9125,N_9105);
or U9217 (N_9217,N_9087,N_9075);
or U9218 (N_9218,N_9017,N_9110);
nor U9219 (N_9219,N_9015,N_9065);
nand U9220 (N_9220,N_9132,N_9050);
or U9221 (N_9221,N_9136,N_9097);
or U9222 (N_9222,N_9064,N_9013);
nand U9223 (N_9223,N_9055,N_9024);
or U9224 (N_9224,N_9112,N_9092);
and U9225 (N_9225,N_9025,N_9065);
nand U9226 (N_9226,N_9023,N_9120);
and U9227 (N_9227,N_9053,N_9079);
or U9228 (N_9228,N_9104,N_9105);
nor U9229 (N_9229,N_9015,N_9074);
or U9230 (N_9230,N_9075,N_9105);
nand U9231 (N_9231,N_9066,N_9078);
xor U9232 (N_9232,N_9059,N_9011);
nor U9233 (N_9233,N_9148,N_9116);
nor U9234 (N_9234,N_9007,N_9103);
nor U9235 (N_9235,N_9119,N_9040);
and U9236 (N_9236,N_9078,N_9124);
and U9237 (N_9237,N_9047,N_9038);
xor U9238 (N_9238,N_9027,N_9141);
nand U9239 (N_9239,N_9023,N_9090);
nand U9240 (N_9240,N_9144,N_9147);
or U9241 (N_9241,N_9109,N_9029);
nand U9242 (N_9242,N_9117,N_9074);
nand U9243 (N_9243,N_9125,N_9142);
and U9244 (N_9244,N_9045,N_9023);
and U9245 (N_9245,N_9026,N_9049);
xnor U9246 (N_9246,N_9101,N_9149);
nor U9247 (N_9247,N_9055,N_9122);
nor U9248 (N_9248,N_9141,N_9093);
or U9249 (N_9249,N_9000,N_9041);
or U9250 (N_9250,N_9096,N_9145);
xor U9251 (N_9251,N_9133,N_9114);
xnor U9252 (N_9252,N_9067,N_9121);
xnor U9253 (N_9253,N_9083,N_9149);
or U9254 (N_9254,N_9142,N_9087);
or U9255 (N_9255,N_9045,N_9098);
nor U9256 (N_9256,N_9096,N_9133);
xor U9257 (N_9257,N_9101,N_9113);
and U9258 (N_9258,N_9058,N_9047);
xor U9259 (N_9259,N_9011,N_9112);
xor U9260 (N_9260,N_9016,N_9106);
xnor U9261 (N_9261,N_9149,N_9119);
or U9262 (N_9262,N_9087,N_9132);
nor U9263 (N_9263,N_9105,N_9137);
nand U9264 (N_9264,N_9030,N_9003);
nor U9265 (N_9265,N_9060,N_9142);
nand U9266 (N_9266,N_9125,N_9048);
nand U9267 (N_9267,N_9121,N_9113);
xnor U9268 (N_9268,N_9106,N_9044);
nor U9269 (N_9269,N_9012,N_9141);
nor U9270 (N_9270,N_9036,N_9020);
nor U9271 (N_9271,N_9028,N_9035);
nand U9272 (N_9272,N_9097,N_9122);
xnor U9273 (N_9273,N_9099,N_9131);
nor U9274 (N_9274,N_9123,N_9124);
and U9275 (N_9275,N_9101,N_9032);
or U9276 (N_9276,N_9140,N_9071);
or U9277 (N_9277,N_9113,N_9074);
or U9278 (N_9278,N_9119,N_9052);
or U9279 (N_9279,N_9052,N_9006);
or U9280 (N_9280,N_9019,N_9015);
nor U9281 (N_9281,N_9082,N_9020);
nor U9282 (N_9282,N_9143,N_9111);
nor U9283 (N_9283,N_9138,N_9036);
and U9284 (N_9284,N_9018,N_9127);
or U9285 (N_9285,N_9127,N_9129);
and U9286 (N_9286,N_9080,N_9010);
nor U9287 (N_9287,N_9011,N_9105);
nor U9288 (N_9288,N_9046,N_9007);
xor U9289 (N_9289,N_9098,N_9102);
nor U9290 (N_9290,N_9054,N_9104);
or U9291 (N_9291,N_9146,N_9080);
nor U9292 (N_9292,N_9140,N_9146);
nor U9293 (N_9293,N_9110,N_9084);
nor U9294 (N_9294,N_9067,N_9143);
nor U9295 (N_9295,N_9137,N_9100);
xnor U9296 (N_9296,N_9092,N_9141);
or U9297 (N_9297,N_9080,N_9060);
nand U9298 (N_9298,N_9009,N_9029);
xnor U9299 (N_9299,N_9112,N_9104);
nand U9300 (N_9300,N_9299,N_9179);
or U9301 (N_9301,N_9254,N_9296);
or U9302 (N_9302,N_9156,N_9242);
xnor U9303 (N_9303,N_9211,N_9250);
nand U9304 (N_9304,N_9199,N_9259);
nand U9305 (N_9305,N_9153,N_9188);
xor U9306 (N_9306,N_9251,N_9298);
or U9307 (N_9307,N_9272,N_9177);
nor U9308 (N_9308,N_9200,N_9249);
nand U9309 (N_9309,N_9245,N_9152);
xnor U9310 (N_9310,N_9190,N_9252);
or U9311 (N_9311,N_9263,N_9180);
nor U9312 (N_9312,N_9162,N_9206);
nand U9313 (N_9313,N_9243,N_9231);
or U9314 (N_9314,N_9170,N_9227);
nand U9315 (N_9315,N_9165,N_9209);
and U9316 (N_9316,N_9262,N_9161);
and U9317 (N_9317,N_9192,N_9213);
and U9318 (N_9318,N_9284,N_9256);
or U9319 (N_9319,N_9225,N_9151);
or U9320 (N_9320,N_9257,N_9277);
and U9321 (N_9321,N_9198,N_9247);
nand U9322 (N_9322,N_9276,N_9289);
nor U9323 (N_9323,N_9197,N_9228);
or U9324 (N_9324,N_9260,N_9282);
and U9325 (N_9325,N_9155,N_9202);
or U9326 (N_9326,N_9232,N_9264);
nor U9327 (N_9327,N_9218,N_9150);
or U9328 (N_9328,N_9295,N_9160);
xnor U9329 (N_9329,N_9196,N_9290);
nor U9330 (N_9330,N_9286,N_9207);
and U9331 (N_9331,N_9287,N_9274);
nand U9332 (N_9332,N_9163,N_9240);
nand U9333 (N_9333,N_9269,N_9195);
or U9334 (N_9334,N_9171,N_9178);
xnor U9335 (N_9335,N_9241,N_9248);
nor U9336 (N_9336,N_9212,N_9278);
nand U9337 (N_9337,N_9221,N_9182);
nor U9338 (N_9338,N_9174,N_9288);
xnor U9339 (N_9339,N_9154,N_9293);
nor U9340 (N_9340,N_9172,N_9253);
nor U9341 (N_9341,N_9261,N_9283);
and U9342 (N_9342,N_9193,N_9235);
or U9343 (N_9343,N_9191,N_9181);
nand U9344 (N_9344,N_9270,N_9271);
or U9345 (N_9345,N_9279,N_9184);
and U9346 (N_9346,N_9268,N_9291);
nand U9347 (N_9347,N_9224,N_9236);
and U9348 (N_9348,N_9208,N_9219);
or U9349 (N_9349,N_9183,N_9275);
xor U9350 (N_9350,N_9297,N_9167);
nor U9351 (N_9351,N_9210,N_9157);
nand U9352 (N_9352,N_9280,N_9158);
or U9353 (N_9353,N_9233,N_9166);
or U9354 (N_9354,N_9168,N_9220);
nand U9355 (N_9355,N_9187,N_9173);
and U9356 (N_9356,N_9217,N_9215);
xor U9357 (N_9357,N_9203,N_9159);
xor U9358 (N_9358,N_9294,N_9204);
xnor U9359 (N_9359,N_9267,N_9273);
nor U9360 (N_9360,N_9234,N_9175);
or U9361 (N_9361,N_9169,N_9186);
nor U9362 (N_9362,N_9292,N_9265);
nand U9363 (N_9363,N_9205,N_9185);
xor U9364 (N_9364,N_9281,N_9201);
xnor U9365 (N_9365,N_9238,N_9266);
nand U9366 (N_9366,N_9229,N_9164);
nand U9367 (N_9367,N_9194,N_9230);
xor U9368 (N_9368,N_9222,N_9189);
or U9369 (N_9369,N_9226,N_9223);
and U9370 (N_9370,N_9244,N_9239);
and U9371 (N_9371,N_9258,N_9285);
nand U9372 (N_9372,N_9216,N_9176);
xor U9373 (N_9373,N_9246,N_9214);
nor U9374 (N_9374,N_9237,N_9255);
and U9375 (N_9375,N_9199,N_9291);
or U9376 (N_9376,N_9280,N_9154);
and U9377 (N_9377,N_9208,N_9252);
and U9378 (N_9378,N_9242,N_9235);
nand U9379 (N_9379,N_9226,N_9184);
nand U9380 (N_9380,N_9277,N_9299);
or U9381 (N_9381,N_9271,N_9185);
nor U9382 (N_9382,N_9239,N_9202);
or U9383 (N_9383,N_9289,N_9176);
xnor U9384 (N_9384,N_9254,N_9176);
nand U9385 (N_9385,N_9153,N_9183);
or U9386 (N_9386,N_9200,N_9267);
xor U9387 (N_9387,N_9188,N_9193);
or U9388 (N_9388,N_9269,N_9268);
nand U9389 (N_9389,N_9254,N_9268);
or U9390 (N_9390,N_9239,N_9283);
nor U9391 (N_9391,N_9241,N_9230);
and U9392 (N_9392,N_9263,N_9251);
nand U9393 (N_9393,N_9258,N_9295);
or U9394 (N_9394,N_9182,N_9201);
xnor U9395 (N_9395,N_9172,N_9247);
nand U9396 (N_9396,N_9248,N_9212);
and U9397 (N_9397,N_9194,N_9250);
or U9398 (N_9398,N_9220,N_9175);
xor U9399 (N_9399,N_9292,N_9256);
nand U9400 (N_9400,N_9229,N_9163);
and U9401 (N_9401,N_9289,N_9250);
or U9402 (N_9402,N_9290,N_9192);
xor U9403 (N_9403,N_9167,N_9161);
or U9404 (N_9404,N_9208,N_9242);
nand U9405 (N_9405,N_9187,N_9294);
or U9406 (N_9406,N_9298,N_9211);
and U9407 (N_9407,N_9226,N_9265);
or U9408 (N_9408,N_9169,N_9166);
or U9409 (N_9409,N_9151,N_9150);
xnor U9410 (N_9410,N_9261,N_9239);
nor U9411 (N_9411,N_9190,N_9171);
nor U9412 (N_9412,N_9250,N_9197);
or U9413 (N_9413,N_9176,N_9279);
nor U9414 (N_9414,N_9226,N_9250);
nand U9415 (N_9415,N_9215,N_9180);
xnor U9416 (N_9416,N_9247,N_9263);
or U9417 (N_9417,N_9224,N_9232);
or U9418 (N_9418,N_9222,N_9181);
xnor U9419 (N_9419,N_9213,N_9282);
nor U9420 (N_9420,N_9240,N_9191);
xnor U9421 (N_9421,N_9280,N_9179);
or U9422 (N_9422,N_9151,N_9212);
and U9423 (N_9423,N_9224,N_9202);
nor U9424 (N_9424,N_9226,N_9217);
or U9425 (N_9425,N_9196,N_9254);
and U9426 (N_9426,N_9218,N_9246);
nand U9427 (N_9427,N_9283,N_9233);
or U9428 (N_9428,N_9204,N_9279);
xor U9429 (N_9429,N_9292,N_9249);
nand U9430 (N_9430,N_9271,N_9212);
nand U9431 (N_9431,N_9276,N_9230);
xnor U9432 (N_9432,N_9178,N_9242);
nor U9433 (N_9433,N_9212,N_9246);
or U9434 (N_9434,N_9196,N_9165);
xnor U9435 (N_9435,N_9188,N_9233);
and U9436 (N_9436,N_9286,N_9195);
and U9437 (N_9437,N_9259,N_9158);
or U9438 (N_9438,N_9282,N_9229);
and U9439 (N_9439,N_9281,N_9217);
and U9440 (N_9440,N_9151,N_9216);
xnor U9441 (N_9441,N_9222,N_9173);
xor U9442 (N_9442,N_9172,N_9234);
nor U9443 (N_9443,N_9231,N_9152);
xor U9444 (N_9444,N_9178,N_9225);
or U9445 (N_9445,N_9262,N_9194);
nand U9446 (N_9446,N_9191,N_9271);
nor U9447 (N_9447,N_9233,N_9214);
or U9448 (N_9448,N_9180,N_9174);
xnor U9449 (N_9449,N_9159,N_9199);
or U9450 (N_9450,N_9406,N_9370);
and U9451 (N_9451,N_9316,N_9407);
nor U9452 (N_9452,N_9385,N_9326);
xor U9453 (N_9453,N_9436,N_9338);
or U9454 (N_9454,N_9303,N_9302);
nand U9455 (N_9455,N_9318,N_9333);
or U9456 (N_9456,N_9317,N_9366);
nand U9457 (N_9457,N_9349,N_9428);
nor U9458 (N_9458,N_9341,N_9367);
nor U9459 (N_9459,N_9330,N_9364);
nand U9460 (N_9460,N_9363,N_9343);
or U9461 (N_9461,N_9380,N_9397);
or U9462 (N_9462,N_9323,N_9305);
or U9463 (N_9463,N_9405,N_9437);
and U9464 (N_9464,N_9427,N_9306);
and U9465 (N_9465,N_9342,N_9379);
or U9466 (N_9466,N_9415,N_9403);
nand U9467 (N_9467,N_9413,N_9314);
xor U9468 (N_9468,N_9441,N_9329);
and U9469 (N_9469,N_9374,N_9391);
nor U9470 (N_9470,N_9371,N_9347);
and U9471 (N_9471,N_9399,N_9402);
xor U9472 (N_9472,N_9320,N_9411);
and U9473 (N_9473,N_9313,N_9445);
nand U9474 (N_9474,N_9408,N_9404);
and U9475 (N_9475,N_9376,N_9440);
xor U9476 (N_9476,N_9373,N_9410);
xnor U9477 (N_9477,N_9360,N_9439);
or U9478 (N_9478,N_9448,N_9421);
nand U9479 (N_9479,N_9310,N_9369);
or U9480 (N_9480,N_9361,N_9429);
xnor U9481 (N_9481,N_9394,N_9426);
or U9482 (N_9482,N_9311,N_9345);
nand U9483 (N_9483,N_9433,N_9396);
nor U9484 (N_9484,N_9356,N_9322);
nand U9485 (N_9485,N_9357,N_9315);
nor U9486 (N_9486,N_9331,N_9355);
nand U9487 (N_9487,N_9312,N_9382);
or U9488 (N_9488,N_9414,N_9434);
or U9489 (N_9489,N_9419,N_9348);
and U9490 (N_9490,N_9446,N_9346);
nand U9491 (N_9491,N_9431,N_9409);
nand U9492 (N_9492,N_9447,N_9359);
xor U9493 (N_9493,N_9335,N_9358);
xnor U9494 (N_9494,N_9351,N_9352);
or U9495 (N_9495,N_9412,N_9368);
and U9496 (N_9496,N_9388,N_9389);
xnor U9497 (N_9497,N_9344,N_9377);
xnor U9498 (N_9498,N_9390,N_9332);
nand U9499 (N_9499,N_9420,N_9386);
nor U9500 (N_9500,N_9325,N_9438);
nor U9501 (N_9501,N_9400,N_9340);
xnor U9502 (N_9502,N_9319,N_9309);
and U9503 (N_9503,N_9304,N_9398);
nor U9504 (N_9504,N_9435,N_9301);
or U9505 (N_9505,N_9430,N_9444);
and U9506 (N_9506,N_9432,N_9353);
xnor U9507 (N_9507,N_9336,N_9328);
xor U9508 (N_9508,N_9378,N_9418);
nor U9509 (N_9509,N_9449,N_9422);
and U9510 (N_9510,N_9416,N_9395);
nand U9511 (N_9511,N_9443,N_9362);
nand U9512 (N_9512,N_9300,N_9375);
and U9513 (N_9513,N_9337,N_9339);
and U9514 (N_9514,N_9393,N_9387);
and U9515 (N_9515,N_9384,N_9334);
xnor U9516 (N_9516,N_9423,N_9383);
nor U9517 (N_9517,N_9442,N_9381);
nand U9518 (N_9518,N_9425,N_9321);
nand U9519 (N_9519,N_9417,N_9324);
nor U9520 (N_9520,N_9350,N_9308);
xnor U9521 (N_9521,N_9372,N_9354);
or U9522 (N_9522,N_9327,N_9424);
and U9523 (N_9523,N_9401,N_9392);
or U9524 (N_9524,N_9365,N_9307);
xor U9525 (N_9525,N_9345,N_9333);
nand U9526 (N_9526,N_9334,N_9342);
nor U9527 (N_9527,N_9376,N_9405);
nor U9528 (N_9528,N_9412,N_9340);
nand U9529 (N_9529,N_9342,N_9365);
and U9530 (N_9530,N_9401,N_9334);
or U9531 (N_9531,N_9316,N_9303);
and U9532 (N_9532,N_9315,N_9310);
and U9533 (N_9533,N_9408,N_9357);
nand U9534 (N_9534,N_9422,N_9361);
xnor U9535 (N_9535,N_9324,N_9323);
nor U9536 (N_9536,N_9358,N_9340);
and U9537 (N_9537,N_9442,N_9309);
and U9538 (N_9538,N_9368,N_9377);
nor U9539 (N_9539,N_9448,N_9396);
and U9540 (N_9540,N_9419,N_9396);
nor U9541 (N_9541,N_9423,N_9387);
nand U9542 (N_9542,N_9409,N_9349);
or U9543 (N_9543,N_9448,N_9443);
xnor U9544 (N_9544,N_9333,N_9404);
and U9545 (N_9545,N_9309,N_9353);
nand U9546 (N_9546,N_9344,N_9433);
xnor U9547 (N_9547,N_9436,N_9346);
nand U9548 (N_9548,N_9343,N_9393);
or U9549 (N_9549,N_9410,N_9437);
nor U9550 (N_9550,N_9387,N_9309);
xnor U9551 (N_9551,N_9322,N_9365);
nand U9552 (N_9552,N_9318,N_9390);
and U9553 (N_9553,N_9372,N_9393);
nand U9554 (N_9554,N_9335,N_9325);
or U9555 (N_9555,N_9333,N_9361);
or U9556 (N_9556,N_9335,N_9322);
xnor U9557 (N_9557,N_9337,N_9426);
xor U9558 (N_9558,N_9333,N_9449);
and U9559 (N_9559,N_9432,N_9308);
nor U9560 (N_9560,N_9332,N_9338);
nand U9561 (N_9561,N_9319,N_9415);
nor U9562 (N_9562,N_9419,N_9403);
nand U9563 (N_9563,N_9353,N_9422);
or U9564 (N_9564,N_9410,N_9350);
xor U9565 (N_9565,N_9368,N_9434);
nor U9566 (N_9566,N_9399,N_9401);
or U9567 (N_9567,N_9414,N_9334);
nor U9568 (N_9568,N_9395,N_9334);
nor U9569 (N_9569,N_9352,N_9444);
nor U9570 (N_9570,N_9430,N_9414);
nor U9571 (N_9571,N_9338,N_9396);
nand U9572 (N_9572,N_9413,N_9349);
or U9573 (N_9573,N_9440,N_9428);
and U9574 (N_9574,N_9417,N_9376);
xor U9575 (N_9575,N_9371,N_9346);
nor U9576 (N_9576,N_9356,N_9408);
and U9577 (N_9577,N_9430,N_9338);
xnor U9578 (N_9578,N_9394,N_9347);
or U9579 (N_9579,N_9398,N_9318);
nor U9580 (N_9580,N_9391,N_9389);
nor U9581 (N_9581,N_9418,N_9302);
and U9582 (N_9582,N_9340,N_9385);
nor U9583 (N_9583,N_9310,N_9441);
xor U9584 (N_9584,N_9354,N_9339);
nand U9585 (N_9585,N_9399,N_9365);
xor U9586 (N_9586,N_9413,N_9447);
nand U9587 (N_9587,N_9414,N_9429);
and U9588 (N_9588,N_9379,N_9367);
or U9589 (N_9589,N_9310,N_9381);
nand U9590 (N_9590,N_9317,N_9335);
nor U9591 (N_9591,N_9350,N_9416);
nand U9592 (N_9592,N_9365,N_9360);
nand U9593 (N_9593,N_9430,N_9440);
and U9594 (N_9594,N_9379,N_9386);
and U9595 (N_9595,N_9399,N_9346);
nand U9596 (N_9596,N_9362,N_9411);
nor U9597 (N_9597,N_9342,N_9438);
and U9598 (N_9598,N_9431,N_9389);
nor U9599 (N_9599,N_9362,N_9393);
nand U9600 (N_9600,N_9526,N_9542);
and U9601 (N_9601,N_9482,N_9459);
xnor U9602 (N_9602,N_9592,N_9519);
nor U9603 (N_9603,N_9552,N_9549);
and U9604 (N_9604,N_9465,N_9537);
xnor U9605 (N_9605,N_9505,N_9568);
nor U9606 (N_9606,N_9518,N_9547);
and U9607 (N_9607,N_9506,N_9462);
and U9608 (N_9608,N_9579,N_9486);
xnor U9609 (N_9609,N_9501,N_9528);
and U9610 (N_9610,N_9450,N_9531);
and U9611 (N_9611,N_9551,N_9540);
or U9612 (N_9612,N_9585,N_9480);
nor U9613 (N_9613,N_9550,N_9455);
nand U9614 (N_9614,N_9458,N_9467);
nor U9615 (N_9615,N_9577,N_9595);
nand U9616 (N_9616,N_9581,N_9495);
nor U9617 (N_9617,N_9536,N_9477);
nand U9618 (N_9618,N_9504,N_9510);
xnor U9619 (N_9619,N_9490,N_9493);
and U9620 (N_9620,N_9523,N_9586);
nand U9621 (N_9621,N_9466,N_9497);
nor U9622 (N_9622,N_9561,N_9451);
nand U9623 (N_9623,N_9529,N_9573);
nor U9624 (N_9624,N_9520,N_9479);
or U9625 (N_9625,N_9464,N_9481);
nor U9626 (N_9626,N_9570,N_9580);
xnor U9627 (N_9627,N_9484,N_9521);
nand U9628 (N_9628,N_9576,N_9475);
nor U9629 (N_9629,N_9457,N_9534);
nor U9630 (N_9630,N_9596,N_9589);
nor U9631 (N_9631,N_9485,N_9583);
nor U9632 (N_9632,N_9500,N_9470);
nand U9633 (N_9633,N_9558,N_9516);
nand U9634 (N_9634,N_9565,N_9548);
or U9635 (N_9635,N_9554,N_9532);
and U9636 (N_9636,N_9511,N_9476);
nand U9637 (N_9637,N_9498,N_9473);
and U9638 (N_9638,N_9572,N_9541);
nand U9639 (N_9639,N_9599,N_9512);
nor U9640 (N_9640,N_9453,N_9488);
nand U9641 (N_9641,N_9525,N_9494);
or U9642 (N_9642,N_9496,N_9574);
or U9643 (N_9643,N_9508,N_9503);
and U9644 (N_9644,N_9492,N_9560);
or U9645 (N_9645,N_9471,N_9489);
xnor U9646 (N_9646,N_9557,N_9566);
and U9647 (N_9647,N_9590,N_9587);
nor U9648 (N_9648,N_9502,N_9460);
xnor U9649 (N_9649,N_9527,N_9571);
xor U9650 (N_9650,N_9517,N_9544);
nand U9651 (N_9651,N_9598,N_9463);
nor U9652 (N_9652,N_9546,N_9564);
xnor U9653 (N_9653,N_9593,N_9509);
or U9654 (N_9654,N_9591,N_9569);
nand U9655 (N_9655,N_9468,N_9538);
nand U9656 (N_9656,N_9578,N_9575);
and U9657 (N_9657,N_9555,N_9515);
nor U9658 (N_9658,N_9584,N_9530);
xnor U9659 (N_9659,N_9478,N_9522);
nor U9660 (N_9660,N_9454,N_9588);
xnor U9661 (N_9661,N_9563,N_9452);
nor U9662 (N_9662,N_9483,N_9594);
or U9663 (N_9663,N_9491,N_9461);
xnor U9664 (N_9664,N_9499,N_9456);
nor U9665 (N_9665,N_9507,N_9567);
and U9666 (N_9666,N_9472,N_9582);
xnor U9667 (N_9667,N_9539,N_9545);
nand U9668 (N_9668,N_9559,N_9553);
nand U9669 (N_9669,N_9514,N_9556);
or U9670 (N_9670,N_9597,N_9524);
or U9671 (N_9671,N_9535,N_9562);
or U9672 (N_9672,N_9487,N_9543);
xor U9673 (N_9673,N_9474,N_9513);
and U9674 (N_9674,N_9533,N_9469);
and U9675 (N_9675,N_9517,N_9524);
nand U9676 (N_9676,N_9591,N_9563);
nand U9677 (N_9677,N_9527,N_9501);
or U9678 (N_9678,N_9470,N_9513);
xor U9679 (N_9679,N_9466,N_9491);
or U9680 (N_9680,N_9565,N_9534);
xor U9681 (N_9681,N_9502,N_9595);
nand U9682 (N_9682,N_9531,N_9524);
or U9683 (N_9683,N_9504,N_9597);
nand U9684 (N_9684,N_9511,N_9467);
and U9685 (N_9685,N_9531,N_9454);
or U9686 (N_9686,N_9509,N_9533);
and U9687 (N_9687,N_9541,N_9537);
nor U9688 (N_9688,N_9534,N_9460);
and U9689 (N_9689,N_9583,N_9475);
or U9690 (N_9690,N_9483,N_9487);
or U9691 (N_9691,N_9523,N_9546);
xor U9692 (N_9692,N_9593,N_9589);
and U9693 (N_9693,N_9561,N_9461);
nor U9694 (N_9694,N_9484,N_9541);
nand U9695 (N_9695,N_9584,N_9451);
or U9696 (N_9696,N_9465,N_9531);
xor U9697 (N_9697,N_9480,N_9536);
xor U9698 (N_9698,N_9454,N_9518);
nand U9699 (N_9699,N_9543,N_9595);
and U9700 (N_9700,N_9509,N_9505);
nor U9701 (N_9701,N_9539,N_9578);
or U9702 (N_9702,N_9522,N_9599);
nand U9703 (N_9703,N_9555,N_9505);
nor U9704 (N_9704,N_9474,N_9473);
nor U9705 (N_9705,N_9484,N_9511);
and U9706 (N_9706,N_9509,N_9574);
and U9707 (N_9707,N_9496,N_9571);
and U9708 (N_9708,N_9578,N_9574);
and U9709 (N_9709,N_9584,N_9498);
nor U9710 (N_9710,N_9524,N_9570);
xnor U9711 (N_9711,N_9518,N_9577);
or U9712 (N_9712,N_9493,N_9506);
nand U9713 (N_9713,N_9564,N_9572);
and U9714 (N_9714,N_9488,N_9588);
xnor U9715 (N_9715,N_9564,N_9569);
or U9716 (N_9716,N_9491,N_9579);
and U9717 (N_9717,N_9455,N_9525);
or U9718 (N_9718,N_9591,N_9514);
and U9719 (N_9719,N_9560,N_9556);
xor U9720 (N_9720,N_9548,N_9526);
nand U9721 (N_9721,N_9466,N_9494);
and U9722 (N_9722,N_9469,N_9454);
nor U9723 (N_9723,N_9510,N_9475);
nand U9724 (N_9724,N_9562,N_9500);
nand U9725 (N_9725,N_9583,N_9535);
xor U9726 (N_9726,N_9460,N_9487);
nand U9727 (N_9727,N_9526,N_9515);
xnor U9728 (N_9728,N_9501,N_9503);
nand U9729 (N_9729,N_9522,N_9509);
nand U9730 (N_9730,N_9469,N_9556);
or U9731 (N_9731,N_9567,N_9531);
or U9732 (N_9732,N_9530,N_9563);
xnor U9733 (N_9733,N_9562,N_9466);
xnor U9734 (N_9734,N_9504,N_9480);
nor U9735 (N_9735,N_9502,N_9485);
and U9736 (N_9736,N_9481,N_9558);
xor U9737 (N_9737,N_9553,N_9571);
xor U9738 (N_9738,N_9552,N_9494);
and U9739 (N_9739,N_9451,N_9465);
or U9740 (N_9740,N_9596,N_9531);
or U9741 (N_9741,N_9549,N_9495);
nor U9742 (N_9742,N_9515,N_9528);
or U9743 (N_9743,N_9476,N_9533);
xor U9744 (N_9744,N_9556,N_9553);
or U9745 (N_9745,N_9451,N_9495);
nor U9746 (N_9746,N_9529,N_9569);
nor U9747 (N_9747,N_9561,N_9525);
nor U9748 (N_9748,N_9501,N_9486);
nand U9749 (N_9749,N_9566,N_9465);
and U9750 (N_9750,N_9692,N_9611);
nand U9751 (N_9751,N_9735,N_9657);
xnor U9752 (N_9752,N_9643,N_9631);
nand U9753 (N_9753,N_9636,N_9629);
and U9754 (N_9754,N_9743,N_9724);
nor U9755 (N_9755,N_9718,N_9617);
and U9756 (N_9756,N_9690,N_9622);
or U9757 (N_9757,N_9600,N_9729);
nor U9758 (N_9758,N_9640,N_9652);
nand U9759 (N_9759,N_9702,N_9659);
and U9760 (N_9760,N_9701,N_9660);
and U9761 (N_9761,N_9608,N_9647);
or U9762 (N_9762,N_9678,N_9684);
or U9763 (N_9763,N_9697,N_9637);
nand U9764 (N_9764,N_9679,N_9700);
and U9765 (N_9765,N_9717,N_9695);
and U9766 (N_9766,N_9723,N_9696);
xor U9767 (N_9767,N_9710,N_9646);
or U9768 (N_9768,N_9747,N_9655);
nor U9769 (N_9769,N_9669,N_9601);
or U9770 (N_9770,N_9681,N_9612);
xor U9771 (N_9771,N_9736,N_9605);
or U9772 (N_9772,N_9653,N_9626);
or U9773 (N_9773,N_9663,N_9706);
nand U9774 (N_9774,N_9742,N_9651);
nand U9775 (N_9775,N_9711,N_9732);
nand U9776 (N_9776,N_9661,N_9650);
xnor U9777 (N_9777,N_9658,N_9606);
nor U9778 (N_9778,N_9632,N_9683);
and U9779 (N_9779,N_9734,N_9746);
nand U9780 (N_9780,N_9676,N_9677);
and U9781 (N_9781,N_9740,N_9728);
and U9782 (N_9782,N_9604,N_9615);
or U9783 (N_9783,N_9628,N_9727);
nor U9784 (N_9784,N_9642,N_9730);
xnor U9785 (N_9785,N_9635,N_9667);
xor U9786 (N_9786,N_9707,N_9733);
nand U9787 (N_9787,N_9648,N_9666);
nand U9788 (N_9788,N_9691,N_9694);
and U9789 (N_9789,N_9641,N_9685);
xor U9790 (N_9790,N_9686,N_9633);
nand U9791 (N_9791,N_9630,N_9712);
nand U9792 (N_9792,N_9720,N_9731);
or U9793 (N_9793,N_9644,N_9623);
xor U9794 (N_9794,N_9614,N_9674);
xor U9795 (N_9795,N_9621,N_9625);
nand U9796 (N_9796,N_9603,N_9680);
or U9797 (N_9797,N_9610,N_9748);
and U9798 (N_9798,N_9638,N_9716);
or U9799 (N_9799,N_9654,N_9639);
xor U9800 (N_9800,N_9616,N_9739);
nand U9801 (N_9801,N_9689,N_9627);
or U9802 (N_9802,N_9656,N_9607);
nor U9803 (N_9803,N_9682,N_9726);
and U9804 (N_9804,N_9725,N_9619);
and U9805 (N_9805,N_9699,N_9609);
and U9806 (N_9806,N_9721,N_9737);
nand U9807 (N_9807,N_9687,N_9704);
xnor U9808 (N_9808,N_9709,N_9645);
xor U9809 (N_9809,N_9719,N_9620);
nand U9810 (N_9810,N_9698,N_9741);
nand U9811 (N_9811,N_9708,N_9670);
nor U9812 (N_9812,N_9673,N_9668);
xnor U9813 (N_9813,N_9613,N_9688);
nand U9814 (N_9814,N_9705,N_9665);
xnor U9815 (N_9815,N_9675,N_9671);
and U9816 (N_9816,N_9672,N_9738);
and U9817 (N_9817,N_9703,N_9649);
or U9818 (N_9818,N_9602,N_9722);
or U9819 (N_9819,N_9713,N_9693);
xor U9820 (N_9820,N_9624,N_9744);
xnor U9821 (N_9821,N_9664,N_9618);
and U9822 (N_9822,N_9715,N_9745);
nor U9823 (N_9823,N_9662,N_9714);
and U9824 (N_9824,N_9749,N_9634);
or U9825 (N_9825,N_9648,N_9735);
and U9826 (N_9826,N_9660,N_9742);
nand U9827 (N_9827,N_9725,N_9739);
xor U9828 (N_9828,N_9606,N_9673);
xor U9829 (N_9829,N_9638,N_9682);
xor U9830 (N_9830,N_9706,N_9689);
nor U9831 (N_9831,N_9622,N_9679);
nand U9832 (N_9832,N_9605,N_9667);
and U9833 (N_9833,N_9623,N_9741);
nand U9834 (N_9834,N_9630,N_9709);
nand U9835 (N_9835,N_9725,N_9661);
and U9836 (N_9836,N_9712,N_9748);
nor U9837 (N_9837,N_9658,N_9731);
nor U9838 (N_9838,N_9742,N_9678);
nor U9839 (N_9839,N_9629,N_9654);
xor U9840 (N_9840,N_9644,N_9703);
and U9841 (N_9841,N_9609,N_9707);
or U9842 (N_9842,N_9618,N_9658);
xnor U9843 (N_9843,N_9689,N_9636);
nor U9844 (N_9844,N_9618,N_9725);
or U9845 (N_9845,N_9702,N_9689);
and U9846 (N_9846,N_9710,N_9602);
and U9847 (N_9847,N_9701,N_9674);
nand U9848 (N_9848,N_9704,N_9746);
or U9849 (N_9849,N_9652,N_9701);
xor U9850 (N_9850,N_9672,N_9625);
nand U9851 (N_9851,N_9715,N_9633);
or U9852 (N_9852,N_9604,N_9638);
nor U9853 (N_9853,N_9714,N_9649);
nand U9854 (N_9854,N_9655,N_9628);
xor U9855 (N_9855,N_9661,N_9678);
xor U9856 (N_9856,N_9673,N_9688);
xor U9857 (N_9857,N_9705,N_9740);
xor U9858 (N_9858,N_9684,N_9706);
nor U9859 (N_9859,N_9705,N_9634);
nor U9860 (N_9860,N_9675,N_9672);
or U9861 (N_9861,N_9720,N_9721);
nor U9862 (N_9862,N_9611,N_9661);
nor U9863 (N_9863,N_9614,N_9695);
or U9864 (N_9864,N_9696,N_9701);
nand U9865 (N_9865,N_9680,N_9704);
nand U9866 (N_9866,N_9644,N_9696);
or U9867 (N_9867,N_9640,N_9741);
and U9868 (N_9868,N_9631,N_9706);
and U9869 (N_9869,N_9707,N_9625);
and U9870 (N_9870,N_9663,N_9674);
xor U9871 (N_9871,N_9732,N_9636);
and U9872 (N_9872,N_9614,N_9640);
nor U9873 (N_9873,N_9717,N_9609);
and U9874 (N_9874,N_9725,N_9672);
and U9875 (N_9875,N_9740,N_9717);
nor U9876 (N_9876,N_9726,N_9639);
nand U9877 (N_9877,N_9622,N_9651);
or U9878 (N_9878,N_9684,N_9640);
and U9879 (N_9879,N_9647,N_9634);
xor U9880 (N_9880,N_9681,N_9719);
nor U9881 (N_9881,N_9626,N_9641);
and U9882 (N_9882,N_9722,N_9747);
nor U9883 (N_9883,N_9713,N_9622);
and U9884 (N_9884,N_9660,N_9680);
or U9885 (N_9885,N_9629,N_9746);
xnor U9886 (N_9886,N_9653,N_9639);
and U9887 (N_9887,N_9671,N_9638);
and U9888 (N_9888,N_9716,N_9608);
nand U9889 (N_9889,N_9652,N_9605);
xor U9890 (N_9890,N_9698,N_9651);
or U9891 (N_9891,N_9615,N_9603);
nor U9892 (N_9892,N_9631,N_9632);
or U9893 (N_9893,N_9671,N_9682);
nand U9894 (N_9894,N_9625,N_9740);
xnor U9895 (N_9895,N_9621,N_9639);
or U9896 (N_9896,N_9690,N_9633);
nand U9897 (N_9897,N_9716,N_9654);
xnor U9898 (N_9898,N_9635,N_9670);
xnor U9899 (N_9899,N_9683,N_9714);
xor U9900 (N_9900,N_9793,N_9829);
and U9901 (N_9901,N_9876,N_9813);
or U9902 (N_9902,N_9766,N_9798);
or U9903 (N_9903,N_9865,N_9868);
nand U9904 (N_9904,N_9825,N_9756);
and U9905 (N_9905,N_9776,N_9787);
or U9906 (N_9906,N_9899,N_9757);
nand U9907 (N_9907,N_9844,N_9788);
nand U9908 (N_9908,N_9781,N_9831);
nor U9909 (N_9909,N_9883,N_9817);
and U9910 (N_9910,N_9786,N_9790);
xor U9911 (N_9911,N_9857,N_9833);
or U9912 (N_9912,N_9862,N_9848);
and U9913 (N_9913,N_9753,N_9889);
xnor U9914 (N_9914,N_9797,N_9860);
nor U9915 (N_9915,N_9871,N_9824);
xor U9916 (N_9916,N_9769,N_9820);
xor U9917 (N_9917,N_9805,N_9891);
or U9918 (N_9918,N_9821,N_9785);
nor U9919 (N_9919,N_9750,N_9783);
nand U9920 (N_9920,N_9878,N_9839);
nor U9921 (N_9921,N_9841,N_9804);
nor U9922 (N_9922,N_9755,N_9775);
xnor U9923 (N_9923,N_9764,N_9855);
nand U9924 (N_9924,N_9759,N_9808);
nor U9925 (N_9925,N_9814,N_9890);
nor U9926 (N_9926,N_9765,N_9854);
nor U9927 (N_9927,N_9838,N_9879);
nand U9928 (N_9928,N_9880,N_9850);
nand U9929 (N_9929,N_9796,N_9751);
nor U9930 (N_9930,N_9898,N_9851);
and U9931 (N_9931,N_9822,N_9837);
nor U9932 (N_9932,N_9806,N_9877);
xor U9933 (N_9933,N_9772,N_9780);
or U9934 (N_9934,N_9810,N_9761);
and U9935 (N_9935,N_9762,N_9847);
nor U9936 (N_9936,N_9778,N_9773);
xor U9937 (N_9937,N_9859,N_9774);
nor U9938 (N_9938,N_9843,N_9894);
and U9939 (N_9939,N_9752,N_9884);
nand U9940 (N_9940,N_9858,N_9849);
and U9941 (N_9941,N_9807,N_9801);
xor U9942 (N_9942,N_9836,N_9770);
and U9943 (N_9943,N_9893,N_9784);
and U9944 (N_9944,N_9830,N_9875);
xor U9945 (N_9945,N_9792,N_9885);
or U9946 (N_9946,N_9867,N_9826);
or U9947 (N_9947,N_9815,N_9768);
and U9948 (N_9948,N_9896,N_9863);
nor U9949 (N_9949,N_9828,N_9779);
or U9950 (N_9950,N_9853,N_9861);
nor U9951 (N_9951,N_9892,N_9811);
nor U9952 (N_9952,N_9887,N_9795);
and U9953 (N_9953,N_9760,N_9818);
xor U9954 (N_9954,N_9881,N_9834);
nand U9955 (N_9955,N_9812,N_9886);
or U9956 (N_9956,N_9895,N_9809);
nand U9957 (N_9957,N_9763,N_9856);
or U9958 (N_9958,N_9800,N_9754);
xor U9959 (N_9959,N_9840,N_9872);
xor U9960 (N_9960,N_9799,N_9767);
nor U9961 (N_9961,N_9827,N_9794);
nand U9962 (N_9962,N_9864,N_9874);
nor U9963 (N_9963,N_9816,N_9777);
nor U9964 (N_9964,N_9802,N_9873);
or U9965 (N_9965,N_9852,N_9842);
nand U9966 (N_9966,N_9888,N_9782);
xor U9967 (N_9967,N_9832,N_9846);
xor U9968 (N_9968,N_9897,N_9758);
and U9969 (N_9969,N_9823,N_9866);
or U9970 (N_9970,N_9803,N_9870);
nor U9971 (N_9971,N_9845,N_9882);
nand U9972 (N_9972,N_9869,N_9789);
or U9973 (N_9973,N_9771,N_9791);
and U9974 (N_9974,N_9819,N_9835);
or U9975 (N_9975,N_9893,N_9771);
xor U9976 (N_9976,N_9799,N_9878);
and U9977 (N_9977,N_9786,N_9894);
or U9978 (N_9978,N_9864,N_9806);
and U9979 (N_9979,N_9837,N_9767);
xor U9980 (N_9980,N_9838,N_9819);
and U9981 (N_9981,N_9890,N_9834);
nor U9982 (N_9982,N_9873,N_9846);
xnor U9983 (N_9983,N_9859,N_9759);
nand U9984 (N_9984,N_9860,N_9771);
nand U9985 (N_9985,N_9823,N_9771);
nand U9986 (N_9986,N_9884,N_9847);
or U9987 (N_9987,N_9799,N_9883);
nand U9988 (N_9988,N_9811,N_9780);
xor U9989 (N_9989,N_9860,N_9866);
or U9990 (N_9990,N_9841,N_9871);
xor U9991 (N_9991,N_9819,N_9757);
xnor U9992 (N_9992,N_9788,N_9837);
or U9993 (N_9993,N_9881,N_9766);
and U9994 (N_9994,N_9773,N_9857);
nand U9995 (N_9995,N_9866,N_9801);
nor U9996 (N_9996,N_9768,N_9804);
nand U9997 (N_9997,N_9821,N_9828);
or U9998 (N_9998,N_9793,N_9759);
xor U9999 (N_9999,N_9788,N_9868);
nor U10000 (N_10000,N_9783,N_9836);
or U10001 (N_10001,N_9834,N_9791);
and U10002 (N_10002,N_9862,N_9813);
xor U10003 (N_10003,N_9782,N_9763);
nor U10004 (N_10004,N_9878,N_9787);
and U10005 (N_10005,N_9860,N_9795);
nor U10006 (N_10006,N_9802,N_9822);
or U10007 (N_10007,N_9812,N_9786);
or U10008 (N_10008,N_9779,N_9777);
nand U10009 (N_10009,N_9867,N_9855);
nand U10010 (N_10010,N_9792,N_9896);
nand U10011 (N_10011,N_9805,N_9896);
nor U10012 (N_10012,N_9823,N_9791);
nand U10013 (N_10013,N_9851,N_9755);
nand U10014 (N_10014,N_9847,N_9841);
or U10015 (N_10015,N_9875,N_9846);
nand U10016 (N_10016,N_9804,N_9874);
nand U10017 (N_10017,N_9896,N_9890);
nand U10018 (N_10018,N_9771,N_9780);
and U10019 (N_10019,N_9801,N_9806);
nand U10020 (N_10020,N_9802,N_9880);
xnor U10021 (N_10021,N_9801,N_9874);
nor U10022 (N_10022,N_9813,N_9761);
or U10023 (N_10023,N_9897,N_9872);
and U10024 (N_10024,N_9841,N_9802);
nand U10025 (N_10025,N_9816,N_9835);
or U10026 (N_10026,N_9756,N_9776);
or U10027 (N_10027,N_9820,N_9892);
nand U10028 (N_10028,N_9796,N_9887);
nor U10029 (N_10029,N_9810,N_9878);
or U10030 (N_10030,N_9815,N_9821);
and U10031 (N_10031,N_9805,N_9768);
and U10032 (N_10032,N_9884,N_9871);
or U10033 (N_10033,N_9764,N_9880);
nand U10034 (N_10034,N_9771,N_9879);
nand U10035 (N_10035,N_9757,N_9837);
or U10036 (N_10036,N_9878,N_9885);
xor U10037 (N_10037,N_9877,N_9895);
or U10038 (N_10038,N_9867,N_9863);
nor U10039 (N_10039,N_9841,N_9882);
xnor U10040 (N_10040,N_9864,N_9750);
or U10041 (N_10041,N_9767,N_9793);
or U10042 (N_10042,N_9815,N_9869);
and U10043 (N_10043,N_9844,N_9870);
or U10044 (N_10044,N_9801,N_9763);
nand U10045 (N_10045,N_9811,N_9857);
nand U10046 (N_10046,N_9752,N_9899);
xnor U10047 (N_10047,N_9792,N_9890);
nand U10048 (N_10048,N_9788,N_9762);
xnor U10049 (N_10049,N_9871,N_9878);
nor U10050 (N_10050,N_9913,N_9919);
nor U10051 (N_10051,N_9923,N_9977);
and U10052 (N_10052,N_10016,N_9989);
nor U10053 (N_10053,N_10034,N_9998);
and U10054 (N_10054,N_9941,N_10004);
xor U10055 (N_10055,N_9980,N_9905);
xor U10056 (N_10056,N_9986,N_10047);
nor U10057 (N_10057,N_9999,N_9908);
nand U10058 (N_10058,N_9962,N_9955);
nand U10059 (N_10059,N_10007,N_10020);
nor U10060 (N_10060,N_9925,N_10026);
nor U10061 (N_10061,N_10039,N_10006);
nand U10062 (N_10062,N_9951,N_9979);
nand U10063 (N_10063,N_10003,N_9964);
or U10064 (N_10064,N_9976,N_9963);
or U10065 (N_10065,N_10048,N_10038);
nand U10066 (N_10066,N_9995,N_9992);
or U10067 (N_10067,N_9982,N_9900);
nor U10068 (N_10068,N_10013,N_9965);
nor U10069 (N_10069,N_9985,N_9969);
or U10070 (N_10070,N_9987,N_10033);
nor U10071 (N_10071,N_9950,N_9944);
or U10072 (N_10072,N_10049,N_9914);
nand U10073 (N_10073,N_9947,N_9931);
xor U10074 (N_10074,N_9935,N_9975);
nor U10075 (N_10075,N_9946,N_9934);
nand U10076 (N_10076,N_9997,N_9983);
and U10077 (N_10077,N_9984,N_9937);
xor U10078 (N_10078,N_9988,N_10043);
or U10079 (N_10079,N_9996,N_9953);
nor U10080 (N_10080,N_10024,N_10015);
nor U10081 (N_10081,N_9970,N_9922);
nor U10082 (N_10082,N_9916,N_9911);
nand U10083 (N_10083,N_10040,N_9904);
nand U10084 (N_10084,N_10008,N_10036);
nand U10085 (N_10085,N_9971,N_9981);
nor U10086 (N_10086,N_10031,N_10005);
nor U10087 (N_10087,N_9939,N_9917);
and U10088 (N_10088,N_9910,N_10042);
nor U10089 (N_10089,N_9943,N_10025);
or U10090 (N_10090,N_9938,N_9952);
nor U10091 (N_10091,N_10023,N_9974);
xor U10092 (N_10092,N_9949,N_9921);
and U10093 (N_10093,N_9991,N_10045);
nand U10094 (N_10094,N_10037,N_9901);
or U10095 (N_10095,N_9993,N_10018);
and U10096 (N_10096,N_10012,N_10027);
or U10097 (N_10097,N_9930,N_9932);
or U10098 (N_10098,N_9928,N_10029);
and U10099 (N_10099,N_10035,N_9994);
and U10100 (N_10100,N_9929,N_9926);
xnor U10101 (N_10101,N_10010,N_9967);
and U10102 (N_10102,N_10041,N_9927);
nor U10103 (N_10103,N_9915,N_10009);
xor U10104 (N_10104,N_9912,N_9902);
nor U10105 (N_10105,N_9966,N_10028);
or U10106 (N_10106,N_10011,N_9978);
or U10107 (N_10107,N_9936,N_9959);
xnor U10108 (N_10108,N_10044,N_9918);
xor U10109 (N_10109,N_10046,N_9924);
nor U10110 (N_10110,N_9954,N_10032);
nor U10111 (N_10111,N_9907,N_10030);
and U10112 (N_10112,N_10001,N_9909);
nand U10113 (N_10113,N_9973,N_9957);
and U10114 (N_10114,N_10021,N_9940);
or U10115 (N_10115,N_9956,N_9903);
and U10116 (N_10116,N_10000,N_9990);
nand U10117 (N_10117,N_9945,N_9972);
nor U10118 (N_10118,N_9906,N_9958);
nor U10119 (N_10119,N_10019,N_9920);
or U10120 (N_10120,N_10017,N_9942);
nor U10121 (N_10121,N_10014,N_9960);
nand U10122 (N_10122,N_9961,N_9948);
and U10123 (N_10123,N_9933,N_10022);
nor U10124 (N_10124,N_9968,N_10002);
nand U10125 (N_10125,N_9990,N_10014);
and U10126 (N_10126,N_10047,N_9930);
xnor U10127 (N_10127,N_9956,N_10018);
and U10128 (N_10128,N_9935,N_10009);
nand U10129 (N_10129,N_9912,N_9900);
nand U10130 (N_10130,N_9950,N_9993);
nor U10131 (N_10131,N_9922,N_9964);
nand U10132 (N_10132,N_9969,N_9949);
nor U10133 (N_10133,N_9930,N_10036);
nand U10134 (N_10134,N_9915,N_9992);
xnor U10135 (N_10135,N_9943,N_9999);
or U10136 (N_10136,N_10018,N_10014);
xor U10137 (N_10137,N_10008,N_9920);
and U10138 (N_10138,N_9917,N_10021);
nand U10139 (N_10139,N_10038,N_10018);
nand U10140 (N_10140,N_9915,N_9974);
nor U10141 (N_10141,N_9969,N_10046);
and U10142 (N_10142,N_9998,N_9932);
or U10143 (N_10143,N_9919,N_10025);
nand U10144 (N_10144,N_10029,N_9993);
nor U10145 (N_10145,N_9920,N_9916);
nor U10146 (N_10146,N_9978,N_9965);
xnor U10147 (N_10147,N_9971,N_10026);
xnor U10148 (N_10148,N_9956,N_9949);
nand U10149 (N_10149,N_9903,N_10002);
and U10150 (N_10150,N_9922,N_9908);
xnor U10151 (N_10151,N_10030,N_9948);
nand U10152 (N_10152,N_9975,N_10038);
nand U10153 (N_10153,N_9917,N_9993);
or U10154 (N_10154,N_9962,N_9989);
nand U10155 (N_10155,N_10002,N_9996);
nand U10156 (N_10156,N_9948,N_10004);
or U10157 (N_10157,N_9996,N_9915);
nand U10158 (N_10158,N_9980,N_9964);
nand U10159 (N_10159,N_9930,N_9951);
nor U10160 (N_10160,N_9987,N_10045);
or U10161 (N_10161,N_10047,N_9936);
xor U10162 (N_10162,N_9920,N_9978);
and U10163 (N_10163,N_9901,N_9933);
and U10164 (N_10164,N_9971,N_10025);
or U10165 (N_10165,N_9922,N_9933);
xor U10166 (N_10166,N_9985,N_9937);
nand U10167 (N_10167,N_9912,N_10004);
nor U10168 (N_10168,N_10034,N_9902);
nand U10169 (N_10169,N_10031,N_10043);
nand U10170 (N_10170,N_9941,N_9969);
or U10171 (N_10171,N_9974,N_10046);
or U10172 (N_10172,N_9979,N_9943);
or U10173 (N_10173,N_10031,N_9977);
or U10174 (N_10174,N_9912,N_9934);
or U10175 (N_10175,N_9973,N_9969);
and U10176 (N_10176,N_9982,N_9937);
and U10177 (N_10177,N_10004,N_9986);
or U10178 (N_10178,N_9959,N_10023);
and U10179 (N_10179,N_9948,N_10045);
or U10180 (N_10180,N_9920,N_10007);
or U10181 (N_10181,N_9971,N_9907);
nor U10182 (N_10182,N_9977,N_9969);
nand U10183 (N_10183,N_10025,N_10000);
xor U10184 (N_10184,N_10011,N_9915);
nand U10185 (N_10185,N_9952,N_9981);
and U10186 (N_10186,N_9994,N_10022);
and U10187 (N_10187,N_9915,N_9967);
nor U10188 (N_10188,N_10038,N_10026);
xor U10189 (N_10189,N_9983,N_9950);
xor U10190 (N_10190,N_10020,N_9926);
nor U10191 (N_10191,N_9989,N_9991);
nand U10192 (N_10192,N_10025,N_10030);
xor U10193 (N_10193,N_10043,N_9967);
nand U10194 (N_10194,N_10004,N_9943);
and U10195 (N_10195,N_9935,N_9945);
nor U10196 (N_10196,N_10048,N_9911);
and U10197 (N_10197,N_9925,N_9958);
nor U10198 (N_10198,N_9964,N_9915);
and U10199 (N_10199,N_9974,N_9971);
nor U10200 (N_10200,N_10085,N_10191);
or U10201 (N_10201,N_10080,N_10193);
nand U10202 (N_10202,N_10093,N_10190);
nor U10203 (N_10203,N_10142,N_10186);
nor U10204 (N_10204,N_10141,N_10130);
nand U10205 (N_10205,N_10172,N_10060);
nor U10206 (N_10206,N_10051,N_10128);
nor U10207 (N_10207,N_10158,N_10167);
nand U10208 (N_10208,N_10148,N_10102);
xnor U10209 (N_10209,N_10137,N_10062);
nor U10210 (N_10210,N_10179,N_10092);
and U10211 (N_10211,N_10090,N_10108);
xor U10212 (N_10212,N_10189,N_10099);
and U10213 (N_10213,N_10112,N_10192);
nand U10214 (N_10214,N_10050,N_10087);
xnor U10215 (N_10215,N_10074,N_10098);
nand U10216 (N_10216,N_10119,N_10175);
xnor U10217 (N_10217,N_10168,N_10089);
or U10218 (N_10218,N_10164,N_10147);
xnor U10219 (N_10219,N_10053,N_10095);
xnor U10220 (N_10220,N_10161,N_10121);
and U10221 (N_10221,N_10066,N_10065);
or U10222 (N_10222,N_10151,N_10071);
nor U10223 (N_10223,N_10133,N_10152);
nand U10224 (N_10224,N_10166,N_10070);
xor U10225 (N_10225,N_10198,N_10083);
or U10226 (N_10226,N_10079,N_10131);
xor U10227 (N_10227,N_10054,N_10059);
nor U10228 (N_10228,N_10123,N_10109);
nor U10229 (N_10229,N_10155,N_10105);
nor U10230 (N_10230,N_10143,N_10110);
nand U10231 (N_10231,N_10063,N_10129);
nand U10232 (N_10232,N_10106,N_10124);
nand U10233 (N_10233,N_10178,N_10185);
nand U10234 (N_10234,N_10165,N_10199);
nand U10235 (N_10235,N_10146,N_10156);
and U10236 (N_10236,N_10180,N_10182);
nor U10237 (N_10237,N_10187,N_10169);
or U10238 (N_10238,N_10118,N_10132);
nor U10239 (N_10239,N_10096,N_10153);
nor U10240 (N_10240,N_10150,N_10068);
xor U10241 (N_10241,N_10086,N_10078);
nor U10242 (N_10242,N_10170,N_10061);
nand U10243 (N_10243,N_10094,N_10177);
nand U10244 (N_10244,N_10072,N_10184);
or U10245 (N_10245,N_10082,N_10136);
or U10246 (N_10246,N_10111,N_10194);
nand U10247 (N_10247,N_10183,N_10107);
xnor U10248 (N_10248,N_10056,N_10076);
nand U10249 (N_10249,N_10181,N_10113);
nand U10250 (N_10250,N_10157,N_10114);
xor U10251 (N_10251,N_10154,N_10067);
or U10252 (N_10252,N_10101,N_10139);
nand U10253 (N_10253,N_10075,N_10162);
nand U10254 (N_10254,N_10116,N_10077);
xnor U10255 (N_10255,N_10149,N_10126);
or U10256 (N_10256,N_10163,N_10055);
or U10257 (N_10257,N_10117,N_10127);
or U10258 (N_10258,N_10073,N_10058);
or U10259 (N_10259,N_10064,N_10174);
nand U10260 (N_10260,N_10138,N_10057);
or U10261 (N_10261,N_10197,N_10091);
xnor U10262 (N_10262,N_10097,N_10052);
or U10263 (N_10263,N_10196,N_10069);
nand U10264 (N_10264,N_10144,N_10171);
nand U10265 (N_10265,N_10125,N_10103);
xnor U10266 (N_10266,N_10195,N_10084);
or U10267 (N_10267,N_10120,N_10115);
nor U10268 (N_10268,N_10122,N_10135);
xor U10269 (N_10269,N_10159,N_10173);
and U10270 (N_10270,N_10140,N_10104);
nand U10271 (N_10271,N_10088,N_10176);
nor U10272 (N_10272,N_10081,N_10100);
and U10273 (N_10273,N_10160,N_10134);
xor U10274 (N_10274,N_10145,N_10188);
and U10275 (N_10275,N_10144,N_10069);
nand U10276 (N_10276,N_10182,N_10093);
nor U10277 (N_10277,N_10193,N_10076);
nor U10278 (N_10278,N_10069,N_10108);
nor U10279 (N_10279,N_10063,N_10147);
nor U10280 (N_10280,N_10182,N_10163);
xnor U10281 (N_10281,N_10110,N_10193);
nand U10282 (N_10282,N_10145,N_10106);
or U10283 (N_10283,N_10057,N_10124);
or U10284 (N_10284,N_10066,N_10097);
and U10285 (N_10285,N_10129,N_10143);
and U10286 (N_10286,N_10102,N_10169);
nand U10287 (N_10287,N_10106,N_10065);
or U10288 (N_10288,N_10073,N_10162);
or U10289 (N_10289,N_10145,N_10068);
nand U10290 (N_10290,N_10181,N_10067);
nand U10291 (N_10291,N_10065,N_10051);
xnor U10292 (N_10292,N_10057,N_10123);
nor U10293 (N_10293,N_10138,N_10142);
nor U10294 (N_10294,N_10151,N_10148);
xnor U10295 (N_10295,N_10143,N_10092);
nor U10296 (N_10296,N_10189,N_10073);
nor U10297 (N_10297,N_10178,N_10069);
nand U10298 (N_10298,N_10183,N_10099);
nor U10299 (N_10299,N_10087,N_10116);
xnor U10300 (N_10300,N_10141,N_10108);
or U10301 (N_10301,N_10124,N_10127);
and U10302 (N_10302,N_10124,N_10101);
nor U10303 (N_10303,N_10147,N_10051);
xor U10304 (N_10304,N_10090,N_10136);
or U10305 (N_10305,N_10147,N_10145);
and U10306 (N_10306,N_10193,N_10138);
xnor U10307 (N_10307,N_10166,N_10098);
nor U10308 (N_10308,N_10182,N_10135);
and U10309 (N_10309,N_10098,N_10185);
xnor U10310 (N_10310,N_10170,N_10135);
nor U10311 (N_10311,N_10066,N_10099);
and U10312 (N_10312,N_10138,N_10085);
and U10313 (N_10313,N_10112,N_10083);
nor U10314 (N_10314,N_10149,N_10073);
xnor U10315 (N_10315,N_10099,N_10156);
nand U10316 (N_10316,N_10088,N_10053);
nand U10317 (N_10317,N_10060,N_10107);
nor U10318 (N_10318,N_10094,N_10153);
and U10319 (N_10319,N_10106,N_10175);
nor U10320 (N_10320,N_10052,N_10086);
and U10321 (N_10321,N_10196,N_10191);
nand U10322 (N_10322,N_10180,N_10194);
nor U10323 (N_10323,N_10105,N_10069);
or U10324 (N_10324,N_10108,N_10175);
nand U10325 (N_10325,N_10085,N_10107);
nand U10326 (N_10326,N_10120,N_10055);
xnor U10327 (N_10327,N_10152,N_10159);
or U10328 (N_10328,N_10076,N_10051);
nor U10329 (N_10329,N_10145,N_10184);
or U10330 (N_10330,N_10149,N_10108);
nand U10331 (N_10331,N_10199,N_10113);
or U10332 (N_10332,N_10171,N_10098);
and U10333 (N_10333,N_10194,N_10147);
or U10334 (N_10334,N_10170,N_10183);
nor U10335 (N_10335,N_10098,N_10102);
xnor U10336 (N_10336,N_10054,N_10100);
nand U10337 (N_10337,N_10168,N_10102);
nor U10338 (N_10338,N_10131,N_10087);
nor U10339 (N_10339,N_10192,N_10109);
xor U10340 (N_10340,N_10075,N_10184);
nand U10341 (N_10341,N_10194,N_10142);
or U10342 (N_10342,N_10192,N_10107);
or U10343 (N_10343,N_10190,N_10118);
nand U10344 (N_10344,N_10190,N_10150);
or U10345 (N_10345,N_10077,N_10173);
xnor U10346 (N_10346,N_10079,N_10182);
xor U10347 (N_10347,N_10144,N_10070);
xnor U10348 (N_10348,N_10124,N_10188);
nor U10349 (N_10349,N_10168,N_10130);
xnor U10350 (N_10350,N_10252,N_10316);
nor U10351 (N_10351,N_10347,N_10245);
nand U10352 (N_10352,N_10265,N_10337);
and U10353 (N_10353,N_10280,N_10209);
nor U10354 (N_10354,N_10247,N_10326);
and U10355 (N_10355,N_10291,N_10306);
nor U10356 (N_10356,N_10323,N_10292);
or U10357 (N_10357,N_10235,N_10324);
nand U10358 (N_10358,N_10257,N_10238);
xnor U10359 (N_10359,N_10312,N_10284);
xor U10360 (N_10360,N_10200,N_10330);
nor U10361 (N_10361,N_10332,N_10283);
nand U10362 (N_10362,N_10253,N_10222);
xnor U10363 (N_10363,N_10258,N_10211);
or U10364 (N_10364,N_10321,N_10214);
xor U10365 (N_10365,N_10242,N_10348);
nor U10366 (N_10366,N_10219,N_10266);
and U10367 (N_10367,N_10307,N_10344);
nor U10368 (N_10368,N_10317,N_10327);
xnor U10369 (N_10369,N_10262,N_10213);
and U10370 (N_10370,N_10338,N_10299);
or U10371 (N_10371,N_10296,N_10276);
nand U10372 (N_10372,N_10304,N_10297);
or U10373 (N_10373,N_10249,N_10237);
nor U10374 (N_10374,N_10232,N_10329);
nand U10375 (N_10375,N_10341,N_10325);
xnor U10376 (N_10376,N_10243,N_10210);
or U10377 (N_10377,N_10349,N_10216);
and U10378 (N_10378,N_10309,N_10225);
nor U10379 (N_10379,N_10202,N_10305);
xnor U10380 (N_10380,N_10293,N_10319);
and U10381 (N_10381,N_10259,N_10256);
xor U10382 (N_10382,N_10346,N_10208);
xnor U10383 (N_10383,N_10205,N_10342);
nand U10384 (N_10384,N_10203,N_10318);
xor U10385 (N_10385,N_10272,N_10302);
nand U10386 (N_10386,N_10333,N_10335);
nand U10387 (N_10387,N_10331,N_10288);
nand U10388 (N_10388,N_10311,N_10201);
nor U10389 (N_10389,N_10287,N_10294);
and U10390 (N_10390,N_10286,N_10269);
nand U10391 (N_10391,N_10345,N_10282);
or U10392 (N_10392,N_10278,N_10221);
and U10393 (N_10393,N_10343,N_10246);
nand U10394 (N_10394,N_10261,N_10298);
nand U10395 (N_10395,N_10223,N_10322);
nand U10396 (N_10396,N_10277,N_10217);
and U10397 (N_10397,N_10239,N_10328);
or U10398 (N_10398,N_10248,N_10264);
xor U10399 (N_10399,N_10206,N_10295);
xnor U10400 (N_10400,N_10241,N_10270);
nand U10401 (N_10401,N_10320,N_10310);
and U10402 (N_10402,N_10336,N_10339);
nor U10403 (N_10403,N_10313,N_10273);
nor U10404 (N_10404,N_10224,N_10274);
and U10405 (N_10405,N_10289,N_10251);
nor U10406 (N_10406,N_10244,N_10229);
nor U10407 (N_10407,N_10303,N_10334);
nand U10408 (N_10408,N_10250,N_10240);
and U10409 (N_10409,N_10263,N_10254);
or U10410 (N_10410,N_10230,N_10260);
and U10411 (N_10411,N_10228,N_10207);
and U10412 (N_10412,N_10308,N_10227);
nand U10413 (N_10413,N_10301,N_10215);
xnor U10414 (N_10414,N_10220,N_10231);
and U10415 (N_10415,N_10314,N_10268);
xnor U10416 (N_10416,N_10285,N_10267);
nand U10417 (N_10417,N_10271,N_10234);
xnor U10418 (N_10418,N_10204,N_10340);
nor U10419 (N_10419,N_10233,N_10275);
and U10420 (N_10420,N_10279,N_10290);
xor U10421 (N_10421,N_10315,N_10300);
nand U10422 (N_10422,N_10236,N_10255);
xor U10423 (N_10423,N_10212,N_10281);
nand U10424 (N_10424,N_10218,N_10226);
and U10425 (N_10425,N_10343,N_10234);
xor U10426 (N_10426,N_10215,N_10209);
or U10427 (N_10427,N_10224,N_10328);
and U10428 (N_10428,N_10218,N_10211);
nand U10429 (N_10429,N_10306,N_10225);
or U10430 (N_10430,N_10333,N_10273);
or U10431 (N_10431,N_10288,N_10340);
or U10432 (N_10432,N_10271,N_10311);
and U10433 (N_10433,N_10281,N_10228);
xnor U10434 (N_10434,N_10346,N_10341);
nand U10435 (N_10435,N_10234,N_10219);
nor U10436 (N_10436,N_10229,N_10315);
nand U10437 (N_10437,N_10328,N_10252);
and U10438 (N_10438,N_10219,N_10308);
or U10439 (N_10439,N_10306,N_10202);
nor U10440 (N_10440,N_10326,N_10273);
nand U10441 (N_10441,N_10321,N_10337);
or U10442 (N_10442,N_10299,N_10206);
nand U10443 (N_10443,N_10256,N_10224);
or U10444 (N_10444,N_10333,N_10313);
nand U10445 (N_10445,N_10338,N_10268);
or U10446 (N_10446,N_10265,N_10289);
and U10447 (N_10447,N_10284,N_10272);
nor U10448 (N_10448,N_10281,N_10252);
and U10449 (N_10449,N_10219,N_10335);
or U10450 (N_10450,N_10278,N_10237);
nor U10451 (N_10451,N_10286,N_10221);
or U10452 (N_10452,N_10302,N_10294);
or U10453 (N_10453,N_10325,N_10281);
nand U10454 (N_10454,N_10300,N_10264);
and U10455 (N_10455,N_10221,N_10265);
nand U10456 (N_10456,N_10316,N_10279);
xnor U10457 (N_10457,N_10302,N_10295);
nor U10458 (N_10458,N_10267,N_10218);
and U10459 (N_10459,N_10222,N_10278);
nor U10460 (N_10460,N_10227,N_10306);
nor U10461 (N_10461,N_10210,N_10236);
nand U10462 (N_10462,N_10316,N_10285);
nor U10463 (N_10463,N_10312,N_10202);
or U10464 (N_10464,N_10214,N_10200);
and U10465 (N_10465,N_10272,N_10253);
xnor U10466 (N_10466,N_10303,N_10247);
nand U10467 (N_10467,N_10201,N_10251);
xor U10468 (N_10468,N_10246,N_10236);
and U10469 (N_10469,N_10268,N_10212);
nor U10470 (N_10470,N_10342,N_10226);
nand U10471 (N_10471,N_10320,N_10296);
and U10472 (N_10472,N_10343,N_10327);
xor U10473 (N_10473,N_10234,N_10241);
nor U10474 (N_10474,N_10287,N_10305);
nand U10475 (N_10475,N_10245,N_10274);
xnor U10476 (N_10476,N_10233,N_10284);
or U10477 (N_10477,N_10270,N_10306);
nand U10478 (N_10478,N_10235,N_10279);
xor U10479 (N_10479,N_10200,N_10250);
nand U10480 (N_10480,N_10265,N_10324);
xor U10481 (N_10481,N_10307,N_10316);
or U10482 (N_10482,N_10249,N_10318);
and U10483 (N_10483,N_10272,N_10331);
nor U10484 (N_10484,N_10220,N_10226);
nor U10485 (N_10485,N_10266,N_10255);
nand U10486 (N_10486,N_10253,N_10291);
xor U10487 (N_10487,N_10254,N_10341);
and U10488 (N_10488,N_10282,N_10283);
or U10489 (N_10489,N_10324,N_10299);
nor U10490 (N_10490,N_10218,N_10306);
and U10491 (N_10491,N_10335,N_10250);
nor U10492 (N_10492,N_10321,N_10326);
and U10493 (N_10493,N_10303,N_10295);
xor U10494 (N_10494,N_10312,N_10263);
and U10495 (N_10495,N_10309,N_10222);
nand U10496 (N_10496,N_10224,N_10290);
nand U10497 (N_10497,N_10341,N_10234);
xor U10498 (N_10498,N_10300,N_10281);
or U10499 (N_10499,N_10212,N_10302);
nand U10500 (N_10500,N_10417,N_10485);
nand U10501 (N_10501,N_10449,N_10453);
xnor U10502 (N_10502,N_10462,N_10472);
nand U10503 (N_10503,N_10437,N_10484);
and U10504 (N_10504,N_10441,N_10412);
and U10505 (N_10505,N_10434,N_10439);
and U10506 (N_10506,N_10460,N_10388);
or U10507 (N_10507,N_10474,N_10487);
nand U10508 (N_10508,N_10406,N_10461);
or U10509 (N_10509,N_10360,N_10433);
or U10510 (N_10510,N_10410,N_10395);
nand U10511 (N_10511,N_10425,N_10436);
and U10512 (N_10512,N_10498,N_10390);
nor U10513 (N_10513,N_10481,N_10483);
or U10514 (N_10514,N_10391,N_10473);
nor U10515 (N_10515,N_10418,N_10414);
and U10516 (N_10516,N_10429,N_10488);
nand U10517 (N_10517,N_10421,N_10468);
or U10518 (N_10518,N_10435,N_10445);
xnor U10519 (N_10519,N_10364,N_10399);
or U10520 (N_10520,N_10374,N_10407);
and U10521 (N_10521,N_10358,N_10448);
nand U10522 (N_10522,N_10478,N_10416);
xor U10523 (N_10523,N_10423,N_10367);
nor U10524 (N_10524,N_10496,N_10464);
nand U10525 (N_10525,N_10394,N_10420);
nand U10526 (N_10526,N_10396,N_10438);
or U10527 (N_10527,N_10353,N_10440);
nor U10528 (N_10528,N_10476,N_10424);
nor U10529 (N_10529,N_10404,N_10446);
xor U10530 (N_10530,N_10432,N_10368);
or U10531 (N_10531,N_10456,N_10465);
and U10532 (N_10532,N_10389,N_10385);
nand U10533 (N_10533,N_10359,N_10492);
nor U10534 (N_10534,N_10370,N_10383);
xnor U10535 (N_10535,N_10379,N_10402);
nor U10536 (N_10536,N_10447,N_10428);
xnor U10537 (N_10537,N_10470,N_10378);
xnor U10538 (N_10538,N_10415,N_10467);
or U10539 (N_10539,N_10362,N_10398);
or U10540 (N_10540,N_10377,N_10463);
nand U10541 (N_10541,N_10422,N_10450);
or U10542 (N_10542,N_10366,N_10430);
xnor U10543 (N_10543,N_10405,N_10486);
or U10544 (N_10544,N_10471,N_10499);
or U10545 (N_10545,N_10451,N_10419);
xnor U10546 (N_10546,N_10427,N_10459);
nand U10547 (N_10547,N_10490,N_10466);
nand U10548 (N_10548,N_10371,N_10452);
or U10549 (N_10549,N_10493,N_10469);
and U10550 (N_10550,N_10477,N_10357);
or U10551 (N_10551,N_10431,N_10455);
or U10552 (N_10552,N_10384,N_10443);
nand U10553 (N_10553,N_10400,N_10403);
nand U10554 (N_10554,N_10475,N_10409);
or U10555 (N_10555,N_10458,N_10392);
xnor U10556 (N_10556,N_10387,N_10376);
nand U10557 (N_10557,N_10386,N_10375);
xnor U10558 (N_10558,N_10401,N_10356);
and U10559 (N_10559,N_10480,N_10369);
nor U10560 (N_10560,N_10381,N_10408);
and U10561 (N_10561,N_10489,N_10363);
xnor U10562 (N_10562,N_10351,N_10380);
nor U10563 (N_10563,N_10393,N_10350);
nand U10564 (N_10564,N_10457,N_10491);
xnor U10565 (N_10565,N_10495,N_10411);
xnor U10566 (N_10566,N_10354,N_10413);
or U10567 (N_10567,N_10361,N_10355);
and U10568 (N_10568,N_10479,N_10444);
xor U10569 (N_10569,N_10494,N_10482);
nor U10570 (N_10570,N_10352,N_10373);
xor U10571 (N_10571,N_10382,N_10372);
nor U10572 (N_10572,N_10497,N_10397);
nor U10573 (N_10573,N_10454,N_10426);
and U10574 (N_10574,N_10442,N_10365);
nand U10575 (N_10575,N_10401,N_10489);
and U10576 (N_10576,N_10497,N_10372);
or U10577 (N_10577,N_10382,N_10450);
nand U10578 (N_10578,N_10358,N_10427);
and U10579 (N_10579,N_10496,N_10404);
nand U10580 (N_10580,N_10483,N_10385);
or U10581 (N_10581,N_10460,N_10435);
and U10582 (N_10582,N_10424,N_10453);
xor U10583 (N_10583,N_10353,N_10370);
nor U10584 (N_10584,N_10364,N_10387);
or U10585 (N_10585,N_10471,N_10442);
xor U10586 (N_10586,N_10448,N_10391);
xor U10587 (N_10587,N_10453,N_10404);
and U10588 (N_10588,N_10440,N_10482);
xor U10589 (N_10589,N_10390,N_10362);
nor U10590 (N_10590,N_10472,N_10449);
or U10591 (N_10591,N_10350,N_10434);
xor U10592 (N_10592,N_10478,N_10377);
nor U10593 (N_10593,N_10440,N_10374);
nor U10594 (N_10594,N_10489,N_10440);
and U10595 (N_10595,N_10360,N_10362);
or U10596 (N_10596,N_10490,N_10454);
xnor U10597 (N_10597,N_10494,N_10459);
nor U10598 (N_10598,N_10431,N_10430);
or U10599 (N_10599,N_10493,N_10474);
xnor U10600 (N_10600,N_10375,N_10439);
nor U10601 (N_10601,N_10444,N_10437);
and U10602 (N_10602,N_10375,N_10354);
xor U10603 (N_10603,N_10480,N_10442);
or U10604 (N_10604,N_10390,N_10478);
nand U10605 (N_10605,N_10468,N_10373);
xnor U10606 (N_10606,N_10434,N_10404);
xnor U10607 (N_10607,N_10425,N_10498);
nand U10608 (N_10608,N_10396,N_10456);
xor U10609 (N_10609,N_10402,N_10458);
or U10610 (N_10610,N_10463,N_10372);
or U10611 (N_10611,N_10389,N_10408);
xor U10612 (N_10612,N_10447,N_10400);
or U10613 (N_10613,N_10428,N_10414);
and U10614 (N_10614,N_10360,N_10492);
nand U10615 (N_10615,N_10443,N_10454);
or U10616 (N_10616,N_10458,N_10394);
nand U10617 (N_10617,N_10494,N_10464);
nand U10618 (N_10618,N_10403,N_10460);
nand U10619 (N_10619,N_10464,N_10379);
and U10620 (N_10620,N_10353,N_10433);
nand U10621 (N_10621,N_10375,N_10369);
or U10622 (N_10622,N_10481,N_10355);
and U10623 (N_10623,N_10358,N_10478);
nor U10624 (N_10624,N_10361,N_10439);
nor U10625 (N_10625,N_10441,N_10388);
xnor U10626 (N_10626,N_10387,N_10412);
and U10627 (N_10627,N_10401,N_10424);
or U10628 (N_10628,N_10447,N_10413);
nand U10629 (N_10629,N_10480,N_10438);
nor U10630 (N_10630,N_10499,N_10373);
and U10631 (N_10631,N_10450,N_10454);
or U10632 (N_10632,N_10442,N_10387);
or U10633 (N_10633,N_10375,N_10484);
and U10634 (N_10634,N_10380,N_10391);
nor U10635 (N_10635,N_10369,N_10363);
or U10636 (N_10636,N_10367,N_10467);
and U10637 (N_10637,N_10470,N_10410);
nor U10638 (N_10638,N_10462,N_10450);
nand U10639 (N_10639,N_10368,N_10379);
nor U10640 (N_10640,N_10482,N_10383);
and U10641 (N_10641,N_10476,N_10426);
nor U10642 (N_10642,N_10418,N_10397);
xor U10643 (N_10643,N_10392,N_10426);
nor U10644 (N_10644,N_10441,N_10462);
and U10645 (N_10645,N_10486,N_10383);
nand U10646 (N_10646,N_10437,N_10400);
nor U10647 (N_10647,N_10404,N_10410);
nor U10648 (N_10648,N_10424,N_10448);
or U10649 (N_10649,N_10415,N_10391);
and U10650 (N_10650,N_10552,N_10558);
xor U10651 (N_10651,N_10576,N_10637);
xor U10652 (N_10652,N_10572,N_10575);
nand U10653 (N_10653,N_10528,N_10557);
and U10654 (N_10654,N_10638,N_10589);
or U10655 (N_10655,N_10596,N_10504);
or U10656 (N_10656,N_10643,N_10644);
xor U10657 (N_10657,N_10615,N_10537);
or U10658 (N_10658,N_10559,N_10619);
nor U10659 (N_10659,N_10505,N_10509);
xnor U10660 (N_10660,N_10533,N_10569);
nor U10661 (N_10661,N_10592,N_10579);
nand U10662 (N_10662,N_10590,N_10609);
or U10663 (N_10663,N_10546,N_10600);
or U10664 (N_10664,N_10525,N_10628);
nand U10665 (N_10665,N_10621,N_10587);
xnor U10666 (N_10666,N_10577,N_10636);
nor U10667 (N_10667,N_10535,N_10648);
and U10668 (N_10668,N_10642,N_10607);
xnor U10669 (N_10669,N_10622,N_10601);
and U10670 (N_10670,N_10503,N_10549);
or U10671 (N_10671,N_10554,N_10624);
nor U10672 (N_10672,N_10581,N_10570);
and U10673 (N_10673,N_10595,N_10632);
and U10674 (N_10674,N_10620,N_10556);
or U10675 (N_10675,N_10594,N_10510);
nor U10676 (N_10676,N_10586,N_10597);
xnor U10677 (N_10677,N_10573,N_10560);
and U10678 (N_10678,N_10611,N_10605);
or U10679 (N_10679,N_10538,N_10530);
nand U10680 (N_10680,N_10531,N_10555);
xor U10681 (N_10681,N_10539,N_10565);
nor U10682 (N_10682,N_10616,N_10629);
or U10683 (N_10683,N_10604,N_10567);
nor U10684 (N_10684,N_10647,N_10522);
nor U10685 (N_10685,N_10519,N_10623);
and U10686 (N_10686,N_10591,N_10610);
nor U10687 (N_10687,N_10551,N_10588);
nand U10688 (N_10688,N_10630,N_10526);
nand U10689 (N_10689,N_10614,N_10548);
nor U10690 (N_10690,N_10512,N_10515);
nor U10691 (N_10691,N_10568,N_10534);
or U10692 (N_10692,N_10529,N_10527);
nor U10693 (N_10693,N_10646,N_10547);
nor U10694 (N_10694,N_10521,N_10608);
or U10695 (N_10695,N_10585,N_10511);
nor U10696 (N_10696,N_10544,N_10541);
nand U10697 (N_10697,N_10625,N_10574);
nand U10698 (N_10698,N_10513,N_10593);
and U10699 (N_10699,N_10536,N_10641);
and U10700 (N_10700,N_10516,N_10550);
and U10701 (N_10701,N_10517,N_10598);
or U10702 (N_10702,N_10520,N_10545);
xor U10703 (N_10703,N_10553,N_10603);
and U10704 (N_10704,N_10501,N_10612);
xor U10705 (N_10705,N_10571,N_10602);
or U10706 (N_10706,N_10508,N_10561);
and U10707 (N_10707,N_10502,N_10532);
or U10708 (N_10708,N_10631,N_10645);
xnor U10709 (N_10709,N_10566,N_10627);
and U10710 (N_10710,N_10562,N_10506);
nand U10711 (N_10711,N_10640,N_10584);
xnor U10712 (N_10712,N_10580,N_10613);
nor U10713 (N_10713,N_10626,N_10563);
or U10714 (N_10714,N_10617,N_10582);
or U10715 (N_10715,N_10543,N_10514);
nand U10716 (N_10716,N_10649,N_10635);
and U10717 (N_10717,N_10606,N_10523);
nand U10718 (N_10718,N_10633,N_10639);
xor U10719 (N_10719,N_10542,N_10564);
or U10720 (N_10720,N_10578,N_10599);
nor U10721 (N_10721,N_10500,N_10518);
nand U10722 (N_10722,N_10540,N_10524);
or U10723 (N_10723,N_10507,N_10618);
or U10724 (N_10724,N_10634,N_10583);
nand U10725 (N_10725,N_10578,N_10554);
nor U10726 (N_10726,N_10539,N_10644);
xor U10727 (N_10727,N_10536,N_10634);
xnor U10728 (N_10728,N_10577,N_10605);
or U10729 (N_10729,N_10535,N_10618);
xor U10730 (N_10730,N_10524,N_10566);
nor U10731 (N_10731,N_10589,N_10503);
nor U10732 (N_10732,N_10563,N_10505);
or U10733 (N_10733,N_10539,N_10648);
or U10734 (N_10734,N_10604,N_10615);
or U10735 (N_10735,N_10500,N_10585);
and U10736 (N_10736,N_10500,N_10620);
xor U10737 (N_10737,N_10540,N_10539);
xnor U10738 (N_10738,N_10629,N_10584);
xnor U10739 (N_10739,N_10580,N_10597);
nand U10740 (N_10740,N_10559,N_10628);
or U10741 (N_10741,N_10618,N_10629);
and U10742 (N_10742,N_10551,N_10613);
or U10743 (N_10743,N_10539,N_10549);
and U10744 (N_10744,N_10586,N_10620);
xor U10745 (N_10745,N_10571,N_10646);
nor U10746 (N_10746,N_10551,N_10635);
xnor U10747 (N_10747,N_10516,N_10517);
nand U10748 (N_10748,N_10501,N_10503);
or U10749 (N_10749,N_10531,N_10525);
xor U10750 (N_10750,N_10635,N_10503);
nor U10751 (N_10751,N_10609,N_10602);
xnor U10752 (N_10752,N_10557,N_10641);
nand U10753 (N_10753,N_10639,N_10638);
xor U10754 (N_10754,N_10647,N_10547);
nand U10755 (N_10755,N_10501,N_10642);
and U10756 (N_10756,N_10554,N_10623);
nor U10757 (N_10757,N_10594,N_10614);
nand U10758 (N_10758,N_10549,N_10508);
nand U10759 (N_10759,N_10557,N_10545);
xor U10760 (N_10760,N_10602,N_10579);
xor U10761 (N_10761,N_10506,N_10513);
nand U10762 (N_10762,N_10598,N_10613);
or U10763 (N_10763,N_10534,N_10502);
or U10764 (N_10764,N_10586,N_10580);
nor U10765 (N_10765,N_10605,N_10502);
nand U10766 (N_10766,N_10636,N_10616);
and U10767 (N_10767,N_10519,N_10535);
xor U10768 (N_10768,N_10533,N_10626);
nand U10769 (N_10769,N_10522,N_10561);
xor U10770 (N_10770,N_10558,N_10546);
xor U10771 (N_10771,N_10515,N_10559);
xnor U10772 (N_10772,N_10556,N_10533);
or U10773 (N_10773,N_10578,N_10648);
xnor U10774 (N_10774,N_10510,N_10561);
or U10775 (N_10775,N_10560,N_10604);
xor U10776 (N_10776,N_10543,N_10571);
nor U10777 (N_10777,N_10501,N_10579);
nand U10778 (N_10778,N_10521,N_10568);
xnor U10779 (N_10779,N_10617,N_10545);
xnor U10780 (N_10780,N_10599,N_10618);
or U10781 (N_10781,N_10522,N_10644);
nor U10782 (N_10782,N_10557,N_10505);
nand U10783 (N_10783,N_10574,N_10532);
xor U10784 (N_10784,N_10559,N_10621);
or U10785 (N_10785,N_10501,N_10566);
nor U10786 (N_10786,N_10646,N_10512);
and U10787 (N_10787,N_10637,N_10577);
or U10788 (N_10788,N_10577,N_10601);
nor U10789 (N_10789,N_10629,N_10619);
and U10790 (N_10790,N_10506,N_10569);
nand U10791 (N_10791,N_10647,N_10549);
or U10792 (N_10792,N_10541,N_10513);
xnor U10793 (N_10793,N_10643,N_10578);
nand U10794 (N_10794,N_10567,N_10558);
or U10795 (N_10795,N_10555,N_10572);
nor U10796 (N_10796,N_10610,N_10503);
nor U10797 (N_10797,N_10638,N_10509);
or U10798 (N_10798,N_10525,N_10615);
nor U10799 (N_10799,N_10535,N_10639);
nor U10800 (N_10800,N_10798,N_10788);
nor U10801 (N_10801,N_10734,N_10762);
nand U10802 (N_10802,N_10696,N_10732);
nand U10803 (N_10803,N_10745,N_10768);
or U10804 (N_10804,N_10786,N_10677);
nor U10805 (N_10805,N_10664,N_10695);
nor U10806 (N_10806,N_10752,N_10766);
and U10807 (N_10807,N_10694,N_10678);
nand U10808 (N_10808,N_10778,N_10785);
nor U10809 (N_10809,N_10708,N_10735);
or U10810 (N_10810,N_10739,N_10757);
nand U10811 (N_10811,N_10730,N_10689);
nor U10812 (N_10812,N_10736,N_10715);
nor U10813 (N_10813,N_10772,N_10775);
nor U10814 (N_10814,N_10780,N_10665);
xor U10815 (N_10815,N_10713,N_10661);
and U10816 (N_10816,N_10748,N_10751);
or U10817 (N_10817,N_10763,N_10783);
or U10818 (N_10818,N_10776,N_10687);
or U10819 (N_10819,N_10784,N_10740);
xor U10820 (N_10820,N_10667,N_10723);
or U10821 (N_10821,N_10765,N_10790);
or U10822 (N_10822,N_10704,N_10685);
nand U10823 (N_10823,N_10753,N_10720);
or U10824 (N_10824,N_10681,N_10705);
nor U10825 (N_10825,N_10682,N_10721);
nand U10826 (N_10826,N_10668,N_10683);
or U10827 (N_10827,N_10794,N_10722);
xor U10828 (N_10828,N_10650,N_10759);
nand U10829 (N_10829,N_10746,N_10737);
nor U10830 (N_10830,N_10669,N_10652);
or U10831 (N_10831,N_10701,N_10719);
or U10832 (N_10832,N_10684,N_10754);
nor U10833 (N_10833,N_10770,N_10771);
or U10834 (N_10834,N_10744,N_10698);
or U10835 (N_10835,N_10797,N_10769);
xnor U10836 (N_10836,N_10699,N_10756);
or U10837 (N_10837,N_10666,N_10660);
nand U10838 (N_10838,N_10654,N_10755);
nand U10839 (N_10839,N_10659,N_10738);
and U10840 (N_10840,N_10706,N_10657);
nor U10841 (N_10841,N_10725,N_10728);
xnor U10842 (N_10842,N_10727,N_10716);
or U10843 (N_10843,N_10764,N_10792);
or U10844 (N_10844,N_10761,N_10747);
nand U10845 (N_10845,N_10658,N_10789);
and U10846 (N_10846,N_10697,N_10714);
and U10847 (N_10847,N_10679,N_10675);
nor U10848 (N_10848,N_10796,N_10782);
or U10849 (N_10849,N_10710,N_10731);
xor U10850 (N_10850,N_10651,N_10767);
nor U10851 (N_10851,N_10676,N_10733);
xnor U10852 (N_10852,N_10717,N_10707);
nor U10853 (N_10853,N_10758,N_10799);
nand U10854 (N_10854,N_10680,N_10703);
nand U10855 (N_10855,N_10691,N_10724);
or U10856 (N_10856,N_10711,N_10779);
nor U10857 (N_10857,N_10655,N_10686);
nor U10858 (N_10858,N_10760,N_10791);
nor U10859 (N_10859,N_10787,N_10673);
nor U10860 (N_10860,N_10749,N_10670);
and U10861 (N_10861,N_10742,N_10656);
and U10862 (N_10862,N_10729,N_10741);
nor U10863 (N_10863,N_10793,N_10690);
or U10864 (N_10864,N_10663,N_10774);
and U10865 (N_10865,N_10672,N_10702);
nor U10866 (N_10866,N_10743,N_10750);
nand U10867 (N_10867,N_10773,N_10662);
or U10868 (N_10868,N_10671,N_10712);
nor U10869 (N_10869,N_10777,N_10726);
or U10870 (N_10870,N_10781,N_10795);
and U10871 (N_10871,N_10700,N_10688);
xnor U10872 (N_10872,N_10692,N_10653);
nand U10873 (N_10873,N_10674,N_10709);
xor U10874 (N_10874,N_10718,N_10693);
nor U10875 (N_10875,N_10759,N_10712);
and U10876 (N_10876,N_10733,N_10670);
nand U10877 (N_10877,N_10757,N_10758);
or U10878 (N_10878,N_10799,N_10702);
xnor U10879 (N_10879,N_10710,N_10701);
nand U10880 (N_10880,N_10672,N_10762);
nand U10881 (N_10881,N_10779,N_10767);
or U10882 (N_10882,N_10799,N_10673);
nand U10883 (N_10883,N_10659,N_10655);
or U10884 (N_10884,N_10657,N_10663);
nand U10885 (N_10885,N_10725,N_10664);
nor U10886 (N_10886,N_10730,N_10672);
xnor U10887 (N_10887,N_10677,N_10780);
and U10888 (N_10888,N_10700,N_10780);
or U10889 (N_10889,N_10669,N_10763);
xor U10890 (N_10890,N_10772,N_10745);
nor U10891 (N_10891,N_10723,N_10776);
and U10892 (N_10892,N_10654,N_10793);
nand U10893 (N_10893,N_10686,N_10674);
and U10894 (N_10894,N_10652,N_10675);
nand U10895 (N_10895,N_10785,N_10701);
or U10896 (N_10896,N_10736,N_10711);
xor U10897 (N_10897,N_10712,N_10743);
nand U10898 (N_10898,N_10767,N_10794);
or U10899 (N_10899,N_10766,N_10693);
or U10900 (N_10900,N_10665,N_10757);
or U10901 (N_10901,N_10786,N_10707);
and U10902 (N_10902,N_10701,N_10680);
and U10903 (N_10903,N_10669,N_10664);
and U10904 (N_10904,N_10744,N_10739);
and U10905 (N_10905,N_10754,N_10706);
or U10906 (N_10906,N_10761,N_10786);
nand U10907 (N_10907,N_10765,N_10705);
xnor U10908 (N_10908,N_10680,N_10711);
and U10909 (N_10909,N_10797,N_10731);
xnor U10910 (N_10910,N_10670,N_10662);
and U10911 (N_10911,N_10710,N_10737);
nor U10912 (N_10912,N_10768,N_10720);
or U10913 (N_10913,N_10737,N_10663);
nor U10914 (N_10914,N_10662,N_10759);
xor U10915 (N_10915,N_10717,N_10740);
nor U10916 (N_10916,N_10737,N_10689);
nor U10917 (N_10917,N_10761,N_10704);
and U10918 (N_10918,N_10675,N_10781);
nand U10919 (N_10919,N_10732,N_10656);
nor U10920 (N_10920,N_10730,N_10702);
xnor U10921 (N_10921,N_10723,N_10686);
and U10922 (N_10922,N_10689,N_10728);
nor U10923 (N_10923,N_10673,N_10671);
or U10924 (N_10924,N_10767,N_10792);
nand U10925 (N_10925,N_10701,N_10741);
or U10926 (N_10926,N_10705,N_10650);
nor U10927 (N_10927,N_10731,N_10746);
nor U10928 (N_10928,N_10674,N_10667);
xnor U10929 (N_10929,N_10792,N_10771);
and U10930 (N_10930,N_10656,N_10751);
nand U10931 (N_10931,N_10754,N_10740);
nor U10932 (N_10932,N_10757,N_10664);
nor U10933 (N_10933,N_10706,N_10715);
and U10934 (N_10934,N_10660,N_10654);
nand U10935 (N_10935,N_10759,N_10778);
xnor U10936 (N_10936,N_10682,N_10799);
nand U10937 (N_10937,N_10737,N_10690);
xor U10938 (N_10938,N_10727,N_10774);
and U10939 (N_10939,N_10739,N_10660);
nor U10940 (N_10940,N_10704,N_10667);
xor U10941 (N_10941,N_10746,N_10680);
nor U10942 (N_10942,N_10752,N_10651);
or U10943 (N_10943,N_10683,N_10777);
nand U10944 (N_10944,N_10736,N_10744);
or U10945 (N_10945,N_10742,N_10752);
nor U10946 (N_10946,N_10682,N_10684);
and U10947 (N_10947,N_10742,N_10654);
nor U10948 (N_10948,N_10678,N_10778);
nand U10949 (N_10949,N_10758,N_10660);
nand U10950 (N_10950,N_10868,N_10894);
nor U10951 (N_10951,N_10943,N_10877);
and U10952 (N_10952,N_10909,N_10862);
nor U10953 (N_10953,N_10929,N_10856);
xor U10954 (N_10954,N_10828,N_10802);
nand U10955 (N_10955,N_10801,N_10916);
nor U10956 (N_10956,N_10865,N_10899);
and U10957 (N_10957,N_10849,N_10942);
xnor U10958 (N_10958,N_10810,N_10923);
nand U10959 (N_10959,N_10816,N_10852);
nor U10960 (N_10960,N_10872,N_10863);
nand U10961 (N_10961,N_10926,N_10815);
nor U10962 (N_10962,N_10891,N_10813);
nand U10963 (N_10963,N_10911,N_10866);
nor U10964 (N_10964,N_10887,N_10913);
nand U10965 (N_10965,N_10915,N_10833);
xnor U10966 (N_10966,N_10857,N_10830);
or U10967 (N_10967,N_10897,N_10914);
nor U10968 (N_10968,N_10859,N_10837);
or U10969 (N_10969,N_10920,N_10807);
nand U10970 (N_10970,N_10876,N_10935);
xnor U10971 (N_10971,N_10917,N_10853);
nand U10972 (N_10972,N_10896,N_10928);
or U10973 (N_10973,N_10886,N_10930);
nor U10974 (N_10974,N_10846,N_10808);
nor U10975 (N_10975,N_10944,N_10947);
or U10976 (N_10976,N_10939,N_10882);
and U10977 (N_10977,N_10925,N_10860);
nor U10978 (N_10978,N_10805,N_10905);
nand U10979 (N_10979,N_10873,N_10812);
nor U10980 (N_10980,N_10848,N_10927);
nand U10981 (N_10981,N_10893,N_10839);
or U10982 (N_10982,N_10821,N_10870);
nand U10983 (N_10983,N_10847,N_10824);
xnor U10984 (N_10984,N_10900,N_10831);
and U10985 (N_10985,N_10888,N_10902);
nor U10986 (N_10986,N_10945,N_10861);
or U10987 (N_10987,N_10921,N_10814);
nor U10988 (N_10988,N_10835,N_10883);
and U10989 (N_10989,N_10910,N_10843);
or U10990 (N_10990,N_10912,N_10803);
and U10991 (N_10991,N_10871,N_10858);
nor U10992 (N_10992,N_10841,N_10885);
nand U10993 (N_10993,N_10949,N_10834);
nand U10994 (N_10994,N_10948,N_10844);
nor U10995 (N_10995,N_10820,N_10881);
nor U10996 (N_10996,N_10937,N_10867);
nor U10997 (N_10997,N_10880,N_10869);
nand U10998 (N_10998,N_10931,N_10879);
or U10999 (N_10999,N_10918,N_10800);
nor U11000 (N_11000,N_10822,N_10832);
and U11001 (N_11001,N_10884,N_10903);
or U11002 (N_11002,N_10850,N_10875);
xnor U11003 (N_11003,N_10818,N_10845);
or U11004 (N_11004,N_10809,N_10936);
or U11005 (N_11005,N_10878,N_10804);
nor U11006 (N_11006,N_10842,N_10901);
xnor U11007 (N_11007,N_10932,N_10940);
xor U11008 (N_11008,N_10836,N_10892);
nand U11009 (N_11009,N_10919,N_10934);
or U11010 (N_11010,N_10906,N_10825);
nand U11011 (N_11011,N_10806,N_10890);
nor U11012 (N_11012,N_10889,N_10907);
or U11013 (N_11013,N_10840,N_10898);
nand U11014 (N_11014,N_10895,N_10933);
and U11015 (N_11015,N_10855,N_10908);
nor U11016 (N_11016,N_10829,N_10811);
and U11017 (N_11017,N_10864,N_10938);
xnor U11018 (N_11018,N_10941,N_10817);
nor U11019 (N_11019,N_10838,N_10819);
nand U11020 (N_11020,N_10924,N_10851);
nor U11021 (N_11021,N_10826,N_10904);
and U11022 (N_11022,N_10946,N_10823);
or U11023 (N_11023,N_10827,N_10922);
nand U11024 (N_11024,N_10854,N_10874);
xor U11025 (N_11025,N_10906,N_10877);
and U11026 (N_11026,N_10852,N_10865);
and U11027 (N_11027,N_10813,N_10876);
and U11028 (N_11028,N_10893,N_10827);
nand U11029 (N_11029,N_10836,N_10876);
nor U11030 (N_11030,N_10817,N_10834);
nor U11031 (N_11031,N_10934,N_10925);
and U11032 (N_11032,N_10863,N_10878);
xnor U11033 (N_11033,N_10922,N_10876);
nand U11034 (N_11034,N_10803,N_10866);
and U11035 (N_11035,N_10927,N_10937);
or U11036 (N_11036,N_10836,N_10841);
and U11037 (N_11037,N_10819,N_10903);
nand U11038 (N_11038,N_10817,N_10930);
xor U11039 (N_11039,N_10859,N_10943);
xor U11040 (N_11040,N_10823,N_10818);
nor U11041 (N_11041,N_10915,N_10935);
nor U11042 (N_11042,N_10928,N_10843);
nor U11043 (N_11043,N_10855,N_10879);
xor U11044 (N_11044,N_10942,N_10817);
nor U11045 (N_11045,N_10924,N_10808);
nand U11046 (N_11046,N_10880,N_10830);
or U11047 (N_11047,N_10882,N_10809);
or U11048 (N_11048,N_10863,N_10862);
nand U11049 (N_11049,N_10948,N_10859);
nor U11050 (N_11050,N_10889,N_10807);
xnor U11051 (N_11051,N_10835,N_10881);
nand U11052 (N_11052,N_10883,N_10847);
and U11053 (N_11053,N_10908,N_10833);
nand U11054 (N_11054,N_10876,N_10917);
nand U11055 (N_11055,N_10854,N_10906);
xnor U11056 (N_11056,N_10865,N_10809);
and U11057 (N_11057,N_10936,N_10833);
and U11058 (N_11058,N_10857,N_10810);
nor U11059 (N_11059,N_10830,N_10940);
nor U11060 (N_11060,N_10829,N_10942);
nand U11061 (N_11061,N_10811,N_10816);
or U11062 (N_11062,N_10933,N_10864);
and U11063 (N_11063,N_10920,N_10868);
nor U11064 (N_11064,N_10898,N_10873);
nand U11065 (N_11065,N_10889,N_10928);
or U11066 (N_11066,N_10939,N_10846);
nor U11067 (N_11067,N_10832,N_10885);
and U11068 (N_11068,N_10852,N_10932);
xnor U11069 (N_11069,N_10905,N_10943);
and U11070 (N_11070,N_10846,N_10871);
nor U11071 (N_11071,N_10904,N_10840);
nand U11072 (N_11072,N_10887,N_10899);
xnor U11073 (N_11073,N_10817,N_10865);
or U11074 (N_11074,N_10807,N_10913);
xor U11075 (N_11075,N_10946,N_10909);
xnor U11076 (N_11076,N_10877,N_10903);
nor U11077 (N_11077,N_10835,N_10873);
and U11078 (N_11078,N_10860,N_10834);
xor U11079 (N_11079,N_10902,N_10883);
and U11080 (N_11080,N_10916,N_10941);
nor U11081 (N_11081,N_10869,N_10926);
or U11082 (N_11082,N_10873,N_10832);
and U11083 (N_11083,N_10931,N_10871);
xor U11084 (N_11084,N_10880,N_10887);
nor U11085 (N_11085,N_10837,N_10826);
nor U11086 (N_11086,N_10916,N_10929);
nor U11087 (N_11087,N_10888,N_10916);
or U11088 (N_11088,N_10911,N_10817);
xnor U11089 (N_11089,N_10932,N_10880);
nand U11090 (N_11090,N_10835,N_10862);
nand U11091 (N_11091,N_10814,N_10827);
xnor U11092 (N_11092,N_10891,N_10830);
nand U11093 (N_11093,N_10851,N_10807);
xnor U11094 (N_11094,N_10928,N_10911);
and U11095 (N_11095,N_10856,N_10822);
xnor U11096 (N_11096,N_10870,N_10876);
xnor U11097 (N_11097,N_10854,N_10905);
and U11098 (N_11098,N_10801,N_10853);
nand U11099 (N_11099,N_10922,N_10904);
or U11100 (N_11100,N_10983,N_10955);
nand U11101 (N_11101,N_11034,N_10962);
xor U11102 (N_11102,N_11085,N_10956);
or U11103 (N_11103,N_10957,N_11020);
nand U11104 (N_11104,N_11006,N_11081);
nand U11105 (N_11105,N_11086,N_10967);
and U11106 (N_11106,N_10976,N_11056);
and U11107 (N_11107,N_11050,N_11030);
or U11108 (N_11108,N_10980,N_11018);
nor U11109 (N_11109,N_10959,N_11047);
nand U11110 (N_11110,N_10981,N_11026);
nand U11111 (N_11111,N_11094,N_10993);
xor U11112 (N_11112,N_11053,N_11046);
or U11113 (N_11113,N_10968,N_11075);
nand U11114 (N_11114,N_11015,N_11093);
xor U11115 (N_11115,N_10974,N_11038);
nand U11116 (N_11116,N_11091,N_10953);
and U11117 (N_11117,N_11089,N_11005);
and U11118 (N_11118,N_11042,N_11088);
and U11119 (N_11119,N_10982,N_11077);
nand U11120 (N_11120,N_10987,N_10973);
and U11121 (N_11121,N_11004,N_11052);
xor U11122 (N_11122,N_11079,N_10994);
and U11123 (N_11123,N_11048,N_10995);
and U11124 (N_11124,N_11043,N_11074);
or U11125 (N_11125,N_11014,N_11098);
nor U11126 (N_11126,N_10965,N_11033);
and U11127 (N_11127,N_11076,N_10966);
nor U11128 (N_11128,N_11008,N_11012);
xnor U11129 (N_11129,N_11057,N_11040);
nand U11130 (N_11130,N_11044,N_11065);
or U11131 (N_11131,N_11095,N_11060);
nand U11132 (N_11132,N_11009,N_11083);
nand U11133 (N_11133,N_10969,N_11017);
or U11134 (N_11134,N_11037,N_11025);
or U11135 (N_11135,N_11059,N_10997);
xor U11136 (N_11136,N_11041,N_10963);
xor U11137 (N_11137,N_11064,N_11031);
nand U11138 (N_11138,N_11067,N_11063);
nor U11139 (N_11139,N_11003,N_11013);
or U11140 (N_11140,N_11035,N_11019);
or U11141 (N_11141,N_10986,N_11016);
nand U11142 (N_11142,N_11082,N_10964);
or U11143 (N_11143,N_10985,N_10961);
nand U11144 (N_11144,N_11027,N_11080);
and U11145 (N_11145,N_10954,N_11087);
and U11146 (N_11146,N_11072,N_11061);
nand U11147 (N_11147,N_10958,N_11010);
or U11148 (N_11148,N_10998,N_11049);
and U11149 (N_11149,N_11023,N_11051);
xnor U11150 (N_11150,N_11007,N_10990);
xor U11151 (N_11151,N_11028,N_11099);
nor U11152 (N_11152,N_10951,N_11036);
xnor U11153 (N_11153,N_10972,N_11021);
or U11154 (N_11154,N_11032,N_11000);
nand U11155 (N_11155,N_11055,N_10996);
xnor U11156 (N_11156,N_10971,N_10991);
or U11157 (N_11157,N_11039,N_11071);
nand U11158 (N_11158,N_10984,N_10979);
and U11159 (N_11159,N_10988,N_11070);
or U11160 (N_11160,N_11078,N_11022);
and U11161 (N_11161,N_11024,N_11029);
and U11162 (N_11162,N_10952,N_11073);
and U11163 (N_11163,N_11096,N_11066);
and U11164 (N_11164,N_11054,N_11011);
nand U11165 (N_11165,N_11058,N_10989);
and U11166 (N_11166,N_11062,N_10999);
and U11167 (N_11167,N_10977,N_11090);
xor U11168 (N_11168,N_10975,N_10950);
or U11169 (N_11169,N_10978,N_11097);
or U11170 (N_11170,N_10970,N_11068);
xnor U11171 (N_11171,N_11092,N_11001);
and U11172 (N_11172,N_11045,N_11002);
nor U11173 (N_11173,N_10992,N_11084);
xnor U11174 (N_11174,N_10960,N_11069);
and U11175 (N_11175,N_11050,N_11044);
nor U11176 (N_11176,N_10974,N_10969);
nand U11177 (N_11177,N_11091,N_11009);
nand U11178 (N_11178,N_10967,N_11044);
and U11179 (N_11179,N_10966,N_11049);
and U11180 (N_11180,N_10955,N_10956);
nor U11181 (N_11181,N_11070,N_10960);
and U11182 (N_11182,N_11095,N_11087);
nand U11183 (N_11183,N_11089,N_11024);
or U11184 (N_11184,N_10963,N_11000);
and U11185 (N_11185,N_11044,N_11064);
nor U11186 (N_11186,N_11003,N_11058);
or U11187 (N_11187,N_11078,N_11013);
or U11188 (N_11188,N_10989,N_10991);
nand U11189 (N_11189,N_11074,N_11099);
nand U11190 (N_11190,N_10986,N_11037);
or U11191 (N_11191,N_11023,N_11030);
nand U11192 (N_11192,N_11001,N_11018);
xor U11193 (N_11193,N_11049,N_10978);
and U11194 (N_11194,N_10959,N_11099);
nor U11195 (N_11195,N_11016,N_10974);
xnor U11196 (N_11196,N_10987,N_11054);
nor U11197 (N_11197,N_10964,N_11071);
nand U11198 (N_11198,N_10980,N_11097);
nor U11199 (N_11199,N_11062,N_10998);
nand U11200 (N_11200,N_11036,N_11086);
xnor U11201 (N_11201,N_11097,N_10966);
nor U11202 (N_11202,N_11075,N_10951);
and U11203 (N_11203,N_11039,N_11038);
xnor U11204 (N_11204,N_11077,N_11031);
xor U11205 (N_11205,N_11044,N_11048);
nand U11206 (N_11206,N_11005,N_11093);
xor U11207 (N_11207,N_11002,N_11043);
nand U11208 (N_11208,N_11081,N_11010);
nor U11209 (N_11209,N_11043,N_11065);
and U11210 (N_11210,N_11011,N_10982);
and U11211 (N_11211,N_11065,N_10957);
xnor U11212 (N_11212,N_11002,N_11023);
and U11213 (N_11213,N_11092,N_10975);
and U11214 (N_11214,N_11052,N_11073);
nor U11215 (N_11215,N_11086,N_11016);
and U11216 (N_11216,N_10955,N_11097);
nor U11217 (N_11217,N_11092,N_11047);
xnor U11218 (N_11218,N_11093,N_11046);
and U11219 (N_11219,N_11082,N_11036);
nor U11220 (N_11220,N_11032,N_10984);
xnor U11221 (N_11221,N_11029,N_11019);
xor U11222 (N_11222,N_10971,N_10984);
and U11223 (N_11223,N_11071,N_11036);
nand U11224 (N_11224,N_11090,N_11004);
or U11225 (N_11225,N_11021,N_11009);
xnor U11226 (N_11226,N_11097,N_11073);
or U11227 (N_11227,N_10981,N_10955);
or U11228 (N_11228,N_11017,N_10989);
xor U11229 (N_11229,N_10976,N_11001);
nor U11230 (N_11230,N_10977,N_11076);
nor U11231 (N_11231,N_11011,N_11006);
and U11232 (N_11232,N_11029,N_11041);
nor U11233 (N_11233,N_10951,N_11017);
and U11234 (N_11234,N_11023,N_11014);
xnor U11235 (N_11235,N_10988,N_11061);
or U11236 (N_11236,N_11034,N_10997);
xnor U11237 (N_11237,N_10969,N_11022);
and U11238 (N_11238,N_10966,N_11041);
nand U11239 (N_11239,N_11086,N_10955);
xor U11240 (N_11240,N_11088,N_11005);
nand U11241 (N_11241,N_11079,N_10950);
nand U11242 (N_11242,N_10975,N_10959);
nor U11243 (N_11243,N_11045,N_11068);
nor U11244 (N_11244,N_11001,N_11088);
nand U11245 (N_11245,N_11009,N_11092);
nand U11246 (N_11246,N_10957,N_11048);
xor U11247 (N_11247,N_11038,N_11095);
and U11248 (N_11248,N_11014,N_10986);
nand U11249 (N_11249,N_10981,N_11043);
nor U11250 (N_11250,N_11120,N_11248);
and U11251 (N_11251,N_11205,N_11113);
and U11252 (N_11252,N_11139,N_11148);
and U11253 (N_11253,N_11202,N_11129);
and U11254 (N_11254,N_11221,N_11117);
nor U11255 (N_11255,N_11230,N_11106);
xnor U11256 (N_11256,N_11153,N_11211);
or U11257 (N_11257,N_11147,N_11224);
xnor U11258 (N_11258,N_11125,N_11116);
nand U11259 (N_11259,N_11157,N_11130);
nor U11260 (N_11260,N_11235,N_11183);
nand U11261 (N_11261,N_11169,N_11100);
or U11262 (N_11262,N_11174,N_11239);
or U11263 (N_11263,N_11191,N_11241);
or U11264 (N_11264,N_11222,N_11114);
nor U11265 (N_11265,N_11236,N_11231);
or U11266 (N_11266,N_11180,N_11170);
nand U11267 (N_11267,N_11247,N_11154);
nor U11268 (N_11268,N_11243,N_11182);
nor U11269 (N_11269,N_11109,N_11223);
or U11270 (N_11270,N_11214,N_11245);
xor U11271 (N_11271,N_11225,N_11187);
and U11272 (N_11272,N_11168,N_11244);
xor U11273 (N_11273,N_11212,N_11156);
or U11274 (N_11274,N_11162,N_11132);
nor U11275 (N_11275,N_11232,N_11186);
nand U11276 (N_11276,N_11220,N_11146);
nor U11277 (N_11277,N_11201,N_11194);
xnor U11278 (N_11278,N_11200,N_11215);
or U11279 (N_11279,N_11122,N_11138);
nor U11280 (N_11280,N_11192,N_11181);
xor U11281 (N_11281,N_11103,N_11121);
nand U11282 (N_11282,N_11137,N_11203);
nand U11283 (N_11283,N_11115,N_11133);
nand U11284 (N_11284,N_11119,N_11190);
nor U11285 (N_11285,N_11185,N_11179);
and U11286 (N_11286,N_11164,N_11126);
xor U11287 (N_11287,N_11166,N_11124);
or U11288 (N_11288,N_11172,N_11135);
and U11289 (N_11289,N_11237,N_11177);
nand U11290 (N_11290,N_11158,N_11151);
and U11291 (N_11291,N_11150,N_11219);
or U11292 (N_11292,N_11217,N_11112);
nor U11293 (N_11293,N_11165,N_11141);
or U11294 (N_11294,N_11171,N_11188);
nor U11295 (N_11295,N_11197,N_11173);
and U11296 (N_11296,N_11195,N_11227);
nor U11297 (N_11297,N_11175,N_11210);
nand U11298 (N_11298,N_11184,N_11206);
xor U11299 (N_11299,N_11143,N_11216);
nand U11300 (N_11300,N_11149,N_11128);
nand U11301 (N_11301,N_11213,N_11198);
xor U11302 (N_11302,N_11140,N_11226);
nor U11303 (N_11303,N_11196,N_11207);
nand U11304 (N_11304,N_11167,N_11240);
or U11305 (N_11305,N_11218,N_11107);
nand U11306 (N_11306,N_11118,N_11228);
xnor U11307 (N_11307,N_11136,N_11189);
nor U11308 (N_11308,N_11127,N_11159);
xnor U11309 (N_11309,N_11199,N_11155);
nor U11310 (N_11310,N_11142,N_11204);
nor U11311 (N_11311,N_11176,N_11229);
or U11312 (N_11312,N_11145,N_11108);
nand U11313 (N_11313,N_11110,N_11160);
nor U11314 (N_11314,N_11242,N_11193);
nand U11315 (N_11315,N_11161,N_11111);
nand U11316 (N_11316,N_11131,N_11144);
or U11317 (N_11317,N_11102,N_11238);
nand U11318 (N_11318,N_11163,N_11208);
or U11319 (N_11319,N_11249,N_11105);
xnor U11320 (N_11320,N_11246,N_11178);
and U11321 (N_11321,N_11152,N_11209);
nand U11322 (N_11322,N_11134,N_11104);
and U11323 (N_11323,N_11234,N_11233);
and U11324 (N_11324,N_11123,N_11101);
xnor U11325 (N_11325,N_11213,N_11108);
or U11326 (N_11326,N_11123,N_11161);
and U11327 (N_11327,N_11227,N_11161);
and U11328 (N_11328,N_11181,N_11221);
nor U11329 (N_11329,N_11210,N_11216);
nand U11330 (N_11330,N_11178,N_11172);
and U11331 (N_11331,N_11183,N_11234);
xor U11332 (N_11332,N_11172,N_11243);
xnor U11333 (N_11333,N_11106,N_11147);
xnor U11334 (N_11334,N_11164,N_11130);
xnor U11335 (N_11335,N_11196,N_11212);
xor U11336 (N_11336,N_11127,N_11229);
and U11337 (N_11337,N_11160,N_11132);
or U11338 (N_11338,N_11160,N_11148);
nand U11339 (N_11339,N_11168,N_11210);
and U11340 (N_11340,N_11229,N_11214);
xor U11341 (N_11341,N_11140,N_11129);
xnor U11342 (N_11342,N_11249,N_11129);
and U11343 (N_11343,N_11240,N_11160);
and U11344 (N_11344,N_11234,N_11176);
xor U11345 (N_11345,N_11178,N_11130);
or U11346 (N_11346,N_11208,N_11168);
nor U11347 (N_11347,N_11116,N_11197);
or U11348 (N_11348,N_11107,N_11207);
or U11349 (N_11349,N_11139,N_11215);
or U11350 (N_11350,N_11101,N_11199);
or U11351 (N_11351,N_11249,N_11179);
or U11352 (N_11352,N_11180,N_11125);
and U11353 (N_11353,N_11236,N_11239);
or U11354 (N_11354,N_11206,N_11231);
and U11355 (N_11355,N_11131,N_11220);
xor U11356 (N_11356,N_11190,N_11174);
xor U11357 (N_11357,N_11152,N_11173);
nor U11358 (N_11358,N_11243,N_11219);
xnor U11359 (N_11359,N_11190,N_11155);
and U11360 (N_11360,N_11187,N_11211);
xnor U11361 (N_11361,N_11128,N_11162);
or U11362 (N_11362,N_11170,N_11130);
xor U11363 (N_11363,N_11234,N_11196);
and U11364 (N_11364,N_11163,N_11193);
nand U11365 (N_11365,N_11105,N_11151);
or U11366 (N_11366,N_11220,N_11218);
or U11367 (N_11367,N_11137,N_11181);
nand U11368 (N_11368,N_11245,N_11117);
or U11369 (N_11369,N_11236,N_11121);
nand U11370 (N_11370,N_11154,N_11225);
and U11371 (N_11371,N_11191,N_11121);
or U11372 (N_11372,N_11158,N_11204);
nand U11373 (N_11373,N_11224,N_11110);
and U11374 (N_11374,N_11213,N_11229);
or U11375 (N_11375,N_11151,N_11223);
nand U11376 (N_11376,N_11134,N_11230);
nor U11377 (N_11377,N_11101,N_11214);
and U11378 (N_11378,N_11109,N_11231);
and U11379 (N_11379,N_11119,N_11225);
nor U11380 (N_11380,N_11171,N_11143);
nand U11381 (N_11381,N_11184,N_11118);
xnor U11382 (N_11382,N_11199,N_11224);
nand U11383 (N_11383,N_11118,N_11146);
nand U11384 (N_11384,N_11249,N_11175);
or U11385 (N_11385,N_11152,N_11174);
xnor U11386 (N_11386,N_11148,N_11246);
or U11387 (N_11387,N_11188,N_11144);
and U11388 (N_11388,N_11222,N_11146);
nand U11389 (N_11389,N_11111,N_11128);
xor U11390 (N_11390,N_11172,N_11125);
nand U11391 (N_11391,N_11169,N_11109);
xnor U11392 (N_11392,N_11116,N_11207);
nor U11393 (N_11393,N_11134,N_11232);
nand U11394 (N_11394,N_11236,N_11104);
nand U11395 (N_11395,N_11113,N_11163);
nand U11396 (N_11396,N_11200,N_11111);
or U11397 (N_11397,N_11249,N_11214);
and U11398 (N_11398,N_11137,N_11132);
xnor U11399 (N_11399,N_11184,N_11120);
nand U11400 (N_11400,N_11370,N_11291);
nand U11401 (N_11401,N_11361,N_11376);
nand U11402 (N_11402,N_11336,N_11290);
and U11403 (N_11403,N_11334,N_11345);
nand U11404 (N_11404,N_11295,N_11342);
or U11405 (N_11405,N_11297,N_11276);
and U11406 (N_11406,N_11310,N_11364);
xor U11407 (N_11407,N_11374,N_11317);
nand U11408 (N_11408,N_11287,N_11350);
or U11409 (N_11409,N_11251,N_11395);
xor U11410 (N_11410,N_11316,N_11378);
and U11411 (N_11411,N_11371,N_11301);
xor U11412 (N_11412,N_11286,N_11302);
nand U11413 (N_11413,N_11323,N_11326);
nand U11414 (N_11414,N_11289,N_11377);
or U11415 (N_11415,N_11389,N_11259);
xnor U11416 (N_11416,N_11281,N_11320);
or U11417 (N_11417,N_11380,N_11294);
nand U11418 (N_11418,N_11348,N_11292);
xor U11419 (N_11419,N_11340,N_11325);
nand U11420 (N_11420,N_11365,N_11314);
xnor U11421 (N_11421,N_11390,N_11283);
xnor U11422 (N_11422,N_11381,N_11332);
or U11423 (N_11423,N_11265,N_11330);
or U11424 (N_11424,N_11299,N_11321);
xnor U11425 (N_11425,N_11254,N_11344);
and U11426 (N_11426,N_11267,N_11360);
xnor U11427 (N_11427,N_11309,N_11272);
and U11428 (N_11428,N_11252,N_11382);
or U11429 (N_11429,N_11392,N_11278);
nand U11430 (N_11430,N_11358,N_11372);
nor U11431 (N_11431,N_11319,N_11305);
and U11432 (N_11432,N_11341,N_11356);
xor U11433 (N_11433,N_11352,N_11394);
xnor U11434 (N_11434,N_11386,N_11318);
and U11435 (N_11435,N_11293,N_11300);
or U11436 (N_11436,N_11282,N_11355);
or U11437 (N_11437,N_11346,N_11391);
nor U11438 (N_11438,N_11328,N_11284);
or U11439 (N_11439,N_11397,N_11322);
or U11440 (N_11440,N_11343,N_11357);
xnor U11441 (N_11441,N_11262,N_11312);
or U11442 (N_11442,N_11315,N_11275);
nand U11443 (N_11443,N_11393,N_11264);
nand U11444 (N_11444,N_11363,N_11384);
nand U11445 (N_11445,N_11270,N_11269);
and U11446 (N_11446,N_11387,N_11338);
nand U11447 (N_11447,N_11308,N_11383);
and U11448 (N_11448,N_11367,N_11324);
xor U11449 (N_11449,N_11398,N_11396);
nand U11450 (N_11450,N_11273,N_11351);
nor U11451 (N_11451,N_11311,N_11253);
or U11452 (N_11452,N_11327,N_11304);
or U11453 (N_11453,N_11277,N_11388);
and U11454 (N_11454,N_11288,N_11353);
nor U11455 (N_11455,N_11373,N_11255);
nor U11456 (N_11456,N_11257,N_11359);
xor U11457 (N_11457,N_11271,N_11366);
and U11458 (N_11458,N_11280,N_11306);
xor U11459 (N_11459,N_11260,N_11335);
nand U11460 (N_11460,N_11331,N_11399);
xor U11461 (N_11461,N_11274,N_11258);
and U11462 (N_11462,N_11354,N_11368);
nand U11463 (N_11463,N_11337,N_11261);
nor U11464 (N_11464,N_11298,N_11339);
xnor U11465 (N_11465,N_11266,N_11303);
xnor U11466 (N_11466,N_11385,N_11279);
or U11467 (N_11467,N_11268,N_11347);
and U11468 (N_11468,N_11296,N_11349);
and U11469 (N_11469,N_11313,N_11329);
nor U11470 (N_11470,N_11263,N_11369);
nor U11471 (N_11471,N_11362,N_11256);
nor U11472 (N_11472,N_11379,N_11307);
nor U11473 (N_11473,N_11285,N_11375);
xnor U11474 (N_11474,N_11333,N_11250);
nand U11475 (N_11475,N_11366,N_11281);
nor U11476 (N_11476,N_11361,N_11394);
or U11477 (N_11477,N_11349,N_11358);
nor U11478 (N_11478,N_11344,N_11276);
and U11479 (N_11479,N_11367,N_11277);
or U11480 (N_11480,N_11361,N_11284);
nand U11481 (N_11481,N_11282,N_11324);
or U11482 (N_11482,N_11335,N_11390);
xor U11483 (N_11483,N_11395,N_11322);
and U11484 (N_11484,N_11311,N_11270);
and U11485 (N_11485,N_11310,N_11383);
and U11486 (N_11486,N_11349,N_11283);
or U11487 (N_11487,N_11386,N_11349);
nor U11488 (N_11488,N_11363,N_11311);
xor U11489 (N_11489,N_11324,N_11365);
or U11490 (N_11490,N_11257,N_11322);
and U11491 (N_11491,N_11385,N_11393);
xor U11492 (N_11492,N_11374,N_11272);
or U11493 (N_11493,N_11288,N_11370);
xnor U11494 (N_11494,N_11338,N_11290);
nor U11495 (N_11495,N_11255,N_11383);
and U11496 (N_11496,N_11254,N_11357);
nand U11497 (N_11497,N_11328,N_11281);
xor U11498 (N_11498,N_11364,N_11284);
and U11499 (N_11499,N_11378,N_11376);
or U11500 (N_11500,N_11310,N_11373);
and U11501 (N_11501,N_11279,N_11397);
nand U11502 (N_11502,N_11382,N_11302);
or U11503 (N_11503,N_11304,N_11369);
nor U11504 (N_11504,N_11285,N_11388);
or U11505 (N_11505,N_11319,N_11392);
and U11506 (N_11506,N_11288,N_11359);
nor U11507 (N_11507,N_11352,N_11319);
or U11508 (N_11508,N_11306,N_11370);
and U11509 (N_11509,N_11274,N_11396);
xor U11510 (N_11510,N_11387,N_11395);
nand U11511 (N_11511,N_11398,N_11312);
nand U11512 (N_11512,N_11391,N_11388);
nor U11513 (N_11513,N_11389,N_11300);
xor U11514 (N_11514,N_11325,N_11287);
nand U11515 (N_11515,N_11347,N_11307);
or U11516 (N_11516,N_11304,N_11389);
and U11517 (N_11517,N_11339,N_11340);
or U11518 (N_11518,N_11250,N_11257);
and U11519 (N_11519,N_11370,N_11332);
xnor U11520 (N_11520,N_11323,N_11385);
nor U11521 (N_11521,N_11310,N_11338);
or U11522 (N_11522,N_11327,N_11331);
xor U11523 (N_11523,N_11313,N_11331);
nor U11524 (N_11524,N_11397,N_11324);
and U11525 (N_11525,N_11346,N_11310);
and U11526 (N_11526,N_11335,N_11333);
or U11527 (N_11527,N_11376,N_11349);
or U11528 (N_11528,N_11281,N_11369);
nor U11529 (N_11529,N_11354,N_11376);
nand U11530 (N_11530,N_11290,N_11334);
or U11531 (N_11531,N_11368,N_11266);
xor U11532 (N_11532,N_11379,N_11370);
or U11533 (N_11533,N_11354,N_11345);
xor U11534 (N_11534,N_11270,N_11377);
or U11535 (N_11535,N_11334,N_11327);
or U11536 (N_11536,N_11307,N_11343);
xor U11537 (N_11537,N_11255,N_11345);
xor U11538 (N_11538,N_11344,N_11391);
or U11539 (N_11539,N_11305,N_11290);
nor U11540 (N_11540,N_11271,N_11313);
nand U11541 (N_11541,N_11385,N_11254);
and U11542 (N_11542,N_11295,N_11380);
or U11543 (N_11543,N_11368,N_11373);
or U11544 (N_11544,N_11354,N_11398);
xnor U11545 (N_11545,N_11294,N_11259);
xnor U11546 (N_11546,N_11293,N_11290);
nor U11547 (N_11547,N_11364,N_11256);
xnor U11548 (N_11548,N_11360,N_11378);
nand U11549 (N_11549,N_11332,N_11268);
xnor U11550 (N_11550,N_11458,N_11538);
xnor U11551 (N_11551,N_11422,N_11514);
nand U11552 (N_11552,N_11469,N_11532);
nand U11553 (N_11553,N_11445,N_11461);
or U11554 (N_11554,N_11515,N_11417);
and U11555 (N_11555,N_11456,N_11475);
xor U11556 (N_11556,N_11471,N_11472);
nand U11557 (N_11557,N_11503,N_11527);
xor U11558 (N_11558,N_11541,N_11505);
nand U11559 (N_11559,N_11473,N_11440);
and U11560 (N_11560,N_11502,N_11518);
or U11561 (N_11561,N_11483,N_11513);
xnor U11562 (N_11562,N_11526,N_11433);
and U11563 (N_11563,N_11412,N_11431);
and U11564 (N_11564,N_11492,N_11524);
and U11565 (N_11565,N_11481,N_11428);
nand U11566 (N_11566,N_11419,N_11522);
nor U11567 (N_11567,N_11537,N_11521);
xnor U11568 (N_11568,N_11465,N_11546);
xor U11569 (N_11569,N_11528,N_11457);
xor U11570 (N_11570,N_11511,N_11549);
nor U11571 (N_11571,N_11426,N_11420);
nor U11572 (N_11572,N_11544,N_11407);
nand U11573 (N_11573,N_11485,N_11450);
and U11574 (N_11574,N_11452,N_11447);
xnor U11575 (N_11575,N_11493,N_11400);
nor U11576 (N_11576,N_11487,N_11545);
or U11577 (N_11577,N_11454,N_11506);
nor U11578 (N_11578,N_11548,N_11476);
nor U11579 (N_11579,N_11509,N_11491);
and U11580 (N_11580,N_11468,N_11444);
nor U11581 (N_11581,N_11543,N_11455);
and U11582 (N_11582,N_11496,N_11427);
nand U11583 (N_11583,N_11448,N_11429);
or U11584 (N_11584,N_11401,N_11520);
nor U11585 (N_11585,N_11478,N_11414);
xor U11586 (N_11586,N_11434,N_11453);
nor U11587 (N_11587,N_11500,N_11531);
nand U11588 (N_11588,N_11542,N_11406);
or U11589 (N_11589,N_11463,N_11533);
or U11590 (N_11590,N_11470,N_11512);
or U11591 (N_11591,N_11446,N_11442);
nand U11592 (N_11592,N_11415,N_11529);
nand U11593 (N_11593,N_11494,N_11525);
or U11594 (N_11594,N_11467,N_11411);
and U11595 (N_11595,N_11477,N_11466);
and U11596 (N_11596,N_11439,N_11449);
xor U11597 (N_11597,N_11443,N_11504);
nand U11598 (N_11598,N_11482,N_11402);
or U11599 (N_11599,N_11418,N_11408);
or U11600 (N_11600,N_11425,N_11480);
xnor U11601 (N_11601,N_11519,N_11409);
and U11602 (N_11602,N_11510,N_11437);
nand U11603 (N_11603,N_11436,N_11438);
nor U11604 (N_11604,N_11416,N_11495);
nor U11605 (N_11605,N_11507,N_11535);
nand U11606 (N_11606,N_11486,N_11462);
or U11607 (N_11607,N_11451,N_11404);
xor U11608 (N_11608,N_11523,N_11464);
or U11609 (N_11609,N_11489,N_11474);
nor U11610 (N_11610,N_11499,N_11435);
nor U11611 (N_11611,N_11424,N_11497);
xnor U11612 (N_11612,N_11536,N_11430);
xor U11613 (N_11613,N_11530,N_11413);
and U11614 (N_11614,N_11421,N_11441);
nor U11615 (N_11615,N_11540,N_11410);
nand U11616 (N_11616,N_11539,N_11490);
or U11617 (N_11617,N_11479,N_11508);
xnor U11618 (N_11618,N_11516,N_11547);
xnor U11619 (N_11619,N_11423,N_11459);
and U11620 (N_11620,N_11403,N_11484);
xnor U11621 (N_11621,N_11432,N_11498);
xor U11622 (N_11622,N_11405,N_11517);
nor U11623 (N_11623,N_11488,N_11501);
nor U11624 (N_11624,N_11534,N_11460);
xnor U11625 (N_11625,N_11504,N_11406);
or U11626 (N_11626,N_11515,N_11470);
and U11627 (N_11627,N_11521,N_11512);
xnor U11628 (N_11628,N_11423,N_11519);
and U11629 (N_11629,N_11433,N_11469);
nor U11630 (N_11630,N_11494,N_11503);
or U11631 (N_11631,N_11502,N_11436);
nor U11632 (N_11632,N_11531,N_11408);
nor U11633 (N_11633,N_11436,N_11513);
xnor U11634 (N_11634,N_11462,N_11517);
or U11635 (N_11635,N_11446,N_11403);
or U11636 (N_11636,N_11424,N_11514);
xor U11637 (N_11637,N_11494,N_11505);
nand U11638 (N_11638,N_11426,N_11471);
xnor U11639 (N_11639,N_11469,N_11528);
nor U11640 (N_11640,N_11478,N_11460);
nor U11641 (N_11641,N_11527,N_11487);
and U11642 (N_11642,N_11439,N_11471);
and U11643 (N_11643,N_11453,N_11467);
or U11644 (N_11644,N_11421,N_11487);
xor U11645 (N_11645,N_11523,N_11531);
nor U11646 (N_11646,N_11549,N_11531);
or U11647 (N_11647,N_11531,N_11489);
or U11648 (N_11648,N_11515,N_11467);
nor U11649 (N_11649,N_11426,N_11430);
nor U11650 (N_11650,N_11440,N_11490);
and U11651 (N_11651,N_11415,N_11469);
or U11652 (N_11652,N_11542,N_11521);
and U11653 (N_11653,N_11489,N_11490);
or U11654 (N_11654,N_11526,N_11534);
or U11655 (N_11655,N_11481,N_11464);
xor U11656 (N_11656,N_11502,N_11453);
nor U11657 (N_11657,N_11473,N_11415);
nand U11658 (N_11658,N_11418,N_11412);
nand U11659 (N_11659,N_11549,N_11538);
or U11660 (N_11660,N_11506,N_11466);
xor U11661 (N_11661,N_11408,N_11433);
or U11662 (N_11662,N_11446,N_11494);
and U11663 (N_11663,N_11476,N_11483);
and U11664 (N_11664,N_11505,N_11468);
and U11665 (N_11665,N_11430,N_11439);
nand U11666 (N_11666,N_11545,N_11522);
or U11667 (N_11667,N_11441,N_11487);
nor U11668 (N_11668,N_11497,N_11433);
or U11669 (N_11669,N_11444,N_11483);
or U11670 (N_11670,N_11514,N_11535);
nor U11671 (N_11671,N_11529,N_11541);
and U11672 (N_11672,N_11492,N_11466);
or U11673 (N_11673,N_11524,N_11463);
and U11674 (N_11674,N_11471,N_11450);
and U11675 (N_11675,N_11548,N_11479);
nand U11676 (N_11676,N_11502,N_11486);
nor U11677 (N_11677,N_11461,N_11528);
nand U11678 (N_11678,N_11524,N_11526);
nor U11679 (N_11679,N_11410,N_11519);
xnor U11680 (N_11680,N_11531,N_11540);
and U11681 (N_11681,N_11498,N_11513);
nor U11682 (N_11682,N_11448,N_11432);
or U11683 (N_11683,N_11418,N_11532);
nor U11684 (N_11684,N_11425,N_11415);
and U11685 (N_11685,N_11467,N_11435);
and U11686 (N_11686,N_11498,N_11473);
xnor U11687 (N_11687,N_11501,N_11518);
or U11688 (N_11688,N_11482,N_11491);
or U11689 (N_11689,N_11520,N_11405);
nand U11690 (N_11690,N_11442,N_11436);
or U11691 (N_11691,N_11540,N_11421);
and U11692 (N_11692,N_11509,N_11546);
nor U11693 (N_11693,N_11524,N_11493);
and U11694 (N_11694,N_11439,N_11410);
nor U11695 (N_11695,N_11458,N_11546);
xnor U11696 (N_11696,N_11511,N_11519);
nor U11697 (N_11697,N_11432,N_11411);
nand U11698 (N_11698,N_11536,N_11427);
nor U11699 (N_11699,N_11415,N_11517);
and U11700 (N_11700,N_11627,N_11590);
xnor U11701 (N_11701,N_11586,N_11670);
or U11702 (N_11702,N_11633,N_11622);
nor U11703 (N_11703,N_11634,N_11550);
nand U11704 (N_11704,N_11635,N_11688);
and U11705 (N_11705,N_11675,N_11566);
nor U11706 (N_11706,N_11589,N_11674);
nand U11707 (N_11707,N_11624,N_11564);
nor U11708 (N_11708,N_11642,N_11603);
and U11709 (N_11709,N_11698,N_11684);
or U11710 (N_11710,N_11647,N_11613);
nor U11711 (N_11711,N_11690,N_11626);
nor U11712 (N_11712,N_11637,N_11617);
and U11713 (N_11713,N_11672,N_11598);
nor U11714 (N_11714,N_11681,N_11588);
nand U11715 (N_11715,N_11665,N_11680);
nand U11716 (N_11716,N_11677,N_11685);
nand U11717 (N_11717,N_11560,N_11636);
and U11718 (N_11718,N_11577,N_11629);
nor U11719 (N_11719,N_11563,N_11667);
and U11720 (N_11720,N_11559,N_11628);
or U11721 (N_11721,N_11692,N_11610);
or U11722 (N_11722,N_11668,N_11679);
or U11723 (N_11723,N_11600,N_11657);
and U11724 (N_11724,N_11693,N_11609);
or U11725 (N_11725,N_11659,N_11654);
and U11726 (N_11726,N_11691,N_11561);
or U11727 (N_11727,N_11594,N_11611);
nand U11728 (N_11728,N_11619,N_11655);
or U11729 (N_11729,N_11696,N_11663);
nor U11730 (N_11730,N_11614,N_11662);
nand U11731 (N_11731,N_11576,N_11682);
nand U11732 (N_11732,N_11631,N_11595);
nand U11733 (N_11733,N_11656,N_11699);
or U11734 (N_11734,N_11676,N_11557);
nand U11735 (N_11735,N_11565,N_11646);
nand U11736 (N_11736,N_11695,N_11621);
and U11737 (N_11737,N_11582,N_11669);
and U11738 (N_11738,N_11570,N_11607);
and U11739 (N_11739,N_11650,N_11639);
or U11740 (N_11740,N_11605,N_11556);
and U11741 (N_11741,N_11683,N_11583);
nand U11742 (N_11742,N_11587,N_11606);
xor U11743 (N_11743,N_11567,N_11579);
nor U11744 (N_11744,N_11616,N_11553);
nor U11745 (N_11745,N_11604,N_11552);
and U11746 (N_11746,N_11568,N_11578);
and U11747 (N_11747,N_11671,N_11593);
or U11748 (N_11748,N_11569,N_11643);
or U11749 (N_11749,N_11649,N_11638);
nand U11750 (N_11750,N_11697,N_11630);
nor U11751 (N_11751,N_11664,N_11584);
nand U11752 (N_11752,N_11660,N_11585);
nor U11753 (N_11753,N_11623,N_11571);
nand U11754 (N_11754,N_11689,N_11572);
nand U11755 (N_11755,N_11661,N_11615);
or U11756 (N_11756,N_11580,N_11562);
or U11757 (N_11757,N_11651,N_11653);
and U11758 (N_11758,N_11555,N_11599);
nand U11759 (N_11759,N_11645,N_11694);
or U11760 (N_11760,N_11592,N_11602);
xnor U11761 (N_11761,N_11573,N_11558);
or U11762 (N_11762,N_11612,N_11652);
and U11763 (N_11763,N_11575,N_11554);
or U11764 (N_11764,N_11641,N_11666);
or U11765 (N_11765,N_11591,N_11551);
xnor U11766 (N_11766,N_11673,N_11640);
and U11767 (N_11767,N_11678,N_11686);
nand U11768 (N_11768,N_11658,N_11601);
or U11769 (N_11769,N_11620,N_11574);
nor U11770 (N_11770,N_11625,N_11581);
and U11771 (N_11771,N_11644,N_11687);
nand U11772 (N_11772,N_11618,N_11596);
nor U11773 (N_11773,N_11597,N_11608);
nand U11774 (N_11774,N_11648,N_11632);
nand U11775 (N_11775,N_11696,N_11635);
xor U11776 (N_11776,N_11579,N_11606);
xor U11777 (N_11777,N_11638,N_11660);
xor U11778 (N_11778,N_11572,N_11576);
nor U11779 (N_11779,N_11693,N_11592);
and U11780 (N_11780,N_11623,N_11558);
or U11781 (N_11781,N_11682,N_11554);
nor U11782 (N_11782,N_11675,N_11559);
and U11783 (N_11783,N_11647,N_11674);
and U11784 (N_11784,N_11637,N_11555);
xor U11785 (N_11785,N_11563,N_11565);
nor U11786 (N_11786,N_11685,N_11586);
xor U11787 (N_11787,N_11593,N_11632);
and U11788 (N_11788,N_11679,N_11574);
xnor U11789 (N_11789,N_11633,N_11692);
nand U11790 (N_11790,N_11633,N_11654);
xnor U11791 (N_11791,N_11659,N_11620);
or U11792 (N_11792,N_11562,N_11576);
or U11793 (N_11793,N_11557,N_11652);
xor U11794 (N_11794,N_11649,N_11614);
nor U11795 (N_11795,N_11617,N_11677);
xor U11796 (N_11796,N_11566,N_11565);
nand U11797 (N_11797,N_11636,N_11649);
nand U11798 (N_11798,N_11660,N_11684);
nand U11799 (N_11799,N_11605,N_11689);
xnor U11800 (N_11800,N_11643,N_11634);
nor U11801 (N_11801,N_11569,N_11681);
xor U11802 (N_11802,N_11647,N_11645);
xnor U11803 (N_11803,N_11555,N_11551);
nor U11804 (N_11804,N_11588,N_11631);
or U11805 (N_11805,N_11675,N_11660);
nand U11806 (N_11806,N_11680,N_11639);
or U11807 (N_11807,N_11555,N_11614);
or U11808 (N_11808,N_11696,N_11561);
nand U11809 (N_11809,N_11691,N_11682);
xor U11810 (N_11810,N_11689,N_11556);
or U11811 (N_11811,N_11663,N_11617);
nand U11812 (N_11812,N_11666,N_11661);
nor U11813 (N_11813,N_11690,N_11631);
nand U11814 (N_11814,N_11695,N_11617);
or U11815 (N_11815,N_11571,N_11604);
nor U11816 (N_11816,N_11579,N_11699);
and U11817 (N_11817,N_11614,N_11587);
and U11818 (N_11818,N_11563,N_11623);
nor U11819 (N_11819,N_11635,N_11572);
nor U11820 (N_11820,N_11657,N_11682);
nor U11821 (N_11821,N_11558,N_11684);
or U11822 (N_11822,N_11599,N_11627);
or U11823 (N_11823,N_11668,N_11619);
and U11824 (N_11824,N_11623,N_11629);
nand U11825 (N_11825,N_11670,N_11606);
xnor U11826 (N_11826,N_11586,N_11595);
nor U11827 (N_11827,N_11689,N_11662);
or U11828 (N_11828,N_11602,N_11603);
nand U11829 (N_11829,N_11594,N_11619);
nand U11830 (N_11830,N_11644,N_11688);
xor U11831 (N_11831,N_11551,N_11682);
nand U11832 (N_11832,N_11671,N_11694);
nand U11833 (N_11833,N_11557,N_11686);
xor U11834 (N_11834,N_11602,N_11677);
and U11835 (N_11835,N_11666,N_11588);
nand U11836 (N_11836,N_11561,N_11697);
nand U11837 (N_11837,N_11623,N_11604);
nor U11838 (N_11838,N_11680,N_11648);
or U11839 (N_11839,N_11608,N_11682);
nor U11840 (N_11840,N_11690,N_11596);
xnor U11841 (N_11841,N_11674,N_11572);
nand U11842 (N_11842,N_11573,N_11600);
and U11843 (N_11843,N_11568,N_11657);
nor U11844 (N_11844,N_11613,N_11616);
nor U11845 (N_11845,N_11562,N_11554);
xnor U11846 (N_11846,N_11614,N_11565);
or U11847 (N_11847,N_11603,N_11624);
or U11848 (N_11848,N_11672,N_11620);
nand U11849 (N_11849,N_11631,N_11681);
or U11850 (N_11850,N_11820,N_11756);
or U11851 (N_11851,N_11751,N_11734);
nor U11852 (N_11852,N_11824,N_11719);
and U11853 (N_11853,N_11737,N_11806);
nor U11854 (N_11854,N_11837,N_11723);
nor U11855 (N_11855,N_11742,N_11821);
nand U11856 (N_11856,N_11709,N_11780);
nor U11857 (N_11857,N_11777,N_11741);
or U11858 (N_11858,N_11828,N_11787);
and U11859 (N_11859,N_11794,N_11749);
nand U11860 (N_11860,N_11710,N_11813);
nand U11861 (N_11861,N_11785,N_11778);
or U11862 (N_11862,N_11711,N_11804);
xor U11863 (N_11863,N_11844,N_11760);
nor U11864 (N_11864,N_11816,N_11765);
nand U11865 (N_11865,N_11838,N_11707);
xor U11866 (N_11866,N_11700,N_11758);
xnor U11867 (N_11867,N_11834,N_11729);
and U11868 (N_11868,N_11803,N_11724);
or U11869 (N_11869,N_11846,N_11745);
and U11870 (N_11870,N_11739,N_11818);
xor U11871 (N_11871,N_11790,N_11800);
nor U11872 (N_11872,N_11799,N_11796);
nor U11873 (N_11873,N_11797,N_11746);
or U11874 (N_11874,N_11802,N_11831);
nand U11875 (N_11875,N_11717,N_11716);
or U11876 (N_11876,N_11830,N_11848);
xnor U11877 (N_11877,N_11793,N_11714);
and U11878 (N_11878,N_11731,N_11779);
nand U11879 (N_11879,N_11792,N_11726);
nand U11880 (N_11880,N_11773,N_11732);
xor U11881 (N_11881,N_11704,N_11825);
nand U11882 (N_11882,N_11771,N_11713);
or U11883 (N_11883,N_11706,N_11827);
xnor U11884 (N_11884,N_11715,N_11769);
xor U11885 (N_11885,N_11738,N_11757);
nor U11886 (N_11886,N_11730,N_11767);
or U11887 (N_11887,N_11798,N_11774);
or U11888 (N_11888,N_11708,N_11843);
xor U11889 (N_11889,N_11705,N_11826);
xnor U11890 (N_11890,N_11743,N_11791);
nor U11891 (N_11891,N_11733,N_11776);
nand U11892 (N_11892,N_11781,N_11783);
nor U11893 (N_11893,N_11811,N_11702);
or U11894 (N_11894,N_11809,N_11839);
and U11895 (N_11895,N_11725,N_11750);
xnor U11896 (N_11896,N_11722,N_11807);
or U11897 (N_11897,N_11748,N_11808);
nor U11898 (N_11898,N_11759,N_11836);
and U11899 (N_11899,N_11701,N_11849);
nand U11900 (N_11900,N_11833,N_11766);
nand U11901 (N_11901,N_11728,N_11770);
xnor U11902 (N_11902,N_11829,N_11764);
nor U11903 (N_11903,N_11819,N_11784);
nand U11904 (N_11904,N_11847,N_11795);
or U11905 (N_11905,N_11720,N_11744);
xor U11906 (N_11906,N_11752,N_11740);
and U11907 (N_11907,N_11823,N_11718);
nor U11908 (N_11908,N_11768,N_11727);
nor U11909 (N_11909,N_11840,N_11822);
nor U11910 (N_11910,N_11753,N_11817);
nor U11911 (N_11911,N_11832,N_11763);
nor U11912 (N_11912,N_11761,N_11712);
or U11913 (N_11913,N_11775,N_11835);
nand U11914 (N_11914,N_11788,N_11842);
xnor U11915 (N_11915,N_11845,N_11801);
nand U11916 (N_11916,N_11735,N_11755);
or U11917 (N_11917,N_11736,N_11782);
nor U11918 (N_11918,N_11812,N_11789);
xnor U11919 (N_11919,N_11762,N_11805);
or U11920 (N_11920,N_11815,N_11810);
or U11921 (N_11921,N_11814,N_11841);
and U11922 (N_11922,N_11747,N_11721);
and U11923 (N_11923,N_11786,N_11772);
and U11924 (N_11924,N_11754,N_11703);
xor U11925 (N_11925,N_11706,N_11845);
or U11926 (N_11926,N_11704,N_11831);
or U11927 (N_11927,N_11715,N_11793);
and U11928 (N_11928,N_11809,N_11749);
xor U11929 (N_11929,N_11835,N_11709);
nor U11930 (N_11930,N_11702,N_11706);
nor U11931 (N_11931,N_11849,N_11707);
or U11932 (N_11932,N_11799,N_11711);
nor U11933 (N_11933,N_11794,N_11747);
xor U11934 (N_11934,N_11819,N_11704);
or U11935 (N_11935,N_11799,N_11735);
nand U11936 (N_11936,N_11745,N_11737);
nor U11937 (N_11937,N_11777,N_11733);
and U11938 (N_11938,N_11796,N_11753);
xor U11939 (N_11939,N_11832,N_11810);
or U11940 (N_11940,N_11816,N_11833);
and U11941 (N_11941,N_11839,N_11778);
nand U11942 (N_11942,N_11787,N_11785);
and U11943 (N_11943,N_11805,N_11780);
or U11944 (N_11944,N_11790,N_11836);
and U11945 (N_11945,N_11782,N_11759);
nor U11946 (N_11946,N_11778,N_11825);
or U11947 (N_11947,N_11712,N_11788);
xnor U11948 (N_11948,N_11777,N_11702);
nor U11949 (N_11949,N_11800,N_11717);
and U11950 (N_11950,N_11804,N_11713);
nand U11951 (N_11951,N_11836,N_11823);
xnor U11952 (N_11952,N_11711,N_11732);
nor U11953 (N_11953,N_11835,N_11710);
xor U11954 (N_11954,N_11784,N_11733);
nor U11955 (N_11955,N_11795,N_11776);
and U11956 (N_11956,N_11808,N_11766);
and U11957 (N_11957,N_11730,N_11750);
nor U11958 (N_11958,N_11749,N_11771);
nand U11959 (N_11959,N_11843,N_11768);
nor U11960 (N_11960,N_11787,N_11731);
xor U11961 (N_11961,N_11831,N_11735);
xor U11962 (N_11962,N_11717,N_11803);
and U11963 (N_11963,N_11843,N_11837);
nor U11964 (N_11964,N_11820,N_11818);
or U11965 (N_11965,N_11785,N_11714);
or U11966 (N_11966,N_11780,N_11797);
nand U11967 (N_11967,N_11719,N_11778);
nor U11968 (N_11968,N_11836,N_11785);
and U11969 (N_11969,N_11725,N_11780);
nand U11970 (N_11970,N_11730,N_11796);
or U11971 (N_11971,N_11735,N_11767);
nand U11972 (N_11972,N_11703,N_11718);
xnor U11973 (N_11973,N_11763,N_11848);
or U11974 (N_11974,N_11827,N_11747);
xor U11975 (N_11975,N_11747,N_11800);
or U11976 (N_11976,N_11848,N_11847);
and U11977 (N_11977,N_11767,N_11834);
and U11978 (N_11978,N_11718,N_11737);
nand U11979 (N_11979,N_11845,N_11724);
nor U11980 (N_11980,N_11758,N_11812);
nand U11981 (N_11981,N_11814,N_11819);
nand U11982 (N_11982,N_11760,N_11774);
or U11983 (N_11983,N_11784,N_11719);
nand U11984 (N_11984,N_11779,N_11788);
xnor U11985 (N_11985,N_11838,N_11767);
xnor U11986 (N_11986,N_11717,N_11743);
and U11987 (N_11987,N_11827,N_11816);
xnor U11988 (N_11988,N_11738,N_11784);
or U11989 (N_11989,N_11816,N_11733);
and U11990 (N_11990,N_11838,N_11826);
nand U11991 (N_11991,N_11718,N_11794);
nor U11992 (N_11992,N_11808,N_11814);
nor U11993 (N_11993,N_11716,N_11727);
nor U11994 (N_11994,N_11777,N_11751);
xor U11995 (N_11995,N_11766,N_11702);
nand U11996 (N_11996,N_11703,N_11839);
xor U11997 (N_11997,N_11738,N_11700);
and U11998 (N_11998,N_11784,N_11796);
or U11999 (N_11999,N_11838,N_11797);
and U12000 (N_12000,N_11917,N_11943);
nand U12001 (N_12001,N_11908,N_11885);
and U12002 (N_12002,N_11884,N_11964);
or U12003 (N_12003,N_11965,N_11871);
and U12004 (N_12004,N_11920,N_11963);
or U12005 (N_12005,N_11967,N_11932);
nand U12006 (N_12006,N_11953,N_11913);
nand U12007 (N_12007,N_11888,N_11882);
nand U12008 (N_12008,N_11983,N_11996);
or U12009 (N_12009,N_11989,N_11931);
nor U12010 (N_12010,N_11880,N_11914);
xor U12011 (N_12011,N_11962,N_11906);
nor U12012 (N_12012,N_11933,N_11993);
or U12013 (N_12013,N_11923,N_11970);
xnor U12014 (N_12014,N_11898,N_11957);
and U12015 (N_12015,N_11975,N_11936);
nor U12016 (N_12016,N_11984,N_11988);
or U12017 (N_12017,N_11903,N_11946);
and U12018 (N_12018,N_11981,N_11948);
and U12019 (N_12019,N_11929,N_11886);
or U12020 (N_12020,N_11941,N_11990);
or U12021 (N_12021,N_11900,N_11955);
and U12022 (N_12022,N_11912,N_11939);
or U12023 (N_12023,N_11907,N_11918);
or U12024 (N_12024,N_11947,N_11887);
or U12025 (N_12025,N_11897,N_11869);
nor U12026 (N_12026,N_11935,N_11873);
or U12027 (N_12027,N_11905,N_11893);
nor U12028 (N_12028,N_11949,N_11919);
xor U12029 (N_12029,N_11892,N_11854);
nand U12030 (N_12030,N_11878,N_11994);
or U12031 (N_12031,N_11977,N_11866);
nand U12032 (N_12032,N_11901,N_11870);
nor U12033 (N_12033,N_11899,N_11868);
xor U12034 (N_12034,N_11863,N_11942);
and U12035 (N_12035,N_11850,N_11934);
or U12036 (N_12036,N_11891,N_11978);
xnor U12037 (N_12037,N_11875,N_11954);
nand U12038 (N_12038,N_11862,N_11979);
xnor U12039 (N_12039,N_11991,N_11950);
and U12040 (N_12040,N_11864,N_11945);
nor U12041 (N_12041,N_11928,N_11937);
nand U12042 (N_12042,N_11976,N_11940);
xnor U12043 (N_12043,N_11971,N_11960);
nand U12044 (N_12044,N_11852,N_11927);
nor U12045 (N_12045,N_11910,N_11915);
and U12046 (N_12046,N_11958,N_11961);
and U12047 (N_12047,N_11980,N_11944);
nand U12048 (N_12048,N_11998,N_11925);
nand U12049 (N_12049,N_11853,N_11890);
xor U12050 (N_12050,N_11872,N_11952);
or U12051 (N_12051,N_11924,N_11982);
nand U12052 (N_12052,N_11930,N_11896);
nor U12053 (N_12053,N_11992,N_11999);
and U12054 (N_12054,N_11861,N_11922);
nand U12055 (N_12055,N_11859,N_11876);
or U12056 (N_12056,N_11926,N_11973);
and U12057 (N_12057,N_11997,N_11956);
nor U12058 (N_12058,N_11916,N_11911);
nand U12059 (N_12059,N_11966,N_11921);
nor U12060 (N_12060,N_11909,N_11857);
and U12061 (N_12061,N_11974,N_11874);
and U12062 (N_12062,N_11969,N_11889);
nor U12063 (N_12063,N_11959,N_11968);
nor U12064 (N_12064,N_11972,N_11985);
and U12065 (N_12065,N_11879,N_11987);
xor U12066 (N_12066,N_11858,N_11894);
and U12067 (N_12067,N_11904,N_11895);
or U12068 (N_12068,N_11877,N_11856);
and U12069 (N_12069,N_11986,N_11883);
nor U12070 (N_12070,N_11938,N_11855);
nand U12071 (N_12071,N_11902,N_11867);
or U12072 (N_12072,N_11881,N_11865);
and U12073 (N_12073,N_11860,N_11851);
xnor U12074 (N_12074,N_11951,N_11995);
or U12075 (N_12075,N_11984,N_11851);
nor U12076 (N_12076,N_11925,N_11907);
xor U12077 (N_12077,N_11887,N_11878);
xor U12078 (N_12078,N_11853,N_11881);
nor U12079 (N_12079,N_11999,N_11908);
and U12080 (N_12080,N_11850,N_11926);
or U12081 (N_12081,N_11926,N_11994);
nor U12082 (N_12082,N_11884,N_11859);
nor U12083 (N_12083,N_11929,N_11881);
nand U12084 (N_12084,N_11913,N_11966);
or U12085 (N_12085,N_11985,N_11875);
nand U12086 (N_12086,N_11854,N_11997);
xor U12087 (N_12087,N_11989,N_11856);
nand U12088 (N_12088,N_11867,N_11964);
or U12089 (N_12089,N_11958,N_11895);
xnor U12090 (N_12090,N_11927,N_11928);
and U12091 (N_12091,N_11878,N_11918);
or U12092 (N_12092,N_11990,N_11922);
and U12093 (N_12093,N_11920,N_11942);
xor U12094 (N_12094,N_11985,N_11994);
and U12095 (N_12095,N_11851,N_11914);
and U12096 (N_12096,N_11896,N_11939);
or U12097 (N_12097,N_11895,N_11877);
nand U12098 (N_12098,N_11998,N_11935);
nor U12099 (N_12099,N_11998,N_11911);
or U12100 (N_12100,N_11861,N_11997);
and U12101 (N_12101,N_11900,N_11989);
and U12102 (N_12102,N_11917,N_11872);
and U12103 (N_12103,N_11890,N_11966);
or U12104 (N_12104,N_11949,N_11857);
nor U12105 (N_12105,N_11853,N_11903);
and U12106 (N_12106,N_11912,N_11899);
or U12107 (N_12107,N_11851,N_11992);
and U12108 (N_12108,N_11911,N_11889);
nor U12109 (N_12109,N_11872,N_11915);
nand U12110 (N_12110,N_11977,N_11967);
nor U12111 (N_12111,N_11981,N_11976);
xor U12112 (N_12112,N_11945,N_11872);
nand U12113 (N_12113,N_11972,N_11903);
nand U12114 (N_12114,N_11955,N_11949);
nand U12115 (N_12115,N_11927,N_11911);
xnor U12116 (N_12116,N_11918,N_11981);
or U12117 (N_12117,N_11985,N_11902);
and U12118 (N_12118,N_11953,N_11940);
xnor U12119 (N_12119,N_11874,N_11879);
nor U12120 (N_12120,N_11875,N_11919);
or U12121 (N_12121,N_11944,N_11988);
or U12122 (N_12122,N_11869,N_11967);
nand U12123 (N_12123,N_11916,N_11884);
and U12124 (N_12124,N_11910,N_11875);
and U12125 (N_12125,N_11924,N_11969);
and U12126 (N_12126,N_11930,N_11913);
nor U12127 (N_12127,N_11996,N_11910);
or U12128 (N_12128,N_11904,N_11931);
and U12129 (N_12129,N_11921,N_11975);
and U12130 (N_12130,N_11899,N_11936);
and U12131 (N_12131,N_11953,N_11952);
or U12132 (N_12132,N_11953,N_11930);
nor U12133 (N_12133,N_11883,N_11983);
nand U12134 (N_12134,N_11998,N_11861);
nand U12135 (N_12135,N_11878,N_11938);
xor U12136 (N_12136,N_11929,N_11868);
nand U12137 (N_12137,N_11997,N_11869);
nor U12138 (N_12138,N_11942,N_11916);
or U12139 (N_12139,N_11909,N_11984);
nor U12140 (N_12140,N_11917,N_11887);
xnor U12141 (N_12141,N_11982,N_11976);
nor U12142 (N_12142,N_11928,N_11866);
and U12143 (N_12143,N_11896,N_11977);
nor U12144 (N_12144,N_11905,N_11874);
nand U12145 (N_12145,N_11991,N_11878);
and U12146 (N_12146,N_11855,N_11985);
nor U12147 (N_12147,N_11860,N_11956);
or U12148 (N_12148,N_11969,N_11886);
nand U12149 (N_12149,N_11980,N_11941);
or U12150 (N_12150,N_12056,N_12144);
nand U12151 (N_12151,N_12114,N_12085);
nand U12152 (N_12152,N_12097,N_12067);
and U12153 (N_12153,N_12108,N_12140);
and U12154 (N_12154,N_12054,N_12104);
xnor U12155 (N_12155,N_12132,N_12095);
or U12156 (N_12156,N_12003,N_12099);
or U12157 (N_12157,N_12063,N_12025);
and U12158 (N_12158,N_12070,N_12051);
or U12159 (N_12159,N_12079,N_12026);
and U12160 (N_12160,N_12135,N_12141);
or U12161 (N_12161,N_12033,N_12064);
nor U12162 (N_12162,N_12058,N_12116);
nor U12163 (N_12163,N_12014,N_12048);
nand U12164 (N_12164,N_12084,N_12069);
and U12165 (N_12165,N_12131,N_12005);
nor U12166 (N_12166,N_12093,N_12136);
or U12167 (N_12167,N_12074,N_12105);
nor U12168 (N_12168,N_12021,N_12027);
and U12169 (N_12169,N_12018,N_12062);
nor U12170 (N_12170,N_12006,N_12077);
or U12171 (N_12171,N_12008,N_12089);
and U12172 (N_12172,N_12013,N_12039);
nor U12173 (N_12173,N_12088,N_12125);
nor U12174 (N_12174,N_12111,N_12129);
and U12175 (N_12175,N_12142,N_12009);
xnor U12176 (N_12176,N_12061,N_12083);
and U12177 (N_12177,N_12107,N_12007);
xnor U12178 (N_12178,N_12115,N_12049);
or U12179 (N_12179,N_12100,N_12012);
or U12180 (N_12180,N_12035,N_12110);
nor U12181 (N_12181,N_12094,N_12134);
xor U12182 (N_12182,N_12038,N_12047);
or U12183 (N_12183,N_12023,N_12148);
nand U12184 (N_12184,N_12113,N_12103);
and U12185 (N_12185,N_12001,N_12045);
or U12186 (N_12186,N_12126,N_12128);
nor U12187 (N_12187,N_12032,N_12091);
xnor U12188 (N_12188,N_12065,N_12127);
xor U12189 (N_12189,N_12092,N_12098);
nor U12190 (N_12190,N_12066,N_12010);
nor U12191 (N_12191,N_12019,N_12090);
or U12192 (N_12192,N_12040,N_12016);
and U12193 (N_12193,N_12015,N_12109);
nand U12194 (N_12194,N_12086,N_12096);
or U12195 (N_12195,N_12137,N_12036);
xnor U12196 (N_12196,N_12020,N_12106);
or U12197 (N_12197,N_12044,N_12138);
nand U12198 (N_12198,N_12043,N_12034);
and U12199 (N_12199,N_12119,N_12011);
or U12200 (N_12200,N_12055,N_12000);
nand U12201 (N_12201,N_12120,N_12146);
xor U12202 (N_12202,N_12143,N_12042);
xnor U12203 (N_12203,N_12124,N_12078);
nor U12204 (N_12204,N_12087,N_12080);
xnor U12205 (N_12205,N_12081,N_12082);
and U12206 (N_12206,N_12057,N_12068);
xnor U12207 (N_12207,N_12053,N_12072);
xor U12208 (N_12208,N_12004,N_12133);
and U12209 (N_12209,N_12002,N_12101);
or U12210 (N_12210,N_12017,N_12117);
nand U12211 (N_12211,N_12030,N_12139);
nor U12212 (N_12212,N_12121,N_12130);
nand U12213 (N_12213,N_12022,N_12118);
and U12214 (N_12214,N_12031,N_12060);
and U12215 (N_12215,N_12145,N_12122);
and U12216 (N_12216,N_12149,N_12046);
and U12217 (N_12217,N_12037,N_12076);
and U12218 (N_12218,N_12050,N_12059);
and U12219 (N_12219,N_12075,N_12147);
or U12220 (N_12220,N_12028,N_12071);
nor U12221 (N_12221,N_12029,N_12112);
or U12222 (N_12222,N_12073,N_12123);
nand U12223 (N_12223,N_12024,N_12102);
nand U12224 (N_12224,N_12041,N_12052);
nor U12225 (N_12225,N_12080,N_12125);
nand U12226 (N_12226,N_12136,N_12036);
nor U12227 (N_12227,N_12026,N_12025);
nand U12228 (N_12228,N_12076,N_12111);
and U12229 (N_12229,N_12132,N_12093);
and U12230 (N_12230,N_12091,N_12025);
and U12231 (N_12231,N_12043,N_12097);
xor U12232 (N_12232,N_12081,N_12117);
or U12233 (N_12233,N_12127,N_12062);
nand U12234 (N_12234,N_12088,N_12022);
nor U12235 (N_12235,N_12001,N_12079);
xnor U12236 (N_12236,N_12042,N_12076);
xnor U12237 (N_12237,N_12099,N_12006);
and U12238 (N_12238,N_12074,N_12034);
and U12239 (N_12239,N_12081,N_12123);
and U12240 (N_12240,N_12048,N_12047);
or U12241 (N_12241,N_12103,N_12063);
and U12242 (N_12242,N_12147,N_12047);
nor U12243 (N_12243,N_12054,N_12133);
xor U12244 (N_12244,N_12132,N_12092);
and U12245 (N_12245,N_12130,N_12046);
nand U12246 (N_12246,N_12044,N_12092);
nor U12247 (N_12247,N_12031,N_12101);
and U12248 (N_12248,N_12074,N_12079);
and U12249 (N_12249,N_12086,N_12089);
nand U12250 (N_12250,N_12079,N_12103);
nand U12251 (N_12251,N_12007,N_12149);
and U12252 (N_12252,N_12007,N_12058);
and U12253 (N_12253,N_12105,N_12066);
nand U12254 (N_12254,N_12143,N_12133);
xor U12255 (N_12255,N_12108,N_12088);
and U12256 (N_12256,N_12105,N_12125);
nor U12257 (N_12257,N_12007,N_12148);
or U12258 (N_12258,N_12132,N_12147);
xor U12259 (N_12259,N_12090,N_12006);
and U12260 (N_12260,N_12099,N_12112);
or U12261 (N_12261,N_12132,N_12004);
xor U12262 (N_12262,N_12100,N_12059);
nor U12263 (N_12263,N_12089,N_12005);
and U12264 (N_12264,N_12069,N_12077);
xor U12265 (N_12265,N_12143,N_12037);
xnor U12266 (N_12266,N_12078,N_12000);
or U12267 (N_12267,N_12111,N_12029);
xor U12268 (N_12268,N_12008,N_12115);
nand U12269 (N_12269,N_12079,N_12124);
nor U12270 (N_12270,N_12136,N_12005);
nand U12271 (N_12271,N_12133,N_12051);
xor U12272 (N_12272,N_12112,N_12063);
nor U12273 (N_12273,N_12104,N_12082);
nor U12274 (N_12274,N_12080,N_12064);
or U12275 (N_12275,N_12024,N_12080);
or U12276 (N_12276,N_12103,N_12119);
and U12277 (N_12277,N_12127,N_12123);
nor U12278 (N_12278,N_12046,N_12017);
xnor U12279 (N_12279,N_12107,N_12023);
nand U12280 (N_12280,N_12036,N_12139);
or U12281 (N_12281,N_12038,N_12069);
and U12282 (N_12282,N_12069,N_12048);
nor U12283 (N_12283,N_12097,N_12143);
nor U12284 (N_12284,N_12138,N_12034);
or U12285 (N_12285,N_12093,N_12000);
or U12286 (N_12286,N_12092,N_12123);
nand U12287 (N_12287,N_12096,N_12133);
or U12288 (N_12288,N_12067,N_12123);
and U12289 (N_12289,N_12108,N_12100);
nor U12290 (N_12290,N_12138,N_12028);
xnor U12291 (N_12291,N_12039,N_12074);
and U12292 (N_12292,N_12051,N_12028);
or U12293 (N_12293,N_12000,N_12146);
or U12294 (N_12294,N_12128,N_12102);
xor U12295 (N_12295,N_12063,N_12109);
and U12296 (N_12296,N_12030,N_12009);
and U12297 (N_12297,N_12022,N_12127);
xor U12298 (N_12298,N_12015,N_12068);
nand U12299 (N_12299,N_12007,N_12085);
or U12300 (N_12300,N_12245,N_12297);
and U12301 (N_12301,N_12284,N_12274);
and U12302 (N_12302,N_12243,N_12267);
or U12303 (N_12303,N_12230,N_12182);
xor U12304 (N_12304,N_12215,N_12269);
nand U12305 (N_12305,N_12293,N_12238);
xnor U12306 (N_12306,N_12291,N_12263);
and U12307 (N_12307,N_12295,N_12199);
nand U12308 (N_12308,N_12173,N_12228);
and U12309 (N_12309,N_12299,N_12162);
or U12310 (N_12310,N_12264,N_12231);
or U12311 (N_12311,N_12201,N_12156);
xnor U12312 (N_12312,N_12247,N_12208);
xnor U12313 (N_12313,N_12285,N_12193);
xor U12314 (N_12314,N_12187,N_12160);
or U12315 (N_12315,N_12229,N_12172);
xnor U12316 (N_12316,N_12197,N_12296);
and U12317 (N_12317,N_12268,N_12218);
and U12318 (N_12318,N_12184,N_12234);
nand U12319 (N_12319,N_12178,N_12248);
and U12320 (N_12320,N_12246,N_12233);
and U12321 (N_12321,N_12158,N_12177);
nor U12322 (N_12322,N_12232,N_12287);
nor U12323 (N_12323,N_12191,N_12249);
xor U12324 (N_12324,N_12235,N_12194);
nor U12325 (N_12325,N_12169,N_12183);
or U12326 (N_12326,N_12276,N_12205);
xor U12327 (N_12327,N_12209,N_12265);
or U12328 (N_12328,N_12161,N_12254);
or U12329 (N_12329,N_12179,N_12251);
xnor U12330 (N_12330,N_12278,N_12151);
xnor U12331 (N_12331,N_12219,N_12255);
nand U12332 (N_12332,N_12239,N_12279);
and U12333 (N_12333,N_12275,N_12206);
xor U12334 (N_12334,N_12250,N_12272);
nor U12335 (N_12335,N_12170,N_12256);
and U12336 (N_12336,N_12286,N_12202);
nor U12337 (N_12337,N_12152,N_12283);
or U12338 (N_12338,N_12280,N_12176);
xnor U12339 (N_12339,N_12240,N_12159);
nor U12340 (N_12340,N_12189,N_12198);
and U12341 (N_12341,N_12259,N_12281);
xnor U12342 (N_12342,N_12174,N_12292);
nand U12343 (N_12343,N_12186,N_12180);
or U12344 (N_12344,N_12195,N_12214);
nand U12345 (N_12345,N_12167,N_12223);
or U12346 (N_12346,N_12273,N_12271);
nor U12347 (N_12347,N_12190,N_12155);
nor U12348 (N_12348,N_12210,N_12192);
nor U12349 (N_12349,N_12282,N_12227);
and U12350 (N_12350,N_12216,N_12252);
nand U12351 (N_12351,N_12241,N_12168);
and U12352 (N_12352,N_12171,N_12266);
nor U12353 (N_12353,N_12277,N_12225);
nor U12354 (N_12354,N_12298,N_12222);
xnor U12355 (N_12355,N_12288,N_12185);
and U12356 (N_12356,N_12242,N_12257);
or U12357 (N_12357,N_12261,N_12181);
xor U12358 (N_12358,N_12207,N_12212);
and U12359 (N_12359,N_12289,N_12220);
nor U12360 (N_12360,N_12211,N_12157);
xnor U12361 (N_12361,N_12154,N_12164);
nor U12362 (N_12362,N_12175,N_12188);
xor U12363 (N_12363,N_12236,N_12150);
xor U12364 (N_12364,N_12253,N_12217);
and U12365 (N_12365,N_12163,N_12270);
and U12366 (N_12366,N_12200,N_12153);
nand U12367 (N_12367,N_12221,N_12213);
xnor U12368 (N_12368,N_12260,N_12294);
nor U12369 (N_12369,N_12166,N_12224);
xor U12370 (N_12370,N_12165,N_12237);
nand U12371 (N_12371,N_12203,N_12244);
or U12372 (N_12372,N_12196,N_12226);
nor U12373 (N_12373,N_12258,N_12204);
nand U12374 (N_12374,N_12262,N_12290);
xor U12375 (N_12375,N_12196,N_12162);
xnor U12376 (N_12376,N_12269,N_12287);
xor U12377 (N_12377,N_12164,N_12171);
or U12378 (N_12378,N_12278,N_12224);
or U12379 (N_12379,N_12293,N_12196);
nor U12380 (N_12380,N_12159,N_12274);
nand U12381 (N_12381,N_12248,N_12171);
nor U12382 (N_12382,N_12273,N_12154);
xor U12383 (N_12383,N_12215,N_12278);
or U12384 (N_12384,N_12236,N_12167);
or U12385 (N_12385,N_12257,N_12215);
nand U12386 (N_12386,N_12233,N_12288);
and U12387 (N_12387,N_12266,N_12280);
nand U12388 (N_12388,N_12257,N_12210);
nor U12389 (N_12389,N_12212,N_12236);
nand U12390 (N_12390,N_12223,N_12267);
xor U12391 (N_12391,N_12187,N_12249);
xnor U12392 (N_12392,N_12288,N_12158);
nor U12393 (N_12393,N_12159,N_12190);
or U12394 (N_12394,N_12268,N_12282);
and U12395 (N_12395,N_12283,N_12175);
xnor U12396 (N_12396,N_12200,N_12159);
nor U12397 (N_12397,N_12185,N_12241);
nor U12398 (N_12398,N_12231,N_12240);
and U12399 (N_12399,N_12263,N_12195);
or U12400 (N_12400,N_12208,N_12243);
nand U12401 (N_12401,N_12204,N_12273);
nand U12402 (N_12402,N_12159,N_12214);
and U12403 (N_12403,N_12175,N_12154);
nor U12404 (N_12404,N_12191,N_12167);
and U12405 (N_12405,N_12153,N_12266);
nand U12406 (N_12406,N_12264,N_12196);
or U12407 (N_12407,N_12287,N_12263);
nand U12408 (N_12408,N_12275,N_12194);
nand U12409 (N_12409,N_12156,N_12165);
and U12410 (N_12410,N_12243,N_12185);
nor U12411 (N_12411,N_12243,N_12236);
nor U12412 (N_12412,N_12260,N_12167);
xor U12413 (N_12413,N_12185,N_12150);
nor U12414 (N_12414,N_12204,N_12226);
and U12415 (N_12415,N_12205,N_12236);
or U12416 (N_12416,N_12259,N_12220);
or U12417 (N_12417,N_12237,N_12263);
and U12418 (N_12418,N_12276,N_12259);
xnor U12419 (N_12419,N_12214,N_12240);
nor U12420 (N_12420,N_12264,N_12235);
xnor U12421 (N_12421,N_12155,N_12205);
or U12422 (N_12422,N_12259,N_12175);
xor U12423 (N_12423,N_12235,N_12223);
nand U12424 (N_12424,N_12177,N_12160);
nand U12425 (N_12425,N_12175,N_12238);
and U12426 (N_12426,N_12184,N_12244);
and U12427 (N_12427,N_12155,N_12179);
or U12428 (N_12428,N_12231,N_12171);
nand U12429 (N_12429,N_12223,N_12219);
or U12430 (N_12430,N_12257,N_12290);
and U12431 (N_12431,N_12282,N_12219);
and U12432 (N_12432,N_12153,N_12209);
xnor U12433 (N_12433,N_12256,N_12227);
or U12434 (N_12434,N_12180,N_12240);
or U12435 (N_12435,N_12291,N_12285);
xor U12436 (N_12436,N_12291,N_12205);
and U12437 (N_12437,N_12299,N_12249);
nand U12438 (N_12438,N_12286,N_12211);
xnor U12439 (N_12439,N_12272,N_12271);
or U12440 (N_12440,N_12213,N_12242);
xnor U12441 (N_12441,N_12257,N_12213);
xnor U12442 (N_12442,N_12171,N_12161);
xnor U12443 (N_12443,N_12203,N_12254);
nand U12444 (N_12444,N_12216,N_12259);
nor U12445 (N_12445,N_12292,N_12271);
xnor U12446 (N_12446,N_12186,N_12185);
xnor U12447 (N_12447,N_12197,N_12282);
nor U12448 (N_12448,N_12152,N_12154);
and U12449 (N_12449,N_12209,N_12282);
or U12450 (N_12450,N_12317,N_12425);
and U12451 (N_12451,N_12313,N_12322);
and U12452 (N_12452,N_12388,N_12347);
xnor U12453 (N_12453,N_12325,N_12382);
nor U12454 (N_12454,N_12436,N_12403);
or U12455 (N_12455,N_12412,N_12316);
nand U12456 (N_12456,N_12390,N_12442);
and U12457 (N_12457,N_12398,N_12417);
and U12458 (N_12458,N_12326,N_12364);
and U12459 (N_12459,N_12427,N_12304);
xor U12460 (N_12460,N_12370,N_12401);
and U12461 (N_12461,N_12335,N_12352);
xor U12462 (N_12462,N_12374,N_12440);
xnor U12463 (N_12463,N_12367,N_12318);
xnor U12464 (N_12464,N_12319,N_12360);
nor U12465 (N_12465,N_12428,N_12324);
xor U12466 (N_12466,N_12345,N_12418);
and U12467 (N_12467,N_12393,N_12310);
and U12468 (N_12468,N_12340,N_12435);
nand U12469 (N_12469,N_12353,N_12355);
nand U12470 (N_12470,N_12331,N_12338);
or U12471 (N_12471,N_12446,N_12387);
xnor U12472 (N_12472,N_12327,N_12375);
nor U12473 (N_12473,N_12311,N_12300);
or U12474 (N_12474,N_12302,N_12426);
xor U12475 (N_12475,N_12429,N_12341);
and U12476 (N_12476,N_12423,N_12408);
and U12477 (N_12477,N_12445,N_12358);
or U12478 (N_12478,N_12373,N_12330);
and U12479 (N_12479,N_12357,N_12447);
or U12480 (N_12480,N_12439,N_12362);
and U12481 (N_12481,N_12348,N_12312);
or U12482 (N_12482,N_12307,N_12350);
nor U12483 (N_12483,N_12306,N_12328);
and U12484 (N_12484,N_12409,N_12421);
or U12485 (N_12485,N_12399,N_12397);
nand U12486 (N_12486,N_12415,N_12379);
xor U12487 (N_12487,N_12321,N_12444);
and U12488 (N_12488,N_12315,N_12380);
or U12489 (N_12489,N_12371,N_12349);
nor U12490 (N_12490,N_12346,N_12422);
or U12491 (N_12491,N_12411,N_12416);
nor U12492 (N_12492,N_12339,N_12424);
or U12493 (N_12493,N_12314,N_12378);
or U12494 (N_12494,N_12431,N_12356);
and U12495 (N_12495,N_12342,N_12301);
or U12496 (N_12496,N_12448,N_12406);
or U12497 (N_12497,N_12396,N_12385);
xnor U12498 (N_12498,N_12363,N_12383);
or U12499 (N_12499,N_12320,N_12365);
nand U12500 (N_12500,N_12392,N_12402);
and U12501 (N_12501,N_12361,N_12323);
xor U12502 (N_12502,N_12343,N_12381);
nor U12503 (N_12503,N_12386,N_12384);
nor U12504 (N_12504,N_12430,N_12432);
and U12505 (N_12505,N_12344,N_12414);
nor U12506 (N_12506,N_12405,N_12351);
nor U12507 (N_12507,N_12333,N_12420);
and U12508 (N_12508,N_12334,N_12443);
and U12509 (N_12509,N_12366,N_12369);
nor U12510 (N_12510,N_12359,N_12441);
nand U12511 (N_12511,N_12449,N_12337);
nor U12512 (N_12512,N_12368,N_12329);
and U12513 (N_12513,N_12309,N_12437);
nor U12514 (N_12514,N_12434,N_12433);
or U12515 (N_12515,N_12308,N_12410);
nor U12516 (N_12516,N_12419,N_12303);
or U12517 (N_12517,N_12354,N_12395);
or U12518 (N_12518,N_12389,N_12376);
nand U12519 (N_12519,N_12305,N_12377);
nor U12520 (N_12520,N_12404,N_12391);
or U12521 (N_12521,N_12413,N_12336);
nand U12522 (N_12522,N_12394,N_12372);
xnor U12523 (N_12523,N_12438,N_12400);
nand U12524 (N_12524,N_12407,N_12332);
xnor U12525 (N_12525,N_12343,N_12411);
nand U12526 (N_12526,N_12437,N_12323);
xor U12527 (N_12527,N_12386,N_12312);
xnor U12528 (N_12528,N_12340,N_12446);
or U12529 (N_12529,N_12323,N_12373);
nor U12530 (N_12530,N_12320,N_12396);
nor U12531 (N_12531,N_12398,N_12439);
nand U12532 (N_12532,N_12351,N_12308);
and U12533 (N_12533,N_12417,N_12353);
and U12534 (N_12534,N_12360,N_12358);
xor U12535 (N_12535,N_12301,N_12348);
and U12536 (N_12536,N_12370,N_12355);
nor U12537 (N_12537,N_12365,N_12324);
nand U12538 (N_12538,N_12415,N_12366);
nand U12539 (N_12539,N_12374,N_12365);
xor U12540 (N_12540,N_12332,N_12371);
or U12541 (N_12541,N_12434,N_12440);
nand U12542 (N_12542,N_12421,N_12358);
nand U12543 (N_12543,N_12380,N_12329);
and U12544 (N_12544,N_12421,N_12360);
or U12545 (N_12545,N_12399,N_12303);
xor U12546 (N_12546,N_12343,N_12309);
nor U12547 (N_12547,N_12361,N_12412);
and U12548 (N_12548,N_12357,N_12441);
nand U12549 (N_12549,N_12392,N_12337);
or U12550 (N_12550,N_12351,N_12345);
xor U12551 (N_12551,N_12349,N_12449);
nor U12552 (N_12552,N_12402,N_12321);
xnor U12553 (N_12553,N_12369,N_12401);
or U12554 (N_12554,N_12312,N_12364);
nor U12555 (N_12555,N_12388,N_12327);
nor U12556 (N_12556,N_12317,N_12378);
nor U12557 (N_12557,N_12373,N_12363);
nand U12558 (N_12558,N_12329,N_12394);
and U12559 (N_12559,N_12303,N_12422);
and U12560 (N_12560,N_12363,N_12407);
and U12561 (N_12561,N_12347,N_12370);
xnor U12562 (N_12562,N_12327,N_12303);
xnor U12563 (N_12563,N_12435,N_12405);
or U12564 (N_12564,N_12348,N_12309);
nor U12565 (N_12565,N_12383,N_12403);
nand U12566 (N_12566,N_12392,N_12390);
and U12567 (N_12567,N_12314,N_12360);
and U12568 (N_12568,N_12423,N_12380);
nor U12569 (N_12569,N_12354,N_12440);
or U12570 (N_12570,N_12323,N_12308);
nor U12571 (N_12571,N_12320,N_12432);
or U12572 (N_12572,N_12365,N_12370);
or U12573 (N_12573,N_12433,N_12307);
nand U12574 (N_12574,N_12356,N_12370);
nor U12575 (N_12575,N_12329,N_12312);
or U12576 (N_12576,N_12425,N_12400);
nand U12577 (N_12577,N_12356,N_12327);
and U12578 (N_12578,N_12372,N_12406);
nor U12579 (N_12579,N_12389,N_12362);
xnor U12580 (N_12580,N_12382,N_12406);
xor U12581 (N_12581,N_12308,N_12439);
nor U12582 (N_12582,N_12339,N_12325);
nor U12583 (N_12583,N_12332,N_12329);
xor U12584 (N_12584,N_12366,N_12359);
nor U12585 (N_12585,N_12423,N_12435);
nor U12586 (N_12586,N_12364,N_12343);
xnor U12587 (N_12587,N_12411,N_12408);
xor U12588 (N_12588,N_12344,N_12326);
nand U12589 (N_12589,N_12431,N_12397);
xor U12590 (N_12590,N_12416,N_12427);
nand U12591 (N_12591,N_12440,N_12376);
xor U12592 (N_12592,N_12341,N_12317);
and U12593 (N_12593,N_12446,N_12390);
nand U12594 (N_12594,N_12426,N_12355);
xnor U12595 (N_12595,N_12344,N_12434);
and U12596 (N_12596,N_12416,N_12406);
or U12597 (N_12597,N_12355,N_12325);
and U12598 (N_12598,N_12353,N_12435);
nand U12599 (N_12599,N_12395,N_12347);
xnor U12600 (N_12600,N_12577,N_12466);
and U12601 (N_12601,N_12459,N_12536);
or U12602 (N_12602,N_12452,N_12499);
and U12603 (N_12603,N_12513,N_12593);
or U12604 (N_12604,N_12565,N_12488);
nor U12605 (N_12605,N_12522,N_12569);
or U12606 (N_12606,N_12542,N_12451);
nor U12607 (N_12607,N_12551,N_12591);
nor U12608 (N_12608,N_12586,N_12579);
or U12609 (N_12609,N_12547,N_12465);
nor U12610 (N_12610,N_12462,N_12599);
xor U12611 (N_12611,N_12523,N_12534);
xor U12612 (N_12612,N_12475,N_12543);
nor U12613 (N_12613,N_12470,N_12487);
nand U12614 (N_12614,N_12507,N_12483);
or U12615 (N_12615,N_12486,N_12587);
nor U12616 (N_12616,N_12588,N_12598);
and U12617 (N_12617,N_12464,N_12566);
and U12618 (N_12618,N_12535,N_12519);
nand U12619 (N_12619,N_12576,N_12479);
or U12620 (N_12620,N_12510,N_12564);
xor U12621 (N_12621,N_12512,N_12578);
and U12622 (N_12622,N_12545,N_12489);
or U12623 (N_12623,N_12456,N_12544);
or U12624 (N_12624,N_12495,N_12532);
and U12625 (N_12625,N_12500,N_12538);
nand U12626 (N_12626,N_12550,N_12469);
or U12627 (N_12627,N_12539,N_12540);
and U12628 (N_12628,N_12580,N_12527);
xnor U12629 (N_12629,N_12570,N_12521);
and U12630 (N_12630,N_12548,N_12557);
xor U12631 (N_12631,N_12582,N_12460);
xor U12632 (N_12632,N_12457,N_12480);
nand U12633 (N_12633,N_12589,N_12455);
xnor U12634 (N_12634,N_12563,N_12514);
or U12635 (N_12635,N_12458,N_12561);
xor U12636 (N_12636,N_12511,N_12506);
nor U12637 (N_12637,N_12516,N_12574);
nand U12638 (N_12638,N_12450,N_12485);
and U12639 (N_12639,N_12491,N_12508);
nand U12640 (N_12640,N_12454,N_12583);
or U12641 (N_12641,N_12472,N_12473);
or U12642 (N_12642,N_12526,N_12471);
nor U12643 (N_12643,N_12501,N_12515);
and U12644 (N_12644,N_12590,N_12559);
nor U12645 (N_12645,N_12585,N_12482);
xor U12646 (N_12646,N_12555,N_12562);
xor U12647 (N_12647,N_12517,N_12572);
or U12648 (N_12648,N_12467,N_12478);
and U12649 (N_12649,N_12584,N_12463);
and U12650 (N_12650,N_12568,N_12481);
nor U12651 (N_12651,N_12531,N_12595);
or U12652 (N_12652,N_12537,N_12529);
or U12653 (N_12653,N_12554,N_12504);
nor U12654 (N_12654,N_12567,N_12571);
and U12655 (N_12655,N_12558,N_12503);
or U12656 (N_12656,N_12530,N_12474);
nor U12657 (N_12657,N_12502,N_12553);
and U12658 (N_12658,N_12520,N_12573);
xor U12659 (N_12659,N_12549,N_12492);
nand U12660 (N_12660,N_12575,N_12546);
or U12661 (N_12661,N_12596,N_12518);
xor U12662 (N_12662,N_12541,N_12597);
xnor U12663 (N_12663,N_12477,N_12524);
nor U12664 (N_12664,N_12533,N_12509);
and U12665 (N_12665,N_12525,N_12581);
or U12666 (N_12666,N_12496,N_12497);
and U12667 (N_12667,N_12556,N_12453);
nand U12668 (N_12668,N_12592,N_12484);
xor U12669 (N_12669,N_12505,N_12461);
and U12670 (N_12670,N_12498,N_12560);
and U12671 (N_12671,N_12594,N_12552);
nand U12672 (N_12672,N_12528,N_12468);
or U12673 (N_12673,N_12494,N_12476);
and U12674 (N_12674,N_12490,N_12493);
nor U12675 (N_12675,N_12463,N_12554);
or U12676 (N_12676,N_12561,N_12588);
xor U12677 (N_12677,N_12507,N_12491);
nand U12678 (N_12678,N_12524,N_12562);
xnor U12679 (N_12679,N_12506,N_12567);
nor U12680 (N_12680,N_12529,N_12505);
nor U12681 (N_12681,N_12455,N_12494);
xor U12682 (N_12682,N_12488,N_12482);
or U12683 (N_12683,N_12464,N_12535);
nand U12684 (N_12684,N_12569,N_12552);
or U12685 (N_12685,N_12503,N_12522);
and U12686 (N_12686,N_12498,N_12539);
xnor U12687 (N_12687,N_12545,N_12517);
and U12688 (N_12688,N_12518,N_12510);
xor U12689 (N_12689,N_12580,N_12464);
nand U12690 (N_12690,N_12590,N_12454);
nor U12691 (N_12691,N_12469,N_12496);
nand U12692 (N_12692,N_12596,N_12472);
and U12693 (N_12693,N_12519,N_12528);
nor U12694 (N_12694,N_12569,N_12462);
nor U12695 (N_12695,N_12553,N_12562);
nand U12696 (N_12696,N_12469,N_12573);
nor U12697 (N_12697,N_12483,N_12560);
xnor U12698 (N_12698,N_12462,N_12556);
nor U12699 (N_12699,N_12591,N_12568);
and U12700 (N_12700,N_12587,N_12565);
xnor U12701 (N_12701,N_12499,N_12533);
xor U12702 (N_12702,N_12535,N_12521);
xnor U12703 (N_12703,N_12559,N_12465);
nor U12704 (N_12704,N_12482,N_12550);
or U12705 (N_12705,N_12576,N_12566);
xor U12706 (N_12706,N_12516,N_12461);
nand U12707 (N_12707,N_12585,N_12491);
or U12708 (N_12708,N_12531,N_12582);
nor U12709 (N_12709,N_12558,N_12550);
nand U12710 (N_12710,N_12519,N_12551);
or U12711 (N_12711,N_12548,N_12572);
or U12712 (N_12712,N_12570,N_12558);
xnor U12713 (N_12713,N_12497,N_12562);
nand U12714 (N_12714,N_12564,N_12521);
or U12715 (N_12715,N_12539,N_12589);
or U12716 (N_12716,N_12560,N_12492);
nand U12717 (N_12717,N_12469,N_12540);
xor U12718 (N_12718,N_12474,N_12556);
and U12719 (N_12719,N_12539,N_12458);
nand U12720 (N_12720,N_12576,N_12548);
nor U12721 (N_12721,N_12549,N_12552);
nand U12722 (N_12722,N_12459,N_12511);
nor U12723 (N_12723,N_12552,N_12450);
nor U12724 (N_12724,N_12540,N_12596);
and U12725 (N_12725,N_12532,N_12584);
xnor U12726 (N_12726,N_12536,N_12558);
nand U12727 (N_12727,N_12519,N_12482);
and U12728 (N_12728,N_12487,N_12523);
xor U12729 (N_12729,N_12568,N_12597);
nand U12730 (N_12730,N_12534,N_12458);
nand U12731 (N_12731,N_12474,N_12571);
and U12732 (N_12732,N_12515,N_12576);
or U12733 (N_12733,N_12497,N_12592);
xnor U12734 (N_12734,N_12563,N_12512);
nand U12735 (N_12735,N_12512,N_12457);
xnor U12736 (N_12736,N_12562,N_12585);
or U12737 (N_12737,N_12561,N_12582);
or U12738 (N_12738,N_12536,N_12470);
nor U12739 (N_12739,N_12487,N_12509);
nand U12740 (N_12740,N_12517,N_12477);
nor U12741 (N_12741,N_12514,N_12520);
nand U12742 (N_12742,N_12537,N_12576);
xor U12743 (N_12743,N_12596,N_12454);
nor U12744 (N_12744,N_12522,N_12529);
and U12745 (N_12745,N_12536,N_12593);
nor U12746 (N_12746,N_12567,N_12530);
nand U12747 (N_12747,N_12478,N_12480);
and U12748 (N_12748,N_12549,N_12461);
xor U12749 (N_12749,N_12489,N_12582);
and U12750 (N_12750,N_12739,N_12681);
xnor U12751 (N_12751,N_12610,N_12747);
and U12752 (N_12752,N_12711,N_12643);
or U12753 (N_12753,N_12665,N_12686);
xor U12754 (N_12754,N_12746,N_12741);
or U12755 (N_12755,N_12647,N_12736);
and U12756 (N_12756,N_12651,N_12669);
and U12757 (N_12757,N_12718,N_12743);
xor U12758 (N_12758,N_12679,N_12659);
and U12759 (N_12759,N_12668,N_12705);
and U12760 (N_12760,N_12616,N_12609);
xnor U12761 (N_12761,N_12708,N_12626);
xor U12762 (N_12762,N_12640,N_12693);
nand U12763 (N_12763,N_12704,N_12694);
or U12764 (N_12764,N_12667,N_12622);
and U12765 (N_12765,N_12723,N_12670);
and U12766 (N_12766,N_12678,N_12676);
nor U12767 (N_12767,N_12638,N_12715);
nand U12768 (N_12768,N_12707,N_12748);
or U12769 (N_12769,N_12688,N_12700);
xor U12770 (N_12770,N_12646,N_12733);
xnor U12771 (N_12771,N_12709,N_12735);
nand U12772 (N_12772,N_12689,N_12619);
and U12773 (N_12773,N_12695,N_12637);
xor U12774 (N_12774,N_12644,N_12682);
nor U12775 (N_12775,N_12677,N_12737);
xnor U12776 (N_12776,N_12714,N_12630);
nand U12777 (N_12777,N_12608,N_12703);
nand U12778 (N_12778,N_12673,N_12639);
xnor U12779 (N_12779,N_12618,N_12604);
xor U12780 (N_12780,N_12740,N_12687);
or U12781 (N_12781,N_12654,N_12690);
or U12782 (N_12782,N_12655,N_12671);
xnor U12783 (N_12783,N_12692,N_12629);
nand U12784 (N_12784,N_12642,N_12738);
or U12785 (N_12785,N_12648,N_12652);
nand U12786 (N_12786,N_12734,N_12620);
nor U12787 (N_12787,N_12658,N_12623);
or U12788 (N_12788,N_12727,N_12613);
or U12789 (N_12789,N_12636,N_12606);
nand U12790 (N_12790,N_12617,N_12600);
or U12791 (N_12791,N_12645,N_12716);
nor U12792 (N_12792,N_12706,N_12656);
and U12793 (N_12793,N_12699,N_12724);
xor U12794 (N_12794,N_12701,N_12663);
xor U12795 (N_12795,N_12691,N_12722);
xor U12796 (N_12796,N_12713,N_12712);
and U12797 (N_12797,N_12614,N_12607);
nand U12798 (N_12798,N_12698,N_12631);
and U12799 (N_12799,N_12702,N_12657);
nand U12800 (N_12800,N_12719,N_12721);
nand U12801 (N_12801,N_12742,N_12732);
or U12802 (N_12802,N_12685,N_12650);
and U12803 (N_12803,N_12649,N_12697);
xnor U12804 (N_12804,N_12729,N_12672);
nor U12805 (N_12805,N_12730,N_12605);
xnor U12806 (N_12806,N_12602,N_12624);
nor U12807 (N_12807,N_12653,N_12627);
nand U12808 (N_12808,N_12625,N_12615);
nand U12809 (N_12809,N_12666,N_12621);
nand U12810 (N_12810,N_12634,N_12641);
nand U12811 (N_12811,N_12745,N_12674);
nand U12812 (N_12812,N_12633,N_12726);
xnor U12813 (N_12813,N_12660,N_12717);
nor U12814 (N_12814,N_12720,N_12725);
and U12815 (N_12815,N_12675,N_12696);
xnor U12816 (N_12816,N_12710,N_12603);
or U12817 (N_12817,N_12632,N_12749);
or U12818 (N_12818,N_12680,N_12635);
nor U12819 (N_12819,N_12664,N_12684);
and U12820 (N_12820,N_12731,N_12601);
nand U12821 (N_12821,N_12662,N_12728);
nand U12822 (N_12822,N_12683,N_12628);
nand U12823 (N_12823,N_12744,N_12611);
and U12824 (N_12824,N_12612,N_12661);
nand U12825 (N_12825,N_12716,N_12647);
nor U12826 (N_12826,N_12713,N_12678);
nand U12827 (N_12827,N_12640,N_12685);
and U12828 (N_12828,N_12708,N_12689);
or U12829 (N_12829,N_12670,N_12692);
xnor U12830 (N_12830,N_12672,N_12635);
and U12831 (N_12831,N_12610,N_12614);
xnor U12832 (N_12832,N_12628,N_12747);
nand U12833 (N_12833,N_12710,N_12741);
nand U12834 (N_12834,N_12684,N_12656);
and U12835 (N_12835,N_12654,N_12631);
nor U12836 (N_12836,N_12670,N_12661);
nand U12837 (N_12837,N_12708,N_12680);
nand U12838 (N_12838,N_12740,N_12678);
xor U12839 (N_12839,N_12667,N_12604);
xnor U12840 (N_12840,N_12621,N_12609);
nand U12841 (N_12841,N_12739,N_12720);
nand U12842 (N_12842,N_12633,N_12719);
xor U12843 (N_12843,N_12706,N_12653);
or U12844 (N_12844,N_12699,N_12681);
xnor U12845 (N_12845,N_12649,N_12627);
xnor U12846 (N_12846,N_12693,N_12647);
xnor U12847 (N_12847,N_12697,N_12655);
and U12848 (N_12848,N_12631,N_12650);
nor U12849 (N_12849,N_12747,N_12670);
and U12850 (N_12850,N_12695,N_12712);
or U12851 (N_12851,N_12624,N_12630);
xor U12852 (N_12852,N_12656,N_12610);
or U12853 (N_12853,N_12742,N_12683);
and U12854 (N_12854,N_12647,N_12708);
and U12855 (N_12855,N_12686,N_12667);
and U12856 (N_12856,N_12636,N_12673);
nor U12857 (N_12857,N_12606,N_12651);
nor U12858 (N_12858,N_12642,N_12736);
and U12859 (N_12859,N_12646,N_12651);
nor U12860 (N_12860,N_12603,N_12707);
and U12861 (N_12861,N_12668,N_12681);
and U12862 (N_12862,N_12698,N_12602);
xor U12863 (N_12863,N_12748,N_12714);
and U12864 (N_12864,N_12725,N_12630);
and U12865 (N_12865,N_12617,N_12730);
and U12866 (N_12866,N_12716,N_12669);
xnor U12867 (N_12867,N_12667,N_12642);
xnor U12868 (N_12868,N_12639,N_12619);
or U12869 (N_12869,N_12643,N_12702);
and U12870 (N_12870,N_12652,N_12634);
xor U12871 (N_12871,N_12664,N_12677);
and U12872 (N_12872,N_12671,N_12601);
nor U12873 (N_12873,N_12688,N_12657);
nand U12874 (N_12874,N_12651,N_12699);
and U12875 (N_12875,N_12611,N_12710);
nor U12876 (N_12876,N_12677,N_12722);
and U12877 (N_12877,N_12632,N_12723);
xor U12878 (N_12878,N_12738,N_12637);
nand U12879 (N_12879,N_12699,N_12734);
xor U12880 (N_12880,N_12677,N_12715);
or U12881 (N_12881,N_12727,N_12737);
nor U12882 (N_12882,N_12645,N_12626);
nand U12883 (N_12883,N_12627,N_12672);
nand U12884 (N_12884,N_12693,N_12748);
or U12885 (N_12885,N_12605,N_12721);
nand U12886 (N_12886,N_12732,N_12727);
nand U12887 (N_12887,N_12636,N_12696);
and U12888 (N_12888,N_12738,N_12614);
xnor U12889 (N_12889,N_12636,N_12706);
xor U12890 (N_12890,N_12621,N_12615);
xor U12891 (N_12891,N_12684,N_12732);
nor U12892 (N_12892,N_12726,N_12681);
nor U12893 (N_12893,N_12664,N_12742);
or U12894 (N_12894,N_12625,N_12636);
nand U12895 (N_12895,N_12666,N_12697);
nand U12896 (N_12896,N_12707,N_12696);
or U12897 (N_12897,N_12708,N_12604);
and U12898 (N_12898,N_12698,N_12654);
nor U12899 (N_12899,N_12674,N_12668);
and U12900 (N_12900,N_12763,N_12890);
nor U12901 (N_12901,N_12859,N_12895);
nand U12902 (N_12902,N_12800,N_12847);
or U12903 (N_12903,N_12863,N_12898);
and U12904 (N_12904,N_12878,N_12880);
and U12905 (N_12905,N_12873,N_12784);
or U12906 (N_12906,N_12777,N_12774);
xnor U12907 (N_12907,N_12810,N_12750);
nor U12908 (N_12908,N_12830,N_12808);
or U12909 (N_12909,N_12821,N_12874);
nor U12910 (N_12910,N_12805,N_12845);
and U12911 (N_12911,N_12759,N_12815);
or U12912 (N_12912,N_12846,N_12771);
nand U12913 (N_12913,N_12892,N_12833);
or U12914 (N_12914,N_12770,N_12764);
xnor U12915 (N_12915,N_12836,N_12844);
nand U12916 (N_12916,N_12769,N_12888);
nand U12917 (N_12917,N_12877,N_12813);
nor U12918 (N_12918,N_12850,N_12885);
nand U12919 (N_12919,N_12818,N_12758);
xor U12920 (N_12920,N_12781,N_12835);
or U12921 (N_12921,N_12761,N_12780);
nand U12922 (N_12922,N_12894,N_12793);
nand U12923 (N_12923,N_12820,N_12767);
and U12924 (N_12924,N_12876,N_12779);
nor U12925 (N_12925,N_12866,N_12807);
or U12926 (N_12926,N_12753,N_12837);
nor U12927 (N_12927,N_12790,N_12857);
or U12928 (N_12928,N_12809,N_12766);
xor U12929 (N_12929,N_12797,N_12801);
nand U12930 (N_12930,N_12896,N_12843);
and U12931 (N_12931,N_12756,N_12760);
or U12932 (N_12932,N_12889,N_12788);
and U12933 (N_12933,N_12861,N_12806);
and U12934 (N_12934,N_12804,N_12768);
nand U12935 (N_12935,N_12839,N_12869);
and U12936 (N_12936,N_12754,N_12841);
or U12937 (N_12937,N_12858,N_12852);
and U12938 (N_12938,N_12787,N_12823);
nand U12939 (N_12939,N_12751,N_12799);
nor U12940 (N_12940,N_12849,N_12824);
xor U12941 (N_12941,N_12840,N_12897);
nor U12942 (N_12942,N_12851,N_12776);
xor U12943 (N_12943,N_12848,N_12811);
nor U12944 (N_12944,N_12884,N_12778);
nor U12945 (N_12945,N_12773,N_12838);
nor U12946 (N_12946,N_12752,N_12831);
and U12947 (N_12947,N_12755,N_12783);
nor U12948 (N_12948,N_12772,N_12855);
and U12949 (N_12949,N_12817,N_12775);
nor U12950 (N_12950,N_12867,N_12757);
nor U12951 (N_12951,N_12795,N_12762);
xnor U12952 (N_12952,N_12862,N_12872);
and U12953 (N_12953,N_12881,N_12853);
nor U12954 (N_12954,N_12825,N_12796);
xor U12955 (N_12955,N_12803,N_12802);
nor U12956 (N_12956,N_12883,N_12832);
or U12957 (N_12957,N_12827,N_12828);
nor U12958 (N_12958,N_12812,N_12886);
and U12959 (N_12959,N_12789,N_12826);
nand U12960 (N_12960,N_12834,N_12882);
xor U12961 (N_12961,N_12854,N_12856);
xor U12962 (N_12962,N_12893,N_12816);
and U12963 (N_12963,N_12814,N_12868);
xnor U12964 (N_12964,N_12794,N_12842);
nand U12965 (N_12965,N_12792,N_12765);
xnor U12966 (N_12966,N_12870,N_12875);
and U12967 (N_12967,N_12782,N_12829);
nand U12968 (N_12968,N_12871,N_12879);
or U12969 (N_12969,N_12822,N_12865);
xor U12970 (N_12970,N_12887,N_12791);
or U12971 (N_12971,N_12798,N_12860);
or U12972 (N_12972,N_12785,N_12819);
and U12973 (N_12973,N_12786,N_12899);
or U12974 (N_12974,N_12864,N_12891);
nor U12975 (N_12975,N_12818,N_12763);
and U12976 (N_12976,N_12880,N_12812);
and U12977 (N_12977,N_12825,N_12828);
and U12978 (N_12978,N_12828,N_12837);
xnor U12979 (N_12979,N_12836,N_12824);
or U12980 (N_12980,N_12887,N_12761);
nand U12981 (N_12981,N_12845,N_12752);
xnor U12982 (N_12982,N_12892,N_12862);
and U12983 (N_12983,N_12840,N_12757);
nand U12984 (N_12984,N_12873,N_12777);
or U12985 (N_12985,N_12882,N_12807);
xor U12986 (N_12986,N_12831,N_12761);
or U12987 (N_12987,N_12766,N_12865);
xor U12988 (N_12988,N_12859,N_12783);
and U12989 (N_12989,N_12827,N_12837);
nor U12990 (N_12990,N_12799,N_12884);
and U12991 (N_12991,N_12860,N_12880);
xor U12992 (N_12992,N_12756,N_12847);
xnor U12993 (N_12993,N_12774,N_12820);
nand U12994 (N_12994,N_12835,N_12850);
or U12995 (N_12995,N_12848,N_12840);
and U12996 (N_12996,N_12824,N_12793);
nand U12997 (N_12997,N_12872,N_12785);
nand U12998 (N_12998,N_12806,N_12754);
nand U12999 (N_12999,N_12812,N_12891);
nand U13000 (N_13000,N_12894,N_12848);
or U13001 (N_13001,N_12800,N_12842);
xor U13002 (N_13002,N_12892,N_12807);
xor U13003 (N_13003,N_12817,N_12779);
xor U13004 (N_13004,N_12881,N_12879);
nor U13005 (N_13005,N_12812,N_12871);
nor U13006 (N_13006,N_12753,N_12806);
nand U13007 (N_13007,N_12778,N_12860);
and U13008 (N_13008,N_12850,N_12883);
nand U13009 (N_13009,N_12841,N_12879);
xor U13010 (N_13010,N_12857,N_12796);
or U13011 (N_13011,N_12771,N_12894);
nor U13012 (N_13012,N_12876,N_12853);
xor U13013 (N_13013,N_12830,N_12800);
nand U13014 (N_13014,N_12812,N_12895);
and U13015 (N_13015,N_12871,N_12839);
nor U13016 (N_13016,N_12807,N_12769);
and U13017 (N_13017,N_12849,N_12783);
nand U13018 (N_13018,N_12776,N_12773);
or U13019 (N_13019,N_12775,N_12784);
nand U13020 (N_13020,N_12864,N_12860);
or U13021 (N_13021,N_12850,N_12846);
xor U13022 (N_13022,N_12790,N_12884);
and U13023 (N_13023,N_12847,N_12792);
or U13024 (N_13024,N_12790,N_12892);
and U13025 (N_13025,N_12803,N_12835);
nor U13026 (N_13026,N_12877,N_12782);
or U13027 (N_13027,N_12807,N_12857);
nor U13028 (N_13028,N_12841,N_12835);
xor U13029 (N_13029,N_12881,N_12787);
and U13030 (N_13030,N_12793,N_12763);
or U13031 (N_13031,N_12857,N_12770);
and U13032 (N_13032,N_12856,N_12779);
nand U13033 (N_13033,N_12759,N_12783);
or U13034 (N_13034,N_12857,N_12795);
and U13035 (N_13035,N_12897,N_12855);
and U13036 (N_13036,N_12884,N_12864);
and U13037 (N_13037,N_12874,N_12826);
nor U13038 (N_13038,N_12854,N_12840);
nor U13039 (N_13039,N_12755,N_12841);
nor U13040 (N_13040,N_12884,N_12870);
and U13041 (N_13041,N_12769,N_12858);
nor U13042 (N_13042,N_12786,N_12784);
xnor U13043 (N_13043,N_12750,N_12807);
or U13044 (N_13044,N_12862,N_12807);
or U13045 (N_13045,N_12808,N_12855);
nand U13046 (N_13046,N_12808,N_12793);
xnor U13047 (N_13047,N_12866,N_12842);
and U13048 (N_13048,N_12823,N_12896);
and U13049 (N_13049,N_12882,N_12890);
nand U13050 (N_13050,N_13031,N_12910);
nand U13051 (N_13051,N_12925,N_12979);
or U13052 (N_13052,N_13048,N_13038);
xnor U13053 (N_13053,N_12937,N_12920);
or U13054 (N_13054,N_13028,N_13019);
or U13055 (N_13055,N_13015,N_12904);
xnor U13056 (N_13056,N_12997,N_12977);
or U13057 (N_13057,N_13035,N_12950);
or U13058 (N_13058,N_13008,N_12981);
and U13059 (N_13059,N_12933,N_12913);
or U13060 (N_13060,N_12941,N_12916);
xnor U13061 (N_13061,N_12949,N_12918);
nand U13062 (N_13062,N_12987,N_13039);
and U13063 (N_13063,N_13002,N_13012);
nor U13064 (N_13064,N_12984,N_12953);
nand U13065 (N_13065,N_12915,N_12988);
and U13066 (N_13066,N_12936,N_12989);
and U13067 (N_13067,N_13042,N_12928);
nand U13068 (N_13068,N_12943,N_12994);
or U13069 (N_13069,N_12959,N_12951);
nand U13070 (N_13070,N_12978,N_12954);
xnor U13071 (N_13071,N_12935,N_12992);
nor U13072 (N_13072,N_12946,N_12964);
xor U13073 (N_13073,N_12995,N_12922);
or U13074 (N_13074,N_12945,N_12930);
or U13075 (N_13075,N_12993,N_12985);
and U13076 (N_13076,N_12944,N_12963);
nor U13077 (N_13077,N_12968,N_12958);
nor U13078 (N_13078,N_13026,N_12932);
nand U13079 (N_13079,N_12952,N_13024);
xnor U13080 (N_13080,N_12905,N_13000);
nand U13081 (N_13081,N_12940,N_12948);
and U13082 (N_13082,N_13021,N_12955);
and U13083 (N_13083,N_13047,N_12926);
xnor U13084 (N_13084,N_13005,N_13036);
and U13085 (N_13085,N_12934,N_13040);
and U13086 (N_13086,N_12911,N_13044);
and U13087 (N_13087,N_13020,N_12919);
nand U13088 (N_13088,N_12900,N_12983);
and U13089 (N_13089,N_12942,N_13007);
nand U13090 (N_13090,N_12996,N_13037);
nor U13091 (N_13091,N_12957,N_12980);
or U13092 (N_13092,N_13009,N_13014);
nand U13093 (N_13093,N_13004,N_13016);
nand U13094 (N_13094,N_12931,N_13011);
or U13095 (N_13095,N_12976,N_13025);
xnor U13096 (N_13096,N_12927,N_13029);
nand U13097 (N_13097,N_13030,N_13001);
and U13098 (N_13098,N_12917,N_12960);
or U13099 (N_13099,N_13034,N_13023);
and U13100 (N_13100,N_13010,N_12906);
and U13101 (N_13101,N_12901,N_12974);
nor U13102 (N_13102,N_13046,N_12956);
and U13103 (N_13103,N_12939,N_12986);
and U13104 (N_13104,N_12914,N_13033);
nor U13105 (N_13105,N_12982,N_12998);
and U13106 (N_13106,N_13017,N_12975);
xnor U13107 (N_13107,N_13032,N_12907);
nor U13108 (N_13108,N_12966,N_13045);
xor U13109 (N_13109,N_12970,N_12967);
xnor U13110 (N_13110,N_12961,N_12923);
nand U13111 (N_13111,N_13043,N_12991);
and U13112 (N_13112,N_12912,N_12999);
and U13113 (N_13113,N_12903,N_13041);
and U13114 (N_13114,N_13018,N_13006);
nand U13115 (N_13115,N_12971,N_13003);
xnor U13116 (N_13116,N_12921,N_12924);
and U13117 (N_13117,N_12938,N_12965);
and U13118 (N_13118,N_12969,N_13013);
and U13119 (N_13119,N_12908,N_12909);
nor U13120 (N_13120,N_12972,N_12947);
nand U13121 (N_13121,N_12973,N_12990);
or U13122 (N_13122,N_13022,N_13027);
nand U13123 (N_13123,N_12902,N_13049);
and U13124 (N_13124,N_12962,N_12929);
and U13125 (N_13125,N_12993,N_13041);
nand U13126 (N_13126,N_13033,N_12993);
xor U13127 (N_13127,N_12986,N_12991);
or U13128 (N_13128,N_12970,N_12960);
or U13129 (N_13129,N_12963,N_13005);
xnor U13130 (N_13130,N_12923,N_13005);
nor U13131 (N_13131,N_13027,N_12951);
and U13132 (N_13132,N_12939,N_12924);
nand U13133 (N_13133,N_13037,N_13017);
nand U13134 (N_13134,N_12990,N_13023);
nor U13135 (N_13135,N_13044,N_12986);
and U13136 (N_13136,N_13044,N_12994);
nor U13137 (N_13137,N_13035,N_12902);
or U13138 (N_13138,N_12939,N_12910);
or U13139 (N_13139,N_13032,N_13025);
or U13140 (N_13140,N_13044,N_13023);
and U13141 (N_13141,N_13036,N_13041);
and U13142 (N_13142,N_12939,N_13041);
nor U13143 (N_13143,N_12911,N_13006);
xor U13144 (N_13144,N_12919,N_12910);
nor U13145 (N_13145,N_12991,N_13033);
nand U13146 (N_13146,N_12976,N_12923);
nor U13147 (N_13147,N_12995,N_13006);
and U13148 (N_13148,N_12901,N_12984);
nor U13149 (N_13149,N_12930,N_13000);
and U13150 (N_13150,N_12982,N_12916);
and U13151 (N_13151,N_12923,N_12934);
nor U13152 (N_13152,N_12927,N_12971);
and U13153 (N_13153,N_13033,N_12998);
nand U13154 (N_13154,N_13009,N_13030);
xnor U13155 (N_13155,N_13046,N_12935);
and U13156 (N_13156,N_12929,N_13048);
nor U13157 (N_13157,N_13047,N_13032);
nor U13158 (N_13158,N_12967,N_13042);
nor U13159 (N_13159,N_13042,N_12996);
or U13160 (N_13160,N_12968,N_12944);
nand U13161 (N_13161,N_12930,N_13014);
nor U13162 (N_13162,N_12934,N_12979);
nor U13163 (N_13163,N_13016,N_12912);
nor U13164 (N_13164,N_13029,N_13040);
or U13165 (N_13165,N_12921,N_13018);
nand U13166 (N_13166,N_12980,N_13022);
and U13167 (N_13167,N_12925,N_12950);
nand U13168 (N_13168,N_12954,N_12920);
or U13169 (N_13169,N_12998,N_13013);
or U13170 (N_13170,N_12927,N_13021);
nand U13171 (N_13171,N_13038,N_12903);
xor U13172 (N_13172,N_12942,N_13032);
xor U13173 (N_13173,N_13030,N_12902);
and U13174 (N_13174,N_12904,N_13004);
nand U13175 (N_13175,N_13033,N_13025);
or U13176 (N_13176,N_12949,N_13003);
and U13177 (N_13177,N_12962,N_12918);
nand U13178 (N_13178,N_12924,N_12946);
nor U13179 (N_13179,N_12917,N_13040);
nor U13180 (N_13180,N_12917,N_12956);
and U13181 (N_13181,N_13014,N_12987);
nor U13182 (N_13182,N_12955,N_12965);
nor U13183 (N_13183,N_12923,N_12987);
nor U13184 (N_13184,N_13039,N_12978);
and U13185 (N_13185,N_12966,N_13048);
nand U13186 (N_13186,N_12922,N_12919);
nand U13187 (N_13187,N_12986,N_12970);
nor U13188 (N_13188,N_12983,N_12905);
and U13189 (N_13189,N_13014,N_12927);
nor U13190 (N_13190,N_12958,N_12979);
or U13191 (N_13191,N_12900,N_12960);
nand U13192 (N_13192,N_13039,N_12965);
and U13193 (N_13193,N_12986,N_13029);
nor U13194 (N_13194,N_12929,N_12921);
and U13195 (N_13195,N_12935,N_12920);
xnor U13196 (N_13196,N_12998,N_12968);
nand U13197 (N_13197,N_12962,N_13008);
xor U13198 (N_13198,N_12922,N_12914);
nand U13199 (N_13199,N_12940,N_13032);
and U13200 (N_13200,N_13162,N_13079);
nand U13201 (N_13201,N_13053,N_13176);
nand U13202 (N_13202,N_13075,N_13094);
nand U13203 (N_13203,N_13187,N_13195);
xor U13204 (N_13204,N_13123,N_13190);
or U13205 (N_13205,N_13168,N_13117);
xnor U13206 (N_13206,N_13148,N_13097);
and U13207 (N_13207,N_13108,N_13183);
nand U13208 (N_13208,N_13104,N_13181);
nand U13209 (N_13209,N_13091,N_13069);
or U13210 (N_13210,N_13198,N_13055);
nand U13211 (N_13211,N_13166,N_13144);
nor U13212 (N_13212,N_13119,N_13184);
nor U13213 (N_13213,N_13150,N_13078);
or U13214 (N_13214,N_13059,N_13131);
nor U13215 (N_13215,N_13191,N_13090);
nor U13216 (N_13216,N_13073,N_13086);
and U13217 (N_13217,N_13118,N_13160);
or U13218 (N_13218,N_13095,N_13057);
nor U13219 (N_13219,N_13120,N_13129);
nor U13220 (N_13220,N_13066,N_13146);
or U13221 (N_13221,N_13138,N_13177);
or U13222 (N_13222,N_13115,N_13098);
xor U13223 (N_13223,N_13064,N_13058);
nand U13224 (N_13224,N_13180,N_13155);
xnor U13225 (N_13225,N_13199,N_13196);
or U13226 (N_13226,N_13134,N_13193);
nand U13227 (N_13227,N_13121,N_13056);
nand U13228 (N_13228,N_13122,N_13145);
or U13229 (N_13229,N_13100,N_13070);
nor U13230 (N_13230,N_13060,N_13151);
nor U13231 (N_13231,N_13105,N_13082);
nand U13232 (N_13232,N_13141,N_13163);
and U13233 (N_13233,N_13167,N_13071);
nand U13234 (N_13234,N_13096,N_13113);
nand U13235 (N_13235,N_13142,N_13172);
xor U13236 (N_13236,N_13174,N_13154);
xnor U13237 (N_13237,N_13067,N_13158);
xnor U13238 (N_13238,N_13085,N_13083);
nor U13239 (N_13239,N_13197,N_13186);
nor U13240 (N_13240,N_13106,N_13099);
nand U13241 (N_13241,N_13124,N_13076);
nor U13242 (N_13242,N_13107,N_13194);
and U13243 (N_13243,N_13084,N_13132);
and U13244 (N_13244,N_13192,N_13152);
xnor U13245 (N_13245,N_13170,N_13110);
and U13246 (N_13246,N_13156,N_13112);
nor U13247 (N_13247,N_13111,N_13114);
nor U13248 (N_13248,N_13101,N_13173);
nor U13249 (N_13249,N_13130,N_13125);
xnor U13250 (N_13250,N_13188,N_13128);
or U13251 (N_13251,N_13102,N_13092);
nand U13252 (N_13252,N_13087,N_13140);
xnor U13253 (N_13253,N_13093,N_13103);
and U13254 (N_13254,N_13153,N_13081);
or U13255 (N_13255,N_13161,N_13147);
and U13256 (N_13256,N_13109,N_13149);
xor U13257 (N_13257,N_13164,N_13143);
nor U13258 (N_13258,N_13072,N_13189);
nor U13259 (N_13259,N_13068,N_13182);
or U13260 (N_13260,N_13127,N_13077);
or U13261 (N_13261,N_13126,N_13054);
or U13262 (N_13262,N_13175,N_13089);
xor U13263 (N_13263,N_13157,N_13050);
xor U13264 (N_13264,N_13052,N_13169);
nand U13265 (N_13265,N_13116,N_13165);
or U13266 (N_13266,N_13062,N_13051);
nor U13267 (N_13267,N_13185,N_13080);
and U13268 (N_13268,N_13171,N_13135);
xnor U13269 (N_13269,N_13061,N_13178);
nand U13270 (N_13270,N_13137,N_13139);
xor U13271 (N_13271,N_13088,N_13133);
nand U13272 (N_13272,N_13065,N_13159);
and U13273 (N_13273,N_13063,N_13074);
or U13274 (N_13274,N_13136,N_13179);
xor U13275 (N_13275,N_13091,N_13181);
or U13276 (N_13276,N_13059,N_13166);
and U13277 (N_13277,N_13131,N_13100);
or U13278 (N_13278,N_13163,N_13109);
nand U13279 (N_13279,N_13059,N_13098);
and U13280 (N_13280,N_13071,N_13191);
nor U13281 (N_13281,N_13085,N_13082);
and U13282 (N_13282,N_13131,N_13187);
nand U13283 (N_13283,N_13165,N_13130);
nand U13284 (N_13284,N_13150,N_13148);
or U13285 (N_13285,N_13163,N_13098);
and U13286 (N_13286,N_13087,N_13078);
nand U13287 (N_13287,N_13197,N_13065);
or U13288 (N_13288,N_13094,N_13188);
nor U13289 (N_13289,N_13143,N_13051);
nor U13290 (N_13290,N_13131,N_13078);
or U13291 (N_13291,N_13188,N_13118);
or U13292 (N_13292,N_13130,N_13187);
or U13293 (N_13293,N_13108,N_13144);
and U13294 (N_13294,N_13154,N_13146);
nand U13295 (N_13295,N_13090,N_13068);
nand U13296 (N_13296,N_13078,N_13135);
xor U13297 (N_13297,N_13157,N_13119);
xnor U13298 (N_13298,N_13136,N_13161);
or U13299 (N_13299,N_13092,N_13176);
or U13300 (N_13300,N_13181,N_13136);
nor U13301 (N_13301,N_13144,N_13167);
nand U13302 (N_13302,N_13167,N_13198);
nand U13303 (N_13303,N_13084,N_13180);
nand U13304 (N_13304,N_13107,N_13126);
xnor U13305 (N_13305,N_13088,N_13178);
nand U13306 (N_13306,N_13052,N_13142);
xor U13307 (N_13307,N_13144,N_13075);
and U13308 (N_13308,N_13171,N_13172);
nor U13309 (N_13309,N_13102,N_13132);
or U13310 (N_13310,N_13199,N_13183);
nand U13311 (N_13311,N_13159,N_13151);
or U13312 (N_13312,N_13167,N_13146);
or U13313 (N_13313,N_13114,N_13067);
xor U13314 (N_13314,N_13194,N_13119);
and U13315 (N_13315,N_13163,N_13190);
nand U13316 (N_13316,N_13164,N_13148);
xnor U13317 (N_13317,N_13113,N_13165);
or U13318 (N_13318,N_13121,N_13153);
and U13319 (N_13319,N_13166,N_13115);
or U13320 (N_13320,N_13179,N_13080);
and U13321 (N_13321,N_13185,N_13157);
xor U13322 (N_13322,N_13161,N_13191);
nor U13323 (N_13323,N_13079,N_13170);
or U13324 (N_13324,N_13183,N_13103);
and U13325 (N_13325,N_13111,N_13051);
xor U13326 (N_13326,N_13149,N_13169);
nand U13327 (N_13327,N_13166,N_13156);
nor U13328 (N_13328,N_13133,N_13159);
xor U13329 (N_13329,N_13107,N_13162);
and U13330 (N_13330,N_13099,N_13129);
nand U13331 (N_13331,N_13194,N_13085);
or U13332 (N_13332,N_13099,N_13083);
and U13333 (N_13333,N_13104,N_13133);
nand U13334 (N_13334,N_13197,N_13093);
and U13335 (N_13335,N_13096,N_13085);
or U13336 (N_13336,N_13127,N_13197);
or U13337 (N_13337,N_13066,N_13109);
nand U13338 (N_13338,N_13098,N_13147);
and U13339 (N_13339,N_13080,N_13138);
or U13340 (N_13340,N_13114,N_13093);
nand U13341 (N_13341,N_13193,N_13099);
and U13342 (N_13342,N_13055,N_13194);
and U13343 (N_13343,N_13075,N_13068);
xnor U13344 (N_13344,N_13052,N_13192);
and U13345 (N_13345,N_13116,N_13129);
nor U13346 (N_13346,N_13161,N_13176);
and U13347 (N_13347,N_13088,N_13083);
nor U13348 (N_13348,N_13064,N_13148);
nand U13349 (N_13349,N_13068,N_13097);
xnor U13350 (N_13350,N_13277,N_13337);
xnor U13351 (N_13351,N_13329,N_13333);
nor U13352 (N_13352,N_13207,N_13324);
xnor U13353 (N_13353,N_13328,N_13260);
nor U13354 (N_13354,N_13244,N_13230);
nand U13355 (N_13355,N_13331,N_13229);
xnor U13356 (N_13356,N_13349,N_13275);
nand U13357 (N_13357,N_13272,N_13286);
nor U13358 (N_13358,N_13208,N_13344);
xnor U13359 (N_13359,N_13338,N_13254);
nand U13360 (N_13360,N_13334,N_13316);
nand U13361 (N_13361,N_13228,N_13330);
nand U13362 (N_13362,N_13278,N_13210);
nor U13363 (N_13363,N_13318,N_13323);
xor U13364 (N_13364,N_13256,N_13282);
nor U13365 (N_13365,N_13243,N_13332);
nand U13366 (N_13366,N_13341,N_13217);
xor U13367 (N_13367,N_13293,N_13250);
nand U13368 (N_13368,N_13271,N_13302);
nand U13369 (N_13369,N_13326,N_13266);
and U13370 (N_13370,N_13346,N_13301);
nor U13371 (N_13371,N_13236,N_13240);
nand U13372 (N_13372,N_13313,N_13252);
xor U13373 (N_13373,N_13213,N_13311);
nand U13374 (N_13374,N_13245,N_13327);
xnor U13375 (N_13375,N_13264,N_13206);
nand U13376 (N_13376,N_13307,N_13291);
nand U13377 (N_13377,N_13283,N_13297);
and U13378 (N_13378,N_13226,N_13200);
nor U13379 (N_13379,N_13241,N_13265);
nor U13380 (N_13380,N_13267,N_13274);
or U13381 (N_13381,N_13246,N_13273);
nor U13382 (N_13382,N_13285,N_13218);
or U13383 (N_13383,N_13221,N_13336);
or U13384 (N_13384,N_13220,N_13232);
xor U13385 (N_13385,N_13234,N_13314);
xor U13386 (N_13386,N_13295,N_13251);
nand U13387 (N_13387,N_13342,N_13340);
and U13388 (N_13388,N_13233,N_13319);
or U13389 (N_13389,N_13255,N_13345);
nand U13390 (N_13390,N_13321,N_13322);
or U13391 (N_13391,N_13253,N_13262);
or U13392 (N_13392,N_13284,N_13270);
nor U13393 (N_13393,N_13247,N_13259);
or U13394 (N_13394,N_13276,N_13203);
or U13395 (N_13395,N_13315,N_13249);
or U13396 (N_13396,N_13202,N_13225);
and U13397 (N_13397,N_13231,N_13237);
or U13398 (N_13398,N_13325,N_13239);
and U13399 (N_13399,N_13235,N_13205);
xor U13400 (N_13400,N_13222,N_13308);
and U13401 (N_13401,N_13312,N_13339);
xor U13402 (N_13402,N_13223,N_13299);
and U13403 (N_13403,N_13347,N_13201);
nand U13404 (N_13404,N_13219,N_13268);
xnor U13405 (N_13405,N_13258,N_13257);
or U13406 (N_13406,N_13261,N_13227);
xnor U13407 (N_13407,N_13279,N_13238);
and U13408 (N_13408,N_13306,N_13317);
xor U13409 (N_13409,N_13305,N_13320);
and U13410 (N_13410,N_13214,N_13289);
nor U13411 (N_13411,N_13292,N_13224);
or U13412 (N_13412,N_13248,N_13216);
or U13413 (N_13413,N_13290,N_13204);
nand U13414 (N_13414,N_13215,N_13303);
xor U13415 (N_13415,N_13298,N_13263);
nor U13416 (N_13416,N_13296,N_13287);
and U13417 (N_13417,N_13242,N_13269);
nor U13418 (N_13418,N_13310,N_13211);
and U13419 (N_13419,N_13212,N_13209);
nor U13420 (N_13420,N_13300,N_13288);
nor U13421 (N_13421,N_13309,N_13281);
nor U13422 (N_13422,N_13294,N_13343);
nand U13423 (N_13423,N_13280,N_13348);
and U13424 (N_13424,N_13304,N_13335);
and U13425 (N_13425,N_13253,N_13217);
nand U13426 (N_13426,N_13303,N_13321);
and U13427 (N_13427,N_13323,N_13295);
or U13428 (N_13428,N_13262,N_13233);
nand U13429 (N_13429,N_13253,N_13342);
or U13430 (N_13430,N_13337,N_13241);
nand U13431 (N_13431,N_13227,N_13299);
nor U13432 (N_13432,N_13223,N_13304);
nand U13433 (N_13433,N_13290,N_13233);
xor U13434 (N_13434,N_13206,N_13284);
xor U13435 (N_13435,N_13320,N_13260);
nand U13436 (N_13436,N_13253,N_13277);
nand U13437 (N_13437,N_13280,N_13247);
nand U13438 (N_13438,N_13290,N_13307);
or U13439 (N_13439,N_13217,N_13301);
or U13440 (N_13440,N_13240,N_13204);
xor U13441 (N_13441,N_13204,N_13226);
nor U13442 (N_13442,N_13241,N_13212);
and U13443 (N_13443,N_13232,N_13269);
and U13444 (N_13444,N_13300,N_13233);
and U13445 (N_13445,N_13278,N_13221);
nand U13446 (N_13446,N_13209,N_13299);
nor U13447 (N_13447,N_13242,N_13276);
nand U13448 (N_13448,N_13203,N_13247);
and U13449 (N_13449,N_13253,N_13292);
xor U13450 (N_13450,N_13226,N_13237);
or U13451 (N_13451,N_13227,N_13326);
nor U13452 (N_13452,N_13242,N_13340);
or U13453 (N_13453,N_13285,N_13211);
and U13454 (N_13454,N_13200,N_13209);
or U13455 (N_13455,N_13300,N_13315);
and U13456 (N_13456,N_13310,N_13263);
or U13457 (N_13457,N_13280,N_13324);
or U13458 (N_13458,N_13265,N_13229);
nand U13459 (N_13459,N_13261,N_13248);
or U13460 (N_13460,N_13269,N_13335);
or U13461 (N_13461,N_13336,N_13273);
nand U13462 (N_13462,N_13308,N_13200);
and U13463 (N_13463,N_13297,N_13321);
nand U13464 (N_13464,N_13205,N_13211);
or U13465 (N_13465,N_13335,N_13320);
nor U13466 (N_13466,N_13334,N_13242);
xnor U13467 (N_13467,N_13259,N_13307);
nand U13468 (N_13468,N_13332,N_13293);
or U13469 (N_13469,N_13305,N_13253);
and U13470 (N_13470,N_13230,N_13218);
or U13471 (N_13471,N_13330,N_13225);
and U13472 (N_13472,N_13281,N_13307);
xnor U13473 (N_13473,N_13241,N_13322);
and U13474 (N_13474,N_13318,N_13334);
or U13475 (N_13475,N_13237,N_13312);
and U13476 (N_13476,N_13224,N_13268);
nor U13477 (N_13477,N_13269,N_13206);
xnor U13478 (N_13478,N_13270,N_13244);
xnor U13479 (N_13479,N_13277,N_13205);
xnor U13480 (N_13480,N_13333,N_13304);
nand U13481 (N_13481,N_13204,N_13284);
xor U13482 (N_13482,N_13208,N_13285);
and U13483 (N_13483,N_13257,N_13241);
xor U13484 (N_13484,N_13213,N_13325);
nand U13485 (N_13485,N_13341,N_13254);
xor U13486 (N_13486,N_13201,N_13218);
nand U13487 (N_13487,N_13327,N_13296);
nor U13488 (N_13488,N_13207,N_13222);
nand U13489 (N_13489,N_13256,N_13228);
nand U13490 (N_13490,N_13318,N_13335);
nor U13491 (N_13491,N_13253,N_13334);
nor U13492 (N_13492,N_13286,N_13331);
xor U13493 (N_13493,N_13221,N_13266);
or U13494 (N_13494,N_13203,N_13222);
nand U13495 (N_13495,N_13279,N_13209);
or U13496 (N_13496,N_13244,N_13323);
and U13497 (N_13497,N_13337,N_13336);
and U13498 (N_13498,N_13274,N_13233);
nand U13499 (N_13499,N_13211,N_13305);
xnor U13500 (N_13500,N_13403,N_13441);
nor U13501 (N_13501,N_13442,N_13458);
and U13502 (N_13502,N_13430,N_13405);
or U13503 (N_13503,N_13409,N_13432);
or U13504 (N_13504,N_13480,N_13490);
and U13505 (N_13505,N_13376,N_13447);
xor U13506 (N_13506,N_13387,N_13357);
xnor U13507 (N_13507,N_13419,N_13439);
nand U13508 (N_13508,N_13494,N_13418);
nand U13509 (N_13509,N_13408,N_13425);
xor U13510 (N_13510,N_13412,N_13469);
and U13511 (N_13511,N_13359,N_13429);
or U13512 (N_13512,N_13371,N_13466);
or U13513 (N_13513,N_13486,N_13406);
xnor U13514 (N_13514,N_13495,N_13421);
nand U13515 (N_13515,N_13400,N_13386);
or U13516 (N_13516,N_13437,N_13448);
or U13517 (N_13517,N_13476,N_13451);
or U13518 (N_13518,N_13392,N_13380);
nand U13519 (N_13519,N_13401,N_13496);
or U13520 (N_13520,N_13453,N_13389);
and U13521 (N_13521,N_13351,N_13384);
and U13522 (N_13522,N_13396,N_13354);
nand U13523 (N_13523,N_13461,N_13365);
and U13524 (N_13524,N_13378,N_13381);
and U13525 (N_13525,N_13445,N_13368);
nor U13526 (N_13526,N_13467,N_13353);
nor U13527 (N_13527,N_13393,N_13352);
nand U13528 (N_13528,N_13350,N_13424);
or U13529 (N_13529,N_13360,N_13383);
and U13530 (N_13530,N_13414,N_13355);
xnor U13531 (N_13531,N_13413,N_13420);
and U13532 (N_13532,N_13394,N_13431);
nor U13533 (N_13533,N_13417,N_13438);
nor U13534 (N_13534,N_13450,N_13398);
and U13535 (N_13535,N_13460,N_13426);
and U13536 (N_13536,N_13385,N_13471);
or U13537 (N_13537,N_13499,N_13475);
and U13538 (N_13538,N_13455,N_13440);
or U13539 (N_13539,N_13372,N_13456);
nor U13540 (N_13540,N_13410,N_13452);
and U13541 (N_13541,N_13464,N_13423);
or U13542 (N_13542,N_13367,N_13358);
nand U13543 (N_13543,N_13375,N_13364);
nor U13544 (N_13544,N_13498,N_13362);
nor U13545 (N_13545,N_13479,N_13474);
or U13546 (N_13546,N_13465,N_13433);
or U13547 (N_13547,N_13434,N_13404);
nand U13548 (N_13548,N_13370,N_13428);
xor U13549 (N_13549,N_13492,N_13415);
xor U13550 (N_13550,N_13435,N_13399);
and U13551 (N_13551,N_13459,N_13457);
nand U13552 (N_13552,N_13373,N_13366);
nand U13553 (N_13553,N_13407,N_13468);
nor U13554 (N_13554,N_13497,N_13454);
nand U13555 (N_13555,N_13374,N_13377);
nor U13556 (N_13556,N_13391,N_13487);
or U13557 (N_13557,N_13379,N_13436);
nand U13558 (N_13558,N_13397,N_13462);
nor U13559 (N_13559,N_13443,N_13422);
xor U13560 (N_13560,N_13491,N_13390);
nor U13561 (N_13561,N_13473,N_13488);
nor U13562 (N_13562,N_13369,N_13477);
nand U13563 (N_13563,N_13481,N_13402);
nor U13564 (N_13564,N_13427,N_13416);
and U13565 (N_13565,N_13485,N_13483);
and U13566 (N_13566,N_13388,N_13382);
or U13567 (N_13567,N_13482,N_13395);
nor U13568 (N_13568,N_13361,N_13446);
xnor U13569 (N_13569,N_13489,N_13493);
or U13570 (N_13570,N_13363,N_13449);
or U13571 (N_13571,N_13444,N_13463);
or U13572 (N_13572,N_13484,N_13356);
and U13573 (N_13573,N_13470,N_13472);
xnor U13574 (N_13574,N_13411,N_13478);
nor U13575 (N_13575,N_13382,N_13451);
nand U13576 (N_13576,N_13430,N_13437);
or U13577 (N_13577,N_13491,N_13473);
nand U13578 (N_13578,N_13399,N_13487);
nand U13579 (N_13579,N_13410,N_13471);
xor U13580 (N_13580,N_13400,N_13447);
or U13581 (N_13581,N_13444,N_13475);
nand U13582 (N_13582,N_13486,N_13391);
nand U13583 (N_13583,N_13403,N_13351);
nor U13584 (N_13584,N_13362,N_13383);
nor U13585 (N_13585,N_13385,N_13419);
or U13586 (N_13586,N_13415,N_13389);
nand U13587 (N_13587,N_13466,N_13402);
nor U13588 (N_13588,N_13387,N_13450);
or U13589 (N_13589,N_13448,N_13454);
or U13590 (N_13590,N_13484,N_13410);
and U13591 (N_13591,N_13484,N_13411);
and U13592 (N_13592,N_13446,N_13355);
or U13593 (N_13593,N_13392,N_13418);
and U13594 (N_13594,N_13496,N_13366);
nor U13595 (N_13595,N_13494,N_13363);
nand U13596 (N_13596,N_13432,N_13356);
nand U13597 (N_13597,N_13429,N_13360);
nand U13598 (N_13598,N_13387,N_13358);
nor U13599 (N_13599,N_13390,N_13470);
and U13600 (N_13600,N_13471,N_13445);
nand U13601 (N_13601,N_13425,N_13393);
xnor U13602 (N_13602,N_13367,N_13475);
nand U13603 (N_13603,N_13482,N_13358);
and U13604 (N_13604,N_13453,N_13442);
nor U13605 (N_13605,N_13366,N_13372);
xnor U13606 (N_13606,N_13419,N_13427);
xor U13607 (N_13607,N_13463,N_13452);
nand U13608 (N_13608,N_13488,N_13350);
xnor U13609 (N_13609,N_13382,N_13406);
xor U13610 (N_13610,N_13355,N_13442);
nand U13611 (N_13611,N_13428,N_13427);
nand U13612 (N_13612,N_13484,N_13442);
nor U13613 (N_13613,N_13449,N_13436);
nor U13614 (N_13614,N_13430,N_13414);
nand U13615 (N_13615,N_13489,N_13357);
or U13616 (N_13616,N_13374,N_13487);
nand U13617 (N_13617,N_13465,N_13387);
nand U13618 (N_13618,N_13362,N_13393);
nor U13619 (N_13619,N_13359,N_13440);
nand U13620 (N_13620,N_13387,N_13435);
or U13621 (N_13621,N_13463,N_13476);
and U13622 (N_13622,N_13406,N_13361);
nor U13623 (N_13623,N_13468,N_13422);
nand U13624 (N_13624,N_13426,N_13456);
xor U13625 (N_13625,N_13488,N_13392);
nand U13626 (N_13626,N_13357,N_13486);
and U13627 (N_13627,N_13493,N_13407);
nand U13628 (N_13628,N_13432,N_13350);
nand U13629 (N_13629,N_13404,N_13428);
or U13630 (N_13630,N_13370,N_13395);
xnor U13631 (N_13631,N_13497,N_13351);
xor U13632 (N_13632,N_13445,N_13392);
nor U13633 (N_13633,N_13462,N_13464);
or U13634 (N_13634,N_13406,N_13366);
nor U13635 (N_13635,N_13460,N_13398);
nor U13636 (N_13636,N_13353,N_13370);
nor U13637 (N_13637,N_13472,N_13458);
xor U13638 (N_13638,N_13373,N_13432);
nor U13639 (N_13639,N_13373,N_13389);
nor U13640 (N_13640,N_13489,N_13407);
or U13641 (N_13641,N_13472,N_13466);
nor U13642 (N_13642,N_13436,N_13396);
nor U13643 (N_13643,N_13460,N_13467);
nand U13644 (N_13644,N_13373,N_13398);
nor U13645 (N_13645,N_13350,N_13391);
and U13646 (N_13646,N_13361,N_13470);
xnor U13647 (N_13647,N_13458,N_13382);
xor U13648 (N_13648,N_13484,N_13489);
nand U13649 (N_13649,N_13481,N_13412);
xor U13650 (N_13650,N_13581,N_13542);
xnor U13651 (N_13651,N_13533,N_13546);
nor U13652 (N_13652,N_13578,N_13556);
nor U13653 (N_13653,N_13547,N_13522);
xnor U13654 (N_13654,N_13637,N_13597);
or U13655 (N_13655,N_13577,N_13591);
and U13656 (N_13656,N_13613,N_13590);
and U13657 (N_13657,N_13570,N_13525);
or U13658 (N_13658,N_13592,N_13609);
xnor U13659 (N_13659,N_13540,N_13505);
and U13660 (N_13660,N_13599,N_13504);
or U13661 (N_13661,N_13610,N_13572);
xnor U13662 (N_13662,N_13523,N_13601);
and U13663 (N_13663,N_13586,N_13524);
and U13664 (N_13664,N_13550,N_13521);
xor U13665 (N_13665,N_13560,N_13568);
or U13666 (N_13666,N_13557,N_13583);
or U13667 (N_13667,N_13573,N_13645);
or U13668 (N_13668,N_13575,N_13537);
nand U13669 (N_13669,N_13565,N_13502);
and U13670 (N_13670,N_13622,N_13614);
xnor U13671 (N_13671,N_13618,N_13519);
nand U13672 (N_13672,N_13602,N_13619);
nand U13673 (N_13673,N_13646,N_13582);
and U13674 (N_13674,N_13563,N_13543);
nor U13675 (N_13675,N_13589,N_13511);
xor U13676 (N_13676,N_13638,N_13640);
and U13677 (N_13677,N_13510,N_13625);
or U13678 (N_13678,N_13594,N_13571);
and U13679 (N_13679,N_13593,N_13629);
nand U13680 (N_13680,N_13567,N_13553);
nor U13681 (N_13681,N_13644,N_13648);
and U13682 (N_13682,N_13503,N_13506);
xnor U13683 (N_13683,N_13635,N_13634);
nor U13684 (N_13684,N_13532,N_13520);
xor U13685 (N_13685,N_13636,N_13580);
xor U13686 (N_13686,N_13544,N_13500);
and U13687 (N_13687,N_13564,N_13512);
or U13688 (N_13688,N_13518,N_13628);
and U13689 (N_13689,N_13536,N_13620);
nand U13690 (N_13690,N_13555,N_13508);
xnor U13691 (N_13691,N_13612,N_13566);
and U13692 (N_13692,N_13551,N_13534);
nand U13693 (N_13693,N_13576,N_13531);
nand U13694 (N_13694,N_13626,N_13608);
and U13695 (N_13695,N_13588,N_13535);
xor U13696 (N_13696,N_13516,N_13643);
xnor U13697 (N_13697,N_13617,N_13595);
xnor U13698 (N_13698,N_13501,N_13587);
nand U13699 (N_13699,N_13517,N_13584);
xnor U13700 (N_13700,N_13603,N_13647);
xnor U13701 (N_13701,N_13574,N_13561);
nand U13702 (N_13702,N_13616,N_13548);
xor U13703 (N_13703,N_13611,N_13598);
and U13704 (N_13704,N_13541,N_13526);
nand U13705 (N_13705,N_13549,N_13545);
and U13706 (N_13706,N_13514,N_13579);
nor U13707 (N_13707,N_13621,N_13641);
xnor U13708 (N_13708,N_13530,N_13539);
nand U13709 (N_13709,N_13515,N_13513);
or U13710 (N_13710,N_13639,N_13596);
xnor U13711 (N_13711,N_13627,N_13559);
and U13712 (N_13712,N_13528,N_13554);
xnor U13713 (N_13713,N_13604,N_13507);
nor U13714 (N_13714,N_13615,N_13630);
nor U13715 (N_13715,N_13552,N_13649);
or U13716 (N_13716,N_13632,N_13569);
nor U13717 (N_13717,N_13562,N_13623);
and U13718 (N_13718,N_13509,N_13600);
xor U13719 (N_13719,N_13538,N_13633);
xnor U13720 (N_13720,N_13527,N_13607);
and U13721 (N_13721,N_13585,N_13624);
and U13722 (N_13722,N_13529,N_13606);
xnor U13723 (N_13723,N_13605,N_13642);
xnor U13724 (N_13724,N_13631,N_13558);
or U13725 (N_13725,N_13520,N_13585);
xor U13726 (N_13726,N_13634,N_13560);
or U13727 (N_13727,N_13602,N_13585);
xor U13728 (N_13728,N_13570,N_13607);
nor U13729 (N_13729,N_13531,N_13600);
xor U13730 (N_13730,N_13567,N_13505);
nand U13731 (N_13731,N_13591,N_13539);
nor U13732 (N_13732,N_13520,N_13608);
or U13733 (N_13733,N_13550,N_13507);
and U13734 (N_13734,N_13508,N_13507);
nor U13735 (N_13735,N_13616,N_13509);
nor U13736 (N_13736,N_13636,N_13549);
xnor U13737 (N_13737,N_13502,N_13616);
nor U13738 (N_13738,N_13557,N_13579);
xnor U13739 (N_13739,N_13616,N_13615);
nand U13740 (N_13740,N_13562,N_13587);
xor U13741 (N_13741,N_13647,N_13563);
and U13742 (N_13742,N_13548,N_13552);
nor U13743 (N_13743,N_13552,N_13589);
or U13744 (N_13744,N_13560,N_13599);
xnor U13745 (N_13745,N_13649,N_13602);
or U13746 (N_13746,N_13533,N_13641);
or U13747 (N_13747,N_13581,N_13565);
or U13748 (N_13748,N_13584,N_13572);
nor U13749 (N_13749,N_13594,N_13586);
nor U13750 (N_13750,N_13526,N_13648);
xnor U13751 (N_13751,N_13506,N_13574);
nor U13752 (N_13752,N_13625,N_13589);
and U13753 (N_13753,N_13535,N_13648);
nand U13754 (N_13754,N_13628,N_13640);
nor U13755 (N_13755,N_13608,N_13569);
xnor U13756 (N_13756,N_13507,N_13573);
nand U13757 (N_13757,N_13636,N_13645);
nand U13758 (N_13758,N_13628,N_13604);
xnor U13759 (N_13759,N_13648,N_13577);
or U13760 (N_13760,N_13567,N_13608);
and U13761 (N_13761,N_13566,N_13514);
and U13762 (N_13762,N_13512,N_13506);
xor U13763 (N_13763,N_13618,N_13528);
xnor U13764 (N_13764,N_13611,N_13515);
xor U13765 (N_13765,N_13622,N_13554);
nor U13766 (N_13766,N_13631,N_13592);
nor U13767 (N_13767,N_13561,N_13571);
and U13768 (N_13768,N_13611,N_13500);
and U13769 (N_13769,N_13623,N_13538);
and U13770 (N_13770,N_13622,N_13589);
and U13771 (N_13771,N_13632,N_13545);
and U13772 (N_13772,N_13616,N_13632);
nor U13773 (N_13773,N_13539,N_13581);
nand U13774 (N_13774,N_13565,N_13541);
xor U13775 (N_13775,N_13567,N_13544);
and U13776 (N_13776,N_13593,N_13649);
and U13777 (N_13777,N_13527,N_13638);
xnor U13778 (N_13778,N_13568,N_13626);
xor U13779 (N_13779,N_13589,N_13547);
or U13780 (N_13780,N_13532,N_13539);
and U13781 (N_13781,N_13528,N_13557);
or U13782 (N_13782,N_13628,N_13647);
nor U13783 (N_13783,N_13649,N_13506);
and U13784 (N_13784,N_13586,N_13555);
nand U13785 (N_13785,N_13550,N_13565);
or U13786 (N_13786,N_13594,N_13612);
and U13787 (N_13787,N_13528,N_13595);
xnor U13788 (N_13788,N_13633,N_13620);
nand U13789 (N_13789,N_13567,N_13618);
nand U13790 (N_13790,N_13612,N_13618);
and U13791 (N_13791,N_13571,N_13643);
xor U13792 (N_13792,N_13589,N_13512);
nor U13793 (N_13793,N_13638,N_13501);
and U13794 (N_13794,N_13560,N_13544);
xnor U13795 (N_13795,N_13649,N_13646);
nand U13796 (N_13796,N_13588,N_13612);
nand U13797 (N_13797,N_13629,N_13597);
or U13798 (N_13798,N_13614,N_13529);
nand U13799 (N_13799,N_13636,N_13519);
nand U13800 (N_13800,N_13793,N_13769);
or U13801 (N_13801,N_13745,N_13724);
or U13802 (N_13802,N_13694,N_13660);
nor U13803 (N_13803,N_13727,N_13767);
and U13804 (N_13804,N_13796,N_13768);
nor U13805 (N_13805,N_13778,N_13704);
or U13806 (N_13806,N_13783,N_13701);
nand U13807 (N_13807,N_13787,N_13653);
and U13808 (N_13808,N_13738,N_13758);
xor U13809 (N_13809,N_13794,N_13772);
xor U13810 (N_13810,N_13795,N_13733);
nor U13811 (N_13811,N_13788,N_13784);
nand U13812 (N_13812,N_13675,N_13756);
or U13813 (N_13813,N_13717,N_13663);
or U13814 (N_13814,N_13687,N_13662);
nand U13815 (N_13815,N_13797,N_13708);
nand U13816 (N_13816,N_13780,N_13755);
nand U13817 (N_13817,N_13760,N_13657);
nor U13818 (N_13818,N_13712,N_13651);
xor U13819 (N_13819,N_13684,N_13765);
or U13820 (N_13820,N_13678,N_13754);
nand U13821 (N_13821,N_13781,N_13693);
xnor U13822 (N_13822,N_13709,N_13688);
nand U13823 (N_13823,N_13764,N_13734);
nand U13824 (N_13824,N_13773,N_13770);
xor U13825 (N_13825,N_13779,N_13707);
nand U13826 (N_13826,N_13757,N_13703);
nand U13827 (N_13827,N_13659,N_13683);
xor U13828 (N_13828,N_13721,N_13751);
nor U13829 (N_13829,N_13785,N_13771);
nor U13830 (N_13830,N_13747,N_13672);
xor U13831 (N_13831,N_13665,N_13689);
or U13832 (N_13832,N_13676,N_13792);
or U13833 (N_13833,N_13731,N_13761);
xnor U13834 (N_13834,N_13695,N_13681);
nand U13835 (N_13835,N_13668,N_13716);
nor U13836 (N_13836,N_13666,N_13697);
xnor U13837 (N_13837,N_13699,N_13669);
nand U13838 (N_13838,N_13710,N_13759);
nand U13839 (N_13839,N_13744,N_13741);
and U13840 (N_13840,N_13735,N_13696);
nand U13841 (N_13841,N_13690,N_13700);
xor U13842 (N_13842,N_13692,N_13762);
nand U13843 (N_13843,N_13671,N_13706);
or U13844 (N_13844,N_13705,N_13691);
nor U13845 (N_13845,N_13674,N_13650);
xor U13846 (N_13846,N_13749,N_13736);
or U13847 (N_13847,N_13763,N_13720);
or U13848 (N_13848,N_13702,N_13658);
xor U13849 (N_13849,N_13742,N_13725);
or U13850 (N_13850,N_13748,N_13774);
xnor U13851 (N_13851,N_13698,N_13686);
nor U13852 (N_13852,N_13753,N_13752);
nand U13853 (N_13853,N_13775,N_13670);
nand U13854 (N_13854,N_13718,N_13715);
nor U13855 (N_13855,N_13790,N_13652);
xnor U13856 (N_13856,N_13782,N_13726);
xor U13857 (N_13857,N_13682,N_13730);
xnor U13858 (N_13858,N_13777,N_13750);
nand U13859 (N_13859,N_13786,N_13728);
nor U13860 (N_13860,N_13746,N_13677);
and U13861 (N_13861,N_13766,N_13711);
nor U13862 (N_13862,N_13673,N_13680);
xor U13863 (N_13863,N_13661,N_13791);
or U13864 (N_13864,N_13776,N_13664);
nor U13865 (N_13865,N_13732,N_13723);
xnor U13866 (N_13866,N_13656,N_13654);
xnor U13867 (N_13867,N_13799,N_13714);
xnor U13868 (N_13868,N_13713,N_13655);
and U13869 (N_13869,N_13798,N_13789);
nand U13870 (N_13870,N_13722,N_13679);
or U13871 (N_13871,N_13719,N_13740);
or U13872 (N_13872,N_13737,N_13667);
and U13873 (N_13873,N_13739,N_13729);
or U13874 (N_13874,N_13743,N_13685);
and U13875 (N_13875,N_13749,N_13742);
xor U13876 (N_13876,N_13694,N_13717);
and U13877 (N_13877,N_13714,N_13681);
nor U13878 (N_13878,N_13791,N_13766);
nand U13879 (N_13879,N_13660,N_13700);
xor U13880 (N_13880,N_13750,N_13761);
nor U13881 (N_13881,N_13706,N_13689);
or U13882 (N_13882,N_13690,N_13742);
nand U13883 (N_13883,N_13782,N_13767);
xor U13884 (N_13884,N_13789,N_13674);
xor U13885 (N_13885,N_13693,N_13761);
nor U13886 (N_13886,N_13689,N_13673);
xnor U13887 (N_13887,N_13770,N_13707);
and U13888 (N_13888,N_13699,N_13751);
and U13889 (N_13889,N_13687,N_13759);
or U13890 (N_13890,N_13726,N_13696);
nand U13891 (N_13891,N_13712,N_13674);
nand U13892 (N_13892,N_13752,N_13675);
and U13893 (N_13893,N_13653,N_13780);
nor U13894 (N_13894,N_13797,N_13688);
or U13895 (N_13895,N_13789,N_13742);
nor U13896 (N_13896,N_13669,N_13740);
nand U13897 (N_13897,N_13712,N_13692);
nor U13898 (N_13898,N_13778,N_13787);
xor U13899 (N_13899,N_13733,N_13706);
nor U13900 (N_13900,N_13695,N_13708);
nand U13901 (N_13901,N_13709,N_13745);
nand U13902 (N_13902,N_13716,N_13703);
nand U13903 (N_13903,N_13679,N_13682);
xor U13904 (N_13904,N_13751,N_13706);
nand U13905 (N_13905,N_13729,N_13685);
or U13906 (N_13906,N_13700,N_13676);
nand U13907 (N_13907,N_13674,N_13777);
or U13908 (N_13908,N_13757,N_13725);
and U13909 (N_13909,N_13652,N_13706);
nor U13910 (N_13910,N_13697,N_13651);
nor U13911 (N_13911,N_13662,N_13675);
and U13912 (N_13912,N_13754,N_13680);
or U13913 (N_13913,N_13651,N_13708);
xor U13914 (N_13914,N_13658,N_13715);
or U13915 (N_13915,N_13700,N_13717);
nor U13916 (N_13916,N_13740,N_13735);
or U13917 (N_13917,N_13787,N_13784);
xnor U13918 (N_13918,N_13655,N_13693);
or U13919 (N_13919,N_13688,N_13741);
nand U13920 (N_13920,N_13712,N_13764);
nand U13921 (N_13921,N_13745,N_13787);
nand U13922 (N_13922,N_13658,N_13785);
and U13923 (N_13923,N_13721,N_13659);
or U13924 (N_13924,N_13668,N_13733);
xor U13925 (N_13925,N_13786,N_13713);
nand U13926 (N_13926,N_13772,N_13669);
xor U13927 (N_13927,N_13716,N_13653);
or U13928 (N_13928,N_13654,N_13671);
nor U13929 (N_13929,N_13679,N_13676);
nand U13930 (N_13930,N_13723,N_13778);
or U13931 (N_13931,N_13745,N_13778);
or U13932 (N_13932,N_13763,N_13742);
and U13933 (N_13933,N_13793,N_13667);
or U13934 (N_13934,N_13787,N_13681);
and U13935 (N_13935,N_13778,N_13740);
or U13936 (N_13936,N_13672,N_13679);
or U13937 (N_13937,N_13768,N_13669);
or U13938 (N_13938,N_13685,N_13765);
nor U13939 (N_13939,N_13733,N_13727);
xnor U13940 (N_13940,N_13719,N_13669);
or U13941 (N_13941,N_13696,N_13740);
and U13942 (N_13942,N_13798,N_13722);
or U13943 (N_13943,N_13797,N_13756);
xnor U13944 (N_13944,N_13665,N_13718);
and U13945 (N_13945,N_13768,N_13775);
and U13946 (N_13946,N_13750,N_13674);
or U13947 (N_13947,N_13714,N_13678);
nor U13948 (N_13948,N_13765,N_13703);
nor U13949 (N_13949,N_13759,N_13742);
xor U13950 (N_13950,N_13879,N_13844);
or U13951 (N_13951,N_13839,N_13875);
or U13952 (N_13952,N_13938,N_13807);
or U13953 (N_13953,N_13815,N_13945);
nor U13954 (N_13954,N_13833,N_13803);
or U13955 (N_13955,N_13863,N_13911);
nand U13956 (N_13956,N_13916,N_13828);
nor U13957 (N_13957,N_13840,N_13846);
and U13958 (N_13958,N_13804,N_13858);
and U13959 (N_13959,N_13872,N_13864);
or U13960 (N_13960,N_13932,N_13886);
nand U13961 (N_13961,N_13907,N_13926);
or U13962 (N_13962,N_13873,N_13816);
or U13963 (N_13963,N_13813,N_13924);
xor U13964 (N_13964,N_13836,N_13852);
and U13965 (N_13965,N_13845,N_13905);
nor U13966 (N_13966,N_13826,N_13920);
nand U13967 (N_13967,N_13820,N_13909);
or U13968 (N_13968,N_13832,N_13933);
nor U13969 (N_13969,N_13812,N_13904);
xor U13970 (N_13970,N_13941,N_13901);
nand U13971 (N_13971,N_13888,N_13925);
or U13972 (N_13972,N_13870,N_13891);
xor U13973 (N_13973,N_13856,N_13835);
nand U13974 (N_13974,N_13889,N_13910);
nor U13975 (N_13975,N_13868,N_13906);
nand U13976 (N_13976,N_13814,N_13881);
xnor U13977 (N_13977,N_13827,N_13854);
nand U13978 (N_13978,N_13940,N_13917);
nor U13979 (N_13979,N_13855,N_13885);
nor U13980 (N_13980,N_13929,N_13802);
or U13981 (N_13981,N_13919,N_13939);
nand U13982 (N_13982,N_13913,N_13850);
or U13983 (N_13983,N_13860,N_13818);
or U13984 (N_13984,N_13805,N_13831);
and U13985 (N_13985,N_13937,N_13918);
xor U13986 (N_13986,N_13942,N_13869);
nor U13987 (N_13987,N_13851,N_13948);
and U13988 (N_13988,N_13834,N_13892);
and U13989 (N_13989,N_13943,N_13822);
or U13990 (N_13990,N_13811,N_13936);
and U13991 (N_13991,N_13922,N_13931);
or U13992 (N_13992,N_13829,N_13876);
nand U13993 (N_13993,N_13946,N_13914);
and U13994 (N_13994,N_13896,N_13912);
nand U13995 (N_13995,N_13823,N_13862);
nand U13996 (N_13996,N_13837,N_13921);
xnor U13997 (N_13997,N_13809,N_13903);
or U13998 (N_13998,N_13865,N_13884);
nand U13999 (N_13999,N_13821,N_13825);
and U14000 (N_14000,N_13949,N_13928);
nand U14001 (N_14001,N_13878,N_13808);
xnor U14002 (N_14002,N_13944,N_13842);
or U14003 (N_14003,N_13890,N_13894);
xnor U14004 (N_14004,N_13897,N_13899);
xnor U14005 (N_14005,N_13923,N_13824);
nor U14006 (N_14006,N_13849,N_13838);
or U14007 (N_14007,N_13915,N_13883);
or U14008 (N_14008,N_13847,N_13817);
xnor U14009 (N_14009,N_13935,N_13882);
or U14010 (N_14010,N_13871,N_13908);
xor U14011 (N_14011,N_13853,N_13880);
and U14012 (N_14012,N_13810,N_13877);
and U14013 (N_14013,N_13895,N_13806);
or U14014 (N_14014,N_13857,N_13887);
or U14015 (N_14015,N_13934,N_13843);
or U14016 (N_14016,N_13947,N_13893);
xnor U14017 (N_14017,N_13866,N_13801);
or U14018 (N_14018,N_13800,N_13898);
nor U14019 (N_14019,N_13927,N_13819);
xor U14020 (N_14020,N_13900,N_13874);
and U14021 (N_14021,N_13867,N_13841);
nand U14022 (N_14022,N_13830,N_13902);
nor U14023 (N_14023,N_13848,N_13861);
and U14024 (N_14024,N_13930,N_13859);
nand U14025 (N_14025,N_13823,N_13927);
nor U14026 (N_14026,N_13826,N_13876);
nor U14027 (N_14027,N_13877,N_13946);
nor U14028 (N_14028,N_13887,N_13900);
xor U14029 (N_14029,N_13806,N_13815);
and U14030 (N_14030,N_13887,N_13848);
or U14031 (N_14031,N_13880,N_13949);
and U14032 (N_14032,N_13850,N_13840);
and U14033 (N_14033,N_13818,N_13881);
or U14034 (N_14034,N_13933,N_13868);
xor U14035 (N_14035,N_13844,N_13915);
nand U14036 (N_14036,N_13933,N_13918);
nor U14037 (N_14037,N_13936,N_13839);
xor U14038 (N_14038,N_13816,N_13826);
or U14039 (N_14039,N_13912,N_13925);
nand U14040 (N_14040,N_13932,N_13843);
xnor U14041 (N_14041,N_13848,N_13853);
xnor U14042 (N_14042,N_13943,N_13844);
or U14043 (N_14043,N_13875,N_13842);
nor U14044 (N_14044,N_13942,N_13849);
nor U14045 (N_14045,N_13855,N_13887);
nand U14046 (N_14046,N_13912,N_13947);
nor U14047 (N_14047,N_13908,N_13862);
nand U14048 (N_14048,N_13888,N_13903);
xor U14049 (N_14049,N_13894,N_13892);
nor U14050 (N_14050,N_13858,N_13940);
or U14051 (N_14051,N_13808,N_13817);
nor U14052 (N_14052,N_13898,N_13852);
nand U14053 (N_14053,N_13934,N_13827);
xnor U14054 (N_14054,N_13813,N_13934);
nand U14055 (N_14055,N_13874,N_13904);
or U14056 (N_14056,N_13915,N_13861);
nor U14057 (N_14057,N_13939,N_13828);
nor U14058 (N_14058,N_13934,N_13826);
nor U14059 (N_14059,N_13924,N_13824);
or U14060 (N_14060,N_13915,N_13932);
and U14061 (N_14061,N_13915,N_13853);
nand U14062 (N_14062,N_13838,N_13820);
and U14063 (N_14063,N_13932,N_13934);
nor U14064 (N_14064,N_13946,N_13921);
or U14065 (N_14065,N_13849,N_13870);
and U14066 (N_14066,N_13877,N_13818);
and U14067 (N_14067,N_13940,N_13870);
nand U14068 (N_14068,N_13884,N_13838);
and U14069 (N_14069,N_13819,N_13856);
nor U14070 (N_14070,N_13864,N_13928);
and U14071 (N_14071,N_13802,N_13829);
nand U14072 (N_14072,N_13942,N_13829);
nand U14073 (N_14073,N_13823,N_13829);
xnor U14074 (N_14074,N_13856,N_13807);
and U14075 (N_14075,N_13832,N_13869);
nand U14076 (N_14076,N_13828,N_13913);
nor U14077 (N_14077,N_13829,N_13938);
and U14078 (N_14078,N_13897,N_13840);
nand U14079 (N_14079,N_13805,N_13810);
nand U14080 (N_14080,N_13861,N_13847);
or U14081 (N_14081,N_13839,N_13886);
nand U14082 (N_14082,N_13895,N_13812);
xnor U14083 (N_14083,N_13826,N_13833);
xor U14084 (N_14084,N_13851,N_13929);
nand U14085 (N_14085,N_13800,N_13872);
nand U14086 (N_14086,N_13913,N_13843);
nor U14087 (N_14087,N_13874,N_13833);
nand U14088 (N_14088,N_13894,N_13837);
nand U14089 (N_14089,N_13804,N_13902);
and U14090 (N_14090,N_13811,N_13944);
nor U14091 (N_14091,N_13932,N_13896);
nor U14092 (N_14092,N_13849,N_13924);
xor U14093 (N_14093,N_13910,N_13918);
nor U14094 (N_14094,N_13845,N_13844);
nand U14095 (N_14095,N_13917,N_13943);
nand U14096 (N_14096,N_13823,N_13913);
xor U14097 (N_14097,N_13907,N_13891);
or U14098 (N_14098,N_13866,N_13896);
or U14099 (N_14099,N_13931,N_13877);
xnor U14100 (N_14100,N_14009,N_13963);
xnor U14101 (N_14101,N_14075,N_14088);
xnor U14102 (N_14102,N_14062,N_13990);
xor U14103 (N_14103,N_13993,N_14061);
and U14104 (N_14104,N_14063,N_14054);
or U14105 (N_14105,N_13975,N_14091);
nand U14106 (N_14106,N_14016,N_13957);
nor U14107 (N_14107,N_13960,N_13958);
xnor U14108 (N_14108,N_13995,N_13985);
xor U14109 (N_14109,N_14085,N_13989);
nand U14110 (N_14110,N_13953,N_13951);
or U14111 (N_14111,N_14028,N_14092);
nand U14112 (N_14112,N_13996,N_14093);
and U14113 (N_14113,N_13983,N_14087);
and U14114 (N_14114,N_14033,N_14090);
xor U14115 (N_14115,N_14025,N_14030);
nor U14116 (N_14116,N_14003,N_13964);
xnor U14117 (N_14117,N_14077,N_14040);
nand U14118 (N_14118,N_13952,N_14052);
nand U14119 (N_14119,N_14037,N_14055);
and U14120 (N_14120,N_13955,N_14060);
xor U14121 (N_14121,N_14023,N_14089);
nor U14122 (N_14122,N_13982,N_13991);
and U14123 (N_14123,N_14038,N_14019);
nor U14124 (N_14124,N_14021,N_14029);
nand U14125 (N_14125,N_14006,N_13980);
nor U14126 (N_14126,N_14053,N_14039);
xnor U14127 (N_14127,N_14031,N_14086);
xnor U14128 (N_14128,N_13977,N_13966);
nand U14129 (N_14129,N_14008,N_13950);
or U14130 (N_14130,N_13992,N_14056);
xnor U14131 (N_14131,N_14080,N_13961);
nor U14132 (N_14132,N_14017,N_14002);
nor U14133 (N_14133,N_14001,N_13968);
and U14134 (N_14134,N_14015,N_13971);
and U14135 (N_14135,N_14066,N_14097);
nand U14136 (N_14136,N_13981,N_14004);
nand U14137 (N_14137,N_14045,N_14076);
and U14138 (N_14138,N_14026,N_13988);
or U14139 (N_14139,N_13962,N_13999);
xor U14140 (N_14140,N_14074,N_14005);
or U14141 (N_14141,N_13956,N_14094);
nor U14142 (N_14142,N_14044,N_14071);
xnor U14143 (N_14143,N_13984,N_14032);
nand U14144 (N_14144,N_14051,N_14027);
or U14145 (N_14145,N_14070,N_14068);
or U14146 (N_14146,N_14046,N_13979);
xor U14147 (N_14147,N_13987,N_14081);
nor U14148 (N_14148,N_13972,N_13959);
or U14149 (N_14149,N_14058,N_14059);
nand U14150 (N_14150,N_14048,N_14065);
xor U14151 (N_14151,N_14095,N_14035);
nand U14152 (N_14152,N_14096,N_13970);
or U14153 (N_14153,N_13976,N_14007);
nand U14154 (N_14154,N_14036,N_14047);
xor U14155 (N_14155,N_14041,N_14012);
nand U14156 (N_14156,N_13978,N_14024);
nand U14157 (N_14157,N_14072,N_14000);
and U14158 (N_14158,N_14082,N_14084);
nor U14159 (N_14159,N_14022,N_14078);
nand U14160 (N_14160,N_14014,N_14064);
xor U14161 (N_14161,N_14043,N_13954);
nor U14162 (N_14162,N_13967,N_14011);
nand U14163 (N_14163,N_14042,N_13965);
and U14164 (N_14164,N_13986,N_14049);
xnor U14165 (N_14165,N_14057,N_14098);
xnor U14166 (N_14166,N_14013,N_13974);
nand U14167 (N_14167,N_14069,N_13994);
or U14168 (N_14168,N_13997,N_13973);
nor U14169 (N_14169,N_13998,N_14083);
nor U14170 (N_14170,N_14073,N_14099);
or U14171 (N_14171,N_14034,N_14067);
nor U14172 (N_14172,N_14018,N_13969);
xor U14173 (N_14173,N_14050,N_14010);
or U14174 (N_14174,N_14020,N_14079);
xnor U14175 (N_14175,N_14058,N_13952);
nor U14176 (N_14176,N_14038,N_14094);
nand U14177 (N_14177,N_13973,N_14069);
nor U14178 (N_14178,N_14009,N_13996);
or U14179 (N_14179,N_14046,N_14068);
nand U14180 (N_14180,N_14028,N_13969);
nor U14181 (N_14181,N_14027,N_14039);
or U14182 (N_14182,N_13984,N_14047);
xor U14183 (N_14183,N_14084,N_13996);
or U14184 (N_14184,N_14000,N_13991);
xor U14185 (N_14185,N_13993,N_14038);
or U14186 (N_14186,N_13964,N_14080);
xnor U14187 (N_14187,N_14088,N_14002);
nand U14188 (N_14188,N_14043,N_14046);
nand U14189 (N_14189,N_13979,N_13950);
and U14190 (N_14190,N_14038,N_13961);
nor U14191 (N_14191,N_14060,N_14037);
or U14192 (N_14192,N_14048,N_14099);
xor U14193 (N_14193,N_14082,N_14064);
nor U14194 (N_14194,N_14007,N_13968);
or U14195 (N_14195,N_14058,N_13997);
or U14196 (N_14196,N_14035,N_14082);
or U14197 (N_14197,N_14055,N_13968);
and U14198 (N_14198,N_14028,N_13982);
or U14199 (N_14199,N_14073,N_14039);
xnor U14200 (N_14200,N_13957,N_14044);
or U14201 (N_14201,N_14095,N_14002);
nand U14202 (N_14202,N_13983,N_14061);
or U14203 (N_14203,N_13995,N_14008);
and U14204 (N_14204,N_14047,N_14044);
nor U14205 (N_14205,N_14039,N_14047);
and U14206 (N_14206,N_13965,N_14016);
nand U14207 (N_14207,N_13991,N_14020);
xor U14208 (N_14208,N_14048,N_14023);
and U14209 (N_14209,N_13989,N_14050);
nand U14210 (N_14210,N_14053,N_14072);
nand U14211 (N_14211,N_14080,N_14028);
nand U14212 (N_14212,N_14072,N_13992);
and U14213 (N_14213,N_14001,N_14046);
nor U14214 (N_14214,N_14082,N_14070);
nand U14215 (N_14215,N_14045,N_14013);
nor U14216 (N_14216,N_13969,N_14013);
or U14217 (N_14217,N_13950,N_14059);
and U14218 (N_14218,N_14036,N_13958);
xor U14219 (N_14219,N_13990,N_13981);
or U14220 (N_14220,N_14069,N_14019);
and U14221 (N_14221,N_14038,N_13980);
nor U14222 (N_14222,N_13991,N_13983);
nor U14223 (N_14223,N_14031,N_13959);
nor U14224 (N_14224,N_14026,N_14095);
or U14225 (N_14225,N_13982,N_14030);
or U14226 (N_14226,N_13966,N_14045);
or U14227 (N_14227,N_14049,N_14042);
or U14228 (N_14228,N_14026,N_14042);
xnor U14229 (N_14229,N_14003,N_13962);
and U14230 (N_14230,N_13964,N_14006);
xor U14231 (N_14231,N_14029,N_14063);
xor U14232 (N_14232,N_14095,N_14060);
nand U14233 (N_14233,N_13991,N_14080);
nand U14234 (N_14234,N_14098,N_13951);
and U14235 (N_14235,N_14015,N_14095);
nand U14236 (N_14236,N_13965,N_14074);
or U14237 (N_14237,N_13978,N_14092);
xnor U14238 (N_14238,N_14099,N_13992);
or U14239 (N_14239,N_14097,N_14070);
or U14240 (N_14240,N_13971,N_14046);
xor U14241 (N_14241,N_13958,N_14047);
nor U14242 (N_14242,N_14020,N_14076);
nand U14243 (N_14243,N_14029,N_14013);
or U14244 (N_14244,N_14031,N_14037);
nor U14245 (N_14245,N_14017,N_14058);
nand U14246 (N_14246,N_14057,N_14093);
nand U14247 (N_14247,N_14017,N_13985);
xnor U14248 (N_14248,N_13955,N_13998);
nor U14249 (N_14249,N_14020,N_14024);
xnor U14250 (N_14250,N_14147,N_14204);
and U14251 (N_14251,N_14196,N_14107);
and U14252 (N_14252,N_14206,N_14217);
nand U14253 (N_14253,N_14186,N_14115);
xor U14254 (N_14254,N_14235,N_14103);
and U14255 (N_14255,N_14202,N_14249);
or U14256 (N_14256,N_14236,N_14237);
xnor U14257 (N_14257,N_14152,N_14219);
xnor U14258 (N_14258,N_14171,N_14157);
xnor U14259 (N_14259,N_14165,N_14230);
and U14260 (N_14260,N_14139,N_14106);
and U14261 (N_14261,N_14129,N_14223);
nor U14262 (N_14262,N_14138,N_14169);
and U14263 (N_14263,N_14172,N_14197);
xor U14264 (N_14264,N_14126,N_14122);
xnor U14265 (N_14265,N_14116,N_14241);
nor U14266 (N_14266,N_14208,N_14212);
nand U14267 (N_14267,N_14140,N_14228);
nor U14268 (N_14268,N_14242,N_14188);
and U14269 (N_14269,N_14160,N_14185);
or U14270 (N_14270,N_14137,N_14229);
xnor U14271 (N_14271,N_14243,N_14112);
or U14272 (N_14272,N_14144,N_14246);
nand U14273 (N_14273,N_14200,N_14199);
nand U14274 (N_14274,N_14234,N_14104);
nor U14275 (N_14275,N_14201,N_14108);
and U14276 (N_14276,N_14216,N_14117);
xor U14277 (N_14277,N_14153,N_14211);
xor U14278 (N_14278,N_14111,N_14183);
nor U14279 (N_14279,N_14105,N_14141);
nand U14280 (N_14280,N_14214,N_14240);
and U14281 (N_14281,N_14119,N_14120);
and U14282 (N_14282,N_14215,N_14248);
or U14283 (N_14283,N_14151,N_14189);
and U14284 (N_14284,N_14166,N_14145);
nand U14285 (N_14285,N_14176,N_14207);
xor U14286 (N_14286,N_14226,N_14187);
and U14287 (N_14287,N_14130,N_14222);
and U14288 (N_14288,N_14158,N_14154);
and U14289 (N_14289,N_14182,N_14168);
xor U14290 (N_14290,N_14156,N_14162);
or U14291 (N_14291,N_14244,N_14150);
nand U14292 (N_14292,N_14180,N_14247);
nand U14293 (N_14293,N_14133,N_14221);
nand U14294 (N_14294,N_14198,N_14102);
xnor U14295 (N_14295,N_14191,N_14110);
or U14296 (N_14296,N_14203,N_14175);
and U14297 (N_14297,N_14155,N_14224);
xor U14298 (N_14298,N_14233,N_14148);
xor U14299 (N_14299,N_14159,N_14113);
or U14300 (N_14300,N_14121,N_14123);
and U14301 (N_14301,N_14125,N_14205);
nor U14302 (N_14302,N_14209,N_14146);
and U14303 (N_14303,N_14149,N_14114);
xnor U14304 (N_14304,N_14132,N_14100);
or U14305 (N_14305,N_14225,N_14179);
nand U14306 (N_14306,N_14194,N_14164);
nand U14307 (N_14307,N_14131,N_14135);
xnor U14308 (N_14308,N_14170,N_14163);
xor U14309 (N_14309,N_14174,N_14142);
and U14310 (N_14310,N_14181,N_14184);
or U14311 (N_14311,N_14220,N_14210);
or U14312 (N_14312,N_14178,N_14239);
xor U14313 (N_14313,N_14128,N_14190);
and U14314 (N_14314,N_14161,N_14238);
and U14315 (N_14315,N_14193,N_14245);
and U14316 (N_14316,N_14195,N_14227);
nor U14317 (N_14317,N_14167,N_14213);
nor U14318 (N_14318,N_14143,N_14218);
or U14319 (N_14319,N_14118,N_14173);
xor U14320 (N_14320,N_14109,N_14136);
or U14321 (N_14321,N_14101,N_14177);
nor U14322 (N_14322,N_14124,N_14232);
and U14323 (N_14323,N_14192,N_14231);
and U14324 (N_14324,N_14134,N_14127);
or U14325 (N_14325,N_14191,N_14179);
xnor U14326 (N_14326,N_14247,N_14198);
nand U14327 (N_14327,N_14123,N_14119);
nor U14328 (N_14328,N_14156,N_14102);
and U14329 (N_14329,N_14159,N_14202);
xnor U14330 (N_14330,N_14128,N_14187);
nor U14331 (N_14331,N_14132,N_14112);
and U14332 (N_14332,N_14213,N_14223);
nor U14333 (N_14333,N_14121,N_14112);
nand U14334 (N_14334,N_14234,N_14194);
xor U14335 (N_14335,N_14130,N_14177);
or U14336 (N_14336,N_14229,N_14112);
nand U14337 (N_14337,N_14196,N_14162);
or U14338 (N_14338,N_14171,N_14222);
xor U14339 (N_14339,N_14190,N_14202);
xor U14340 (N_14340,N_14109,N_14181);
nand U14341 (N_14341,N_14104,N_14166);
xor U14342 (N_14342,N_14104,N_14214);
nor U14343 (N_14343,N_14148,N_14202);
nand U14344 (N_14344,N_14190,N_14247);
xnor U14345 (N_14345,N_14249,N_14134);
or U14346 (N_14346,N_14136,N_14198);
nor U14347 (N_14347,N_14188,N_14106);
or U14348 (N_14348,N_14131,N_14230);
xor U14349 (N_14349,N_14249,N_14205);
nor U14350 (N_14350,N_14109,N_14183);
or U14351 (N_14351,N_14177,N_14141);
nor U14352 (N_14352,N_14192,N_14204);
xnor U14353 (N_14353,N_14212,N_14177);
nor U14354 (N_14354,N_14128,N_14108);
or U14355 (N_14355,N_14168,N_14100);
or U14356 (N_14356,N_14122,N_14234);
nor U14357 (N_14357,N_14218,N_14147);
nor U14358 (N_14358,N_14126,N_14145);
nor U14359 (N_14359,N_14181,N_14155);
and U14360 (N_14360,N_14221,N_14168);
or U14361 (N_14361,N_14246,N_14231);
nor U14362 (N_14362,N_14158,N_14119);
and U14363 (N_14363,N_14180,N_14133);
nand U14364 (N_14364,N_14238,N_14242);
nand U14365 (N_14365,N_14225,N_14155);
nand U14366 (N_14366,N_14224,N_14162);
nand U14367 (N_14367,N_14158,N_14177);
nand U14368 (N_14368,N_14212,N_14108);
xor U14369 (N_14369,N_14195,N_14242);
xnor U14370 (N_14370,N_14106,N_14138);
nor U14371 (N_14371,N_14120,N_14189);
or U14372 (N_14372,N_14197,N_14137);
nand U14373 (N_14373,N_14221,N_14100);
nand U14374 (N_14374,N_14171,N_14132);
xnor U14375 (N_14375,N_14144,N_14162);
xnor U14376 (N_14376,N_14227,N_14101);
or U14377 (N_14377,N_14232,N_14178);
or U14378 (N_14378,N_14175,N_14185);
and U14379 (N_14379,N_14221,N_14130);
nor U14380 (N_14380,N_14129,N_14105);
and U14381 (N_14381,N_14158,N_14153);
nand U14382 (N_14382,N_14235,N_14166);
or U14383 (N_14383,N_14245,N_14231);
or U14384 (N_14384,N_14204,N_14212);
or U14385 (N_14385,N_14239,N_14224);
nor U14386 (N_14386,N_14239,N_14169);
xnor U14387 (N_14387,N_14157,N_14131);
xor U14388 (N_14388,N_14237,N_14208);
and U14389 (N_14389,N_14213,N_14191);
nand U14390 (N_14390,N_14222,N_14242);
and U14391 (N_14391,N_14195,N_14114);
nor U14392 (N_14392,N_14102,N_14143);
xnor U14393 (N_14393,N_14158,N_14155);
and U14394 (N_14394,N_14109,N_14138);
and U14395 (N_14395,N_14132,N_14202);
and U14396 (N_14396,N_14121,N_14124);
nand U14397 (N_14397,N_14177,N_14222);
or U14398 (N_14398,N_14247,N_14107);
and U14399 (N_14399,N_14195,N_14174);
nand U14400 (N_14400,N_14253,N_14356);
or U14401 (N_14401,N_14316,N_14343);
xnor U14402 (N_14402,N_14315,N_14364);
and U14403 (N_14403,N_14276,N_14374);
or U14404 (N_14404,N_14360,N_14377);
xor U14405 (N_14405,N_14286,N_14296);
xor U14406 (N_14406,N_14345,N_14370);
nor U14407 (N_14407,N_14301,N_14342);
nand U14408 (N_14408,N_14382,N_14307);
nor U14409 (N_14409,N_14303,N_14346);
nand U14410 (N_14410,N_14275,N_14349);
and U14411 (N_14411,N_14381,N_14273);
xor U14412 (N_14412,N_14271,N_14262);
xnor U14413 (N_14413,N_14395,N_14363);
and U14414 (N_14414,N_14387,N_14366);
or U14415 (N_14415,N_14338,N_14327);
xor U14416 (N_14416,N_14298,N_14388);
xor U14417 (N_14417,N_14294,N_14281);
nand U14418 (N_14418,N_14354,N_14329);
xor U14419 (N_14419,N_14277,N_14267);
nand U14420 (N_14420,N_14257,N_14309);
xnor U14421 (N_14421,N_14268,N_14306);
nand U14422 (N_14422,N_14384,N_14335);
and U14423 (N_14423,N_14317,N_14337);
or U14424 (N_14424,N_14287,N_14270);
xnor U14425 (N_14425,N_14368,N_14279);
xor U14426 (N_14426,N_14280,N_14269);
or U14427 (N_14427,N_14393,N_14259);
and U14428 (N_14428,N_14341,N_14369);
nand U14429 (N_14429,N_14310,N_14305);
nor U14430 (N_14430,N_14260,N_14302);
nor U14431 (N_14431,N_14394,N_14290);
and U14432 (N_14432,N_14375,N_14320);
and U14433 (N_14433,N_14376,N_14297);
nand U14434 (N_14434,N_14348,N_14261);
nor U14435 (N_14435,N_14398,N_14312);
or U14436 (N_14436,N_14359,N_14344);
nand U14437 (N_14437,N_14386,N_14373);
nand U14438 (N_14438,N_14380,N_14385);
xnor U14439 (N_14439,N_14254,N_14371);
xnor U14440 (N_14440,N_14391,N_14266);
and U14441 (N_14441,N_14331,N_14361);
nor U14442 (N_14442,N_14263,N_14383);
nor U14443 (N_14443,N_14340,N_14278);
and U14444 (N_14444,N_14326,N_14293);
and U14445 (N_14445,N_14399,N_14378);
and U14446 (N_14446,N_14292,N_14333);
nor U14447 (N_14447,N_14285,N_14283);
xnor U14448 (N_14448,N_14324,N_14265);
and U14449 (N_14449,N_14339,N_14289);
or U14450 (N_14450,N_14313,N_14252);
nor U14451 (N_14451,N_14336,N_14367);
and U14452 (N_14452,N_14350,N_14355);
nor U14453 (N_14453,N_14372,N_14322);
nor U14454 (N_14454,N_14250,N_14300);
nor U14455 (N_14455,N_14332,N_14379);
nor U14456 (N_14456,N_14295,N_14314);
xnor U14457 (N_14457,N_14288,N_14389);
nor U14458 (N_14458,N_14299,N_14334);
or U14459 (N_14459,N_14351,N_14258);
nor U14460 (N_14460,N_14392,N_14330);
and U14461 (N_14461,N_14311,N_14396);
nor U14462 (N_14462,N_14353,N_14321);
and U14463 (N_14463,N_14328,N_14319);
xnor U14464 (N_14464,N_14397,N_14357);
or U14465 (N_14465,N_14255,N_14347);
and U14466 (N_14466,N_14308,N_14352);
nand U14467 (N_14467,N_14274,N_14358);
nor U14468 (N_14468,N_14323,N_14304);
and U14469 (N_14469,N_14365,N_14256);
nand U14470 (N_14470,N_14325,N_14362);
xnor U14471 (N_14471,N_14272,N_14284);
nor U14472 (N_14472,N_14390,N_14291);
nor U14473 (N_14473,N_14251,N_14318);
nand U14474 (N_14474,N_14264,N_14282);
and U14475 (N_14475,N_14364,N_14254);
or U14476 (N_14476,N_14305,N_14302);
and U14477 (N_14477,N_14260,N_14387);
xnor U14478 (N_14478,N_14384,N_14286);
or U14479 (N_14479,N_14309,N_14357);
nor U14480 (N_14480,N_14306,N_14348);
xor U14481 (N_14481,N_14285,N_14357);
or U14482 (N_14482,N_14278,N_14391);
or U14483 (N_14483,N_14264,N_14356);
or U14484 (N_14484,N_14306,N_14256);
nor U14485 (N_14485,N_14292,N_14305);
and U14486 (N_14486,N_14297,N_14288);
and U14487 (N_14487,N_14384,N_14289);
nor U14488 (N_14488,N_14361,N_14295);
nand U14489 (N_14489,N_14250,N_14362);
or U14490 (N_14490,N_14334,N_14395);
nand U14491 (N_14491,N_14336,N_14388);
nor U14492 (N_14492,N_14308,N_14298);
xnor U14493 (N_14493,N_14366,N_14307);
xnor U14494 (N_14494,N_14274,N_14365);
xnor U14495 (N_14495,N_14335,N_14389);
nor U14496 (N_14496,N_14328,N_14274);
nand U14497 (N_14497,N_14353,N_14305);
or U14498 (N_14498,N_14309,N_14371);
nand U14499 (N_14499,N_14256,N_14352);
nand U14500 (N_14500,N_14288,N_14292);
or U14501 (N_14501,N_14343,N_14257);
xnor U14502 (N_14502,N_14275,N_14365);
and U14503 (N_14503,N_14292,N_14310);
and U14504 (N_14504,N_14263,N_14280);
nand U14505 (N_14505,N_14275,N_14359);
and U14506 (N_14506,N_14297,N_14363);
nand U14507 (N_14507,N_14332,N_14390);
and U14508 (N_14508,N_14273,N_14306);
nor U14509 (N_14509,N_14355,N_14374);
and U14510 (N_14510,N_14350,N_14348);
nand U14511 (N_14511,N_14256,N_14375);
xor U14512 (N_14512,N_14260,N_14314);
xor U14513 (N_14513,N_14274,N_14385);
and U14514 (N_14514,N_14284,N_14365);
nand U14515 (N_14515,N_14259,N_14390);
or U14516 (N_14516,N_14283,N_14369);
nor U14517 (N_14517,N_14260,N_14276);
xor U14518 (N_14518,N_14358,N_14357);
nand U14519 (N_14519,N_14343,N_14368);
nor U14520 (N_14520,N_14291,N_14396);
nand U14521 (N_14521,N_14331,N_14395);
and U14522 (N_14522,N_14265,N_14377);
and U14523 (N_14523,N_14275,N_14279);
nor U14524 (N_14524,N_14343,N_14282);
nand U14525 (N_14525,N_14368,N_14278);
nand U14526 (N_14526,N_14286,N_14368);
nand U14527 (N_14527,N_14321,N_14349);
or U14528 (N_14528,N_14258,N_14334);
nor U14529 (N_14529,N_14363,N_14318);
nand U14530 (N_14530,N_14381,N_14357);
nand U14531 (N_14531,N_14282,N_14292);
nand U14532 (N_14532,N_14342,N_14395);
nor U14533 (N_14533,N_14267,N_14306);
or U14534 (N_14534,N_14280,N_14345);
nand U14535 (N_14535,N_14325,N_14363);
nand U14536 (N_14536,N_14360,N_14319);
nand U14537 (N_14537,N_14373,N_14299);
xnor U14538 (N_14538,N_14306,N_14388);
or U14539 (N_14539,N_14387,N_14327);
and U14540 (N_14540,N_14315,N_14323);
xnor U14541 (N_14541,N_14340,N_14383);
or U14542 (N_14542,N_14315,N_14280);
nand U14543 (N_14543,N_14397,N_14332);
nand U14544 (N_14544,N_14292,N_14325);
nand U14545 (N_14545,N_14352,N_14372);
and U14546 (N_14546,N_14372,N_14324);
xnor U14547 (N_14547,N_14328,N_14350);
xor U14548 (N_14548,N_14265,N_14263);
and U14549 (N_14549,N_14362,N_14355);
xor U14550 (N_14550,N_14524,N_14462);
nand U14551 (N_14551,N_14461,N_14490);
xnor U14552 (N_14552,N_14460,N_14499);
or U14553 (N_14553,N_14546,N_14534);
xor U14554 (N_14554,N_14440,N_14401);
or U14555 (N_14555,N_14527,N_14530);
or U14556 (N_14556,N_14424,N_14452);
nand U14557 (N_14557,N_14526,N_14548);
nand U14558 (N_14558,N_14518,N_14541);
and U14559 (N_14559,N_14488,N_14400);
and U14560 (N_14560,N_14442,N_14409);
xnor U14561 (N_14561,N_14431,N_14445);
and U14562 (N_14562,N_14477,N_14480);
nor U14563 (N_14563,N_14498,N_14545);
or U14564 (N_14564,N_14422,N_14485);
nor U14565 (N_14565,N_14497,N_14408);
or U14566 (N_14566,N_14463,N_14509);
xor U14567 (N_14567,N_14467,N_14456);
nor U14568 (N_14568,N_14474,N_14435);
nor U14569 (N_14569,N_14532,N_14496);
and U14570 (N_14570,N_14507,N_14468);
and U14571 (N_14571,N_14418,N_14453);
and U14572 (N_14572,N_14495,N_14514);
xnor U14573 (N_14573,N_14448,N_14472);
nor U14574 (N_14574,N_14484,N_14406);
or U14575 (N_14575,N_14520,N_14522);
or U14576 (N_14576,N_14417,N_14427);
nor U14577 (N_14577,N_14403,N_14523);
and U14578 (N_14578,N_14420,N_14421);
nor U14579 (N_14579,N_14471,N_14503);
or U14580 (N_14580,N_14439,N_14482);
and U14581 (N_14581,N_14419,N_14457);
nor U14582 (N_14582,N_14434,N_14525);
xor U14583 (N_14583,N_14493,N_14405);
or U14584 (N_14584,N_14429,N_14455);
or U14585 (N_14585,N_14505,N_14458);
and U14586 (N_14586,N_14410,N_14447);
or U14587 (N_14587,N_14411,N_14483);
and U14588 (N_14588,N_14451,N_14416);
and U14589 (N_14589,N_14539,N_14504);
nor U14590 (N_14590,N_14531,N_14478);
nor U14591 (N_14591,N_14492,N_14487);
nand U14592 (N_14592,N_14481,N_14540);
or U14593 (N_14593,N_14533,N_14430);
xnor U14594 (N_14594,N_14512,N_14432);
nand U14595 (N_14595,N_14538,N_14508);
nand U14596 (N_14596,N_14469,N_14446);
and U14597 (N_14597,N_14426,N_14402);
nor U14598 (N_14598,N_14414,N_14511);
nand U14599 (N_14599,N_14513,N_14506);
and U14600 (N_14600,N_14491,N_14515);
and U14601 (N_14601,N_14516,N_14412);
and U14602 (N_14602,N_14537,N_14437);
or U14603 (N_14603,N_14413,N_14510);
nor U14604 (N_14604,N_14501,N_14544);
or U14605 (N_14605,N_14517,N_14549);
xnor U14606 (N_14606,N_14433,N_14536);
xor U14607 (N_14607,N_14529,N_14479);
nor U14608 (N_14608,N_14438,N_14441);
or U14609 (N_14609,N_14459,N_14423);
and U14610 (N_14610,N_14547,N_14444);
xnor U14611 (N_14611,N_14407,N_14425);
and U14612 (N_14612,N_14443,N_14428);
nor U14613 (N_14613,N_14473,N_14475);
and U14614 (N_14614,N_14494,N_14465);
and U14615 (N_14615,N_14486,N_14519);
or U14616 (N_14616,N_14489,N_14502);
xnor U14617 (N_14617,N_14521,N_14450);
nand U14618 (N_14618,N_14454,N_14404);
xor U14619 (N_14619,N_14415,N_14535);
or U14620 (N_14620,N_14436,N_14449);
nand U14621 (N_14621,N_14543,N_14528);
or U14622 (N_14622,N_14500,N_14476);
and U14623 (N_14623,N_14464,N_14470);
and U14624 (N_14624,N_14466,N_14542);
or U14625 (N_14625,N_14513,N_14452);
and U14626 (N_14626,N_14531,N_14451);
xnor U14627 (N_14627,N_14485,N_14488);
nor U14628 (N_14628,N_14439,N_14492);
or U14629 (N_14629,N_14488,N_14530);
xor U14630 (N_14630,N_14506,N_14478);
or U14631 (N_14631,N_14475,N_14511);
nor U14632 (N_14632,N_14400,N_14459);
or U14633 (N_14633,N_14422,N_14546);
or U14634 (N_14634,N_14491,N_14489);
or U14635 (N_14635,N_14537,N_14411);
xnor U14636 (N_14636,N_14547,N_14449);
xor U14637 (N_14637,N_14453,N_14402);
and U14638 (N_14638,N_14415,N_14525);
nor U14639 (N_14639,N_14412,N_14477);
and U14640 (N_14640,N_14520,N_14473);
nor U14641 (N_14641,N_14517,N_14413);
xor U14642 (N_14642,N_14476,N_14526);
nor U14643 (N_14643,N_14481,N_14537);
and U14644 (N_14644,N_14446,N_14413);
nand U14645 (N_14645,N_14518,N_14539);
or U14646 (N_14646,N_14455,N_14513);
and U14647 (N_14647,N_14408,N_14480);
or U14648 (N_14648,N_14543,N_14429);
and U14649 (N_14649,N_14519,N_14507);
nand U14650 (N_14650,N_14441,N_14481);
nand U14651 (N_14651,N_14495,N_14441);
xor U14652 (N_14652,N_14494,N_14467);
and U14653 (N_14653,N_14419,N_14411);
and U14654 (N_14654,N_14523,N_14535);
xor U14655 (N_14655,N_14508,N_14468);
or U14656 (N_14656,N_14457,N_14414);
xor U14657 (N_14657,N_14498,N_14451);
nand U14658 (N_14658,N_14401,N_14445);
nor U14659 (N_14659,N_14491,N_14412);
or U14660 (N_14660,N_14451,N_14435);
or U14661 (N_14661,N_14504,N_14474);
nor U14662 (N_14662,N_14506,N_14481);
xor U14663 (N_14663,N_14427,N_14548);
nor U14664 (N_14664,N_14433,N_14443);
nor U14665 (N_14665,N_14465,N_14523);
or U14666 (N_14666,N_14516,N_14506);
or U14667 (N_14667,N_14406,N_14483);
nand U14668 (N_14668,N_14442,N_14402);
and U14669 (N_14669,N_14451,N_14406);
and U14670 (N_14670,N_14482,N_14514);
or U14671 (N_14671,N_14480,N_14518);
or U14672 (N_14672,N_14443,N_14548);
and U14673 (N_14673,N_14500,N_14408);
xnor U14674 (N_14674,N_14433,N_14518);
nand U14675 (N_14675,N_14532,N_14464);
and U14676 (N_14676,N_14413,N_14505);
nand U14677 (N_14677,N_14442,N_14492);
nor U14678 (N_14678,N_14416,N_14456);
xnor U14679 (N_14679,N_14458,N_14541);
nand U14680 (N_14680,N_14485,N_14406);
nand U14681 (N_14681,N_14486,N_14416);
and U14682 (N_14682,N_14519,N_14425);
nor U14683 (N_14683,N_14403,N_14448);
nor U14684 (N_14684,N_14464,N_14466);
xor U14685 (N_14685,N_14429,N_14479);
nand U14686 (N_14686,N_14420,N_14469);
nand U14687 (N_14687,N_14434,N_14532);
nor U14688 (N_14688,N_14446,N_14417);
nor U14689 (N_14689,N_14478,N_14412);
nand U14690 (N_14690,N_14540,N_14548);
nand U14691 (N_14691,N_14512,N_14430);
xnor U14692 (N_14692,N_14450,N_14522);
nand U14693 (N_14693,N_14526,N_14411);
nand U14694 (N_14694,N_14425,N_14402);
xor U14695 (N_14695,N_14483,N_14480);
xnor U14696 (N_14696,N_14472,N_14547);
nand U14697 (N_14697,N_14516,N_14419);
xor U14698 (N_14698,N_14467,N_14462);
nand U14699 (N_14699,N_14496,N_14481);
nand U14700 (N_14700,N_14608,N_14607);
and U14701 (N_14701,N_14657,N_14621);
xor U14702 (N_14702,N_14590,N_14639);
xor U14703 (N_14703,N_14673,N_14580);
nor U14704 (N_14704,N_14612,N_14651);
and U14705 (N_14705,N_14640,N_14596);
xor U14706 (N_14706,N_14664,N_14584);
nor U14707 (N_14707,N_14647,N_14571);
and U14708 (N_14708,N_14659,N_14609);
nor U14709 (N_14709,N_14595,N_14698);
xor U14710 (N_14710,N_14672,N_14574);
nor U14711 (N_14711,N_14560,N_14598);
xor U14712 (N_14712,N_14601,N_14551);
xnor U14713 (N_14713,N_14565,N_14628);
or U14714 (N_14714,N_14645,N_14615);
nor U14715 (N_14715,N_14666,N_14685);
or U14716 (N_14716,N_14634,N_14654);
and U14717 (N_14717,N_14695,N_14658);
xnor U14718 (N_14718,N_14688,N_14569);
nand U14719 (N_14719,N_14644,N_14681);
nand U14720 (N_14720,N_14680,N_14573);
nor U14721 (N_14721,N_14694,N_14655);
xor U14722 (N_14722,N_14610,N_14564);
xor U14723 (N_14723,N_14567,N_14589);
and U14724 (N_14724,N_14669,N_14617);
nand U14725 (N_14725,N_14618,N_14559);
xnor U14726 (N_14726,N_14582,N_14587);
and U14727 (N_14727,N_14662,N_14667);
nand U14728 (N_14728,N_14638,N_14578);
xor U14729 (N_14729,N_14653,N_14576);
and U14730 (N_14730,N_14632,N_14699);
xnor U14731 (N_14731,N_14668,N_14629);
and U14732 (N_14732,N_14661,N_14679);
and U14733 (N_14733,N_14689,N_14620);
nor U14734 (N_14734,N_14597,N_14665);
and U14735 (N_14735,N_14622,N_14557);
nand U14736 (N_14736,N_14562,N_14627);
nand U14737 (N_14737,N_14693,N_14624);
nand U14738 (N_14738,N_14630,N_14561);
or U14739 (N_14739,N_14563,N_14697);
nor U14740 (N_14740,N_14619,N_14660);
or U14741 (N_14741,N_14604,N_14550);
and U14742 (N_14742,N_14623,N_14682);
nand U14743 (N_14743,N_14686,N_14570);
or U14744 (N_14744,N_14599,N_14646);
nand U14745 (N_14745,N_14674,N_14684);
xor U14746 (N_14746,N_14579,N_14677);
xnor U14747 (N_14747,N_14588,N_14663);
or U14748 (N_14748,N_14552,N_14671);
nor U14749 (N_14749,N_14648,N_14613);
nand U14750 (N_14750,N_14633,N_14649);
nor U14751 (N_14751,N_14636,N_14637);
or U14752 (N_14752,N_14583,N_14670);
xnor U14753 (N_14753,N_14683,N_14642);
nor U14754 (N_14754,N_14650,N_14553);
and U14755 (N_14755,N_14605,N_14594);
xnor U14756 (N_14756,N_14575,N_14606);
nand U14757 (N_14757,N_14592,N_14631);
or U14758 (N_14758,N_14678,N_14614);
or U14759 (N_14759,N_14616,N_14602);
nand U14760 (N_14760,N_14572,N_14585);
xnor U14761 (N_14761,N_14568,N_14691);
and U14762 (N_14762,N_14696,N_14591);
xor U14763 (N_14763,N_14635,N_14626);
nor U14764 (N_14764,N_14556,N_14643);
xnor U14765 (N_14765,N_14656,N_14611);
xnor U14766 (N_14766,N_14625,N_14555);
nand U14767 (N_14767,N_14600,N_14676);
nor U14768 (N_14768,N_14593,N_14692);
and U14769 (N_14769,N_14603,N_14558);
or U14770 (N_14770,N_14554,N_14566);
and U14771 (N_14771,N_14586,N_14652);
or U14772 (N_14772,N_14675,N_14581);
or U14773 (N_14773,N_14641,N_14687);
nand U14774 (N_14774,N_14577,N_14690);
or U14775 (N_14775,N_14603,N_14587);
nand U14776 (N_14776,N_14660,N_14685);
and U14777 (N_14777,N_14608,N_14695);
nor U14778 (N_14778,N_14557,N_14683);
nor U14779 (N_14779,N_14662,N_14590);
xor U14780 (N_14780,N_14679,N_14671);
xor U14781 (N_14781,N_14604,N_14648);
or U14782 (N_14782,N_14625,N_14639);
nor U14783 (N_14783,N_14658,N_14697);
nand U14784 (N_14784,N_14550,N_14625);
and U14785 (N_14785,N_14667,N_14595);
and U14786 (N_14786,N_14597,N_14655);
and U14787 (N_14787,N_14564,N_14699);
nor U14788 (N_14788,N_14678,N_14603);
xor U14789 (N_14789,N_14637,N_14695);
xnor U14790 (N_14790,N_14616,N_14563);
and U14791 (N_14791,N_14551,N_14630);
or U14792 (N_14792,N_14583,N_14673);
nor U14793 (N_14793,N_14690,N_14553);
nor U14794 (N_14794,N_14562,N_14652);
nor U14795 (N_14795,N_14640,N_14622);
xor U14796 (N_14796,N_14552,N_14694);
or U14797 (N_14797,N_14674,N_14568);
or U14798 (N_14798,N_14674,N_14629);
xnor U14799 (N_14799,N_14666,N_14690);
nand U14800 (N_14800,N_14555,N_14586);
xnor U14801 (N_14801,N_14607,N_14580);
nand U14802 (N_14802,N_14573,N_14674);
nor U14803 (N_14803,N_14606,N_14623);
nand U14804 (N_14804,N_14696,N_14676);
xor U14805 (N_14805,N_14550,N_14569);
and U14806 (N_14806,N_14598,N_14695);
nand U14807 (N_14807,N_14644,N_14696);
xnor U14808 (N_14808,N_14597,N_14673);
and U14809 (N_14809,N_14690,N_14582);
and U14810 (N_14810,N_14639,N_14552);
nor U14811 (N_14811,N_14637,N_14649);
or U14812 (N_14812,N_14645,N_14556);
xor U14813 (N_14813,N_14621,N_14613);
or U14814 (N_14814,N_14678,N_14680);
or U14815 (N_14815,N_14580,N_14637);
xor U14816 (N_14816,N_14649,N_14630);
nor U14817 (N_14817,N_14575,N_14668);
xor U14818 (N_14818,N_14671,N_14592);
xor U14819 (N_14819,N_14597,N_14642);
and U14820 (N_14820,N_14595,N_14558);
xnor U14821 (N_14821,N_14606,N_14611);
nor U14822 (N_14822,N_14664,N_14573);
and U14823 (N_14823,N_14665,N_14687);
and U14824 (N_14824,N_14617,N_14678);
or U14825 (N_14825,N_14571,N_14641);
and U14826 (N_14826,N_14572,N_14673);
nor U14827 (N_14827,N_14551,N_14618);
nor U14828 (N_14828,N_14697,N_14583);
or U14829 (N_14829,N_14595,N_14659);
or U14830 (N_14830,N_14605,N_14648);
or U14831 (N_14831,N_14644,N_14698);
xor U14832 (N_14832,N_14697,N_14698);
xnor U14833 (N_14833,N_14554,N_14642);
nand U14834 (N_14834,N_14563,N_14682);
nor U14835 (N_14835,N_14683,N_14619);
and U14836 (N_14836,N_14637,N_14635);
nor U14837 (N_14837,N_14562,N_14586);
nor U14838 (N_14838,N_14617,N_14571);
xnor U14839 (N_14839,N_14672,N_14580);
or U14840 (N_14840,N_14590,N_14561);
or U14841 (N_14841,N_14550,N_14690);
nor U14842 (N_14842,N_14639,N_14671);
and U14843 (N_14843,N_14621,N_14674);
and U14844 (N_14844,N_14595,N_14569);
nand U14845 (N_14845,N_14605,N_14682);
nor U14846 (N_14846,N_14550,N_14695);
nand U14847 (N_14847,N_14639,N_14661);
or U14848 (N_14848,N_14687,N_14599);
xnor U14849 (N_14849,N_14699,N_14621);
nor U14850 (N_14850,N_14786,N_14706);
nor U14851 (N_14851,N_14811,N_14801);
xnor U14852 (N_14852,N_14732,N_14803);
or U14853 (N_14853,N_14826,N_14814);
nor U14854 (N_14854,N_14719,N_14807);
or U14855 (N_14855,N_14737,N_14756);
and U14856 (N_14856,N_14717,N_14813);
or U14857 (N_14857,N_14795,N_14753);
or U14858 (N_14858,N_14718,N_14789);
and U14859 (N_14859,N_14782,N_14778);
xnor U14860 (N_14860,N_14735,N_14781);
nor U14861 (N_14861,N_14741,N_14798);
nand U14862 (N_14862,N_14791,N_14708);
nor U14863 (N_14863,N_14834,N_14823);
nand U14864 (N_14864,N_14759,N_14771);
nand U14865 (N_14865,N_14747,N_14724);
and U14866 (N_14866,N_14775,N_14780);
xnor U14867 (N_14867,N_14772,N_14704);
xor U14868 (N_14868,N_14725,N_14808);
nand U14869 (N_14869,N_14822,N_14769);
nand U14870 (N_14870,N_14832,N_14714);
xnor U14871 (N_14871,N_14793,N_14846);
or U14872 (N_14872,N_14757,N_14796);
xor U14873 (N_14873,N_14847,N_14707);
nor U14874 (N_14874,N_14820,N_14844);
nand U14875 (N_14875,N_14797,N_14710);
and U14876 (N_14876,N_14767,N_14827);
xor U14877 (N_14877,N_14831,N_14788);
nor U14878 (N_14878,N_14815,N_14709);
xor U14879 (N_14879,N_14729,N_14766);
xor U14880 (N_14880,N_14721,N_14758);
xnor U14881 (N_14881,N_14702,N_14754);
or U14882 (N_14882,N_14806,N_14761);
nand U14883 (N_14883,N_14700,N_14787);
nor U14884 (N_14884,N_14727,N_14792);
or U14885 (N_14885,N_14731,N_14752);
or U14886 (N_14886,N_14734,N_14768);
xor U14887 (N_14887,N_14836,N_14711);
xnor U14888 (N_14888,N_14739,N_14712);
xor U14889 (N_14889,N_14805,N_14736);
or U14890 (N_14890,N_14819,N_14728);
nor U14891 (N_14891,N_14777,N_14743);
xnor U14892 (N_14892,N_14829,N_14722);
xnor U14893 (N_14893,N_14749,N_14713);
nand U14894 (N_14894,N_14705,N_14738);
xnor U14895 (N_14895,N_14848,N_14776);
nand U14896 (N_14896,N_14701,N_14849);
xor U14897 (N_14897,N_14785,N_14716);
nor U14898 (N_14898,N_14760,N_14750);
xnor U14899 (N_14899,N_14830,N_14802);
xnor U14900 (N_14900,N_14804,N_14824);
nand U14901 (N_14901,N_14812,N_14821);
and U14902 (N_14902,N_14703,N_14840);
nor U14903 (N_14903,N_14765,N_14809);
nand U14904 (N_14904,N_14762,N_14748);
nand U14905 (N_14905,N_14764,N_14733);
xor U14906 (N_14906,N_14839,N_14818);
or U14907 (N_14907,N_14835,N_14817);
and U14908 (N_14908,N_14740,N_14838);
and U14909 (N_14909,N_14720,N_14755);
xnor U14910 (N_14910,N_14837,N_14726);
xor U14911 (N_14911,N_14730,N_14833);
nand U14912 (N_14912,N_14828,N_14746);
nor U14913 (N_14913,N_14751,N_14800);
or U14914 (N_14914,N_14745,N_14773);
or U14915 (N_14915,N_14842,N_14770);
nand U14916 (N_14916,N_14794,N_14843);
and U14917 (N_14917,N_14784,N_14841);
nand U14918 (N_14918,N_14744,N_14723);
and U14919 (N_14919,N_14783,N_14810);
xor U14920 (N_14920,N_14799,N_14779);
and U14921 (N_14921,N_14825,N_14845);
or U14922 (N_14922,N_14715,N_14742);
nor U14923 (N_14923,N_14816,N_14790);
xor U14924 (N_14924,N_14763,N_14774);
xor U14925 (N_14925,N_14771,N_14794);
and U14926 (N_14926,N_14837,N_14702);
or U14927 (N_14927,N_14792,N_14843);
xnor U14928 (N_14928,N_14823,N_14724);
and U14929 (N_14929,N_14824,N_14810);
or U14930 (N_14930,N_14765,N_14716);
or U14931 (N_14931,N_14791,N_14839);
nand U14932 (N_14932,N_14742,N_14724);
or U14933 (N_14933,N_14733,N_14703);
xnor U14934 (N_14934,N_14836,N_14847);
or U14935 (N_14935,N_14791,N_14785);
or U14936 (N_14936,N_14823,N_14705);
nand U14937 (N_14937,N_14746,N_14795);
and U14938 (N_14938,N_14756,N_14841);
nand U14939 (N_14939,N_14790,N_14776);
or U14940 (N_14940,N_14775,N_14808);
xor U14941 (N_14941,N_14703,N_14715);
xor U14942 (N_14942,N_14783,N_14773);
xor U14943 (N_14943,N_14808,N_14776);
nor U14944 (N_14944,N_14826,N_14711);
xnor U14945 (N_14945,N_14776,N_14778);
and U14946 (N_14946,N_14768,N_14730);
or U14947 (N_14947,N_14812,N_14837);
nor U14948 (N_14948,N_14716,N_14806);
and U14949 (N_14949,N_14832,N_14740);
xnor U14950 (N_14950,N_14793,N_14751);
nand U14951 (N_14951,N_14755,N_14761);
nor U14952 (N_14952,N_14731,N_14736);
nor U14953 (N_14953,N_14756,N_14740);
xor U14954 (N_14954,N_14704,N_14757);
and U14955 (N_14955,N_14740,N_14806);
xnor U14956 (N_14956,N_14717,N_14718);
or U14957 (N_14957,N_14843,N_14752);
and U14958 (N_14958,N_14715,N_14810);
or U14959 (N_14959,N_14769,N_14714);
xor U14960 (N_14960,N_14827,N_14718);
nand U14961 (N_14961,N_14845,N_14743);
nor U14962 (N_14962,N_14809,N_14719);
nor U14963 (N_14963,N_14716,N_14700);
xnor U14964 (N_14964,N_14721,N_14737);
or U14965 (N_14965,N_14749,N_14818);
nor U14966 (N_14966,N_14827,N_14720);
and U14967 (N_14967,N_14753,N_14818);
nand U14968 (N_14968,N_14799,N_14787);
or U14969 (N_14969,N_14707,N_14848);
nand U14970 (N_14970,N_14726,N_14802);
nor U14971 (N_14971,N_14704,N_14830);
xor U14972 (N_14972,N_14842,N_14834);
or U14973 (N_14973,N_14717,N_14774);
xnor U14974 (N_14974,N_14716,N_14825);
or U14975 (N_14975,N_14834,N_14770);
nand U14976 (N_14976,N_14733,N_14788);
or U14977 (N_14977,N_14784,N_14808);
and U14978 (N_14978,N_14847,N_14704);
and U14979 (N_14979,N_14847,N_14832);
nor U14980 (N_14980,N_14767,N_14749);
nor U14981 (N_14981,N_14764,N_14756);
or U14982 (N_14982,N_14722,N_14798);
nand U14983 (N_14983,N_14826,N_14748);
nor U14984 (N_14984,N_14754,N_14824);
and U14985 (N_14985,N_14753,N_14712);
and U14986 (N_14986,N_14794,N_14819);
or U14987 (N_14987,N_14841,N_14754);
or U14988 (N_14988,N_14808,N_14701);
nor U14989 (N_14989,N_14848,N_14731);
and U14990 (N_14990,N_14726,N_14811);
nand U14991 (N_14991,N_14835,N_14848);
nor U14992 (N_14992,N_14801,N_14769);
nor U14993 (N_14993,N_14734,N_14716);
and U14994 (N_14994,N_14740,N_14834);
nand U14995 (N_14995,N_14742,N_14743);
nor U14996 (N_14996,N_14768,N_14760);
nand U14997 (N_14997,N_14702,N_14785);
nand U14998 (N_14998,N_14816,N_14767);
or U14999 (N_14999,N_14761,N_14751);
or UO_0 (O_0,N_14892,N_14986);
nand UO_1 (O_1,N_14999,N_14995);
xor UO_2 (O_2,N_14926,N_14988);
and UO_3 (O_3,N_14877,N_14985);
or UO_4 (O_4,N_14897,N_14982);
xor UO_5 (O_5,N_14972,N_14946);
and UO_6 (O_6,N_14851,N_14886);
or UO_7 (O_7,N_14983,N_14978);
nor UO_8 (O_8,N_14887,N_14980);
nand UO_9 (O_9,N_14992,N_14885);
and UO_10 (O_10,N_14975,N_14915);
and UO_11 (O_11,N_14906,N_14940);
xor UO_12 (O_12,N_14894,N_14949);
or UO_13 (O_13,N_14878,N_14909);
and UO_14 (O_14,N_14908,N_14859);
nand UO_15 (O_15,N_14873,N_14930);
xor UO_16 (O_16,N_14854,N_14962);
or UO_17 (O_17,N_14852,N_14967);
nand UO_18 (O_18,N_14900,N_14960);
xnor UO_19 (O_19,N_14958,N_14903);
or UO_20 (O_20,N_14996,N_14914);
xnor UO_21 (O_21,N_14884,N_14876);
and UO_22 (O_22,N_14959,N_14923);
or UO_23 (O_23,N_14860,N_14969);
and UO_24 (O_24,N_14895,N_14905);
xnor UO_25 (O_25,N_14870,N_14868);
nand UO_26 (O_26,N_14856,N_14997);
xor UO_27 (O_27,N_14981,N_14970);
nor UO_28 (O_28,N_14998,N_14932);
or UO_29 (O_29,N_14866,N_14971);
and UO_30 (O_30,N_14936,N_14913);
nand UO_31 (O_31,N_14979,N_14910);
xnor UO_32 (O_32,N_14948,N_14867);
and UO_33 (O_33,N_14955,N_14974);
xor UO_34 (O_34,N_14987,N_14991);
xnor UO_35 (O_35,N_14963,N_14850);
or UO_36 (O_36,N_14920,N_14916);
or UO_37 (O_37,N_14872,N_14950);
and UO_38 (O_38,N_14947,N_14954);
nor UO_39 (O_39,N_14862,N_14889);
xnor UO_40 (O_40,N_14935,N_14994);
nor UO_41 (O_41,N_14941,N_14888);
nand UO_42 (O_42,N_14939,N_14864);
or UO_43 (O_43,N_14976,N_14953);
nand UO_44 (O_44,N_14956,N_14928);
xor UO_45 (O_45,N_14890,N_14858);
nand UO_46 (O_46,N_14933,N_14945);
nor UO_47 (O_47,N_14904,N_14931);
or UO_48 (O_48,N_14977,N_14857);
xor UO_49 (O_49,N_14938,N_14925);
and UO_50 (O_50,N_14882,N_14961);
or UO_51 (O_51,N_14927,N_14891);
nand UO_52 (O_52,N_14896,N_14869);
or UO_53 (O_53,N_14861,N_14880);
and UO_54 (O_54,N_14943,N_14951);
or UO_55 (O_55,N_14973,N_14879);
or UO_56 (O_56,N_14901,N_14907);
nor UO_57 (O_57,N_14990,N_14965);
or UO_58 (O_58,N_14952,N_14853);
xnor UO_59 (O_59,N_14912,N_14929);
nand UO_60 (O_60,N_14898,N_14893);
nor UO_61 (O_61,N_14944,N_14865);
xnor UO_62 (O_62,N_14984,N_14871);
or UO_63 (O_63,N_14917,N_14881);
and UO_64 (O_64,N_14934,N_14968);
and UO_65 (O_65,N_14919,N_14911);
nor UO_66 (O_66,N_14902,N_14964);
nand UO_67 (O_67,N_14921,N_14989);
nor UO_68 (O_68,N_14937,N_14918);
nor UO_69 (O_69,N_14875,N_14863);
or UO_70 (O_70,N_14874,N_14899);
nor UO_71 (O_71,N_14966,N_14942);
or UO_72 (O_72,N_14957,N_14883);
nor UO_73 (O_73,N_14855,N_14924);
and UO_74 (O_74,N_14993,N_14922);
and UO_75 (O_75,N_14877,N_14963);
xnor UO_76 (O_76,N_14917,N_14955);
or UO_77 (O_77,N_14943,N_14940);
or UO_78 (O_78,N_14896,N_14979);
nand UO_79 (O_79,N_14861,N_14867);
or UO_80 (O_80,N_14986,N_14996);
or UO_81 (O_81,N_14966,N_14927);
or UO_82 (O_82,N_14851,N_14983);
nand UO_83 (O_83,N_14903,N_14963);
nor UO_84 (O_84,N_14893,N_14941);
nor UO_85 (O_85,N_14923,N_14951);
nor UO_86 (O_86,N_14999,N_14971);
or UO_87 (O_87,N_14862,N_14961);
xor UO_88 (O_88,N_14878,N_14882);
nor UO_89 (O_89,N_14870,N_14961);
and UO_90 (O_90,N_14904,N_14882);
and UO_91 (O_91,N_14969,N_14997);
nor UO_92 (O_92,N_14932,N_14948);
xor UO_93 (O_93,N_14854,N_14943);
nor UO_94 (O_94,N_14926,N_14995);
and UO_95 (O_95,N_14909,N_14944);
or UO_96 (O_96,N_14871,N_14937);
or UO_97 (O_97,N_14851,N_14970);
xnor UO_98 (O_98,N_14858,N_14884);
nor UO_99 (O_99,N_14860,N_14981);
nand UO_100 (O_100,N_14851,N_14978);
nand UO_101 (O_101,N_14991,N_14951);
and UO_102 (O_102,N_14948,N_14859);
nor UO_103 (O_103,N_14976,N_14872);
nand UO_104 (O_104,N_14871,N_14869);
and UO_105 (O_105,N_14964,N_14907);
nor UO_106 (O_106,N_14960,N_14991);
xor UO_107 (O_107,N_14934,N_14920);
nor UO_108 (O_108,N_14993,N_14975);
or UO_109 (O_109,N_14984,N_14853);
xnor UO_110 (O_110,N_14953,N_14889);
nor UO_111 (O_111,N_14974,N_14905);
nand UO_112 (O_112,N_14970,N_14859);
or UO_113 (O_113,N_14950,N_14946);
and UO_114 (O_114,N_14964,N_14912);
nor UO_115 (O_115,N_14955,N_14879);
and UO_116 (O_116,N_14899,N_14895);
or UO_117 (O_117,N_14887,N_14942);
or UO_118 (O_118,N_14877,N_14911);
or UO_119 (O_119,N_14881,N_14909);
nor UO_120 (O_120,N_14935,N_14992);
nand UO_121 (O_121,N_14982,N_14956);
or UO_122 (O_122,N_14949,N_14860);
nand UO_123 (O_123,N_14996,N_14942);
nor UO_124 (O_124,N_14882,N_14941);
xor UO_125 (O_125,N_14932,N_14879);
nand UO_126 (O_126,N_14965,N_14886);
or UO_127 (O_127,N_14908,N_14934);
or UO_128 (O_128,N_14967,N_14857);
nand UO_129 (O_129,N_14899,N_14985);
nor UO_130 (O_130,N_14894,N_14979);
xnor UO_131 (O_131,N_14899,N_14931);
or UO_132 (O_132,N_14943,N_14957);
or UO_133 (O_133,N_14951,N_14857);
or UO_134 (O_134,N_14961,N_14993);
nand UO_135 (O_135,N_14997,N_14987);
or UO_136 (O_136,N_14892,N_14851);
and UO_137 (O_137,N_14967,N_14863);
nor UO_138 (O_138,N_14879,N_14935);
and UO_139 (O_139,N_14938,N_14918);
xor UO_140 (O_140,N_14891,N_14956);
nand UO_141 (O_141,N_14949,N_14942);
nand UO_142 (O_142,N_14961,N_14984);
nor UO_143 (O_143,N_14972,N_14974);
xor UO_144 (O_144,N_14981,N_14902);
nand UO_145 (O_145,N_14896,N_14878);
or UO_146 (O_146,N_14892,N_14958);
or UO_147 (O_147,N_14894,N_14885);
xor UO_148 (O_148,N_14893,N_14951);
xnor UO_149 (O_149,N_14923,N_14913);
nor UO_150 (O_150,N_14985,N_14980);
xor UO_151 (O_151,N_14881,N_14918);
and UO_152 (O_152,N_14985,N_14894);
and UO_153 (O_153,N_14892,N_14954);
nor UO_154 (O_154,N_14960,N_14908);
nor UO_155 (O_155,N_14903,N_14906);
xnor UO_156 (O_156,N_14939,N_14858);
or UO_157 (O_157,N_14923,N_14895);
or UO_158 (O_158,N_14991,N_14920);
or UO_159 (O_159,N_14926,N_14989);
nand UO_160 (O_160,N_14960,N_14976);
nor UO_161 (O_161,N_14872,N_14961);
nand UO_162 (O_162,N_14998,N_14986);
or UO_163 (O_163,N_14897,N_14917);
nor UO_164 (O_164,N_14889,N_14867);
or UO_165 (O_165,N_14909,N_14886);
nor UO_166 (O_166,N_14891,N_14895);
or UO_167 (O_167,N_14922,N_14990);
nand UO_168 (O_168,N_14884,N_14956);
or UO_169 (O_169,N_14871,N_14996);
nor UO_170 (O_170,N_14961,N_14891);
nand UO_171 (O_171,N_14856,N_14890);
and UO_172 (O_172,N_14884,N_14932);
xnor UO_173 (O_173,N_14952,N_14907);
and UO_174 (O_174,N_14930,N_14950);
nand UO_175 (O_175,N_14957,N_14980);
xnor UO_176 (O_176,N_14985,N_14942);
and UO_177 (O_177,N_14924,N_14872);
or UO_178 (O_178,N_14895,N_14882);
nand UO_179 (O_179,N_14991,N_14899);
nand UO_180 (O_180,N_14853,N_14928);
or UO_181 (O_181,N_14923,N_14896);
nor UO_182 (O_182,N_14858,N_14949);
and UO_183 (O_183,N_14897,N_14895);
or UO_184 (O_184,N_14962,N_14996);
nor UO_185 (O_185,N_14869,N_14977);
or UO_186 (O_186,N_14951,N_14927);
and UO_187 (O_187,N_14949,N_14998);
and UO_188 (O_188,N_14916,N_14985);
xor UO_189 (O_189,N_14895,N_14983);
nor UO_190 (O_190,N_14965,N_14863);
and UO_191 (O_191,N_14904,N_14934);
and UO_192 (O_192,N_14892,N_14873);
nand UO_193 (O_193,N_14951,N_14850);
and UO_194 (O_194,N_14916,N_14922);
nand UO_195 (O_195,N_14870,N_14905);
nand UO_196 (O_196,N_14869,N_14870);
nor UO_197 (O_197,N_14900,N_14986);
nand UO_198 (O_198,N_14973,N_14869);
nor UO_199 (O_199,N_14919,N_14955);
or UO_200 (O_200,N_14925,N_14917);
xnor UO_201 (O_201,N_14855,N_14877);
nand UO_202 (O_202,N_14929,N_14867);
xor UO_203 (O_203,N_14860,N_14882);
or UO_204 (O_204,N_14901,N_14905);
or UO_205 (O_205,N_14856,N_14854);
xor UO_206 (O_206,N_14948,N_14922);
or UO_207 (O_207,N_14883,N_14934);
and UO_208 (O_208,N_14928,N_14951);
xor UO_209 (O_209,N_14916,N_14994);
and UO_210 (O_210,N_14922,N_14979);
nor UO_211 (O_211,N_14984,N_14898);
or UO_212 (O_212,N_14913,N_14880);
xor UO_213 (O_213,N_14958,N_14973);
or UO_214 (O_214,N_14857,N_14978);
or UO_215 (O_215,N_14930,N_14865);
or UO_216 (O_216,N_14982,N_14880);
and UO_217 (O_217,N_14948,N_14944);
nand UO_218 (O_218,N_14855,N_14853);
or UO_219 (O_219,N_14987,N_14979);
xnor UO_220 (O_220,N_14966,N_14861);
nor UO_221 (O_221,N_14917,N_14995);
xnor UO_222 (O_222,N_14910,N_14965);
or UO_223 (O_223,N_14860,N_14945);
nor UO_224 (O_224,N_14930,N_14986);
nand UO_225 (O_225,N_14978,N_14907);
xnor UO_226 (O_226,N_14940,N_14983);
nand UO_227 (O_227,N_14876,N_14971);
xor UO_228 (O_228,N_14901,N_14992);
or UO_229 (O_229,N_14959,N_14871);
nor UO_230 (O_230,N_14990,N_14930);
nor UO_231 (O_231,N_14912,N_14907);
and UO_232 (O_232,N_14891,N_14877);
and UO_233 (O_233,N_14955,N_14929);
nand UO_234 (O_234,N_14910,N_14963);
nor UO_235 (O_235,N_14868,N_14950);
and UO_236 (O_236,N_14902,N_14865);
nand UO_237 (O_237,N_14994,N_14871);
xnor UO_238 (O_238,N_14985,N_14961);
nand UO_239 (O_239,N_14930,N_14895);
xnor UO_240 (O_240,N_14984,N_14986);
xnor UO_241 (O_241,N_14925,N_14939);
nor UO_242 (O_242,N_14892,N_14991);
or UO_243 (O_243,N_14927,N_14920);
or UO_244 (O_244,N_14883,N_14984);
nor UO_245 (O_245,N_14942,N_14948);
nor UO_246 (O_246,N_14889,N_14876);
xnor UO_247 (O_247,N_14955,N_14965);
xnor UO_248 (O_248,N_14922,N_14878);
or UO_249 (O_249,N_14972,N_14985);
and UO_250 (O_250,N_14895,N_14904);
nor UO_251 (O_251,N_14854,N_14980);
nor UO_252 (O_252,N_14868,N_14968);
or UO_253 (O_253,N_14914,N_14857);
nand UO_254 (O_254,N_14995,N_14984);
xnor UO_255 (O_255,N_14889,N_14908);
and UO_256 (O_256,N_14864,N_14994);
nand UO_257 (O_257,N_14936,N_14889);
and UO_258 (O_258,N_14871,N_14974);
and UO_259 (O_259,N_14981,N_14850);
or UO_260 (O_260,N_14906,N_14961);
nand UO_261 (O_261,N_14868,N_14872);
or UO_262 (O_262,N_14926,N_14943);
and UO_263 (O_263,N_14930,N_14948);
nor UO_264 (O_264,N_14939,N_14877);
and UO_265 (O_265,N_14920,N_14895);
and UO_266 (O_266,N_14861,N_14958);
nand UO_267 (O_267,N_14886,N_14994);
nand UO_268 (O_268,N_14867,N_14931);
nand UO_269 (O_269,N_14992,N_14944);
nor UO_270 (O_270,N_14933,N_14858);
and UO_271 (O_271,N_14926,N_14932);
and UO_272 (O_272,N_14867,N_14961);
and UO_273 (O_273,N_14863,N_14893);
nor UO_274 (O_274,N_14937,N_14892);
xnor UO_275 (O_275,N_14905,N_14906);
xnor UO_276 (O_276,N_14866,N_14929);
nand UO_277 (O_277,N_14968,N_14875);
nand UO_278 (O_278,N_14901,N_14865);
nor UO_279 (O_279,N_14935,N_14859);
or UO_280 (O_280,N_14969,N_14948);
nor UO_281 (O_281,N_14983,N_14889);
nand UO_282 (O_282,N_14899,N_14888);
or UO_283 (O_283,N_14919,N_14988);
or UO_284 (O_284,N_14900,N_14918);
nand UO_285 (O_285,N_14959,N_14983);
xnor UO_286 (O_286,N_14890,N_14916);
xor UO_287 (O_287,N_14868,N_14951);
and UO_288 (O_288,N_14944,N_14981);
and UO_289 (O_289,N_14922,N_14857);
xor UO_290 (O_290,N_14904,N_14987);
nand UO_291 (O_291,N_14853,N_14923);
and UO_292 (O_292,N_14946,N_14882);
xor UO_293 (O_293,N_14857,N_14874);
or UO_294 (O_294,N_14878,N_14875);
nor UO_295 (O_295,N_14888,N_14996);
xnor UO_296 (O_296,N_14937,N_14855);
xor UO_297 (O_297,N_14949,N_14940);
nand UO_298 (O_298,N_14850,N_14969);
or UO_299 (O_299,N_14885,N_14948);
or UO_300 (O_300,N_14896,N_14930);
or UO_301 (O_301,N_14993,N_14980);
nor UO_302 (O_302,N_14962,N_14991);
and UO_303 (O_303,N_14948,N_14857);
nor UO_304 (O_304,N_14996,N_14931);
and UO_305 (O_305,N_14852,N_14937);
nand UO_306 (O_306,N_14942,N_14852);
xnor UO_307 (O_307,N_14856,N_14960);
or UO_308 (O_308,N_14889,N_14892);
nand UO_309 (O_309,N_14962,N_14915);
xor UO_310 (O_310,N_14978,N_14935);
and UO_311 (O_311,N_14934,N_14984);
nor UO_312 (O_312,N_14947,N_14921);
or UO_313 (O_313,N_14916,N_14941);
or UO_314 (O_314,N_14974,N_14897);
and UO_315 (O_315,N_14949,N_14960);
xor UO_316 (O_316,N_14921,N_14887);
and UO_317 (O_317,N_14890,N_14973);
or UO_318 (O_318,N_14963,N_14990);
nand UO_319 (O_319,N_14948,N_14884);
nand UO_320 (O_320,N_14935,N_14997);
or UO_321 (O_321,N_14860,N_14913);
nand UO_322 (O_322,N_14926,N_14913);
nand UO_323 (O_323,N_14944,N_14910);
nor UO_324 (O_324,N_14861,N_14924);
nand UO_325 (O_325,N_14936,N_14981);
or UO_326 (O_326,N_14862,N_14863);
xnor UO_327 (O_327,N_14943,N_14920);
nor UO_328 (O_328,N_14962,N_14992);
xnor UO_329 (O_329,N_14974,N_14919);
and UO_330 (O_330,N_14958,N_14930);
and UO_331 (O_331,N_14882,N_14899);
xor UO_332 (O_332,N_14918,N_14855);
or UO_333 (O_333,N_14921,N_14892);
or UO_334 (O_334,N_14898,N_14995);
or UO_335 (O_335,N_14983,N_14898);
nand UO_336 (O_336,N_14935,N_14955);
nor UO_337 (O_337,N_14925,N_14898);
nand UO_338 (O_338,N_14993,N_14920);
or UO_339 (O_339,N_14918,N_14892);
nand UO_340 (O_340,N_14960,N_14946);
nand UO_341 (O_341,N_14900,N_14944);
or UO_342 (O_342,N_14937,N_14912);
nand UO_343 (O_343,N_14955,N_14995);
and UO_344 (O_344,N_14878,N_14873);
xnor UO_345 (O_345,N_14971,N_14850);
xor UO_346 (O_346,N_14961,N_14962);
nand UO_347 (O_347,N_14859,N_14876);
and UO_348 (O_348,N_14973,N_14974);
nand UO_349 (O_349,N_14909,N_14859);
xor UO_350 (O_350,N_14951,N_14880);
and UO_351 (O_351,N_14943,N_14859);
and UO_352 (O_352,N_14906,N_14994);
and UO_353 (O_353,N_14916,N_14935);
nor UO_354 (O_354,N_14879,N_14863);
and UO_355 (O_355,N_14957,N_14996);
nand UO_356 (O_356,N_14963,N_14895);
nand UO_357 (O_357,N_14975,N_14992);
nor UO_358 (O_358,N_14953,N_14900);
xor UO_359 (O_359,N_14933,N_14865);
nand UO_360 (O_360,N_14955,N_14947);
and UO_361 (O_361,N_14912,N_14985);
or UO_362 (O_362,N_14950,N_14889);
nor UO_363 (O_363,N_14956,N_14911);
xnor UO_364 (O_364,N_14861,N_14988);
xnor UO_365 (O_365,N_14979,N_14999);
or UO_366 (O_366,N_14971,N_14944);
nand UO_367 (O_367,N_14970,N_14871);
nor UO_368 (O_368,N_14863,N_14914);
nor UO_369 (O_369,N_14893,N_14860);
or UO_370 (O_370,N_14902,N_14854);
or UO_371 (O_371,N_14856,N_14932);
and UO_372 (O_372,N_14962,N_14988);
nand UO_373 (O_373,N_14956,N_14960);
xnor UO_374 (O_374,N_14970,N_14969);
xor UO_375 (O_375,N_14912,N_14872);
nand UO_376 (O_376,N_14884,N_14879);
nand UO_377 (O_377,N_14915,N_14977);
and UO_378 (O_378,N_14938,N_14889);
xor UO_379 (O_379,N_14858,N_14997);
nand UO_380 (O_380,N_14862,N_14948);
nand UO_381 (O_381,N_14971,N_14889);
nand UO_382 (O_382,N_14861,N_14900);
or UO_383 (O_383,N_14861,N_14906);
or UO_384 (O_384,N_14918,N_14916);
xor UO_385 (O_385,N_14989,N_14920);
and UO_386 (O_386,N_14906,N_14960);
and UO_387 (O_387,N_14948,N_14929);
xor UO_388 (O_388,N_14890,N_14918);
and UO_389 (O_389,N_14894,N_14905);
and UO_390 (O_390,N_14966,N_14997);
and UO_391 (O_391,N_14904,N_14920);
nand UO_392 (O_392,N_14871,N_14898);
nor UO_393 (O_393,N_14997,N_14957);
xnor UO_394 (O_394,N_14877,N_14996);
nor UO_395 (O_395,N_14889,N_14967);
nor UO_396 (O_396,N_14961,N_14950);
nand UO_397 (O_397,N_14870,N_14883);
xor UO_398 (O_398,N_14880,N_14888);
nand UO_399 (O_399,N_14912,N_14984);
xor UO_400 (O_400,N_14851,N_14929);
or UO_401 (O_401,N_14856,N_14957);
or UO_402 (O_402,N_14883,N_14911);
or UO_403 (O_403,N_14891,N_14957);
xor UO_404 (O_404,N_14872,N_14891);
xnor UO_405 (O_405,N_14978,N_14917);
xnor UO_406 (O_406,N_14934,N_14959);
nand UO_407 (O_407,N_14979,N_14928);
nor UO_408 (O_408,N_14894,N_14941);
or UO_409 (O_409,N_14889,N_14970);
and UO_410 (O_410,N_14858,N_14992);
and UO_411 (O_411,N_14903,N_14868);
nor UO_412 (O_412,N_14986,N_14890);
nor UO_413 (O_413,N_14929,N_14998);
or UO_414 (O_414,N_14975,N_14896);
and UO_415 (O_415,N_14859,N_14889);
nand UO_416 (O_416,N_14946,N_14964);
and UO_417 (O_417,N_14949,N_14990);
and UO_418 (O_418,N_14916,N_14951);
xnor UO_419 (O_419,N_14992,N_14889);
nor UO_420 (O_420,N_14941,N_14901);
or UO_421 (O_421,N_14892,N_14931);
nand UO_422 (O_422,N_14865,N_14935);
nand UO_423 (O_423,N_14960,N_14994);
nand UO_424 (O_424,N_14964,N_14872);
nand UO_425 (O_425,N_14950,N_14967);
xor UO_426 (O_426,N_14976,N_14876);
nor UO_427 (O_427,N_14881,N_14955);
or UO_428 (O_428,N_14931,N_14942);
nand UO_429 (O_429,N_14876,N_14931);
nor UO_430 (O_430,N_14856,N_14913);
nor UO_431 (O_431,N_14877,N_14917);
or UO_432 (O_432,N_14926,N_14884);
nand UO_433 (O_433,N_14902,N_14861);
nor UO_434 (O_434,N_14995,N_14878);
or UO_435 (O_435,N_14984,N_14957);
xnor UO_436 (O_436,N_14911,N_14954);
or UO_437 (O_437,N_14885,N_14906);
or UO_438 (O_438,N_14856,N_14969);
nand UO_439 (O_439,N_14900,N_14911);
nand UO_440 (O_440,N_14888,N_14930);
and UO_441 (O_441,N_14872,N_14982);
nand UO_442 (O_442,N_14976,N_14966);
and UO_443 (O_443,N_14967,N_14926);
or UO_444 (O_444,N_14902,N_14903);
or UO_445 (O_445,N_14952,N_14968);
nand UO_446 (O_446,N_14973,N_14872);
nor UO_447 (O_447,N_14987,N_14892);
nor UO_448 (O_448,N_14873,N_14903);
xnor UO_449 (O_449,N_14900,N_14948);
nor UO_450 (O_450,N_14972,N_14927);
nor UO_451 (O_451,N_14929,N_14878);
xor UO_452 (O_452,N_14887,N_14865);
nor UO_453 (O_453,N_14853,N_14932);
and UO_454 (O_454,N_14954,N_14877);
or UO_455 (O_455,N_14964,N_14970);
and UO_456 (O_456,N_14987,N_14857);
and UO_457 (O_457,N_14996,N_14895);
and UO_458 (O_458,N_14867,N_14884);
nand UO_459 (O_459,N_14974,N_14900);
and UO_460 (O_460,N_14938,N_14958);
nor UO_461 (O_461,N_14893,N_14958);
nand UO_462 (O_462,N_14866,N_14979);
nor UO_463 (O_463,N_14959,N_14916);
or UO_464 (O_464,N_14931,N_14959);
xor UO_465 (O_465,N_14939,N_14878);
nor UO_466 (O_466,N_14864,N_14919);
xor UO_467 (O_467,N_14914,N_14904);
and UO_468 (O_468,N_14947,N_14863);
xor UO_469 (O_469,N_14917,N_14905);
nor UO_470 (O_470,N_14883,N_14859);
nor UO_471 (O_471,N_14893,N_14980);
nor UO_472 (O_472,N_14944,N_14987);
xnor UO_473 (O_473,N_14867,N_14928);
and UO_474 (O_474,N_14957,N_14897);
nor UO_475 (O_475,N_14901,N_14967);
and UO_476 (O_476,N_14986,N_14912);
nor UO_477 (O_477,N_14891,N_14932);
nor UO_478 (O_478,N_14997,N_14878);
nand UO_479 (O_479,N_14996,N_14990);
nand UO_480 (O_480,N_14861,N_14892);
xnor UO_481 (O_481,N_14859,N_14994);
and UO_482 (O_482,N_14957,N_14940);
nor UO_483 (O_483,N_14861,N_14852);
xnor UO_484 (O_484,N_14908,N_14854);
nor UO_485 (O_485,N_14858,N_14913);
nand UO_486 (O_486,N_14912,N_14997);
or UO_487 (O_487,N_14952,N_14970);
nor UO_488 (O_488,N_14888,N_14972);
xnor UO_489 (O_489,N_14891,N_14993);
nor UO_490 (O_490,N_14939,N_14903);
xnor UO_491 (O_491,N_14997,N_14890);
nand UO_492 (O_492,N_14852,N_14907);
and UO_493 (O_493,N_14904,N_14955);
nor UO_494 (O_494,N_14978,N_14928);
nand UO_495 (O_495,N_14875,N_14862);
nand UO_496 (O_496,N_14850,N_14860);
xor UO_497 (O_497,N_14909,N_14974);
xor UO_498 (O_498,N_14975,N_14879);
nor UO_499 (O_499,N_14914,N_14954);
or UO_500 (O_500,N_14916,N_14924);
nand UO_501 (O_501,N_14929,N_14962);
nor UO_502 (O_502,N_14862,N_14855);
xor UO_503 (O_503,N_14943,N_14988);
and UO_504 (O_504,N_14976,N_14933);
nor UO_505 (O_505,N_14873,N_14995);
and UO_506 (O_506,N_14907,N_14869);
and UO_507 (O_507,N_14910,N_14957);
xor UO_508 (O_508,N_14999,N_14902);
and UO_509 (O_509,N_14992,N_14904);
and UO_510 (O_510,N_14928,N_14919);
and UO_511 (O_511,N_14965,N_14963);
and UO_512 (O_512,N_14914,N_14949);
nand UO_513 (O_513,N_14902,N_14882);
or UO_514 (O_514,N_14900,N_14945);
or UO_515 (O_515,N_14926,N_14859);
and UO_516 (O_516,N_14992,N_14902);
and UO_517 (O_517,N_14870,N_14882);
and UO_518 (O_518,N_14916,N_14986);
and UO_519 (O_519,N_14892,N_14865);
nor UO_520 (O_520,N_14873,N_14883);
and UO_521 (O_521,N_14924,N_14900);
or UO_522 (O_522,N_14850,N_14901);
nor UO_523 (O_523,N_14913,N_14998);
nor UO_524 (O_524,N_14974,N_14881);
nand UO_525 (O_525,N_14865,N_14889);
nand UO_526 (O_526,N_14965,N_14991);
xnor UO_527 (O_527,N_14925,N_14890);
xnor UO_528 (O_528,N_14885,N_14924);
xnor UO_529 (O_529,N_14926,N_14982);
and UO_530 (O_530,N_14912,N_14918);
and UO_531 (O_531,N_14905,N_14879);
xnor UO_532 (O_532,N_14974,N_14983);
xor UO_533 (O_533,N_14927,N_14947);
xor UO_534 (O_534,N_14917,N_14967);
and UO_535 (O_535,N_14882,N_14876);
xnor UO_536 (O_536,N_14995,N_14862);
nand UO_537 (O_537,N_14981,N_14874);
and UO_538 (O_538,N_14958,N_14920);
and UO_539 (O_539,N_14850,N_14869);
or UO_540 (O_540,N_14959,N_14940);
xnor UO_541 (O_541,N_14876,N_14998);
nor UO_542 (O_542,N_14861,N_14956);
and UO_543 (O_543,N_14887,N_14945);
or UO_544 (O_544,N_14925,N_14906);
xor UO_545 (O_545,N_14976,N_14850);
or UO_546 (O_546,N_14974,N_14993);
xnor UO_547 (O_547,N_14911,N_14995);
xnor UO_548 (O_548,N_14893,N_14919);
or UO_549 (O_549,N_14960,N_14876);
and UO_550 (O_550,N_14970,N_14856);
nor UO_551 (O_551,N_14917,N_14982);
nand UO_552 (O_552,N_14890,N_14920);
nor UO_553 (O_553,N_14897,N_14900);
and UO_554 (O_554,N_14966,N_14961);
or UO_555 (O_555,N_14884,N_14998);
nand UO_556 (O_556,N_14856,N_14877);
nand UO_557 (O_557,N_14992,N_14995);
and UO_558 (O_558,N_14917,N_14972);
nor UO_559 (O_559,N_14997,N_14962);
nand UO_560 (O_560,N_14945,N_14976);
nor UO_561 (O_561,N_14955,N_14928);
nor UO_562 (O_562,N_14881,N_14896);
nand UO_563 (O_563,N_14951,N_14965);
and UO_564 (O_564,N_14942,N_14925);
and UO_565 (O_565,N_14943,N_14882);
nand UO_566 (O_566,N_14865,N_14999);
nor UO_567 (O_567,N_14976,N_14956);
nor UO_568 (O_568,N_14991,N_14977);
or UO_569 (O_569,N_14879,N_14907);
and UO_570 (O_570,N_14996,N_14894);
or UO_571 (O_571,N_14922,N_14898);
or UO_572 (O_572,N_14959,N_14928);
and UO_573 (O_573,N_14923,N_14866);
and UO_574 (O_574,N_14961,N_14910);
xnor UO_575 (O_575,N_14967,N_14958);
and UO_576 (O_576,N_14859,N_14996);
nand UO_577 (O_577,N_14868,N_14883);
xor UO_578 (O_578,N_14954,N_14915);
and UO_579 (O_579,N_14968,N_14900);
nor UO_580 (O_580,N_14911,N_14945);
nand UO_581 (O_581,N_14935,N_14899);
or UO_582 (O_582,N_14936,N_14892);
nor UO_583 (O_583,N_14946,N_14945);
nor UO_584 (O_584,N_14893,N_14916);
nor UO_585 (O_585,N_14956,N_14880);
and UO_586 (O_586,N_14970,N_14995);
xnor UO_587 (O_587,N_14850,N_14949);
and UO_588 (O_588,N_14978,N_14998);
nor UO_589 (O_589,N_14912,N_14978);
nand UO_590 (O_590,N_14934,N_14994);
xor UO_591 (O_591,N_14925,N_14964);
or UO_592 (O_592,N_14933,N_14869);
nor UO_593 (O_593,N_14961,N_14967);
xnor UO_594 (O_594,N_14990,N_14903);
and UO_595 (O_595,N_14917,N_14930);
nand UO_596 (O_596,N_14859,N_14964);
and UO_597 (O_597,N_14858,N_14934);
and UO_598 (O_598,N_14859,N_14898);
and UO_599 (O_599,N_14950,N_14944);
or UO_600 (O_600,N_14961,N_14957);
nor UO_601 (O_601,N_14884,N_14901);
nor UO_602 (O_602,N_14854,N_14993);
xnor UO_603 (O_603,N_14970,N_14867);
or UO_604 (O_604,N_14949,N_14890);
xnor UO_605 (O_605,N_14923,N_14967);
nor UO_606 (O_606,N_14950,N_14974);
nand UO_607 (O_607,N_14873,N_14871);
or UO_608 (O_608,N_14940,N_14860);
xor UO_609 (O_609,N_14962,N_14873);
and UO_610 (O_610,N_14862,N_14932);
and UO_611 (O_611,N_14895,N_14911);
nand UO_612 (O_612,N_14980,N_14964);
or UO_613 (O_613,N_14934,N_14860);
nor UO_614 (O_614,N_14902,N_14993);
nor UO_615 (O_615,N_14975,N_14874);
xnor UO_616 (O_616,N_14854,N_14938);
and UO_617 (O_617,N_14969,N_14893);
xnor UO_618 (O_618,N_14921,N_14960);
xnor UO_619 (O_619,N_14917,N_14862);
nand UO_620 (O_620,N_14903,N_14922);
nand UO_621 (O_621,N_14913,N_14990);
and UO_622 (O_622,N_14887,N_14960);
nand UO_623 (O_623,N_14967,N_14983);
or UO_624 (O_624,N_14974,N_14924);
and UO_625 (O_625,N_14958,N_14950);
xor UO_626 (O_626,N_14980,N_14919);
nor UO_627 (O_627,N_14974,N_14874);
xnor UO_628 (O_628,N_14912,N_14909);
or UO_629 (O_629,N_14978,N_14880);
xor UO_630 (O_630,N_14877,N_14906);
or UO_631 (O_631,N_14938,N_14879);
and UO_632 (O_632,N_14894,N_14968);
and UO_633 (O_633,N_14974,N_14995);
nor UO_634 (O_634,N_14971,N_14968);
or UO_635 (O_635,N_14938,N_14940);
nor UO_636 (O_636,N_14874,N_14852);
and UO_637 (O_637,N_14942,N_14970);
nand UO_638 (O_638,N_14953,N_14999);
and UO_639 (O_639,N_14951,N_14971);
nand UO_640 (O_640,N_14968,N_14927);
and UO_641 (O_641,N_14977,N_14962);
or UO_642 (O_642,N_14903,N_14852);
nor UO_643 (O_643,N_14927,N_14885);
nand UO_644 (O_644,N_14920,N_14957);
nor UO_645 (O_645,N_14989,N_14889);
and UO_646 (O_646,N_14898,N_14882);
xnor UO_647 (O_647,N_14887,N_14948);
nor UO_648 (O_648,N_14992,N_14896);
nand UO_649 (O_649,N_14944,N_14853);
xor UO_650 (O_650,N_14933,N_14982);
nor UO_651 (O_651,N_14940,N_14979);
or UO_652 (O_652,N_14982,N_14860);
and UO_653 (O_653,N_14963,N_14904);
nor UO_654 (O_654,N_14933,N_14907);
nor UO_655 (O_655,N_14979,N_14963);
or UO_656 (O_656,N_14948,N_14973);
nand UO_657 (O_657,N_14988,N_14980);
nand UO_658 (O_658,N_14924,N_14896);
and UO_659 (O_659,N_14864,N_14933);
and UO_660 (O_660,N_14871,N_14927);
nand UO_661 (O_661,N_14935,N_14968);
nand UO_662 (O_662,N_14925,N_14994);
or UO_663 (O_663,N_14856,N_14947);
or UO_664 (O_664,N_14897,N_14869);
or UO_665 (O_665,N_14977,N_14873);
or UO_666 (O_666,N_14979,N_14937);
and UO_667 (O_667,N_14959,N_14979);
or UO_668 (O_668,N_14873,N_14897);
nand UO_669 (O_669,N_14927,N_14894);
xor UO_670 (O_670,N_14932,N_14929);
or UO_671 (O_671,N_14934,N_14917);
nand UO_672 (O_672,N_14970,N_14968);
nor UO_673 (O_673,N_14957,N_14939);
or UO_674 (O_674,N_14880,N_14983);
nor UO_675 (O_675,N_14933,N_14953);
or UO_676 (O_676,N_14977,N_14903);
nand UO_677 (O_677,N_14920,N_14896);
xor UO_678 (O_678,N_14880,N_14903);
nor UO_679 (O_679,N_14963,N_14865);
and UO_680 (O_680,N_14884,N_14945);
nand UO_681 (O_681,N_14856,N_14880);
or UO_682 (O_682,N_14991,N_14866);
nand UO_683 (O_683,N_14859,N_14990);
nand UO_684 (O_684,N_14981,N_14855);
or UO_685 (O_685,N_14905,N_14972);
nand UO_686 (O_686,N_14877,N_14935);
or UO_687 (O_687,N_14927,N_14907);
and UO_688 (O_688,N_14995,N_14954);
nor UO_689 (O_689,N_14901,N_14924);
or UO_690 (O_690,N_14874,N_14918);
or UO_691 (O_691,N_14881,N_14932);
or UO_692 (O_692,N_14931,N_14861);
nand UO_693 (O_693,N_14970,N_14927);
xor UO_694 (O_694,N_14915,N_14866);
or UO_695 (O_695,N_14890,N_14938);
or UO_696 (O_696,N_14851,N_14941);
and UO_697 (O_697,N_14942,N_14895);
nand UO_698 (O_698,N_14896,N_14990);
or UO_699 (O_699,N_14978,N_14942);
nand UO_700 (O_700,N_14930,N_14991);
or UO_701 (O_701,N_14954,N_14959);
nor UO_702 (O_702,N_14955,N_14903);
or UO_703 (O_703,N_14855,N_14957);
and UO_704 (O_704,N_14949,N_14897);
nand UO_705 (O_705,N_14928,N_14968);
xnor UO_706 (O_706,N_14938,N_14979);
or UO_707 (O_707,N_14929,N_14965);
nand UO_708 (O_708,N_14896,N_14925);
nand UO_709 (O_709,N_14917,N_14921);
and UO_710 (O_710,N_14951,N_14947);
xnor UO_711 (O_711,N_14920,N_14851);
xor UO_712 (O_712,N_14991,N_14912);
nand UO_713 (O_713,N_14949,N_14973);
nor UO_714 (O_714,N_14933,N_14909);
or UO_715 (O_715,N_14870,N_14886);
nand UO_716 (O_716,N_14921,N_14983);
nand UO_717 (O_717,N_14964,N_14904);
or UO_718 (O_718,N_14917,N_14891);
and UO_719 (O_719,N_14991,N_14908);
xnor UO_720 (O_720,N_14970,N_14908);
nor UO_721 (O_721,N_14991,N_14999);
nor UO_722 (O_722,N_14878,N_14960);
xnor UO_723 (O_723,N_14903,N_14874);
nor UO_724 (O_724,N_14997,N_14934);
or UO_725 (O_725,N_14909,N_14966);
and UO_726 (O_726,N_14873,N_14958);
or UO_727 (O_727,N_14978,N_14941);
xnor UO_728 (O_728,N_14935,N_14971);
nand UO_729 (O_729,N_14859,N_14995);
and UO_730 (O_730,N_14851,N_14874);
or UO_731 (O_731,N_14980,N_14933);
nor UO_732 (O_732,N_14926,N_14887);
nor UO_733 (O_733,N_14946,N_14953);
xnor UO_734 (O_734,N_14964,N_14889);
and UO_735 (O_735,N_14950,N_14853);
or UO_736 (O_736,N_14972,N_14914);
and UO_737 (O_737,N_14921,N_14994);
and UO_738 (O_738,N_14931,N_14966);
nor UO_739 (O_739,N_14929,N_14961);
xnor UO_740 (O_740,N_14997,N_14854);
nor UO_741 (O_741,N_14953,N_14940);
and UO_742 (O_742,N_14897,N_14973);
xor UO_743 (O_743,N_14978,N_14856);
or UO_744 (O_744,N_14983,N_14987);
xnor UO_745 (O_745,N_14933,N_14946);
xnor UO_746 (O_746,N_14907,N_14891);
or UO_747 (O_747,N_14976,N_14874);
xnor UO_748 (O_748,N_14913,N_14989);
xor UO_749 (O_749,N_14881,N_14927);
nand UO_750 (O_750,N_14877,N_14853);
nor UO_751 (O_751,N_14931,N_14989);
or UO_752 (O_752,N_14857,N_14991);
xor UO_753 (O_753,N_14936,N_14915);
or UO_754 (O_754,N_14930,N_14997);
and UO_755 (O_755,N_14901,N_14978);
xnor UO_756 (O_756,N_14957,N_14966);
and UO_757 (O_757,N_14957,N_14998);
nor UO_758 (O_758,N_14924,N_14943);
xor UO_759 (O_759,N_14963,N_14962);
nand UO_760 (O_760,N_14865,N_14953);
or UO_761 (O_761,N_14881,N_14850);
or UO_762 (O_762,N_14958,N_14872);
nand UO_763 (O_763,N_14909,N_14873);
and UO_764 (O_764,N_14867,N_14918);
or UO_765 (O_765,N_14964,N_14879);
xnor UO_766 (O_766,N_14997,N_14880);
xor UO_767 (O_767,N_14885,N_14873);
nor UO_768 (O_768,N_14920,N_14983);
or UO_769 (O_769,N_14852,N_14913);
nor UO_770 (O_770,N_14877,N_14982);
and UO_771 (O_771,N_14988,N_14878);
xnor UO_772 (O_772,N_14886,N_14957);
nor UO_773 (O_773,N_14957,N_14971);
and UO_774 (O_774,N_14924,N_14882);
xnor UO_775 (O_775,N_14941,N_14952);
nor UO_776 (O_776,N_14930,N_14960);
xnor UO_777 (O_777,N_14901,N_14936);
and UO_778 (O_778,N_14857,N_14873);
xor UO_779 (O_779,N_14971,N_14946);
and UO_780 (O_780,N_14993,N_14878);
nand UO_781 (O_781,N_14873,N_14884);
nor UO_782 (O_782,N_14938,N_14876);
xnor UO_783 (O_783,N_14893,N_14963);
or UO_784 (O_784,N_14991,N_14938);
and UO_785 (O_785,N_14920,N_14962);
and UO_786 (O_786,N_14897,N_14859);
nand UO_787 (O_787,N_14970,N_14949);
or UO_788 (O_788,N_14984,N_14943);
xor UO_789 (O_789,N_14993,N_14874);
nor UO_790 (O_790,N_14978,N_14913);
xnor UO_791 (O_791,N_14991,N_14996);
and UO_792 (O_792,N_14893,N_14971);
xnor UO_793 (O_793,N_14985,N_14979);
nand UO_794 (O_794,N_14989,N_14853);
nor UO_795 (O_795,N_14948,N_14939);
nor UO_796 (O_796,N_14937,N_14861);
xnor UO_797 (O_797,N_14893,N_14989);
nor UO_798 (O_798,N_14984,N_14930);
nor UO_799 (O_799,N_14854,N_14898);
and UO_800 (O_800,N_14883,N_14914);
and UO_801 (O_801,N_14866,N_14985);
and UO_802 (O_802,N_14936,N_14945);
nand UO_803 (O_803,N_14964,N_14906);
nand UO_804 (O_804,N_14925,N_14956);
nor UO_805 (O_805,N_14868,N_14905);
nand UO_806 (O_806,N_14931,N_14915);
or UO_807 (O_807,N_14960,N_14884);
or UO_808 (O_808,N_14886,N_14985);
or UO_809 (O_809,N_14878,N_14856);
xnor UO_810 (O_810,N_14867,N_14910);
and UO_811 (O_811,N_14922,N_14869);
xnor UO_812 (O_812,N_14999,N_14909);
nor UO_813 (O_813,N_14926,N_14907);
nand UO_814 (O_814,N_14985,N_14897);
nand UO_815 (O_815,N_14901,N_14916);
and UO_816 (O_816,N_14964,N_14895);
and UO_817 (O_817,N_14938,N_14944);
nand UO_818 (O_818,N_14889,N_14986);
or UO_819 (O_819,N_14995,N_14994);
xnor UO_820 (O_820,N_14868,N_14936);
or UO_821 (O_821,N_14908,N_14927);
xor UO_822 (O_822,N_14920,N_14862);
or UO_823 (O_823,N_14920,N_14866);
and UO_824 (O_824,N_14913,N_14981);
nand UO_825 (O_825,N_14983,N_14963);
nand UO_826 (O_826,N_14868,N_14939);
nor UO_827 (O_827,N_14987,N_14917);
xor UO_828 (O_828,N_14955,N_14898);
nand UO_829 (O_829,N_14990,N_14984);
or UO_830 (O_830,N_14950,N_14920);
nor UO_831 (O_831,N_14854,N_14866);
nor UO_832 (O_832,N_14986,N_14940);
xor UO_833 (O_833,N_14886,N_14885);
or UO_834 (O_834,N_14998,N_14900);
xnor UO_835 (O_835,N_14863,N_14889);
nand UO_836 (O_836,N_14917,N_14928);
and UO_837 (O_837,N_14873,N_14975);
and UO_838 (O_838,N_14926,N_14897);
nand UO_839 (O_839,N_14980,N_14952);
nor UO_840 (O_840,N_14886,N_14941);
nor UO_841 (O_841,N_14879,N_14855);
and UO_842 (O_842,N_14929,N_14899);
or UO_843 (O_843,N_14914,N_14908);
and UO_844 (O_844,N_14855,N_14851);
nor UO_845 (O_845,N_14980,N_14884);
or UO_846 (O_846,N_14984,N_14938);
or UO_847 (O_847,N_14855,N_14961);
nor UO_848 (O_848,N_14898,N_14993);
xor UO_849 (O_849,N_14908,N_14884);
nor UO_850 (O_850,N_14905,N_14860);
and UO_851 (O_851,N_14900,N_14985);
nor UO_852 (O_852,N_14920,N_14953);
and UO_853 (O_853,N_14875,N_14983);
and UO_854 (O_854,N_14967,N_14867);
and UO_855 (O_855,N_14991,N_14953);
nor UO_856 (O_856,N_14972,N_14898);
and UO_857 (O_857,N_14930,N_14913);
and UO_858 (O_858,N_14857,N_14963);
or UO_859 (O_859,N_14920,N_14898);
and UO_860 (O_860,N_14901,N_14986);
nand UO_861 (O_861,N_14968,N_14953);
nor UO_862 (O_862,N_14942,N_14896);
or UO_863 (O_863,N_14872,N_14937);
xor UO_864 (O_864,N_14877,N_14929);
and UO_865 (O_865,N_14993,N_14856);
xor UO_866 (O_866,N_14962,N_14899);
nand UO_867 (O_867,N_14975,N_14910);
and UO_868 (O_868,N_14977,N_14928);
nand UO_869 (O_869,N_14989,N_14950);
nand UO_870 (O_870,N_14919,N_14865);
xor UO_871 (O_871,N_14900,N_14866);
nor UO_872 (O_872,N_14950,N_14994);
nand UO_873 (O_873,N_14980,N_14905);
nor UO_874 (O_874,N_14868,N_14892);
nor UO_875 (O_875,N_14999,N_14959);
nor UO_876 (O_876,N_14861,N_14894);
xor UO_877 (O_877,N_14945,N_14956);
or UO_878 (O_878,N_14908,N_14928);
nor UO_879 (O_879,N_14884,N_14994);
xor UO_880 (O_880,N_14938,N_14917);
or UO_881 (O_881,N_14994,N_14959);
nor UO_882 (O_882,N_14876,N_14878);
xor UO_883 (O_883,N_14976,N_14926);
xnor UO_884 (O_884,N_14982,N_14890);
xor UO_885 (O_885,N_14925,N_14944);
nand UO_886 (O_886,N_14861,N_14870);
nor UO_887 (O_887,N_14865,N_14880);
nand UO_888 (O_888,N_14989,N_14900);
nand UO_889 (O_889,N_14908,N_14878);
nor UO_890 (O_890,N_14850,N_14952);
nor UO_891 (O_891,N_14904,N_14891);
and UO_892 (O_892,N_14927,N_14943);
or UO_893 (O_893,N_14869,N_14879);
or UO_894 (O_894,N_14877,N_14886);
nand UO_895 (O_895,N_14924,N_14852);
nand UO_896 (O_896,N_14857,N_14923);
nor UO_897 (O_897,N_14852,N_14954);
nor UO_898 (O_898,N_14874,N_14856);
nand UO_899 (O_899,N_14934,N_14938);
nand UO_900 (O_900,N_14946,N_14998);
and UO_901 (O_901,N_14956,N_14917);
xnor UO_902 (O_902,N_14915,N_14955);
xor UO_903 (O_903,N_14984,N_14866);
and UO_904 (O_904,N_14911,N_14943);
and UO_905 (O_905,N_14972,N_14891);
xnor UO_906 (O_906,N_14976,N_14962);
or UO_907 (O_907,N_14872,N_14944);
or UO_908 (O_908,N_14929,N_14939);
or UO_909 (O_909,N_14983,N_14935);
and UO_910 (O_910,N_14964,N_14967);
xnor UO_911 (O_911,N_14887,N_14992);
nor UO_912 (O_912,N_14947,N_14930);
and UO_913 (O_913,N_14943,N_14856);
nor UO_914 (O_914,N_14967,N_14979);
nand UO_915 (O_915,N_14859,N_14933);
and UO_916 (O_916,N_14910,N_14882);
and UO_917 (O_917,N_14918,N_14926);
nand UO_918 (O_918,N_14961,N_14894);
or UO_919 (O_919,N_14999,N_14931);
xor UO_920 (O_920,N_14920,N_14990);
and UO_921 (O_921,N_14958,N_14982);
nand UO_922 (O_922,N_14917,N_14964);
or UO_923 (O_923,N_14876,N_14902);
and UO_924 (O_924,N_14890,N_14927);
xnor UO_925 (O_925,N_14884,N_14854);
or UO_926 (O_926,N_14993,N_14910);
and UO_927 (O_927,N_14928,N_14937);
xor UO_928 (O_928,N_14956,N_14858);
or UO_929 (O_929,N_14884,N_14989);
or UO_930 (O_930,N_14894,N_14864);
nor UO_931 (O_931,N_14946,N_14872);
and UO_932 (O_932,N_14883,N_14916);
or UO_933 (O_933,N_14938,N_14993);
nor UO_934 (O_934,N_14931,N_14851);
or UO_935 (O_935,N_14913,N_14964);
nor UO_936 (O_936,N_14926,N_14850);
or UO_937 (O_937,N_14901,N_14990);
nand UO_938 (O_938,N_14998,N_14915);
and UO_939 (O_939,N_14870,N_14947);
nand UO_940 (O_940,N_14911,N_14896);
nor UO_941 (O_941,N_14887,N_14858);
nor UO_942 (O_942,N_14930,N_14853);
nand UO_943 (O_943,N_14969,N_14949);
xor UO_944 (O_944,N_14976,N_14854);
nor UO_945 (O_945,N_14892,N_14972);
nor UO_946 (O_946,N_14873,N_14986);
and UO_947 (O_947,N_14890,N_14893);
xnor UO_948 (O_948,N_14891,N_14945);
nand UO_949 (O_949,N_14991,N_14984);
or UO_950 (O_950,N_14919,N_14998);
nor UO_951 (O_951,N_14937,N_14962);
xnor UO_952 (O_952,N_14888,N_14874);
nor UO_953 (O_953,N_14999,N_14904);
and UO_954 (O_954,N_14912,N_14889);
nor UO_955 (O_955,N_14960,N_14880);
and UO_956 (O_956,N_14988,N_14870);
nand UO_957 (O_957,N_14939,N_14991);
nor UO_958 (O_958,N_14995,N_14883);
nor UO_959 (O_959,N_14905,N_14924);
xnor UO_960 (O_960,N_14947,N_14901);
nor UO_961 (O_961,N_14903,N_14986);
nand UO_962 (O_962,N_14945,N_14856);
nand UO_963 (O_963,N_14894,N_14851);
xnor UO_964 (O_964,N_14941,N_14968);
nand UO_965 (O_965,N_14868,N_14893);
or UO_966 (O_966,N_14991,N_14881);
xnor UO_967 (O_967,N_14915,N_14867);
nand UO_968 (O_968,N_14948,N_14923);
nor UO_969 (O_969,N_14926,N_14972);
nand UO_970 (O_970,N_14994,N_14856);
or UO_971 (O_971,N_14851,N_14986);
nand UO_972 (O_972,N_14929,N_14908);
and UO_973 (O_973,N_14866,N_14871);
nand UO_974 (O_974,N_14851,N_14955);
and UO_975 (O_975,N_14968,N_14994);
nor UO_976 (O_976,N_14874,N_14988);
and UO_977 (O_977,N_14989,N_14988);
xnor UO_978 (O_978,N_14882,N_14888);
or UO_979 (O_979,N_14872,N_14926);
nand UO_980 (O_980,N_14902,N_14985);
and UO_981 (O_981,N_14979,N_14878);
and UO_982 (O_982,N_14978,N_14954);
nor UO_983 (O_983,N_14940,N_14878);
xor UO_984 (O_984,N_14974,N_14920);
nand UO_985 (O_985,N_14943,N_14874);
or UO_986 (O_986,N_14871,N_14853);
xnor UO_987 (O_987,N_14934,N_14881);
and UO_988 (O_988,N_14998,N_14958);
or UO_989 (O_989,N_14995,N_14949);
or UO_990 (O_990,N_14930,N_14956);
or UO_991 (O_991,N_14925,N_14971);
or UO_992 (O_992,N_14937,N_14991);
xnor UO_993 (O_993,N_14980,N_14970);
or UO_994 (O_994,N_14941,N_14957);
or UO_995 (O_995,N_14887,N_14989);
nand UO_996 (O_996,N_14944,N_14965);
xnor UO_997 (O_997,N_14952,N_14940);
or UO_998 (O_998,N_14883,N_14875);
or UO_999 (O_999,N_14925,N_14977);
or UO_1000 (O_1000,N_14981,N_14857);
or UO_1001 (O_1001,N_14918,N_14923);
nand UO_1002 (O_1002,N_14874,N_14985);
or UO_1003 (O_1003,N_14987,N_14871);
or UO_1004 (O_1004,N_14916,N_14937);
or UO_1005 (O_1005,N_14861,N_14996);
nand UO_1006 (O_1006,N_14928,N_14868);
and UO_1007 (O_1007,N_14974,N_14864);
nand UO_1008 (O_1008,N_14869,N_14949);
nor UO_1009 (O_1009,N_14931,N_14929);
and UO_1010 (O_1010,N_14966,N_14988);
and UO_1011 (O_1011,N_14980,N_14900);
nor UO_1012 (O_1012,N_14864,N_14963);
xnor UO_1013 (O_1013,N_14878,N_14871);
or UO_1014 (O_1014,N_14905,N_14968);
and UO_1015 (O_1015,N_14865,N_14938);
and UO_1016 (O_1016,N_14956,N_14935);
nor UO_1017 (O_1017,N_14927,N_14868);
nor UO_1018 (O_1018,N_14916,N_14960);
or UO_1019 (O_1019,N_14895,N_14862);
nor UO_1020 (O_1020,N_14974,N_14970);
xnor UO_1021 (O_1021,N_14898,N_14880);
nor UO_1022 (O_1022,N_14965,N_14947);
nand UO_1023 (O_1023,N_14990,N_14880);
or UO_1024 (O_1024,N_14913,N_14872);
nor UO_1025 (O_1025,N_14866,N_14914);
nand UO_1026 (O_1026,N_14916,N_14936);
or UO_1027 (O_1027,N_14940,N_14937);
and UO_1028 (O_1028,N_14997,N_14906);
nor UO_1029 (O_1029,N_14871,N_14855);
xnor UO_1030 (O_1030,N_14922,N_14987);
nor UO_1031 (O_1031,N_14855,N_14872);
xor UO_1032 (O_1032,N_14987,N_14980);
nand UO_1033 (O_1033,N_14876,N_14928);
and UO_1034 (O_1034,N_14865,N_14989);
and UO_1035 (O_1035,N_14989,N_14881);
nand UO_1036 (O_1036,N_14875,N_14966);
or UO_1037 (O_1037,N_14931,N_14919);
nor UO_1038 (O_1038,N_14938,N_14892);
nor UO_1039 (O_1039,N_14908,N_14941);
xor UO_1040 (O_1040,N_14979,N_14885);
nor UO_1041 (O_1041,N_14926,N_14994);
or UO_1042 (O_1042,N_14865,N_14884);
or UO_1043 (O_1043,N_14854,N_14955);
xor UO_1044 (O_1044,N_14994,N_14887);
and UO_1045 (O_1045,N_14861,N_14961);
xnor UO_1046 (O_1046,N_14893,N_14929);
nor UO_1047 (O_1047,N_14931,N_14906);
nor UO_1048 (O_1048,N_14850,N_14858);
and UO_1049 (O_1049,N_14991,N_14972);
nor UO_1050 (O_1050,N_14975,N_14908);
and UO_1051 (O_1051,N_14939,N_14937);
xor UO_1052 (O_1052,N_14987,N_14925);
or UO_1053 (O_1053,N_14945,N_14941);
nor UO_1054 (O_1054,N_14970,N_14907);
xor UO_1055 (O_1055,N_14958,N_14974);
xnor UO_1056 (O_1056,N_14888,N_14933);
or UO_1057 (O_1057,N_14867,N_14858);
xor UO_1058 (O_1058,N_14903,N_14997);
or UO_1059 (O_1059,N_14852,N_14936);
and UO_1060 (O_1060,N_14869,N_14886);
nor UO_1061 (O_1061,N_14872,N_14880);
xnor UO_1062 (O_1062,N_14994,N_14941);
and UO_1063 (O_1063,N_14911,N_14990);
or UO_1064 (O_1064,N_14903,N_14901);
and UO_1065 (O_1065,N_14982,N_14927);
nand UO_1066 (O_1066,N_14888,N_14988);
xnor UO_1067 (O_1067,N_14915,N_14888);
or UO_1068 (O_1068,N_14943,N_14987);
nor UO_1069 (O_1069,N_14969,N_14979);
xnor UO_1070 (O_1070,N_14921,N_14936);
or UO_1071 (O_1071,N_14928,N_14966);
xnor UO_1072 (O_1072,N_14924,N_14956);
and UO_1073 (O_1073,N_14902,N_14901);
nor UO_1074 (O_1074,N_14959,N_14953);
and UO_1075 (O_1075,N_14930,N_14863);
nor UO_1076 (O_1076,N_14993,N_14865);
nor UO_1077 (O_1077,N_14887,N_14975);
xnor UO_1078 (O_1078,N_14973,N_14997);
and UO_1079 (O_1079,N_14944,N_14866);
and UO_1080 (O_1080,N_14883,N_14997);
and UO_1081 (O_1081,N_14961,N_14895);
nand UO_1082 (O_1082,N_14884,N_14963);
xnor UO_1083 (O_1083,N_14897,N_14909);
or UO_1084 (O_1084,N_14914,N_14951);
nor UO_1085 (O_1085,N_14906,N_14864);
nand UO_1086 (O_1086,N_14910,N_14992);
or UO_1087 (O_1087,N_14939,N_14919);
nor UO_1088 (O_1088,N_14994,N_14928);
or UO_1089 (O_1089,N_14974,N_14935);
nor UO_1090 (O_1090,N_14923,N_14862);
nand UO_1091 (O_1091,N_14935,N_14989);
nor UO_1092 (O_1092,N_14948,N_14926);
nor UO_1093 (O_1093,N_14957,N_14927);
nor UO_1094 (O_1094,N_14939,N_14927);
xor UO_1095 (O_1095,N_14975,N_14984);
or UO_1096 (O_1096,N_14890,N_14882);
and UO_1097 (O_1097,N_14875,N_14911);
or UO_1098 (O_1098,N_14920,N_14995);
and UO_1099 (O_1099,N_14883,N_14951);
nand UO_1100 (O_1100,N_14876,N_14989);
xnor UO_1101 (O_1101,N_14979,N_14911);
nor UO_1102 (O_1102,N_14921,N_14933);
xnor UO_1103 (O_1103,N_14863,N_14910);
and UO_1104 (O_1104,N_14863,N_14898);
nor UO_1105 (O_1105,N_14950,N_14982);
or UO_1106 (O_1106,N_14977,N_14893);
and UO_1107 (O_1107,N_14909,N_14962);
nand UO_1108 (O_1108,N_14974,N_14882);
xor UO_1109 (O_1109,N_14946,N_14884);
nand UO_1110 (O_1110,N_14965,N_14878);
and UO_1111 (O_1111,N_14956,N_14957);
xnor UO_1112 (O_1112,N_14920,N_14885);
nand UO_1113 (O_1113,N_14912,N_14993);
or UO_1114 (O_1114,N_14961,N_14859);
xor UO_1115 (O_1115,N_14902,N_14851);
or UO_1116 (O_1116,N_14866,N_14874);
nand UO_1117 (O_1117,N_14972,N_14910);
xor UO_1118 (O_1118,N_14879,N_14982);
nand UO_1119 (O_1119,N_14938,N_14956);
and UO_1120 (O_1120,N_14985,N_14876);
or UO_1121 (O_1121,N_14904,N_14877);
xnor UO_1122 (O_1122,N_14875,N_14953);
xnor UO_1123 (O_1123,N_14882,N_14893);
nand UO_1124 (O_1124,N_14873,N_14933);
nand UO_1125 (O_1125,N_14948,N_14912);
nor UO_1126 (O_1126,N_14943,N_14915);
and UO_1127 (O_1127,N_14912,N_14862);
and UO_1128 (O_1128,N_14882,N_14958);
xnor UO_1129 (O_1129,N_14922,N_14902);
nand UO_1130 (O_1130,N_14998,N_14872);
xor UO_1131 (O_1131,N_14997,N_14970);
and UO_1132 (O_1132,N_14880,N_14928);
and UO_1133 (O_1133,N_14946,N_14913);
or UO_1134 (O_1134,N_14873,N_14900);
or UO_1135 (O_1135,N_14898,N_14853);
and UO_1136 (O_1136,N_14909,N_14860);
nor UO_1137 (O_1137,N_14979,N_14913);
nor UO_1138 (O_1138,N_14907,N_14889);
or UO_1139 (O_1139,N_14859,N_14911);
nor UO_1140 (O_1140,N_14939,N_14886);
and UO_1141 (O_1141,N_14957,N_14970);
nor UO_1142 (O_1142,N_14882,N_14864);
and UO_1143 (O_1143,N_14928,N_14915);
or UO_1144 (O_1144,N_14918,N_14884);
and UO_1145 (O_1145,N_14933,N_14993);
or UO_1146 (O_1146,N_14896,N_14905);
xnor UO_1147 (O_1147,N_14920,N_14944);
or UO_1148 (O_1148,N_14972,N_14975);
or UO_1149 (O_1149,N_14948,N_14951);
or UO_1150 (O_1150,N_14951,N_14865);
xor UO_1151 (O_1151,N_14867,N_14859);
and UO_1152 (O_1152,N_14948,N_14940);
or UO_1153 (O_1153,N_14992,N_14928);
and UO_1154 (O_1154,N_14875,N_14985);
nor UO_1155 (O_1155,N_14874,N_14867);
and UO_1156 (O_1156,N_14968,N_14865);
xor UO_1157 (O_1157,N_14916,N_14865);
xnor UO_1158 (O_1158,N_14915,N_14978);
and UO_1159 (O_1159,N_14858,N_14903);
nor UO_1160 (O_1160,N_14901,N_14968);
nand UO_1161 (O_1161,N_14962,N_14979);
or UO_1162 (O_1162,N_14984,N_14857);
nand UO_1163 (O_1163,N_14895,N_14871);
and UO_1164 (O_1164,N_14883,N_14988);
nand UO_1165 (O_1165,N_14855,N_14869);
nand UO_1166 (O_1166,N_14877,N_14884);
or UO_1167 (O_1167,N_14950,N_14936);
xnor UO_1168 (O_1168,N_14956,N_14899);
xor UO_1169 (O_1169,N_14945,N_14867);
or UO_1170 (O_1170,N_14886,N_14871);
nand UO_1171 (O_1171,N_14933,N_14970);
and UO_1172 (O_1172,N_14986,N_14985);
xnor UO_1173 (O_1173,N_14876,N_14944);
xnor UO_1174 (O_1174,N_14853,N_14886);
nor UO_1175 (O_1175,N_14991,N_14913);
nor UO_1176 (O_1176,N_14890,N_14851);
and UO_1177 (O_1177,N_14979,N_14915);
and UO_1178 (O_1178,N_14876,N_14939);
or UO_1179 (O_1179,N_14863,N_14961);
xnor UO_1180 (O_1180,N_14928,N_14861);
or UO_1181 (O_1181,N_14995,N_14909);
or UO_1182 (O_1182,N_14960,N_14879);
nor UO_1183 (O_1183,N_14860,N_14929);
or UO_1184 (O_1184,N_14887,N_14889);
and UO_1185 (O_1185,N_14864,N_14914);
and UO_1186 (O_1186,N_14925,N_14892);
nor UO_1187 (O_1187,N_14975,N_14967);
nand UO_1188 (O_1188,N_14901,N_14870);
nand UO_1189 (O_1189,N_14864,N_14890);
nor UO_1190 (O_1190,N_14967,N_14998);
xnor UO_1191 (O_1191,N_14942,N_14891);
xnor UO_1192 (O_1192,N_14985,N_14915);
nor UO_1193 (O_1193,N_14910,N_14990);
nor UO_1194 (O_1194,N_14927,N_14960);
nor UO_1195 (O_1195,N_14921,N_14950);
or UO_1196 (O_1196,N_14965,N_14918);
and UO_1197 (O_1197,N_14925,N_14878);
or UO_1198 (O_1198,N_14923,N_14878);
or UO_1199 (O_1199,N_14961,N_14885);
and UO_1200 (O_1200,N_14994,N_14902);
nand UO_1201 (O_1201,N_14870,N_14893);
and UO_1202 (O_1202,N_14903,N_14883);
and UO_1203 (O_1203,N_14993,N_14862);
xnor UO_1204 (O_1204,N_14934,N_14894);
or UO_1205 (O_1205,N_14894,N_14955);
or UO_1206 (O_1206,N_14985,N_14920);
or UO_1207 (O_1207,N_14930,N_14976);
and UO_1208 (O_1208,N_14947,N_14992);
and UO_1209 (O_1209,N_14937,N_14982);
nand UO_1210 (O_1210,N_14936,N_14967);
nand UO_1211 (O_1211,N_14946,N_14853);
and UO_1212 (O_1212,N_14903,N_14953);
or UO_1213 (O_1213,N_14952,N_14953);
nand UO_1214 (O_1214,N_14959,N_14930);
xnor UO_1215 (O_1215,N_14907,N_14981);
and UO_1216 (O_1216,N_14901,N_14908);
xnor UO_1217 (O_1217,N_14910,N_14932);
and UO_1218 (O_1218,N_14923,N_14890);
nor UO_1219 (O_1219,N_14882,N_14884);
or UO_1220 (O_1220,N_14887,N_14892);
nor UO_1221 (O_1221,N_14877,N_14940);
or UO_1222 (O_1222,N_14995,N_14934);
or UO_1223 (O_1223,N_14926,N_14949);
nor UO_1224 (O_1224,N_14954,N_14929);
and UO_1225 (O_1225,N_14869,N_14917);
xnor UO_1226 (O_1226,N_14875,N_14901);
and UO_1227 (O_1227,N_14869,N_14952);
or UO_1228 (O_1228,N_14883,N_14858);
and UO_1229 (O_1229,N_14901,N_14930);
nor UO_1230 (O_1230,N_14880,N_14855);
and UO_1231 (O_1231,N_14898,N_14861);
and UO_1232 (O_1232,N_14873,N_14860);
and UO_1233 (O_1233,N_14913,N_14931);
or UO_1234 (O_1234,N_14863,N_14986);
or UO_1235 (O_1235,N_14897,N_14886);
nor UO_1236 (O_1236,N_14857,N_14869);
and UO_1237 (O_1237,N_14964,N_14935);
nor UO_1238 (O_1238,N_14978,N_14852);
nand UO_1239 (O_1239,N_14864,N_14941);
nor UO_1240 (O_1240,N_14947,N_14974);
nand UO_1241 (O_1241,N_14856,N_14863);
and UO_1242 (O_1242,N_14969,N_14881);
and UO_1243 (O_1243,N_14992,N_14892);
xnor UO_1244 (O_1244,N_14895,N_14960);
nor UO_1245 (O_1245,N_14936,N_14914);
nor UO_1246 (O_1246,N_14945,N_14925);
nor UO_1247 (O_1247,N_14986,N_14990);
nand UO_1248 (O_1248,N_14963,N_14927);
or UO_1249 (O_1249,N_14851,N_14888);
nand UO_1250 (O_1250,N_14975,N_14962);
or UO_1251 (O_1251,N_14976,N_14863);
nor UO_1252 (O_1252,N_14856,N_14853);
or UO_1253 (O_1253,N_14891,N_14871);
nor UO_1254 (O_1254,N_14860,N_14936);
nor UO_1255 (O_1255,N_14907,N_14906);
or UO_1256 (O_1256,N_14863,N_14881);
xnor UO_1257 (O_1257,N_14864,N_14952);
nand UO_1258 (O_1258,N_14884,N_14996);
nand UO_1259 (O_1259,N_14967,N_14880);
nor UO_1260 (O_1260,N_14953,N_14855);
nor UO_1261 (O_1261,N_14876,N_14940);
xnor UO_1262 (O_1262,N_14967,N_14921);
or UO_1263 (O_1263,N_14877,N_14984);
and UO_1264 (O_1264,N_14938,N_14972);
or UO_1265 (O_1265,N_14959,N_14929);
or UO_1266 (O_1266,N_14978,N_14933);
nor UO_1267 (O_1267,N_14914,N_14939);
and UO_1268 (O_1268,N_14974,N_14851);
or UO_1269 (O_1269,N_14870,N_14917);
xnor UO_1270 (O_1270,N_14897,N_14901);
and UO_1271 (O_1271,N_14988,N_14927);
or UO_1272 (O_1272,N_14868,N_14867);
nor UO_1273 (O_1273,N_14986,N_14886);
nor UO_1274 (O_1274,N_14925,N_14927);
xor UO_1275 (O_1275,N_14959,N_14859);
xor UO_1276 (O_1276,N_14954,N_14958);
nand UO_1277 (O_1277,N_14870,N_14957);
xnor UO_1278 (O_1278,N_14891,N_14998);
nand UO_1279 (O_1279,N_14975,N_14920);
and UO_1280 (O_1280,N_14854,N_14889);
xnor UO_1281 (O_1281,N_14994,N_14891);
nor UO_1282 (O_1282,N_14971,N_14937);
nor UO_1283 (O_1283,N_14913,N_14993);
nor UO_1284 (O_1284,N_14962,N_14989);
and UO_1285 (O_1285,N_14990,N_14897);
nor UO_1286 (O_1286,N_14905,N_14940);
xnor UO_1287 (O_1287,N_14879,N_14950);
xor UO_1288 (O_1288,N_14913,N_14878);
nand UO_1289 (O_1289,N_14990,N_14883);
and UO_1290 (O_1290,N_14860,N_14863);
nor UO_1291 (O_1291,N_14928,N_14914);
and UO_1292 (O_1292,N_14971,N_14976);
nor UO_1293 (O_1293,N_14953,N_14918);
nor UO_1294 (O_1294,N_14862,N_14928);
and UO_1295 (O_1295,N_14881,N_14941);
or UO_1296 (O_1296,N_14942,N_14917);
or UO_1297 (O_1297,N_14888,N_14919);
or UO_1298 (O_1298,N_14964,N_14920);
and UO_1299 (O_1299,N_14976,N_14905);
nor UO_1300 (O_1300,N_14857,N_14886);
xor UO_1301 (O_1301,N_14999,N_14918);
nand UO_1302 (O_1302,N_14858,N_14944);
xnor UO_1303 (O_1303,N_14918,N_14974);
or UO_1304 (O_1304,N_14956,N_14907);
nor UO_1305 (O_1305,N_14963,N_14907);
and UO_1306 (O_1306,N_14864,N_14912);
nand UO_1307 (O_1307,N_14925,N_14851);
or UO_1308 (O_1308,N_14934,N_14933);
xnor UO_1309 (O_1309,N_14955,N_14975);
nand UO_1310 (O_1310,N_14990,N_14943);
nand UO_1311 (O_1311,N_14927,N_14959);
xnor UO_1312 (O_1312,N_14851,N_14959);
xor UO_1313 (O_1313,N_14858,N_14916);
nand UO_1314 (O_1314,N_14894,N_14868);
nand UO_1315 (O_1315,N_14926,N_14892);
nor UO_1316 (O_1316,N_14977,N_14875);
or UO_1317 (O_1317,N_14999,N_14940);
nor UO_1318 (O_1318,N_14865,N_14928);
nand UO_1319 (O_1319,N_14912,N_14961);
and UO_1320 (O_1320,N_14853,N_14995);
and UO_1321 (O_1321,N_14891,N_14928);
or UO_1322 (O_1322,N_14978,N_14946);
or UO_1323 (O_1323,N_14870,N_14858);
and UO_1324 (O_1324,N_14988,N_14856);
and UO_1325 (O_1325,N_14942,N_14892);
xor UO_1326 (O_1326,N_14948,N_14994);
or UO_1327 (O_1327,N_14924,N_14997);
xnor UO_1328 (O_1328,N_14977,N_14887);
nor UO_1329 (O_1329,N_14891,N_14952);
nor UO_1330 (O_1330,N_14908,N_14892);
and UO_1331 (O_1331,N_14886,N_14884);
and UO_1332 (O_1332,N_14864,N_14900);
or UO_1333 (O_1333,N_14985,N_14908);
nand UO_1334 (O_1334,N_14972,N_14937);
nand UO_1335 (O_1335,N_14971,N_14863);
nand UO_1336 (O_1336,N_14976,N_14894);
nor UO_1337 (O_1337,N_14984,N_14974);
nor UO_1338 (O_1338,N_14952,N_14934);
and UO_1339 (O_1339,N_14904,N_14988);
nand UO_1340 (O_1340,N_14918,N_14858);
nor UO_1341 (O_1341,N_14881,N_14900);
or UO_1342 (O_1342,N_14885,N_14971);
nor UO_1343 (O_1343,N_14976,N_14856);
nand UO_1344 (O_1344,N_14979,N_14995);
and UO_1345 (O_1345,N_14922,N_14982);
or UO_1346 (O_1346,N_14852,N_14938);
nand UO_1347 (O_1347,N_14862,N_14907);
or UO_1348 (O_1348,N_14888,N_14913);
or UO_1349 (O_1349,N_14960,N_14901);
nand UO_1350 (O_1350,N_14870,N_14952);
nand UO_1351 (O_1351,N_14873,N_14875);
xnor UO_1352 (O_1352,N_14857,N_14958);
nand UO_1353 (O_1353,N_14869,N_14899);
or UO_1354 (O_1354,N_14998,N_14902);
and UO_1355 (O_1355,N_14981,N_14929);
xnor UO_1356 (O_1356,N_14921,N_14959);
xnor UO_1357 (O_1357,N_14967,N_14886);
and UO_1358 (O_1358,N_14964,N_14900);
xnor UO_1359 (O_1359,N_14907,N_14896);
or UO_1360 (O_1360,N_14915,N_14914);
nand UO_1361 (O_1361,N_14993,N_14988);
and UO_1362 (O_1362,N_14975,N_14863);
nand UO_1363 (O_1363,N_14856,N_14909);
or UO_1364 (O_1364,N_14950,N_14996);
xnor UO_1365 (O_1365,N_14983,N_14964);
xnor UO_1366 (O_1366,N_14933,N_14903);
xnor UO_1367 (O_1367,N_14922,N_14884);
xor UO_1368 (O_1368,N_14881,N_14971);
or UO_1369 (O_1369,N_14930,N_14922);
and UO_1370 (O_1370,N_14983,N_14941);
nand UO_1371 (O_1371,N_14899,N_14934);
xnor UO_1372 (O_1372,N_14952,N_14948);
xnor UO_1373 (O_1373,N_14920,N_14889);
nand UO_1374 (O_1374,N_14968,N_14974);
nand UO_1375 (O_1375,N_14888,N_14863);
xor UO_1376 (O_1376,N_14960,N_14933);
or UO_1377 (O_1377,N_14995,N_14899);
or UO_1378 (O_1378,N_14855,N_14977);
and UO_1379 (O_1379,N_14936,N_14862);
or UO_1380 (O_1380,N_14921,N_14930);
or UO_1381 (O_1381,N_14954,N_14996);
nor UO_1382 (O_1382,N_14882,N_14906);
and UO_1383 (O_1383,N_14956,N_14856);
and UO_1384 (O_1384,N_14986,N_14869);
nand UO_1385 (O_1385,N_14920,N_14853);
xor UO_1386 (O_1386,N_14947,N_14854);
nor UO_1387 (O_1387,N_14892,N_14961);
nand UO_1388 (O_1388,N_14936,N_14910);
or UO_1389 (O_1389,N_14944,N_14962);
nand UO_1390 (O_1390,N_14967,N_14872);
xor UO_1391 (O_1391,N_14973,N_14960);
xnor UO_1392 (O_1392,N_14994,N_14900);
nand UO_1393 (O_1393,N_14922,N_14942);
nand UO_1394 (O_1394,N_14878,N_14937);
nor UO_1395 (O_1395,N_14880,N_14943);
nor UO_1396 (O_1396,N_14870,N_14857);
nand UO_1397 (O_1397,N_14964,N_14928);
or UO_1398 (O_1398,N_14962,N_14877);
or UO_1399 (O_1399,N_14966,N_14908);
nand UO_1400 (O_1400,N_14852,N_14983);
nor UO_1401 (O_1401,N_14871,N_14922);
nand UO_1402 (O_1402,N_14978,N_14984);
or UO_1403 (O_1403,N_14881,N_14916);
xor UO_1404 (O_1404,N_14954,N_14919);
nor UO_1405 (O_1405,N_14875,N_14951);
nor UO_1406 (O_1406,N_14965,N_14957);
and UO_1407 (O_1407,N_14997,N_14865);
and UO_1408 (O_1408,N_14861,N_14895);
nand UO_1409 (O_1409,N_14931,N_14950);
nor UO_1410 (O_1410,N_14854,N_14899);
nor UO_1411 (O_1411,N_14956,N_14997);
xnor UO_1412 (O_1412,N_14958,N_14876);
or UO_1413 (O_1413,N_14880,N_14914);
or UO_1414 (O_1414,N_14908,N_14945);
or UO_1415 (O_1415,N_14904,N_14947);
nor UO_1416 (O_1416,N_14876,N_14918);
and UO_1417 (O_1417,N_14910,N_14869);
nor UO_1418 (O_1418,N_14936,N_14954);
nor UO_1419 (O_1419,N_14874,N_14977);
xnor UO_1420 (O_1420,N_14941,N_14988);
and UO_1421 (O_1421,N_14890,N_14878);
nor UO_1422 (O_1422,N_14973,N_14939);
and UO_1423 (O_1423,N_14977,N_14881);
xnor UO_1424 (O_1424,N_14871,N_14875);
or UO_1425 (O_1425,N_14933,N_14867);
xor UO_1426 (O_1426,N_14860,N_14896);
and UO_1427 (O_1427,N_14901,N_14882);
nand UO_1428 (O_1428,N_14865,N_14878);
or UO_1429 (O_1429,N_14885,N_14990);
nand UO_1430 (O_1430,N_14931,N_14921);
xnor UO_1431 (O_1431,N_14945,N_14977);
and UO_1432 (O_1432,N_14913,N_14881);
and UO_1433 (O_1433,N_14865,N_14912);
or UO_1434 (O_1434,N_14876,N_14915);
or UO_1435 (O_1435,N_14867,N_14983);
nor UO_1436 (O_1436,N_14922,N_14850);
nor UO_1437 (O_1437,N_14870,N_14962);
nor UO_1438 (O_1438,N_14946,N_14859);
nand UO_1439 (O_1439,N_14985,N_14952);
nand UO_1440 (O_1440,N_14881,N_14952);
and UO_1441 (O_1441,N_14951,N_14864);
xor UO_1442 (O_1442,N_14912,N_14992);
nor UO_1443 (O_1443,N_14885,N_14902);
nand UO_1444 (O_1444,N_14988,N_14905);
and UO_1445 (O_1445,N_14879,N_14850);
xnor UO_1446 (O_1446,N_14867,N_14891);
nand UO_1447 (O_1447,N_14997,N_14885);
nor UO_1448 (O_1448,N_14920,N_14938);
xor UO_1449 (O_1449,N_14982,N_14961);
or UO_1450 (O_1450,N_14872,N_14980);
nand UO_1451 (O_1451,N_14961,N_14873);
xnor UO_1452 (O_1452,N_14884,N_14966);
nand UO_1453 (O_1453,N_14875,N_14850);
and UO_1454 (O_1454,N_14961,N_14986);
and UO_1455 (O_1455,N_14888,N_14960);
or UO_1456 (O_1456,N_14995,N_14868);
or UO_1457 (O_1457,N_14972,N_14944);
nand UO_1458 (O_1458,N_14985,N_14937);
xor UO_1459 (O_1459,N_14910,N_14904);
nor UO_1460 (O_1460,N_14901,N_14891);
xor UO_1461 (O_1461,N_14916,N_14895);
nor UO_1462 (O_1462,N_14898,N_14957);
nor UO_1463 (O_1463,N_14890,N_14913);
xor UO_1464 (O_1464,N_14940,N_14942);
nor UO_1465 (O_1465,N_14925,N_14965);
and UO_1466 (O_1466,N_14956,N_14881);
xor UO_1467 (O_1467,N_14935,N_14913);
nand UO_1468 (O_1468,N_14940,N_14974);
or UO_1469 (O_1469,N_14957,N_14959);
nor UO_1470 (O_1470,N_14875,N_14906);
xor UO_1471 (O_1471,N_14957,N_14999);
nor UO_1472 (O_1472,N_14902,N_14888);
and UO_1473 (O_1473,N_14889,N_14903);
nor UO_1474 (O_1474,N_14923,N_14964);
xor UO_1475 (O_1475,N_14855,N_14979);
and UO_1476 (O_1476,N_14928,N_14940);
nand UO_1477 (O_1477,N_14908,N_14857);
nor UO_1478 (O_1478,N_14907,N_14936);
and UO_1479 (O_1479,N_14920,N_14877);
nor UO_1480 (O_1480,N_14885,N_14863);
nand UO_1481 (O_1481,N_14897,N_14945);
or UO_1482 (O_1482,N_14912,N_14954);
xnor UO_1483 (O_1483,N_14961,N_14932);
nor UO_1484 (O_1484,N_14917,N_14989);
or UO_1485 (O_1485,N_14885,N_14866);
xor UO_1486 (O_1486,N_14869,N_14905);
nor UO_1487 (O_1487,N_14918,N_14861);
and UO_1488 (O_1488,N_14876,N_14965);
nor UO_1489 (O_1489,N_14893,N_14878);
nor UO_1490 (O_1490,N_14896,N_14969);
xnor UO_1491 (O_1491,N_14910,N_14971);
or UO_1492 (O_1492,N_14925,N_14996);
xor UO_1493 (O_1493,N_14922,N_14861);
xnor UO_1494 (O_1494,N_14866,N_14881);
nand UO_1495 (O_1495,N_14992,N_14866);
nand UO_1496 (O_1496,N_14999,N_14911);
nand UO_1497 (O_1497,N_14882,N_14852);
and UO_1498 (O_1498,N_14939,N_14930);
nor UO_1499 (O_1499,N_14894,N_14919);
xnor UO_1500 (O_1500,N_14976,N_14989);
xor UO_1501 (O_1501,N_14852,N_14905);
nor UO_1502 (O_1502,N_14936,N_14861);
nor UO_1503 (O_1503,N_14865,N_14859);
and UO_1504 (O_1504,N_14957,N_14958);
nor UO_1505 (O_1505,N_14883,N_14912);
or UO_1506 (O_1506,N_14850,N_14947);
or UO_1507 (O_1507,N_14881,N_14957);
nor UO_1508 (O_1508,N_14889,N_14935);
and UO_1509 (O_1509,N_14930,N_14900);
nand UO_1510 (O_1510,N_14879,N_14945);
xor UO_1511 (O_1511,N_14974,N_14916);
or UO_1512 (O_1512,N_14940,N_14934);
nor UO_1513 (O_1513,N_14852,N_14856);
and UO_1514 (O_1514,N_14855,N_14903);
nor UO_1515 (O_1515,N_14938,N_14926);
nor UO_1516 (O_1516,N_14876,N_14912);
and UO_1517 (O_1517,N_14946,N_14938);
xnor UO_1518 (O_1518,N_14941,N_14925);
nor UO_1519 (O_1519,N_14865,N_14869);
nand UO_1520 (O_1520,N_14853,N_14943);
and UO_1521 (O_1521,N_14980,N_14976);
and UO_1522 (O_1522,N_14937,N_14922);
nand UO_1523 (O_1523,N_14978,N_14966);
nor UO_1524 (O_1524,N_14860,N_14967);
and UO_1525 (O_1525,N_14990,N_14929);
nor UO_1526 (O_1526,N_14865,N_14925);
xor UO_1527 (O_1527,N_14984,N_14968);
nand UO_1528 (O_1528,N_14864,N_14942);
and UO_1529 (O_1529,N_14962,N_14950);
or UO_1530 (O_1530,N_14884,N_14911);
nor UO_1531 (O_1531,N_14991,N_14988);
and UO_1532 (O_1532,N_14979,N_14889);
and UO_1533 (O_1533,N_14914,N_14938);
and UO_1534 (O_1534,N_14878,N_14915);
and UO_1535 (O_1535,N_14945,N_14957);
nand UO_1536 (O_1536,N_14946,N_14850);
or UO_1537 (O_1537,N_14852,N_14955);
or UO_1538 (O_1538,N_14906,N_14927);
nor UO_1539 (O_1539,N_14912,N_14927);
and UO_1540 (O_1540,N_14908,N_14997);
or UO_1541 (O_1541,N_14906,N_14867);
and UO_1542 (O_1542,N_14966,N_14854);
or UO_1543 (O_1543,N_14939,N_14954);
and UO_1544 (O_1544,N_14866,N_14910);
nand UO_1545 (O_1545,N_14935,N_14948);
nor UO_1546 (O_1546,N_14988,N_14959);
and UO_1547 (O_1547,N_14915,N_14889);
or UO_1548 (O_1548,N_14980,N_14972);
and UO_1549 (O_1549,N_14959,N_14958);
nor UO_1550 (O_1550,N_14932,N_14864);
nor UO_1551 (O_1551,N_14938,N_14909);
xor UO_1552 (O_1552,N_14904,N_14862);
or UO_1553 (O_1553,N_14990,N_14868);
nand UO_1554 (O_1554,N_14883,N_14922);
xor UO_1555 (O_1555,N_14964,N_14950);
and UO_1556 (O_1556,N_14856,N_14971);
xor UO_1557 (O_1557,N_14982,N_14920);
xnor UO_1558 (O_1558,N_14965,N_14877);
nand UO_1559 (O_1559,N_14901,N_14913);
and UO_1560 (O_1560,N_14996,N_14928);
and UO_1561 (O_1561,N_14989,N_14856);
nor UO_1562 (O_1562,N_14983,N_14890);
nand UO_1563 (O_1563,N_14904,N_14985);
nor UO_1564 (O_1564,N_14946,N_14934);
nand UO_1565 (O_1565,N_14891,N_14990);
xor UO_1566 (O_1566,N_14890,N_14995);
nand UO_1567 (O_1567,N_14860,N_14954);
or UO_1568 (O_1568,N_14931,N_14995);
nand UO_1569 (O_1569,N_14904,N_14872);
and UO_1570 (O_1570,N_14906,N_14979);
nand UO_1571 (O_1571,N_14988,N_14908);
xnor UO_1572 (O_1572,N_14992,N_14869);
or UO_1573 (O_1573,N_14969,N_14995);
and UO_1574 (O_1574,N_14990,N_14862);
xor UO_1575 (O_1575,N_14925,N_14970);
nor UO_1576 (O_1576,N_14963,N_14939);
or UO_1577 (O_1577,N_14920,N_14918);
nand UO_1578 (O_1578,N_14890,N_14892);
nor UO_1579 (O_1579,N_14910,N_14955);
xnor UO_1580 (O_1580,N_14975,N_14988);
nor UO_1581 (O_1581,N_14876,N_14871);
nand UO_1582 (O_1582,N_14955,N_14906);
and UO_1583 (O_1583,N_14956,N_14962);
or UO_1584 (O_1584,N_14884,N_14961);
xor UO_1585 (O_1585,N_14941,N_14877);
xor UO_1586 (O_1586,N_14890,N_14996);
nand UO_1587 (O_1587,N_14988,N_14920);
nand UO_1588 (O_1588,N_14998,N_14933);
nor UO_1589 (O_1589,N_14850,N_14892);
or UO_1590 (O_1590,N_14886,N_14977);
xnor UO_1591 (O_1591,N_14933,N_14891);
nor UO_1592 (O_1592,N_14885,N_14896);
xnor UO_1593 (O_1593,N_14907,N_14874);
and UO_1594 (O_1594,N_14931,N_14887);
xor UO_1595 (O_1595,N_14925,N_14931);
or UO_1596 (O_1596,N_14985,N_14931);
and UO_1597 (O_1597,N_14912,N_14963);
and UO_1598 (O_1598,N_14880,N_14904);
nand UO_1599 (O_1599,N_14899,N_14978);
or UO_1600 (O_1600,N_14953,N_14862);
or UO_1601 (O_1601,N_14937,N_14941);
or UO_1602 (O_1602,N_14910,N_14995);
and UO_1603 (O_1603,N_14909,N_14883);
or UO_1604 (O_1604,N_14943,N_14978);
and UO_1605 (O_1605,N_14972,N_14928);
nand UO_1606 (O_1606,N_14873,N_14971);
nand UO_1607 (O_1607,N_14864,N_14909);
nand UO_1608 (O_1608,N_14986,N_14997);
or UO_1609 (O_1609,N_14919,N_14902);
nor UO_1610 (O_1610,N_14930,N_14941);
nand UO_1611 (O_1611,N_14967,N_14909);
or UO_1612 (O_1612,N_14978,N_14873);
xor UO_1613 (O_1613,N_14939,N_14938);
and UO_1614 (O_1614,N_14916,N_14977);
nor UO_1615 (O_1615,N_14948,N_14861);
nor UO_1616 (O_1616,N_14924,N_14933);
xor UO_1617 (O_1617,N_14956,N_14876);
xnor UO_1618 (O_1618,N_14893,N_14883);
nand UO_1619 (O_1619,N_14892,N_14963);
xor UO_1620 (O_1620,N_14899,N_14942);
xor UO_1621 (O_1621,N_14971,N_14943);
and UO_1622 (O_1622,N_14868,N_14884);
nand UO_1623 (O_1623,N_14878,N_14903);
xor UO_1624 (O_1624,N_14926,N_14893);
and UO_1625 (O_1625,N_14895,N_14926);
nor UO_1626 (O_1626,N_14887,N_14922);
and UO_1627 (O_1627,N_14994,N_14912);
or UO_1628 (O_1628,N_14969,N_14930);
or UO_1629 (O_1629,N_14990,N_14982);
xor UO_1630 (O_1630,N_14917,N_14871);
nor UO_1631 (O_1631,N_14861,N_14885);
xnor UO_1632 (O_1632,N_14949,N_14997);
nand UO_1633 (O_1633,N_14896,N_14921);
nor UO_1634 (O_1634,N_14857,N_14928);
nand UO_1635 (O_1635,N_14948,N_14874);
and UO_1636 (O_1636,N_14918,N_14932);
nand UO_1637 (O_1637,N_14913,N_14937);
or UO_1638 (O_1638,N_14988,N_14895);
and UO_1639 (O_1639,N_14985,N_14981);
and UO_1640 (O_1640,N_14855,N_14931);
nor UO_1641 (O_1641,N_14942,N_14916);
and UO_1642 (O_1642,N_14874,N_14937);
xnor UO_1643 (O_1643,N_14908,N_14906);
nand UO_1644 (O_1644,N_14922,N_14880);
nand UO_1645 (O_1645,N_14930,N_14871);
and UO_1646 (O_1646,N_14953,N_14890);
and UO_1647 (O_1647,N_14888,N_14953);
xnor UO_1648 (O_1648,N_14972,N_14976);
nor UO_1649 (O_1649,N_14930,N_14982);
or UO_1650 (O_1650,N_14985,N_14959);
xor UO_1651 (O_1651,N_14889,N_14947);
or UO_1652 (O_1652,N_14854,N_14983);
or UO_1653 (O_1653,N_14899,N_14873);
nand UO_1654 (O_1654,N_14909,N_14898);
xor UO_1655 (O_1655,N_14944,N_14936);
nor UO_1656 (O_1656,N_14877,N_14975);
xnor UO_1657 (O_1657,N_14858,N_14984);
nand UO_1658 (O_1658,N_14853,N_14918);
and UO_1659 (O_1659,N_14915,N_14960);
or UO_1660 (O_1660,N_14960,N_14965);
or UO_1661 (O_1661,N_14874,N_14957);
or UO_1662 (O_1662,N_14971,N_14939);
or UO_1663 (O_1663,N_14873,N_14901);
or UO_1664 (O_1664,N_14900,N_14868);
or UO_1665 (O_1665,N_14873,N_14896);
nand UO_1666 (O_1666,N_14991,N_14957);
xnor UO_1667 (O_1667,N_14943,N_14875);
nand UO_1668 (O_1668,N_14883,N_14921);
and UO_1669 (O_1669,N_14985,N_14879);
xnor UO_1670 (O_1670,N_14920,N_14893);
and UO_1671 (O_1671,N_14917,N_14979);
nand UO_1672 (O_1672,N_14962,N_14994);
nor UO_1673 (O_1673,N_14862,N_14930);
nand UO_1674 (O_1674,N_14939,N_14851);
nor UO_1675 (O_1675,N_14967,N_14883);
xor UO_1676 (O_1676,N_14954,N_14917);
nor UO_1677 (O_1677,N_14878,N_14968);
and UO_1678 (O_1678,N_14898,N_14965);
and UO_1679 (O_1679,N_14950,N_14856);
xor UO_1680 (O_1680,N_14998,N_14959);
xor UO_1681 (O_1681,N_14903,N_14866);
xnor UO_1682 (O_1682,N_14945,N_14882);
nand UO_1683 (O_1683,N_14867,N_14866);
or UO_1684 (O_1684,N_14855,N_14899);
and UO_1685 (O_1685,N_14916,N_14944);
nand UO_1686 (O_1686,N_14882,N_14877);
nor UO_1687 (O_1687,N_14943,N_14983);
xor UO_1688 (O_1688,N_14895,N_14990);
xnor UO_1689 (O_1689,N_14890,N_14989);
and UO_1690 (O_1690,N_14975,N_14966);
nor UO_1691 (O_1691,N_14994,N_14881);
nor UO_1692 (O_1692,N_14996,N_14987);
nand UO_1693 (O_1693,N_14881,N_14855);
nand UO_1694 (O_1694,N_14988,N_14867);
or UO_1695 (O_1695,N_14926,N_14983);
nor UO_1696 (O_1696,N_14860,N_14973);
or UO_1697 (O_1697,N_14999,N_14851);
nand UO_1698 (O_1698,N_14953,N_14990);
xnor UO_1699 (O_1699,N_14938,N_14962);
nand UO_1700 (O_1700,N_14977,N_14981);
xnor UO_1701 (O_1701,N_14857,N_14877);
and UO_1702 (O_1702,N_14917,N_14948);
xor UO_1703 (O_1703,N_14981,N_14960);
and UO_1704 (O_1704,N_14858,N_14960);
or UO_1705 (O_1705,N_14969,N_14866);
and UO_1706 (O_1706,N_14868,N_14895);
nor UO_1707 (O_1707,N_14970,N_14862);
xnor UO_1708 (O_1708,N_14990,N_14875);
nand UO_1709 (O_1709,N_14952,N_14867);
nor UO_1710 (O_1710,N_14906,N_14899);
xor UO_1711 (O_1711,N_14869,N_14902);
nand UO_1712 (O_1712,N_14911,N_14894);
nor UO_1713 (O_1713,N_14853,N_14931);
nand UO_1714 (O_1714,N_14876,N_14854);
nor UO_1715 (O_1715,N_14968,N_14892);
nand UO_1716 (O_1716,N_14926,N_14998);
xnor UO_1717 (O_1717,N_14988,N_14901);
nand UO_1718 (O_1718,N_14984,N_14997);
or UO_1719 (O_1719,N_14910,N_14924);
xnor UO_1720 (O_1720,N_14872,N_14994);
and UO_1721 (O_1721,N_14866,N_14987);
xnor UO_1722 (O_1722,N_14931,N_14883);
or UO_1723 (O_1723,N_14926,N_14886);
xor UO_1724 (O_1724,N_14972,N_14930);
and UO_1725 (O_1725,N_14890,N_14861);
xnor UO_1726 (O_1726,N_14996,N_14926);
or UO_1727 (O_1727,N_14924,N_14930);
nand UO_1728 (O_1728,N_14945,N_14988);
or UO_1729 (O_1729,N_14939,N_14862);
xor UO_1730 (O_1730,N_14941,N_14915);
xnor UO_1731 (O_1731,N_14907,N_14917);
nand UO_1732 (O_1732,N_14859,N_14903);
or UO_1733 (O_1733,N_14887,N_14856);
nand UO_1734 (O_1734,N_14882,N_14889);
and UO_1735 (O_1735,N_14998,N_14979);
or UO_1736 (O_1736,N_14998,N_14855);
and UO_1737 (O_1737,N_14921,N_14876);
nand UO_1738 (O_1738,N_14883,N_14992);
nor UO_1739 (O_1739,N_14997,N_14866);
and UO_1740 (O_1740,N_14859,N_14991);
and UO_1741 (O_1741,N_14996,N_14984);
xor UO_1742 (O_1742,N_14995,N_14939);
xor UO_1743 (O_1743,N_14944,N_14908);
or UO_1744 (O_1744,N_14930,N_14968);
xnor UO_1745 (O_1745,N_14899,N_14884);
nor UO_1746 (O_1746,N_14966,N_14876);
xnor UO_1747 (O_1747,N_14962,N_14968);
nand UO_1748 (O_1748,N_14909,N_14863);
nand UO_1749 (O_1749,N_14992,N_14979);
xnor UO_1750 (O_1750,N_14946,N_14878);
xnor UO_1751 (O_1751,N_14893,N_14881);
and UO_1752 (O_1752,N_14919,N_14906);
xnor UO_1753 (O_1753,N_14896,N_14966);
nor UO_1754 (O_1754,N_14912,N_14868);
nand UO_1755 (O_1755,N_14981,N_14973);
or UO_1756 (O_1756,N_14969,N_14890);
xnor UO_1757 (O_1757,N_14984,N_14967);
or UO_1758 (O_1758,N_14906,N_14863);
xor UO_1759 (O_1759,N_14858,N_14854);
or UO_1760 (O_1760,N_14908,N_14979);
nor UO_1761 (O_1761,N_14967,N_14992);
or UO_1762 (O_1762,N_14900,N_14973);
xor UO_1763 (O_1763,N_14975,N_14929);
nor UO_1764 (O_1764,N_14869,N_14873);
or UO_1765 (O_1765,N_14899,N_14992);
and UO_1766 (O_1766,N_14964,N_14993);
and UO_1767 (O_1767,N_14882,N_14925);
or UO_1768 (O_1768,N_14884,N_14969);
or UO_1769 (O_1769,N_14943,N_14897);
nor UO_1770 (O_1770,N_14962,N_14914);
or UO_1771 (O_1771,N_14916,N_14964);
nor UO_1772 (O_1772,N_14900,N_14959);
and UO_1773 (O_1773,N_14932,N_14905);
and UO_1774 (O_1774,N_14969,N_14975);
or UO_1775 (O_1775,N_14950,N_14983);
nor UO_1776 (O_1776,N_14937,N_14923);
nor UO_1777 (O_1777,N_14907,N_14923);
and UO_1778 (O_1778,N_14946,N_14871);
nor UO_1779 (O_1779,N_14993,N_14944);
nand UO_1780 (O_1780,N_14880,N_14974);
nand UO_1781 (O_1781,N_14870,N_14993);
xnor UO_1782 (O_1782,N_14851,N_14951);
xnor UO_1783 (O_1783,N_14905,N_14903);
and UO_1784 (O_1784,N_14929,N_14989);
xnor UO_1785 (O_1785,N_14956,N_14955);
nor UO_1786 (O_1786,N_14913,N_14984);
nor UO_1787 (O_1787,N_14937,N_14964);
nor UO_1788 (O_1788,N_14966,N_14885);
or UO_1789 (O_1789,N_14933,N_14963);
nor UO_1790 (O_1790,N_14946,N_14852);
nand UO_1791 (O_1791,N_14876,N_14860);
xnor UO_1792 (O_1792,N_14983,N_14999);
and UO_1793 (O_1793,N_14974,N_14954);
nand UO_1794 (O_1794,N_14950,N_14939);
xnor UO_1795 (O_1795,N_14862,N_14900);
nor UO_1796 (O_1796,N_14974,N_14887);
xnor UO_1797 (O_1797,N_14939,N_14941);
and UO_1798 (O_1798,N_14878,N_14992);
nand UO_1799 (O_1799,N_14907,N_14920);
and UO_1800 (O_1800,N_14876,N_14952);
or UO_1801 (O_1801,N_14912,N_14939);
nand UO_1802 (O_1802,N_14859,N_14984);
and UO_1803 (O_1803,N_14965,N_14870);
nor UO_1804 (O_1804,N_14922,N_14999);
and UO_1805 (O_1805,N_14916,N_14913);
nand UO_1806 (O_1806,N_14854,N_14920);
nand UO_1807 (O_1807,N_14875,N_14877);
nand UO_1808 (O_1808,N_14995,N_14981);
xor UO_1809 (O_1809,N_14890,N_14935);
nand UO_1810 (O_1810,N_14983,N_14962);
and UO_1811 (O_1811,N_14867,N_14902);
nor UO_1812 (O_1812,N_14860,N_14916);
xnor UO_1813 (O_1813,N_14975,N_14911);
and UO_1814 (O_1814,N_14966,N_14901);
xnor UO_1815 (O_1815,N_14921,N_14944);
or UO_1816 (O_1816,N_14911,N_14944);
or UO_1817 (O_1817,N_14926,N_14873);
nand UO_1818 (O_1818,N_14893,N_14866);
nand UO_1819 (O_1819,N_14900,N_14929);
nand UO_1820 (O_1820,N_14934,N_14916);
nor UO_1821 (O_1821,N_14893,N_14884);
and UO_1822 (O_1822,N_14922,N_14958);
nand UO_1823 (O_1823,N_14974,N_14917);
nor UO_1824 (O_1824,N_14993,N_14965);
xor UO_1825 (O_1825,N_14964,N_14881);
nand UO_1826 (O_1826,N_14932,N_14990);
xnor UO_1827 (O_1827,N_14963,N_14999);
and UO_1828 (O_1828,N_14871,N_14950);
xor UO_1829 (O_1829,N_14902,N_14874);
or UO_1830 (O_1830,N_14899,N_14924);
nand UO_1831 (O_1831,N_14959,N_14952);
and UO_1832 (O_1832,N_14931,N_14955);
and UO_1833 (O_1833,N_14899,N_14949);
nor UO_1834 (O_1834,N_14914,N_14950);
nor UO_1835 (O_1835,N_14936,N_14966);
xor UO_1836 (O_1836,N_14964,N_14957);
or UO_1837 (O_1837,N_14877,N_14863);
nand UO_1838 (O_1838,N_14860,N_14889);
or UO_1839 (O_1839,N_14992,N_14972);
xor UO_1840 (O_1840,N_14892,N_14880);
or UO_1841 (O_1841,N_14934,N_14886);
and UO_1842 (O_1842,N_14944,N_14978);
nor UO_1843 (O_1843,N_14977,N_14988);
nand UO_1844 (O_1844,N_14857,N_14889);
nand UO_1845 (O_1845,N_14879,N_14981);
or UO_1846 (O_1846,N_14875,N_14914);
nand UO_1847 (O_1847,N_14893,N_14879);
or UO_1848 (O_1848,N_14982,N_14895);
and UO_1849 (O_1849,N_14968,N_14851);
or UO_1850 (O_1850,N_14864,N_14916);
and UO_1851 (O_1851,N_14883,N_14879);
nor UO_1852 (O_1852,N_14938,N_14998);
and UO_1853 (O_1853,N_14869,N_14945);
nor UO_1854 (O_1854,N_14885,N_14937);
and UO_1855 (O_1855,N_14904,N_14879);
nor UO_1856 (O_1856,N_14954,N_14873);
or UO_1857 (O_1857,N_14873,N_14929);
or UO_1858 (O_1858,N_14850,N_14925);
or UO_1859 (O_1859,N_14921,N_14980);
nor UO_1860 (O_1860,N_14889,N_14954);
nand UO_1861 (O_1861,N_14890,N_14911);
and UO_1862 (O_1862,N_14885,N_14911);
nand UO_1863 (O_1863,N_14853,N_14982);
nand UO_1864 (O_1864,N_14909,N_14941);
and UO_1865 (O_1865,N_14959,N_14948);
or UO_1866 (O_1866,N_14917,N_14886);
nand UO_1867 (O_1867,N_14895,N_14914);
or UO_1868 (O_1868,N_14904,N_14945);
and UO_1869 (O_1869,N_14884,N_14914);
xor UO_1870 (O_1870,N_14861,N_14917);
nor UO_1871 (O_1871,N_14975,N_14953);
or UO_1872 (O_1872,N_14928,N_14974);
and UO_1873 (O_1873,N_14964,N_14959);
and UO_1874 (O_1874,N_14969,N_14953);
xnor UO_1875 (O_1875,N_14982,N_14995);
or UO_1876 (O_1876,N_14937,N_14911);
xor UO_1877 (O_1877,N_14922,N_14932);
xor UO_1878 (O_1878,N_14892,N_14886);
xnor UO_1879 (O_1879,N_14906,N_14948);
nand UO_1880 (O_1880,N_14960,N_14920);
xnor UO_1881 (O_1881,N_14967,N_14987);
or UO_1882 (O_1882,N_14932,N_14970);
xor UO_1883 (O_1883,N_14995,N_14855);
and UO_1884 (O_1884,N_14941,N_14872);
and UO_1885 (O_1885,N_14947,N_14881);
and UO_1886 (O_1886,N_14958,N_14991);
nand UO_1887 (O_1887,N_14901,N_14954);
or UO_1888 (O_1888,N_14944,N_14886);
and UO_1889 (O_1889,N_14861,N_14897);
nand UO_1890 (O_1890,N_14962,N_14891);
nor UO_1891 (O_1891,N_14933,N_14851);
nor UO_1892 (O_1892,N_14904,N_14866);
or UO_1893 (O_1893,N_14973,N_14877);
or UO_1894 (O_1894,N_14979,N_14905);
nand UO_1895 (O_1895,N_14934,N_14914);
or UO_1896 (O_1896,N_14943,N_14969);
nand UO_1897 (O_1897,N_14889,N_14939);
nor UO_1898 (O_1898,N_14866,N_14983);
xnor UO_1899 (O_1899,N_14929,N_14881);
and UO_1900 (O_1900,N_14878,N_14884);
xor UO_1901 (O_1901,N_14979,N_14859);
xor UO_1902 (O_1902,N_14967,N_14993);
nor UO_1903 (O_1903,N_14988,N_14923);
or UO_1904 (O_1904,N_14861,N_14990);
nand UO_1905 (O_1905,N_14940,N_14977);
or UO_1906 (O_1906,N_14891,N_14879);
and UO_1907 (O_1907,N_14916,N_14868);
nand UO_1908 (O_1908,N_14993,N_14860);
nor UO_1909 (O_1909,N_14964,N_14890);
nor UO_1910 (O_1910,N_14987,N_14952);
or UO_1911 (O_1911,N_14980,N_14892);
nand UO_1912 (O_1912,N_14887,N_14873);
nor UO_1913 (O_1913,N_14851,N_14985);
and UO_1914 (O_1914,N_14918,N_14921);
nor UO_1915 (O_1915,N_14894,N_14993);
and UO_1916 (O_1916,N_14952,N_14922);
xor UO_1917 (O_1917,N_14855,N_14974);
nand UO_1918 (O_1918,N_14879,N_14940);
xor UO_1919 (O_1919,N_14930,N_14851);
and UO_1920 (O_1920,N_14991,N_14919);
xnor UO_1921 (O_1921,N_14965,N_14996);
nor UO_1922 (O_1922,N_14863,N_14942);
nand UO_1923 (O_1923,N_14894,N_14921);
and UO_1924 (O_1924,N_14975,N_14859);
and UO_1925 (O_1925,N_14990,N_14997);
nand UO_1926 (O_1926,N_14963,N_14890);
nor UO_1927 (O_1927,N_14997,N_14860);
nor UO_1928 (O_1928,N_14943,N_14949);
nand UO_1929 (O_1929,N_14896,N_14895);
and UO_1930 (O_1930,N_14914,N_14991);
or UO_1931 (O_1931,N_14981,N_14871);
and UO_1932 (O_1932,N_14932,N_14930);
and UO_1933 (O_1933,N_14980,N_14852);
nor UO_1934 (O_1934,N_14948,N_14890);
and UO_1935 (O_1935,N_14921,N_14889);
or UO_1936 (O_1936,N_14922,N_14882);
or UO_1937 (O_1937,N_14968,N_14982);
and UO_1938 (O_1938,N_14882,N_14999);
and UO_1939 (O_1939,N_14897,N_14882);
or UO_1940 (O_1940,N_14947,N_14994);
nor UO_1941 (O_1941,N_14914,N_14853);
nor UO_1942 (O_1942,N_14885,N_14994);
or UO_1943 (O_1943,N_14855,N_14965);
and UO_1944 (O_1944,N_14900,N_14982);
nor UO_1945 (O_1945,N_14925,N_14923);
xnor UO_1946 (O_1946,N_14991,N_14923);
and UO_1947 (O_1947,N_14896,N_14926);
xor UO_1948 (O_1948,N_14910,N_14918);
or UO_1949 (O_1949,N_14925,N_14930);
nand UO_1950 (O_1950,N_14959,N_14989);
nor UO_1951 (O_1951,N_14900,N_14975);
xnor UO_1952 (O_1952,N_14856,N_14967);
nand UO_1953 (O_1953,N_14949,N_14855);
or UO_1954 (O_1954,N_14922,N_14943);
and UO_1955 (O_1955,N_14915,N_14912);
and UO_1956 (O_1956,N_14886,N_14925);
and UO_1957 (O_1957,N_14933,N_14874);
or UO_1958 (O_1958,N_14922,N_14889);
or UO_1959 (O_1959,N_14931,N_14935);
nand UO_1960 (O_1960,N_14869,N_14951);
nor UO_1961 (O_1961,N_14926,N_14905);
nor UO_1962 (O_1962,N_14903,N_14909);
nand UO_1963 (O_1963,N_14962,N_14959);
xnor UO_1964 (O_1964,N_14880,N_14952);
nor UO_1965 (O_1965,N_14913,N_14892);
xor UO_1966 (O_1966,N_14951,N_14959);
xor UO_1967 (O_1967,N_14992,N_14942);
and UO_1968 (O_1968,N_14864,N_14855);
or UO_1969 (O_1969,N_14887,N_14859);
or UO_1970 (O_1970,N_14999,N_14937);
xor UO_1971 (O_1971,N_14934,N_14989);
and UO_1972 (O_1972,N_14942,N_14964);
or UO_1973 (O_1973,N_14905,N_14930);
and UO_1974 (O_1974,N_14980,N_14866);
and UO_1975 (O_1975,N_14983,N_14868);
xor UO_1976 (O_1976,N_14877,N_14981);
and UO_1977 (O_1977,N_14916,N_14995);
or UO_1978 (O_1978,N_14877,N_14927);
or UO_1979 (O_1979,N_14873,N_14910);
or UO_1980 (O_1980,N_14999,N_14945);
nand UO_1981 (O_1981,N_14923,N_14945);
or UO_1982 (O_1982,N_14997,N_14882);
or UO_1983 (O_1983,N_14988,N_14955);
nor UO_1984 (O_1984,N_14852,N_14878);
xnor UO_1985 (O_1985,N_14852,N_14880);
or UO_1986 (O_1986,N_14930,N_14973);
and UO_1987 (O_1987,N_14938,N_14931);
and UO_1988 (O_1988,N_14926,N_14925);
nor UO_1989 (O_1989,N_14931,N_14930);
nor UO_1990 (O_1990,N_14988,N_14937);
and UO_1991 (O_1991,N_14894,N_14957);
nor UO_1992 (O_1992,N_14917,N_14950);
or UO_1993 (O_1993,N_14890,N_14859);
xnor UO_1994 (O_1994,N_14967,N_14873);
and UO_1995 (O_1995,N_14902,N_14937);
nand UO_1996 (O_1996,N_14889,N_14944);
and UO_1997 (O_1997,N_14883,N_14908);
nor UO_1998 (O_1998,N_14855,N_14945);
nor UO_1999 (O_1999,N_14952,N_14961);
endmodule