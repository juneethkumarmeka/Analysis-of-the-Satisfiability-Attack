module basic_3000_30000_3500_150_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1868,In_2615);
nor U1 (N_1,In_1370,In_1482);
xnor U2 (N_2,In_1806,In_86);
nand U3 (N_3,In_1171,In_527);
nand U4 (N_4,In_2827,In_1466);
nand U5 (N_5,In_1195,In_43);
or U6 (N_6,In_1376,In_1265);
or U7 (N_7,In_1676,In_97);
nand U8 (N_8,In_210,In_631);
nand U9 (N_9,In_1323,In_1608);
or U10 (N_10,In_1349,In_2217);
xnor U11 (N_11,In_758,In_1991);
xor U12 (N_12,In_1659,In_1109);
xor U13 (N_13,In_622,In_1428);
nand U14 (N_14,In_1933,In_2856);
xnor U15 (N_15,In_2697,In_789);
or U16 (N_16,In_921,In_2720);
xnor U17 (N_17,In_2554,In_768);
or U18 (N_18,In_505,In_1776);
nor U19 (N_19,In_1277,In_18);
or U20 (N_20,In_1408,In_2786);
nor U21 (N_21,In_1320,In_1845);
nor U22 (N_22,In_56,In_590);
nor U23 (N_23,In_909,In_540);
xor U24 (N_24,In_1753,In_246);
and U25 (N_25,In_2934,In_962);
nand U26 (N_26,In_1346,In_305);
nor U27 (N_27,In_2654,In_16);
nand U28 (N_28,In_1434,In_1145);
or U29 (N_29,In_1141,In_1152);
and U30 (N_30,In_355,In_2830);
xnor U31 (N_31,In_1936,In_990);
and U32 (N_32,In_1289,In_876);
or U33 (N_33,In_1382,In_2987);
nor U34 (N_34,In_2738,In_1138);
and U35 (N_35,In_2941,In_933);
nor U36 (N_36,In_2629,In_1628);
xor U37 (N_37,In_35,In_2557);
xnor U38 (N_38,In_2811,In_1083);
xnor U39 (N_39,In_2081,In_2463);
nand U40 (N_40,In_2219,In_2608);
xor U41 (N_41,In_277,In_1554);
xnor U42 (N_42,In_2973,In_1588);
and U43 (N_43,In_2621,In_166);
nor U44 (N_44,In_154,In_754);
and U45 (N_45,In_717,In_2240);
or U46 (N_46,In_176,In_1662);
xnor U47 (N_47,In_2848,In_2622);
xor U48 (N_48,In_2341,In_2668);
xor U49 (N_49,In_552,In_1122);
nand U50 (N_50,In_2017,In_808);
or U51 (N_51,In_2316,In_1194);
xnor U52 (N_52,In_1941,In_1945);
or U53 (N_53,In_2584,In_157);
and U54 (N_54,In_1810,In_1736);
and U55 (N_55,In_2072,In_766);
nor U56 (N_56,In_844,In_2914);
xor U57 (N_57,In_1520,In_1779);
xnor U58 (N_58,In_244,In_1594);
nor U59 (N_59,In_2768,In_680);
and U60 (N_60,In_498,In_2018);
xor U61 (N_61,In_2395,In_1484);
and U62 (N_62,In_987,In_1538);
or U63 (N_63,In_2809,In_2465);
nand U64 (N_64,In_1982,In_175);
and U65 (N_65,In_288,In_256);
and U66 (N_66,In_2873,In_2489);
nor U67 (N_67,In_1282,In_2055);
nand U68 (N_68,In_1177,In_2574);
or U69 (N_69,In_1273,In_2047);
nor U70 (N_70,In_2184,In_551);
and U71 (N_71,In_2705,In_376);
nand U72 (N_72,In_1759,In_863);
xor U73 (N_73,In_2690,In_2958);
or U74 (N_74,In_2276,In_1723);
nand U75 (N_75,In_636,In_129);
xor U76 (N_76,In_1768,In_76);
or U77 (N_77,In_1727,In_1703);
nor U78 (N_78,In_1773,In_1497);
or U79 (N_79,In_1340,In_270);
and U80 (N_80,In_2991,In_1997);
and U81 (N_81,In_2211,In_1039);
nand U82 (N_82,In_2863,In_1355);
nand U83 (N_83,In_2933,In_1262);
xnor U84 (N_84,In_2294,In_373);
nand U85 (N_85,In_1331,In_2226);
and U86 (N_86,In_2338,In_1133);
xnor U87 (N_87,In_661,In_2053);
xnor U88 (N_88,In_2050,In_1948);
xnor U89 (N_89,In_2486,In_753);
xor U90 (N_90,In_1386,In_115);
nor U91 (N_91,In_49,In_2521);
xor U92 (N_92,In_1964,In_140);
nor U93 (N_93,In_2661,In_2459);
or U94 (N_94,In_452,In_2603);
nor U95 (N_95,In_426,In_1867);
or U96 (N_96,In_2350,In_476);
or U97 (N_97,In_2004,In_19);
and U98 (N_98,In_936,In_707);
and U99 (N_99,In_940,In_2028);
nand U100 (N_100,In_2441,In_785);
or U101 (N_101,In_870,In_821);
xor U102 (N_102,In_671,In_2069);
nand U103 (N_103,In_1001,In_1284);
xnor U104 (N_104,In_1011,In_1319);
or U105 (N_105,In_2602,In_388);
nand U106 (N_106,In_2852,In_2037);
nand U107 (N_107,In_61,In_2426);
xnor U108 (N_108,In_994,In_1257);
and U109 (N_109,In_1527,In_1616);
and U110 (N_110,In_1837,In_2742);
nor U111 (N_111,In_2439,In_2974);
xor U112 (N_112,In_461,In_2052);
xnor U113 (N_113,In_51,In_1657);
and U114 (N_114,In_2836,In_1111);
and U115 (N_115,In_1942,In_73);
nand U116 (N_116,In_1770,In_682);
or U117 (N_117,In_2168,In_958);
nand U118 (N_118,In_1215,In_1454);
xor U119 (N_119,In_1605,In_2216);
or U120 (N_120,In_2516,In_513);
or U121 (N_121,In_189,In_2701);
or U122 (N_122,In_2887,In_1623);
and U123 (N_123,In_2386,In_2548);
xor U124 (N_124,In_1557,In_646);
and U125 (N_125,In_1275,In_1621);
xnor U126 (N_126,In_1696,In_137);
nand U127 (N_127,In_917,In_2212);
nand U128 (N_128,In_2903,In_2594);
and U129 (N_129,In_1387,In_1949);
nand U130 (N_130,In_2106,In_687);
xnor U131 (N_131,In_1153,In_2203);
nand U132 (N_132,In_727,In_1430);
and U133 (N_133,In_964,In_2562);
or U134 (N_134,In_2745,In_2101);
nor U135 (N_135,In_1227,In_1451);
nand U136 (N_136,In_460,In_1615);
nand U137 (N_137,In_110,In_977);
xnor U138 (N_138,In_2062,In_2385);
xnor U139 (N_139,In_33,In_2267);
or U140 (N_140,In_975,In_2096);
or U141 (N_141,In_1298,In_1857);
nor U142 (N_142,In_1782,In_2715);
or U143 (N_143,In_2538,In_403);
nand U144 (N_144,In_2826,In_1611);
nand U145 (N_145,In_2948,In_94);
or U146 (N_146,In_664,In_2209);
and U147 (N_147,In_1007,In_2039);
nor U148 (N_148,In_493,In_1720);
xnor U149 (N_149,In_1128,In_2077);
and U150 (N_150,In_2404,In_1180);
and U151 (N_151,In_1673,In_2483);
and U152 (N_152,In_834,In_2503);
xnor U153 (N_153,In_1899,In_932);
and U154 (N_154,In_2589,In_599);
and U155 (N_155,In_1020,In_30);
and U156 (N_156,In_1286,In_143);
nor U157 (N_157,In_1730,In_1105);
and U158 (N_158,In_1000,In_740);
or U159 (N_159,In_1804,In_445);
nand U160 (N_160,In_1062,In_516);
xnor U161 (N_161,In_2894,In_1901);
nor U162 (N_162,In_2539,In_421);
and U163 (N_163,In_2814,In_2921);
nand U164 (N_164,In_1552,In_2191);
xnor U165 (N_165,In_1792,In_2130);
nand U166 (N_166,In_1025,In_2712);
nor U167 (N_167,In_2900,In_912);
xor U168 (N_168,In_603,In_2136);
xnor U169 (N_169,In_262,In_914);
xnor U170 (N_170,In_1926,In_2396);
nand U171 (N_171,In_2936,In_2422);
xnor U172 (N_172,In_356,In_385);
xnor U173 (N_173,In_692,In_69);
and U174 (N_174,In_1296,In_533);
nor U175 (N_175,In_1073,In_2955);
nor U176 (N_176,In_2617,In_2803);
or U177 (N_177,In_616,In_894);
xor U178 (N_178,In_2799,In_827);
xor U179 (N_179,In_1276,In_2074);
nor U180 (N_180,In_1668,In_5);
xor U181 (N_181,In_2778,In_2949);
or U182 (N_182,In_2840,In_547);
and U183 (N_183,In_79,In_2808);
nand U184 (N_184,In_1456,In_2205);
or U185 (N_185,In_406,In_1854);
nor U186 (N_186,In_2869,In_1710);
nand U187 (N_187,In_1504,In_2499);
nand U188 (N_188,In_325,In_575);
nand U189 (N_189,In_2733,In_1999);
xor U190 (N_190,In_359,In_744);
nor U191 (N_191,In_1783,In_119);
and U192 (N_192,In_2369,In_399);
xnor U193 (N_193,In_1789,In_2336);
or U194 (N_194,In_2012,In_594);
nor U195 (N_195,In_1494,In_1738);
nand U196 (N_196,In_128,In_2227);
nand U197 (N_197,In_1674,In_2692);
nor U198 (N_198,In_1785,In_1190);
or U199 (N_199,In_435,In_2542);
xnor U200 (N_200,In_2549,In_454);
nor U201 (N_201,In_2902,In_479);
nor U202 (N_202,In_459,In_453);
and U203 (N_203,In_1835,In_2561);
or U204 (N_204,In_2149,In_2569);
nor U205 (N_205,In_2084,In_923);
nor U206 (N_206,In_44,In_647);
nand U207 (N_207,In_586,In_2695);
or U208 (N_208,In_1102,In_730);
or U209 (N_209,In_1803,In_1700);
or U210 (N_210,In_2148,In_167);
xor U211 (N_211,In_2639,In_2671);
and U212 (N_212,In_2880,In_2323);
nor U213 (N_213,In_1909,In_474);
nand U214 (N_214,In_1050,In_2765);
xor U215 (N_215,In_2927,In_22);
or U216 (N_216,In_2597,In_2930);
nor U217 (N_217,N_196,In_1415);
and U218 (N_218,In_2837,In_793);
or U219 (N_219,In_2423,In_2382);
and U220 (N_220,In_1536,In_855);
and U221 (N_221,In_2364,In_1071);
or U222 (N_222,In_978,In_2245);
and U223 (N_223,In_2107,In_2753);
or U224 (N_224,In_850,In_1158);
nor U225 (N_225,In_1653,N_51);
nor U226 (N_226,In_12,In_1938);
and U227 (N_227,In_1404,In_980);
xor U228 (N_228,In_2740,In_322);
and U229 (N_229,In_87,In_285);
xnor U230 (N_230,In_641,In_1980);
or U231 (N_231,In_319,In_218);
nand U232 (N_232,In_2056,In_2694);
nand U233 (N_233,In_637,In_786);
nor U234 (N_234,In_1435,In_265);
and U235 (N_235,N_88,In_787);
or U236 (N_236,In_190,In_743);
nand U237 (N_237,In_2756,In_2270);
xnor U238 (N_238,In_718,In_1241);
xnor U239 (N_239,In_2755,In_1017);
xor U240 (N_240,In_1612,In_1357);
and U241 (N_241,In_1869,In_338);
nand U242 (N_242,N_181,In_2221);
or U243 (N_243,In_236,In_612);
or U244 (N_244,In_694,In_122);
or U245 (N_245,In_396,In_1755);
xnor U246 (N_246,In_2181,In_1216);
nand U247 (N_247,In_2759,In_1206);
and U248 (N_248,In_1729,In_693);
nor U249 (N_249,In_497,In_2078);
or U250 (N_250,In_2114,In_2648);
and U251 (N_251,In_556,N_100);
or U252 (N_252,In_469,In_2126);
or U253 (N_253,In_503,In_2131);
nand U254 (N_254,In_1266,In_2901);
or U255 (N_255,In_2075,In_2073);
nor U256 (N_256,In_1255,N_115);
nand U257 (N_257,In_2978,In_324);
xnor U258 (N_258,In_833,In_679);
and U259 (N_259,N_117,In_2804);
and U260 (N_260,N_133,In_2817);
nand U261 (N_261,In_2616,In_2770);
or U262 (N_262,In_114,N_50);
and U263 (N_263,In_529,In_838);
or U264 (N_264,In_941,In_643);
xnor U265 (N_265,In_111,In_2523);
nor U266 (N_266,In_1704,In_872);
nor U267 (N_267,In_1272,In_2407);
nor U268 (N_268,In_1389,In_1246);
nor U269 (N_269,In_2854,In_1896);
nand U270 (N_270,In_1392,In_1101);
xor U271 (N_271,In_1442,N_3);
nor U272 (N_272,In_1147,In_14);
or U273 (N_273,In_1965,In_106);
xor U274 (N_274,In_1048,In_1607);
or U275 (N_275,In_2912,In_1908);
nor U276 (N_276,In_714,In_1418);
xnor U277 (N_277,In_2058,In_197);
or U278 (N_278,In_2059,In_1400);
or U279 (N_279,In_2448,In_1577);
xnor U280 (N_280,In_653,In_2286);
nand U281 (N_281,In_1781,In_1469);
or U282 (N_282,In_2882,In_2156);
xnor U283 (N_283,N_30,In_251);
nand U284 (N_284,In_413,In_1975);
xnor U285 (N_285,In_1108,In_587);
xor U286 (N_286,In_1429,In_2438);
nand U287 (N_287,In_1204,In_609);
and U288 (N_288,In_1439,In_625);
xnor U289 (N_289,In_1299,In_967);
and U290 (N_290,In_924,In_2736);
nor U291 (N_291,In_1658,In_1372);
nand U292 (N_292,In_1597,In_2905);
nand U293 (N_293,In_25,In_1064);
xnor U294 (N_294,In_550,In_233);
nand U295 (N_295,In_132,In_1316);
and U296 (N_296,N_118,In_2578);
and U297 (N_297,In_1848,In_689);
nor U298 (N_298,In_37,In_2783);
xor U299 (N_299,In_614,In_2189);
or U300 (N_300,In_955,In_2992);
xnor U301 (N_301,In_1827,In_2689);
or U302 (N_302,In_1790,In_966);
xnor U303 (N_303,In_2174,In_2479);
nand U304 (N_304,In_1546,In_2784);
nand U305 (N_305,In_2528,In_1572);
or U306 (N_306,In_2747,In_2916);
xnor U307 (N_307,In_862,In_794);
and U308 (N_308,In_1795,In_2729);
or U309 (N_309,In_2853,In_1207);
or U310 (N_310,In_2042,In_1365);
nand U311 (N_311,In_588,In_88);
nor U312 (N_312,In_1740,In_302);
xnor U313 (N_313,In_1369,N_194);
nor U314 (N_314,In_241,In_2274);
xor U315 (N_315,In_2278,In_2116);
nor U316 (N_316,In_2986,In_2665);
or U317 (N_317,In_2327,In_485);
xnor U318 (N_318,In_1966,In_2527);
nand U319 (N_319,In_2779,In_2966);
or U320 (N_320,In_1927,In_829);
or U321 (N_321,In_790,In_1721);
or U322 (N_322,In_428,In_2865);
nor U323 (N_323,In_1422,In_1799);
and U324 (N_324,In_2345,In_1447);
nor U325 (N_325,In_2206,In_32);
nand U326 (N_326,In_568,In_971);
nand U327 (N_327,In_2904,In_537);
nor U328 (N_328,In_2476,In_2080);
nand U329 (N_329,In_394,In_2922);
xor U330 (N_330,In_1661,In_2046);
nand U331 (N_331,In_2187,In_1120);
and U332 (N_332,In_567,In_70);
or U333 (N_333,In_276,In_1513);
nand U334 (N_334,In_2435,In_1496);
nand U335 (N_335,In_925,In_734);
nand U336 (N_336,In_1741,In_1411);
or U337 (N_337,In_2436,In_1664);
xnor U338 (N_338,In_2368,In_458);
nand U339 (N_339,In_517,In_2822);
and U340 (N_340,In_2041,In_318);
or U341 (N_341,In_2526,In_2924);
and U342 (N_342,In_816,In_2734);
xor U343 (N_343,N_59,In_311);
or U344 (N_344,In_2913,In_96);
nand U345 (N_345,In_1051,N_180);
nor U346 (N_346,In_2835,In_271);
xor U347 (N_347,In_2496,In_1014);
or U348 (N_348,In_699,In_887);
and U349 (N_349,In_729,In_2506);
and U350 (N_350,In_769,In_830);
nand U351 (N_351,In_1726,In_706);
nor U352 (N_352,In_2908,In_2253);
or U353 (N_353,In_854,In_2911);
nand U354 (N_354,In_2113,In_2129);
nand U355 (N_355,In_436,In_2564);
or U356 (N_356,In_1211,In_2248);
and U357 (N_357,In_736,In_328);
and U358 (N_358,In_1477,In_2192);
nand U359 (N_359,In_2682,In_528);
and U360 (N_360,In_1794,In_2741);
or U361 (N_361,In_767,In_2727);
xor U362 (N_362,In_2285,In_168);
and U363 (N_363,In_951,In_1023);
and U364 (N_364,In_1090,In_716);
xnor U365 (N_365,In_2363,In_247);
or U366 (N_366,In_759,In_722);
xnor U367 (N_367,In_2588,N_179);
nor U368 (N_368,In_741,N_173);
xor U369 (N_369,In_2885,In_1562);
and U370 (N_370,In_2683,In_948);
nor U371 (N_371,In_2821,In_532);
xor U372 (N_372,In_1327,In_1687);
and U373 (N_373,In_613,In_1238);
nor U374 (N_374,In_1961,N_70);
and U375 (N_375,In_1842,In_922);
xnor U376 (N_376,In_1754,In_2618);
or U377 (N_377,In_1943,In_2630);
or U378 (N_378,In_1465,In_2525);
nor U379 (N_379,In_2030,In_108);
nand U380 (N_380,In_1191,In_1749);
nand U381 (N_381,In_690,In_1135);
and U382 (N_382,In_371,In_2289);
or U383 (N_383,In_1591,In_2667);
or U384 (N_384,In_1267,In_2421);
nor U385 (N_385,In_1468,In_472);
nor U386 (N_386,In_774,In_606);
and U387 (N_387,In_1470,In_673);
and U388 (N_388,In_2434,In_2071);
or U389 (N_389,In_2984,N_12);
nand U390 (N_390,In_457,In_1885);
or U391 (N_391,In_2167,In_2619);
nand U392 (N_392,In_1167,In_1677);
nand U393 (N_393,N_57,In_520);
nand U394 (N_394,In_1449,In_1954);
or U395 (N_395,In_1622,In_1306);
xor U396 (N_396,In_755,In_101);
and U397 (N_397,In_2068,In_1902);
or U398 (N_398,In_2318,In_216);
nand U399 (N_399,In_2321,In_502);
or U400 (N_400,In_1718,In_2038);
nor U401 (N_401,In_2021,In_2023);
xor U402 (N_402,N_192,In_230);
nand U403 (N_403,In_1502,In_196);
or U404 (N_404,In_380,In_919);
or U405 (N_405,N_263,In_1526);
and U406 (N_406,In_1940,In_135);
and U407 (N_407,In_1922,In_611);
or U408 (N_408,In_581,In_253);
or U409 (N_409,In_363,In_2699);
nand U410 (N_410,In_970,In_286);
nor U411 (N_411,In_1987,In_2983);
xor U412 (N_412,In_2876,In_1092);
nor U413 (N_413,In_7,N_348);
nand U414 (N_414,In_965,N_278);
xnor U415 (N_415,In_2754,In_1935);
and U416 (N_416,In_2674,In_420);
nand U417 (N_417,N_69,In_2634);
nor U418 (N_418,In_2592,N_153);
nor U419 (N_419,N_312,In_1419);
and U420 (N_420,In_1582,In_507);
and U421 (N_421,In_864,In_2054);
or U422 (N_422,In_261,In_1570);
or U423 (N_423,In_2511,In_407);
xor U424 (N_424,In_2324,In_465);
xor U425 (N_425,N_257,In_2165);
and U426 (N_426,In_2851,In_1501);
nor U427 (N_427,In_2086,In_2560);
and U428 (N_428,In_2233,In_1473);
xnor U429 (N_429,In_1745,In_492);
xor U430 (N_430,In_843,In_2320);
or U431 (N_431,In_772,In_867);
xnor U432 (N_432,In_2782,In_949);
nor U433 (N_433,In_2633,In_2706);
xor U434 (N_434,In_317,In_398);
nor U435 (N_435,In_1840,In_2354);
or U436 (N_436,In_1956,In_2582);
or U437 (N_437,In_579,In_1891);
and U438 (N_438,In_956,In_2259);
nor U439 (N_439,In_1722,In_1706);
or U440 (N_440,In_1463,In_2601);
nand U441 (N_441,In_1127,In_548);
nor U442 (N_442,In_165,N_98);
and U443 (N_443,N_186,In_2802);
nor U444 (N_444,In_1679,In_1855);
or U445 (N_445,In_1029,N_246);
and U446 (N_446,In_2393,In_2210);
xor U447 (N_447,In_1412,In_1441);
or U448 (N_448,In_738,In_2631);
nand U449 (N_449,In_2339,N_11);
or U450 (N_450,In_1563,In_28);
or U451 (N_451,In_370,In_2892);
nor U452 (N_452,In_187,In_213);
xnor U453 (N_453,In_1038,In_2310);
and U454 (N_454,In_2299,In_224);
nor U455 (N_455,N_86,In_1878);
nor U456 (N_456,In_957,In_1436);
or U457 (N_457,N_107,In_2134);
xor U458 (N_458,In_2420,In_487);
and U459 (N_459,In_2684,In_367);
xnor U460 (N_460,N_135,In_2829);
nand U461 (N_461,N_296,In_2875);
nor U462 (N_462,In_1523,In_1317);
nand U463 (N_463,In_2996,In_2474);
nor U464 (N_464,In_1274,N_280);
and U465 (N_465,N_78,In_818);
or U466 (N_466,N_244,In_2330);
xnor U467 (N_467,N_350,In_859);
xor U468 (N_468,In_884,In_2300);
and U469 (N_469,N_182,In_998);
xnor U470 (N_470,N_14,In_2242);
xnor U471 (N_471,N_235,In_67);
nor U472 (N_472,In_2611,In_1506);
or U473 (N_473,N_300,In_1595);
nor U474 (N_474,In_2939,In_2306);
nor U475 (N_475,In_2246,In_1042);
nand U476 (N_476,In_1196,In_2031);
nand U477 (N_477,In_1031,In_2025);
nor U478 (N_478,In_2298,In_2995);
or U479 (N_479,In_381,In_2891);
nand U480 (N_480,In_885,In_1801);
nor U481 (N_481,In_2144,In_2361);
or U482 (N_482,In_1149,In_2954);
nand U483 (N_483,In_2651,In_2977);
and U484 (N_484,In_1617,In_17);
and U485 (N_485,In_666,In_257);
nand U486 (N_486,In_1312,In_2590);
and U487 (N_487,In_1446,In_953);
or U488 (N_488,N_227,In_2952);
nor U489 (N_489,N_237,In_565);
and U490 (N_490,In_1131,In_2142);
and U491 (N_491,In_1383,In_800);
xor U492 (N_492,In_1126,In_1519);
xor U493 (N_493,In_446,N_79);
and U494 (N_494,In_2470,In_874);
xnor U495 (N_495,In_2491,In_214);
or U496 (N_496,In_1480,In_907);
nand U497 (N_497,In_235,In_1012);
and U498 (N_498,N_343,N_81);
nand U499 (N_499,In_2416,In_1348);
nand U500 (N_500,In_2504,N_333);
and U501 (N_501,In_63,N_82);
nand U502 (N_502,In_2640,In_1872);
xor U503 (N_503,In_1334,In_2766);
nand U504 (N_504,In_2159,In_1959);
xnor U505 (N_505,In_1558,In_1181);
xnor U506 (N_506,In_2965,In_1567);
xnor U507 (N_507,In_1485,In_1989);
and U508 (N_508,In_1560,In_2263);
nor U509 (N_509,In_2596,In_1213);
nor U510 (N_510,In_2367,N_331);
nand U511 (N_511,N_308,In_2005);
and U512 (N_512,In_1680,N_281);
or U513 (N_513,In_2374,In_1224);
xnor U514 (N_514,In_708,In_663);
or U515 (N_515,In_1522,In_1757);
and U516 (N_516,In_2570,N_386);
and U517 (N_517,In_2502,In_2514);
xnor U518 (N_518,In_2850,In_1828);
and U519 (N_519,In_275,In_2365);
nand U520 (N_520,In_2175,In_258);
nor U521 (N_521,N_239,In_1823);
or U522 (N_522,In_1178,In_1015);
and U523 (N_523,In_1321,In_220);
nor U524 (N_524,In_899,N_336);
and U525 (N_525,In_2871,In_2166);
nand U526 (N_526,N_255,In_1549);
nand U527 (N_527,In_1395,In_688);
xnor U528 (N_528,In_1829,N_27);
or U529 (N_529,In_1307,In_2452);
or U530 (N_530,In_1187,In_849);
nand U531 (N_531,In_875,In_2961);
and U532 (N_532,In_194,In_2985);
nor U533 (N_533,In_0,In_908);
xnor U534 (N_534,In_287,In_151);
or U535 (N_535,In_1457,In_915);
xnor U536 (N_536,In_2394,In_2687);
and U537 (N_537,In_112,N_193);
or U538 (N_538,In_486,In_2657);
and U539 (N_539,In_127,In_170);
nand U540 (N_540,In_1974,N_241);
xnor U541 (N_541,In_2632,In_2645);
nand U542 (N_542,In_660,In_1688);
xnor U543 (N_543,In_2737,In_1398);
or U544 (N_544,In_147,In_267);
nor U545 (N_545,In_1278,In_1825);
xnor U546 (N_546,In_2581,In_797);
or U547 (N_547,In_2585,In_1243);
nand U548 (N_548,N_325,In_2117);
nor U549 (N_549,In_880,N_335);
xnor U550 (N_550,N_184,In_1330);
xor U551 (N_551,In_1689,N_114);
nand U552 (N_552,In_1675,In_284);
nand U553 (N_553,In_2214,In_1385);
or U554 (N_554,In_185,In_1103);
nand U555 (N_555,In_691,In_219);
nor U556 (N_556,In_1871,In_2331);
nor U557 (N_557,In_323,In_2680);
and U558 (N_558,In_518,In_2988);
xor U559 (N_559,In_2636,In_2262);
xnor U560 (N_560,In_205,In_2472);
xnor U561 (N_561,In_2432,In_2029);
nor U562 (N_562,In_1097,In_1946);
xnor U563 (N_563,In_2497,In_571);
nand U564 (N_564,In_2898,In_563);
nor U565 (N_565,In_1113,N_183);
nor U566 (N_566,In_303,In_438);
and U567 (N_567,In_1547,In_2845);
and U568 (N_568,N_146,In_521);
or U569 (N_569,In_1368,In_1667);
and U570 (N_570,In_602,In_1640);
xnor U571 (N_571,In_207,In_604);
nor U572 (N_572,In_2664,N_0);
nand U573 (N_573,In_1453,In_703);
nand U574 (N_574,In_2714,N_217);
and U575 (N_575,In_566,In_748);
xnor U576 (N_576,In_1905,In_2419);
nor U577 (N_577,In_2928,In_2412);
xor U578 (N_578,In_20,In_1746);
xnor U579 (N_579,N_206,In_1148);
or U580 (N_580,N_58,In_494);
or U581 (N_581,In_2317,In_440);
or U582 (N_582,In_91,In_2447);
and U583 (N_583,N_250,In_1865);
xnor U584 (N_584,N_142,N_96);
and U585 (N_585,In_301,In_2110);
nand U586 (N_586,In_2045,In_1929);
xor U587 (N_587,In_2137,In_2446);
or U588 (N_588,In_1471,N_279);
or U589 (N_589,In_2931,N_313);
and U590 (N_590,In_1049,In_2893);
nand U591 (N_591,In_1498,N_268);
nand U592 (N_592,In_984,In_238);
nor U593 (N_593,In_745,In_1921);
nor U594 (N_594,In_886,In_2151);
and U595 (N_595,In_2842,In_1360);
nor U596 (N_596,In_133,In_2805);
and U597 (N_597,In_2587,In_1765);
nand U598 (N_598,In_1897,In_943);
xnor U599 (N_599,In_243,In_2063);
nand U600 (N_600,In_1691,In_1047);
nand U601 (N_601,In_710,In_1831);
and U602 (N_602,N_508,In_2138);
or U603 (N_603,In_2410,In_1358);
or U604 (N_604,In_2243,In_1491);
nor U605 (N_605,In_2796,In_2670);
and U606 (N_606,In_1003,In_2767);
or U607 (N_607,In_1489,In_2943);
xnor U608 (N_608,In_1367,In_2340);
xnor U609 (N_609,In_13,In_709);
nand U610 (N_610,N_467,In_1493);
nand U611 (N_611,N_535,In_2810);
nor U612 (N_612,In_2907,In_1472);
or U613 (N_613,In_2353,In_2241);
nor U614 (N_614,In_2430,In_182);
or U615 (N_615,N_585,In_1670);
and U616 (N_616,In_1550,In_1205);
xnor U617 (N_617,In_1217,In_1214);
nand U618 (N_618,In_1960,In_2855);
and U619 (N_619,N_178,In_468);
xnor U620 (N_620,In_702,In_386);
and U621 (N_621,In_1347,N_23);
xor U622 (N_622,In_455,In_2007);
nor U623 (N_623,N_355,In_1962);
nand U624 (N_624,N_318,N_164);
or U625 (N_625,N_556,In_1458);
xor U626 (N_626,N_320,In_2200);
and U627 (N_627,In_2573,In_633);
and U628 (N_628,In_2079,In_1892);
xnor U629 (N_629,N_62,In_2170);
xnor U630 (N_630,In_297,In_1672);
and U631 (N_631,In_1843,N_225);
nand U632 (N_632,N_570,In_570);
or U633 (N_633,In_333,In_1235);
nand U634 (N_634,In_2377,N_495);
nor U635 (N_635,In_2723,N_55);
nor U636 (N_636,In_350,In_2610);
or U637 (N_637,N_547,In_773);
nor U638 (N_638,In_2313,In_742);
xor U639 (N_639,In_2095,In_1189);
xnor U640 (N_640,In_2906,In_1796);
and U641 (N_641,In_751,In_1985);
and U642 (N_642,N_226,In_1088);
and U643 (N_643,In_1598,In_1524);
or U644 (N_644,In_466,In_2971);
nand U645 (N_645,N_382,In_1583);
xnor U646 (N_646,In_961,N_459);
xnor U647 (N_647,In_1631,In_593);
nor U648 (N_648,In_638,In_650);
nor U649 (N_649,In_760,N_371);
nand U650 (N_650,N_67,In_2372);
xor U651 (N_651,N_526,In_535);
or U652 (N_652,N_532,In_1531);
nor U653 (N_653,In_316,N_573);
and U654 (N_654,N_529,N_460);
xor U655 (N_655,N_478,In_491);
and U656 (N_656,In_573,In_585);
xnor U657 (N_657,In_644,In_2256);
or U658 (N_658,In_1059,In_2960);
and U659 (N_659,In_2360,In_105);
or U660 (N_660,In_1958,In_1836);
and U661 (N_661,In_2577,In_1361);
and U662 (N_662,In_27,N_97);
nand U663 (N_663,N_406,In_1752);
nand U664 (N_664,In_903,In_2172);
nor U665 (N_665,In_1626,N_6);
and U666 (N_666,In_1862,In_424);
and U667 (N_667,In_2819,In_2193);
nand U668 (N_668,In_422,In_2322);
and U669 (N_669,N_384,In_430);
and U670 (N_670,N_576,In_2725);
xnor U671 (N_671,In_1483,In_2297);
and U672 (N_672,In_1271,In_1708);
nand U673 (N_673,In_405,In_610);
nand U674 (N_674,In_2566,In_2864);
or U675 (N_675,In_2743,In_1313);
xor U676 (N_676,In_1256,In_1318);
nor U677 (N_677,In_2724,In_2510);
nand U678 (N_678,In_2899,N_540);
nand U679 (N_679,In_600,In_423);
or U680 (N_680,In_780,In_434);
nand U681 (N_681,In_1130,N_380);
xor U682 (N_682,In_1774,In_897);
xnor U683 (N_683,In_665,N_10);
and U684 (N_684,In_358,In_1585);
xnor U685 (N_685,In_390,In_2579);
nor U686 (N_686,N_473,In_1393);
nand U687 (N_687,In_1144,In_1414);
and U688 (N_688,In_186,In_1183);
nand U689 (N_689,N_518,In_1510);
and U690 (N_690,In_2644,In_2307);
and U691 (N_691,N_358,N_44);
xor U692 (N_692,In_448,In_2373);
and U693 (N_693,In_1032,In_2083);
xor U694 (N_694,In_2006,N_357);
and U695 (N_695,In_2462,In_2464);
or U696 (N_696,In_2093,In_1881);
xor U697 (N_697,In_2196,In_2838);
or U698 (N_698,In_621,In_763);
and U699 (N_699,In_942,N_537);
nor U700 (N_700,N_506,In_534);
and U701 (N_701,In_1838,In_656);
or U702 (N_702,In_1443,N_172);
or U703 (N_703,In_310,In_2388);
or U704 (N_704,N_489,N_212);
xor U705 (N_705,N_104,In_1920);
or U706 (N_706,N_456,N_233);
nand U707 (N_707,In_1907,In_1028);
and U708 (N_708,In_416,N_28);
nor U709 (N_709,N_511,In_721);
and U710 (N_710,In_1561,In_1870);
nor U711 (N_711,In_1259,N_391);
nand U712 (N_712,In_1553,In_1918);
nor U713 (N_713,In_2735,In_1476);
and U714 (N_714,In_1176,N_247);
and U715 (N_715,N_65,N_54);
nand U716 (N_716,In_2679,N_407);
nand U717 (N_717,In_368,In_1821);
nor U718 (N_718,In_1169,In_339);
xor U719 (N_719,In_447,In_576);
nor U720 (N_720,In_1565,In_1326);
or U721 (N_721,In_47,In_1786);
nor U722 (N_722,In_2659,In_2268);
xnor U723 (N_723,In_2399,In_2160);
nor U724 (N_724,In_1300,In_2010);
nand U725 (N_725,In_107,In_130);
and U726 (N_726,In_2501,In_1761);
xnor U727 (N_727,In_2337,In_2405);
nor U728 (N_728,In_981,In_473);
xnor U729 (N_729,In_572,N_116);
or U730 (N_730,N_149,N_499);
and U731 (N_731,In_1643,In_496);
xnor U732 (N_732,N_530,In_2188);
xnor U733 (N_733,In_336,N_201);
and U734 (N_734,N_123,In_2551);
or U735 (N_735,In_598,N_75);
xor U736 (N_736,In_1619,In_676);
nand U737 (N_737,In_2620,In_477);
nand U738 (N_738,In_2238,N_131);
nand U739 (N_739,In_1402,In_163);
nand U740 (N_740,N_363,In_784);
or U741 (N_741,In_1249,N_121);
nor U742 (N_742,N_39,In_2326);
and U743 (N_743,N_589,In_1290);
nor U744 (N_744,In_242,N_474);
or U745 (N_745,In_2797,N_29);
nor U746 (N_746,N_411,N_25);
and U747 (N_747,In_2195,In_441);
or U748 (N_748,In_2231,In_796);
and U749 (N_749,In_2301,In_2953);
xor U750 (N_750,In_1006,In_1394);
and U751 (N_751,In_1787,N_191);
xor U752 (N_752,N_322,In_2658);
nand U753 (N_753,In_149,In_2469);
and U754 (N_754,In_2379,In_1030);
nor U755 (N_755,In_2923,In_2455);
and U756 (N_756,In_728,In_1894);
nand U757 (N_757,In_1735,In_2009);
xnor U758 (N_758,N_457,In_963);
xor U759 (N_759,In_1118,In_444);
nand U760 (N_760,In_1618,In_2543);
or U761 (N_761,N_575,In_2150);
and U762 (N_762,N_120,In_183);
nand U763 (N_763,In_2787,In_2972);
and U764 (N_764,N_137,In_1095);
or U765 (N_765,In_1281,In_2281);
nand U766 (N_766,N_436,In_1895);
or U767 (N_767,In_1877,In_2993);
and U768 (N_768,N_162,In_805);
xor U769 (N_769,In_369,In_2771);
nand U770 (N_770,N_63,In_2591);
and U771 (N_771,In_1225,In_478);
nor U772 (N_772,In_1534,N_367);
or U773 (N_773,In_2874,N_71);
xor U774 (N_774,In_651,In_280);
xnor U775 (N_775,N_222,N_45);
nand U776 (N_776,N_292,In_2153);
and U777 (N_777,In_1809,In_986);
nand U778 (N_778,In_2271,In_2351);
nand U779 (N_779,N_372,In_2381);
or U780 (N_780,In_1986,N_215);
xnor U781 (N_781,N_344,N_471);
and U782 (N_782,In_1579,N_36);
or U783 (N_783,N_454,N_40);
or U784 (N_784,In_1807,In_443);
nand U785 (N_785,In_484,In_2546);
nand U786 (N_786,In_2342,In_2000);
and U787 (N_787,In_42,N_476);
nand U788 (N_788,N_496,In_1163);
nand U789 (N_789,In_2378,In_2490);
or U790 (N_790,In_968,In_409);
xor U791 (N_791,In_1694,In_720);
nor U792 (N_792,In_2508,In_1251);
xnor U793 (N_793,In_1288,In_2598);
nand U794 (N_794,In_387,N_577);
and U795 (N_795,In_2335,In_2349);
or U796 (N_796,In_2065,N_269);
nor U797 (N_797,In_1715,In_749);
and U798 (N_798,In_223,In_145);
or U799 (N_799,In_1237,In_2704);
nand U800 (N_800,N_479,In_1543);
and U801 (N_801,In_2176,N_398);
and U802 (N_802,In_2409,In_2925);
nor U803 (N_803,N_53,N_776);
xor U804 (N_804,In_871,In_698);
and U805 (N_805,In_2494,In_2411);
or U806 (N_806,In_1075,N_252);
xnor U807 (N_807,In_2612,N_417);
nand U808 (N_808,In_1230,N_316);
and U809 (N_809,N_642,In_2282);
nor U810 (N_810,N_176,In_1788);
and U811 (N_811,In_539,In_2325);
and U812 (N_812,N_742,In_1401);
or U813 (N_813,N_639,In_2868);
and U814 (N_814,In_2273,In_1541);
and U815 (N_815,In_2115,N_578);
nand U816 (N_816,In_1709,In_264);
nand U817 (N_817,In_2157,In_123);
nand U818 (N_818,In_1832,In_2935);
or U819 (N_819,In_152,In_960);
nor U820 (N_820,In_1384,In_1648);
and U821 (N_821,In_1044,In_726);
nand U822 (N_822,In_1248,In_988);
nor U823 (N_823,In_2750,In_1208);
nor U824 (N_824,In_1188,In_248);
nor U825 (N_825,In_68,N_762);
xnor U826 (N_826,In_254,In_269);
and U827 (N_827,In_2505,N_490);
and U828 (N_828,N_303,N_670);
nor U829 (N_829,In_1645,In_1967);
or U830 (N_830,N_715,In_1589);
and U831 (N_831,N_721,In_530);
and U832 (N_832,In_375,In_2442);
xor U833 (N_833,N_49,In_1143);
or U834 (N_834,In_1969,N_161);
nand U835 (N_835,In_1352,In_2182);
nor U836 (N_836,In_713,N_775);
nor U837 (N_837,In_2094,In_2014);
nand U838 (N_838,In_1155,In_227);
and U839 (N_839,N_442,N_310);
nand U840 (N_840,In_462,N_691);
nor U841 (N_841,In_1104,In_2152);
nand U842 (N_842,N_199,In_1258);
or U843 (N_843,N_141,N_758);
nor U844 (N_844,In_944,In_1146);
nor U845 (N_845,N_550,In_1525);
nor U846 (N_846,N_795,In_1808);
xor U847 (N_847,N_332,In_639);
nand U848 (N_848,In_1342,In_640);
and U849 (N_849,In_1888,In_1601);
and U850 (N_850,In_2183,N_681);
xor U851 (N_851,N_746,In_2097);
and U852 (N_852,N_466,In_93);
or U853 (N_853,In_628,In_999);
and U854 (N_854,N_453,In_1571);
or U855 (N_855,In_542,In_1410);
xnor U856 (N_856,In_1481,N_720);
or U857 (N_857,N_469,In_658);
nand U858 (N_858,In_1228,In_522);
nand U859 (N_859,In_670,In_2606);
and U860 (N_860,In_1724,N_446);
or U861 (N_861,In_138,N_311);
or U862 (N_862,In_2638,In_848);
and U863 (N_863,In_481,In_1223);
nor U864 (N_864,In_1699,In_471);
nor U865 (N_865,In_952,N_688);
and U866 (N_866,In_1530,In_2757);
and U867 (N_867,In_1096,In_2926);
nor U868 (N_868,In_159,In_2477);
nand U869 (N_869,N_764,In_2730);
xnor U870 (N_870,In_996,N_784);
or U871 (N_871,In_1199,In_2862);
xnor U872 (N_872,N_749,N_788);
nor U873 (N_873,N_728,N_420);
or U874 (N_874,In_2002,In_391);
and U875 (N_875,N_101,In_2831);
and U876 (N_876,In_1043,In_1060);
or U877 (N_877,In_1115,In_1548);
and U878 (N_878,In_2344,In_290);
nand U879 (N_879,N_592,N_705);
xor U880 (N_880,In_501,In_2312);
nand U881 (N_881,In_1351,N_37);
nor U882 (N_882,In_1972,In_2764);
xor U883 (N_883,In_2355,In_2125);
xnor U884 (N_884,In_783,In_1495);
and U885 (N_885,N_409,In_2964);
nand U886 (N_886,In_2710,N_47);
nor U887 (N_887,N_607,N_763);
nand U888 (N_888,N_32,N_452);
xor U889 (N_889,In_2485,In_1666);
and U890 (N_890,In_2158,In_799);
and U891 (N_891,N_455,In_1822);
nand U892 (N_892,In_2102,N_433);
or U893 (N_893,In_1624,N_368);
nor U894 (N_894,In_404,In_2744);
nor U895 (N_895,N_359,In_81);
xnor U896 (N_896,In_2718,In_332);
nand U897 (N_897,In_1655,In_1568);
or U898 (N_898,N_475,In_822);
or U899 (N_899,N_219,In_2303);
nand U900 (N_900,In_2329,In_21);
nand U901 (N_901,In_1005,N_435);
nor U902 (N_902,N_22,In_1335);
nand U903 (N_903,In_1973,In_1683);
xnor U904 (N_904,In_1066,N_277);
nor U905 (N_905,N_349,In_506);
nand U906 (N_906,N_725,In_557);
nand U907 (N_907,In_2180,N_744);
and U908 (N_908,In_1627,In_2082);
and U909 (N_909,In_2540,In_2957);
and U910 (N_910,N_687,In_2719);
nor U911 (N_911,In_395,In_2449);
nor U912 (N_912,In_1040,N_224);
and U913 (N_913,In_2642,In_2275);
xor U914 (N_914,In_1712,In_2794);
and U915 (N_915,N_501,In_2976);
or U916 (N_916,In_657,In_1170);
and U917 (N_917,In_2979,In_2531);
xor U918 (N_918,N_797,In_901);
nand U919 (N_919,In_1344,N_523);
or U920 (N_920,N_498,In_2785);
nor U921 (N_921,In_1106,In_2825);
nand U922 (N_922,In_1990,In_814);
and U923 (N_923,In_2968,In_234);
and U924 (N_924,In_2194,N_590);
and U925 (N_925,In_771,In_1297);
xnor U926 (N_926,In_71,N_793);
nor U927 (N_927,In_2473,In_526);
nor U928 (N_928,In_2660,N_422);
or U929 (N_929,In_377,N_159);
nand U930 (N_930,In_38,N_752);
and U931 (N_931,In_976,N_160);
or U932 (N_932,In_648,N_195);
xnor U933 (N_933,In_1253,In_2387);
nor U934 (N_934,In_308,In_2481);
xnor U935 (N_935,In_674,In_1518);
nand U936 (N_936,In_2858,In_1853);
xnor U937 (N_937,In_1240,In_1609);
xnor U938 (N_938,N_122,N_262);
nor U939 (N_939,In_2247,N_392);
nor U940 (N_940,In_1569,In_2234);
or U941 (N_941,In_1375,In_1811);
or U942 (N_942,In_2019,In_1399);
nand U943 (N_943,In_2033,In_934);
xor U944 (N_944,In_1911,In_347);
xnor U945 (N_945,N_291,In_868);
or U946 (N_946,In_2940,In_2752);
nor U947 (N_947,N_696,N_611);
and U948 (N_948,In_150,In_1269);
nor U949 (N_949,N_42,N_470);
xnor U950 (N_950,In_543,N_521);
or U951 (N_951,In_1156,N_794);
or U952 (N_952,N_561,In_2509);
or U953 (N_953,N_485,N_492);
xor U954 (N_954,In_2726,In_2040);
xor U955 (N_955,In_411,In_1229);
or U956 (N_956,In_2352,In_1338);
xor U957 (N_957,In_429,In_857);
or U958 (N_958,In_1026,In_1198);
nor U959 (N_959,In_1604,In_202);
nand U960 (N_960,In_1345,In_624);
xor U961 (N_961,In_1184,N_361);
nor U962 (N_962,In_681,N_669);
xnor U963 (N_963,In_1702,In_561);
or U964 (N_964,N_628,In_2773);
nand U965 (N_965,In_2413,N_780);
nand U966 (N_966,N_610,N_289);
xor U967 (N_967,N_772,In_342);
xnor U968 (N_968,In_2944,In_508);
xor U969 (N_969,In_1937,In_991);
or U970 (N_970,In_2015,In_1998);
xor U971 (N_971,In_2290,In_538);
nand U972 (N_972,In_1970,N_68);
xnor U973 (N_973,In_1339,N_1);
nand U974 (N_974,In_2625,In_1174);
xor U975 (N_975,N_649,In_615);
nor U976 (N_976,In_74,N_798);
nand U977 (N_977,In_191,N_594);
and U978 (N_978,In_1165,In_2541);
xnor U979 (N_979,N_674,N_127);
or U980 (N_980,N_240,N_216);
nor U981 (N_981,In_495,In_2909);
xnor U982 (N_982,N_144,In_2512);
nor U983 (N_983,N_77,N_557);
xnor U984 (N_984,N_761,N_574);
or U985 (N_985,N_444,In_1875);
or U986 (N_986,In_1309,In_1841);
nor U987 (N_987,In_158,N_500);
and U988 (N_988,In_1322,In_2495);
xor U989 (N_989,In_2026,N_315);
nand U990 (N_990,In_146,In_553);
xnor U991 (N_991,N_481,In_866);
nand U992 (N_992,N_527,N_364);
xnor U993 (N_993,N_522,In_1440);
or U994 (N_994,N_560,In_29);
nor U995 (N_995,N_638,In_1873);
nor U996 (N_996,In_1580,In_2507);
nor U997 (N_997,In_184,In_2563);
nor U998 (N_998,N_41,In_2036);
nand U999 (N_999,In_2066,In_2709);
nand U1000 (N_1000,In_719,In_620);
xnor U1001 (N_1001,In_1590,In_217);
nand U1002 (N_1002,In_2201,In_2020);
and U1003 (N_1003,In_2389,N_549);
and U1004 (N_1004,In_2146,In_1515);
nor U1005 (N_1005,In_2185,In_1992);
nand U1006 (N_1006,N_260,N_889);
and U1007 (N_1007,In_1652,In_1731);
nor U1008 (N_1008,N_947,In_1529);
or U1009 (N_1009,N_203,In_2555);
and U1010 (N_1010,In_2397,N_493);
nand U1011 (N_1011,In_2346,In_1533);
xnor U1012 (N_1012,In_2164,N_713);
or U1013 (N_1013,N_397,In_2204);
and U1014 (N_1014,In_2828,N_445);
or U1015 (N_1015,N_309,In_2202);
nand U1016 (N_1016,In_201,In_2109);
or U1017 (N_1017,In_60,In_357);
or U1018 (N_1018,In_2044,In_2571);
nand U1019 (N_1019,In_1654,N_555);
nand U1020 (N_1020,In_1833,N_593);
nand U1021 (N_1021,In_902,N_404);
nand U1022 (N_1022,In_102,N_913);
nor U1023 (N_1023,In_2140,N_820);
or U1024 (N_1024,In_2798,In_178);
nor U1025 (N_1025,In_155,In_1913);
and U1026 (N_1026,In_1333,N_379);
and U1027 (N_1027,In_2266,In_451);
and U1028 (N_1028,In_337,In_2917);
nand U1029 (N_1029,In_1304,In_812);
nand U1030 (N_1030,In_1381,N_341);
and U1031 (N_1031,N_686,N_329);
nor U1032 (N_1032,In_938,In_1864);
and U1033 (N_1033,In_2776,In_1634);
nor U1034 (N_1034,N_253,In_1900);
xor U1035 (N_1035,N_232,N_988);
nand U1036 (N_1036,In_1082,In_188);
nand U1037 (N_1037,N_591,In_861);
and U1038 (N_1038,In_1182,N_321);
and U1039 (N_1039,In_2609,In_879);
nor U1040 (N_1040,N_884,In_2091);
and U1041 (N_1041,N_629,N_274);
and U1042 (N_1042,In_1824,In_2677);
xor U1043 (N_1043,In_225,N_839);
or U1044 (N_1044,N_324,In_2866);
xnor U1045 (N_1045,In_2647,In_1542);
nand U1046 (N_1046,N_74,In_1445);
xor U1047 (N_1047,In_512,In_1425);
and U1048 (N_1048,N_826,In_1424);
or U1049 (N_1049,N_158,In_1988);
nor U1050 (N_1050,N_234,In_1036);
xor U1051 (N_1051,In_266,N_242);
or U1052 (N_1052,In_2663,In_2524);
xnor U1053 (N_1053,N_138,N_157);
or U1054 (N_1054,In_2179,In_515);
or U1055 (N_1055,N_722,N_957);
xor U1056 (N_1056,In_239,N_937);
and U1057 (N_1057,N_297,In_2681);
xnor U1058 (N_1058,In_937,N_72);
nor U1059 (N_1059,N_271,In_1260);
or U1060 (N_1060,In_832,In_294);
or U1061 (N_1061,In_1291,N_846);
xnor U1062 (N_1062,N_128,In_11);
nand U1063 (N_1063,In_1311,N_385);
nor U1064 (N_1064,In_1054,In_2104);
nand U1065 (N_1065,N_534,In_2376);
xnor U1066 (N_1066,In_463,In_2793);
or U1067 (N_1067,In_142,N_437);
or U1068 (N_1068,N_356,In_2550);
nor U1069 (N_1069,N_563,In_635);
nand U1070 (N_1070,N_622,In_439);
nor U1071 (N_1071,N_129,In_2224);
or U1072 (N_1072,N_941,In_696);
and U1073 (N_1073,In_2583,In_788);
xor U1074 (N_1074,In_1705,N_757);
and U1075 (N_1075,N_258,N_602);
nor U1076 (N_1076,In_807,N_80);
nand U1077 (N_1077,In_1685,In_559);
xor U1078 (N_1078,In_2565,In_2108);
nand U1079 (N_1079,In_2103,In_2424);
and U1080 (N_1080,N_814,N_971);
xnor U1081 (N_1081,In_2711,In_1976);
nand U1082 (N_1082,In_2553,N_626);
nand U1083 (N_1083,In_1350,In_299);
xor U1084 (N_1084,N_514,In_1994);
xnor U1085 (N_1085,N_582,In_40);
and U1086 (N_1086,In_2781,In_888);
xor U1087 (N_1087,N_400,N_66);
xnor U1088 (N_1088,N_497,N_841);
nor U1089 (N_1089,In_2696,N_87);
xor U1090 (N_1090,In_1763,In_1630);
nor U1091 (N_1091,In_2833,In_2127);
or U1092 (N_1092,N_676,N_932);
nor U1093 (N_1093,In_2249,In_2839);
or U1094 (N_1094,N_963,N_709);
nand U1095 (N_1095,N_650,N_636);
or U1096 (N_1096,N_92,In_842);
or U1097 (N_1097,In_1771,In_1887);
and U1098 (N_1098,In_2897,In_1947);
or U1099 (N_1099,In_226,In_1791);
and U1100 (N_1100,N_850,In_950);
xor U1101 (N_1101,In_2945,In_475);
nor U1102 (N_1102,In_555,N_995);
nand U1103 (N_1103,N_282,In_2237);
or U1104 (N_1104,N_414,In_2795);
or U1105 (N_1105,In_1802,In_1117);
xnor U1106 (N_1106,In_1880,In_1532);
xor U1107 (N_1107,In_1035,N_218);
xnor U1108 (N_1108,N_756,In_554);
or U1109 (N_1109,N_633,In_1478);
and U1110 (N_1110,In_2011,In_608);
xor U1111 (N_1111,N_860,In_121);
and U1112 (N_1112,N_559,In_1315);
nand U1113 (N_1113,In_910,N_229);
xor U1114 (N_1114,N_621,N_685);
or U1115 (N_1115,N_606,N_680);
or U1116 (N_1116,In_2099,In_1008);
xnor U1117 (N_1117,In_2652,In_2356);
or U1118 (N_1118,N_858,In_1057);
xnor U1119 (N_1119,N_419,N_805);
or U1120 (N_1120,In_2453,In_2112);
or U1121 (N_1121,In_732,In_2628);
or U1122 (N_1122,In_747,In_1041);
or U1123 (N_1123,N_739,In_2593);
nor U1124 (N_1124,In_920,N_402);
nand U1125 (N_1125,N_507,In_1728);
xor U1126 (N_1126,N_586,N_553);
and U1127 (N_1127,In_1061,N_926);
or U1128 (N_1128,In_2800,N_736);
nand U1129 (N_1129,In_2938,In_2208);
xor U1130 (N_1130,In_272,N_996);
nor U1131 (N_1131,In_136,N_981);
or U1132 (N_1132,N_125,N_283);
or U1133 (N_1133,N_410,In_2761);
or U1134 (N_1134,In_2252,N_838);
and U1135 (N_1135,N_15,N_922);
xnor U1136 (N_1136,N_245,N_430);
or U1137 (N_1137,In_2600,In_2119);
nor U1138 (N_1138,N_284,In_1100);
or U1139 (N_1139,In_1686,N_921);
nor U1140 (N_1140,In_39,In_1302);
or U1141 (N_1141,In_1978,In_2688);
or U1142 (N_1142,In_2418,N_155);
and U1143 (N_1143,In_1068,In_177);
xor U1144 (N_1144,In_245,N_907);
and U1145 (N_1145,In_1021,N_934);
and U1146 (N_1146,N_869,In_2482);
or U1147 (N_1147,In_1509,In_1939);
and U1148 (N_1148,In_304,N_188);
or U1149 (N_1149,N_632,N_347);
nor U1150 (N_1150,In_2357,N_958);
xor U1151 (N_1151,In_1756,In_2762);
xor U1152 (N_1152,N_565,N_668);
nand U1153 (N_1153,N_878,In_1814);
nor U1154 (N_1154,In_1592,In_2849);
nand U1155 (N_1155,In_1487,In_2143);
or U1156 (N_1156,N_623,In_1775);
or U1157 (N_1157,N_351,N_866);
nand U1158 (N_1158,In_1625,N_615);
and U1159 (N_1159,In_2751,In_2951);
nand U1160 (N_1160,In_410,N_458);
or U1161 (N_1161,N_657,N_874);
and U1162 (N_1162,In_2454,In_2034);
nor U1163 (N_1163,N_787,N_825);
xnor U1164 (N_1164,In_2260,In_2098);
nand U1165 (N_1165,In_1168,In_1280);
nand U1166 (N_1166,In_2818,In_156);
xnor U1167 (N_1167,In_2547,N_461);
nand U1168 (N_1168,N_533,N_671);
nor U1169 (N_1169,N_774,N_551);
nand U1170 (N_1170,In_623,N_865);
nor U1171 (N_1171,N_450,In_2641);
and U1172 (N_1172,N_377,In_906);
and U1173 (N_1173,In_1053,In_1110);
and U1174 (N_1174,N_723,In_2076);
and U1175 (N_1175,N_151,In_2650);
nor U1176 (N_1176,In_66,In_75);
nor U1177 (N_1177,In_2500,In_1179);
or U1178 (N_1178,N_509,N_675);
nand U1179 (N_1179,N_727,In_1359);
nor U1180 (N_1180,In_2867,In_1681);
nor U1181 (N_1181,In_2769,In_1748);
xor U1182 (N_1182,In_401,N_896);
nand U1183 (N_1183,In_2746,In_2178);
xnor U1184 (N_1184,In_4,In_1697);
and U1185 (N_1185,In_2693,N_148);
nor U1186 (N_1186,In_2643,In_2791);
nor U1187 (N_1187,N_991,N_729);
xor U1188 (N_1188,N_596,N_524);
nand U1189 (N_1189,N_248,In_2824);
nand U1190 (N_1190,In_41,In_2998);
nand U1191 (N_1191,In_1744,In_2177);
nand U1192 (N_1192,N_544,N_304);
and U1193 (N_1193,In_1018,In_55);
nand U1194 (N_1194,In_1606,In_1737);
and U1195 (N_1195,N_525,In_330);
or U1196 (N_1196,N_111,In_2788);
nand U1197 (N_1197,In_2315,In_2806);
nor U1198 (N_1198,In_2649,In_1863);
xor U1199 (N_1199,N_482,N_401);
xor U1200 (N_1200,N_726,N_604);
or U1201 (N_1201,N_1006,N_754);
nor U1202 (N_1202,N_427,N_1180);
nand U1203 (N_1203,N_1011,In_1239);
xnor U1204 (N_1204,In_1951,In_2197);
nor U1205 (N_1205,In_2843,N_1170);
or U1206 (N_1206,In_148,N_1054);
nor U1207 (N_1207,N_719,N_1161);
xnor U1208 (N_1208,N_613,In_1161);
xnor U1209 (N_1209,N_900,In_2132);
nand U1210 (N_1210,In_1629,In_2728);
and U1211 (N_1211,N_868,In_629);
or U1212 (N_1212,In_2884,In_1390);
or U1213 (N_1213,In_2881,N_38);
or U1214 (N_1214,N_288,In_1866);
and U1215 (N_1215,In_904,In_2890);
nor U1216 (N_1216,In_589,In_700);
xnor U1217 (N_1217,In_544,N_969);
or U1218 (N_1218,In_362,N_334);
and U1219 (N_1219,In_360,In_2488);
or U1220 (N_1220,In_1671,In_273);
or U1221 (N_1221,N_584,N_480);
nand U1222 (N_1222,In_841,N_989);
or U1223 (N_1223,N_956,In_1045);
or U1224 (N_1224,In_697,In_124);
xnor U1225 (N_1225,In_2518,In_1879);
xnor U1226 (N_1226,In_1244,N_634);
and U1227 (N_1227,N_684,N_942);
xor U1228 (N_1228,In_2218,N_890);
and U1229 (N_1229,N_943,In_100);
nor U1230 (N_1230,In_62,In_2141);
and U1231 (N_1231,N_1064,In_1739);
xor U1232 (N_1232,In_1164,In_372);
or U1233 (N_1233,In_141,In_2676);
xnor U1234 (N_1234,N_513,In_2440);
nor U1235 (N_1235,In_892,In_959);
and U1236 (N_1236,In_1134,N_955);
nor U1237 (N_1237,N_464,N_365);
xor U1238 (N_1238,N_809,In_1151);
nand U1239 (N_1239,In_675,In_1004);
nor U1240 (N_1240,In_1172,In_2604);
xor U1241 (N_1241,N_1155,In_2626);
xor U1242 (N_1242,In_1852,In_164);
or U1243 (N_1243,In_2967,In_1417);
xnor U1244 (N_1244,N_512,In_2427);
nand U1245 (N_1245,In_291,In_2003);
xor U1246 (N_1246,N_783,N_1152);
nand U1247 (N_1247,In_578,In_2559);
nand U1248 (N_1248,In_583,N_609);
nor U1249 (N_1249,In_249,In_2383);
or U1250 (N_1250,In_645,In_1461);
nand U1251 (N_1251,In_1928,In_334);
nand U1252 (N_1252,In_2220,N_1126);
or U1253 (N_1253,N_1158,In_2213);
xor U1254 (N_1254,In_2515,In_104);
xnor U1255 (N_1255,In_2279,N_103);
nor U1256 (N_1256,In_1413,In_1555);
nor U1257 (N_1257,In_26,In_231);
and U1258 (N_1258,N_275,In_889);
nor U1259 (N_1259,N_975,In_591);
xor U1260 (N_1260,In_2920,In_1027);
xor U1261 (N_1261,In_882,In_2556);
and U1262 (N_1262,In_1521,In_1971);
and U1263 (N_1263,In_2302,In_57);
nand U1264 (N_1264,In_1586,In_634);
or U1265 (N_1265,N_24,N_569);
and U1266 (N_1266,N_849,In_746);
or U1267 (N_1267,In_2981,N_202);
and U1268 (N_1268,In_881,In_1077);
nand U1269 (N_1269,In_2982,In_1034);
nand U1270 (N_1270,N_1061,In_1584);
xor U1271 (N_1271,N_89,In_836);
or U1272 (N_1272,In_804,In_511);
nand U1273 (N_1273,In_883,In_1682);
xor U1274 (N_1274,In_819,N_541);
xor U1275 (N_1275,N_378,N_993);
xor U1276 (N_1276,In_2635,N_645);
xnor U1277 (N_1277,N_905,In_1963);
nor U1278 (N_1278,In_53,In_2291);
xnor U1279 (N_1279,In_597,In_2758);
xor U1280 (N_1280,N_375,N_1191);
nor U1281 (N_1281,In_2672,N_747);
or U1282 (N_1282,In_900,In_954);
nand U1283 (N_1283,N_735,In_449);
nor U1284 (N_1284,N_338,In_1925);
nor U1285 (N_1285,N_486,In_1137);
xnor U1286 (N_1286,N_1123,In_630);
or U1287 (N_1287,N_786,In_1263);
nor U1288 (N_1288,In_482,In_500);
nand U1289 (N_1289,N_682,N_935);
nand U1290 (N_1290,N_833,N_1140);
or U1291 (N_1291,N_307,N_821);
and U1292 (N_1292,N_249,In_672);
and U1293 (N_1293,In_831,N_1039);
and U1294 (N_1294,N_76,N_702);
xnor U1295 (N_1295,In_309,In_2816);
nand U1296 (N_1296,In_1644,In_1665);
or U1297 (N_1297,N_83,In_2359);
xor U1298 (N_1298,In_2334,In_1093);
or U1299 (N_1299,N_773,In_1613);
and U1300 (N_1300,N_1034,In_2371);
xnor U1301 (N_1301,In_2467,In_1578);
xor U1302 (N_1302,N_983,In_34);
nand U1303 (N_1303,N_902,N_1085);
or U1304 (N_1304,In_860,N_978);
nand U1305 (N_1305,N_1066,N_765);
xor U1306 (N_1306,In_2437,In_2064);
nand U1307 (N_1307,In_1136,In_1638);
or U1308 (N_1308,In_2962,N_236);
nand U1309 (N_1309,In_939,N_1082);
nor U1310 (N_1310,N_661,In_1233);
nor U1311 (N_1311,In_346,In_1893);
nand U1312 (N_1312,In_777,In_649);
or U1313 (N_1313,In_1380,In_2963);
or U1314 (N_1314,In_278,N_538);
nor U1315 (N_1315,N_314,In_1232);
or U1316 (N_1316,In_281,In_2163);
nor U1317 (N_1317,N_1097,In_2915);
or U1318 (N_1318,N_126,N_1124);
or U1319 (N_1319,N_997,N_1037);
and U1320 (N_1320,N_264,N_302);
nor U1321 (N_1321,In_1910,In_1423);
and U1322 (N_1322,In_169,In_1283);
nand U1323 (N_1323,N_734,N_697);
or U1324 (N_1324,N_46,In_1698);
xnor U1325 (N_1325,N_915,In_2222);
nor U1326 (N_1326,In_2024,In_869);
or U1327 (N_1327,In_354,In_1641);
nor U1328 (N_1328,N_383,In_1388);
and U1329 (N_1329,In_809,N_1112);
nor U1330 (N_1330,N_804,N_64);
nand U1331 (N_1331,In_930,In_418);
xor U1332 (N_1332,N_1033,In_577);
nand U1333 (N_1333,In_1264,N_405);
and U1334 (N_1334,N_1030,N_1089);
and U1335 (N_1335,N_990,N_885);
nand U1336 (N_1336,In_2169,In_1197);
or U1337 (N_1337,In_1343,In_2215);
or U1338 (N_1338,N_416,In_2691);
or U1339 (N_1339,In_781,N_26);
xnor U1340 (N_1340,N_5,N_962);
or U1341 (N_1341,N_919,In_2403);
and U1342 (N_1342,N_168,In_823);
or U1343 (N_1343,In_2305,N_1125);
nor U1344 (N_1344,N_294,In_2133);
xnor U1345 (N_1345,N_1195,N_431);
and U1346 (N_1346,In_2155,In_761);
and U1347 (N_1347,N_1048,In_1448);
xor U1348 (N_1348,In_1373,In_1142);
nand U1349 (N_1349,In_820,In_329);
or U1350 (N_1350,N_1168,In_992);
nand U1351 (N_1351,In_2959,In_2487);
and U1352 (N_1352,In_1116,In_348);
nand U1353 (N_1353,In_1085,In_705);
and U1354 (N_1354,N_778,N_429);
nand U1355 (N_1355,N_503,In_2311);
nand U1356 (N_1356,N_876,In_255);
and U1357 (N_1357,In_2128,In_1793);
or U1358 (N_1358,N_1086,In_378);
nand U1359 (N_1359,In_65,In_1438);
or U1360 (N_1360,N_1004,In_1944);
nor U1361 (N_1361,In_2519,N_462);
or U1362 (N_1362,N_85,N_679);
xnor U1363 (N_1363,N_730,In_1636);
xor U1364 (N_1364,In_2859,In_351);
nor U1365 (N_1365,N_689,In_1587);
nor U1366 (N_1366,N_434,In_1656);
xor U1367 (N_1367,N_910,N_653);
nor U1368 (N_1368,In_619,In_2456);
nor U1369 (N_1369,In_1159,In_212);
and U1370 (N_1370,In_2254,In_2319);
xnor U1371 (N_1371,In_2445,In_353);
nand U1372 (N_1372,N_588,In_935);
nor U1373 (N_1373,N_598,N_617);
nand U1374 (N_1374,In_1747,N_48);
nor U1375 (N_1375,In_1222,In_2530);
and U1376 (N_1376,In_268,In_2251);
and U1377 (N_1377,In_525,In_1934);
or U1378 (N_1378,N_387,N_920);
nand U1379 (N_1379,In_2070,In_1431);
xor U1380 (N_1380,In_2277,In_24);
or U1381 (N_1381,In_2118,N_918);
or U1382 (N_1382,N_1111,In_6);
xnor U1383 (N_1383,N_295,In_2517);
or U1384 (N_1384,N_1084,In_2846);
nor U1385 (N_1385,In_617,N_695);
nand U1386 (N_1386,N_1107,In_1742);
or U1387 (N_1387,In_221,N_109);
or U1388 (N_1388,N_655,In_1231);
nor U1389 (N_1389,In_2333,In_2314);
xor U1390 (N_1390,In_2027,In_1341);
xnor U1391 (N_1391,In_1984,N_899);
and U1392 (N_1392,In_1078,In_837);
xnor U1393 (N_1393,N_543,In_2296);
and U1394 (N_1394,N_223,N_91);
xnor U1395 (N_1395,In_523,N_873);
and U1396 (N_1396,N_1129,In_584);
and U1397 (N_1397,N_982,In_364);
nand U1398 (N_1398,N_1079,In_1488);
or U1399 (N_1399,In_1750,In_1663);
nand U1400 (N_1400,N_1334,N_672);
or U1401 (N_1401,In_878,In_2946);
xor U1402 (N_1402,N_1251,In_383);
or U1403 (N_1403,N_1344,In_846);
nand U1404 (N_1404,In_2380,N_1184);
nand U1405 (N_1405,In_1486,N_1120);
and U1406 (N_1406,N_977,N_425);
or U1407 (N_1407,In_1693,N_1270);
xnor U1408 (N_1408,In_1437,In_1444);
xor U1409 (N_1409,In_2100,N_408);
or U1410 (N_1410,N_953,N_1370);
or U1411 (N_1411,In_782,N_654);
and U1412 (N_1412,N_1072,In_480);
xnor U1413 (N_1413,N_520,N_306);
or U1414 (N_1414,In_1219,In_973);
xor U1415 (N_1415,N_834,N_931);
nor U1416 (N_1416,N_273,In_1474);
nand U1417 (N_1417,In_2425,N_197);
or U1418 (N_1418,N_1185,N_1256);
and U1419 (N_1419,In_1234,N_644);
nand U1420 (N_1420,N_799,In_2586);
and U1421 (N_1421,N_1024,N_298);
nand U1422 (N_1422,In_1995,N_1153);
and U1423 (N_1423,N_13,N_1174);
nor U1424 (N_1424,In_1079,In_564);
and U1425 (N_1425,N_711,In_292);
and U1426 (N_1426,N_1076,In_307);
and U1427 (N_1427,In_139,In_2384);
xor U1428 (N_1428,N_785,In_2760);
and U1429 (N_1429,N_1252,N_1200);
nand U1430 (N_1430,N_1187,N_1088);
and U1431 (N_1431,N_976,In_1162);
and U1432 (N_1432,N_1134,N_1214);
nor U1433 (N_1433,N_1032,N_1386);
nand U1434 (N_1434,In_2390,N_587);
xor U1435 (N_1435,In_2228,N_892);
xor U1436 (N_1436,In_1086,N_1058);
xor U1437 (N_1437,N_810,In_1074);
nor U1438 (N_1438,N_1141,N_1283);
xor U1439 (N_1439,N_1343,In_1517);
nor U1440 (N_1440,In_1221,In_2721);
nand U1441 (N_1441,N_154,N_984);
xor U1442 (N_1442,N_393,In_1890);
or U1443 (N_1443,N_903,In_1743);
and U1444 (N_1444,In_335,N_1130);
nand U1445 (N_1445,In_1581,In_596);
and U1446 (N_1446,N_595,In_2471);
nor U1447 (N_1447,In_2790,N_1190);
nor U1448 (N_1448,In_510,In_1834);
nand U1449 (N_1449,In_2857,N_651);
or U1450 (N_1450,N_740,N_1063);
nand U1451 (N_1451,In_1800,N_1363);
nor U1452 (N_1452,In_1125,In_31);
xnor U1453 (N_1453,N_1382,N_1249);
nand U1454 (N_1454,In_1993,N_1166);
xnor U1455 (N_1455,N_1068,In_715);
nand U1456 (N_1456,N_1319,In_2370);
xor U1457 (N_1457,In_1815,In_1511);
nand U1458 (N_1458,In_1226,N_204);
xnor U1459 (N_1459,In_82,N_1257);
and U1460 (N_1460,In_1957,In_464);
xnor U1461 (N_1461,In_2605,N_871);
and U1462 (N_1462,In_1839,N_1188);
xnor U1463 (N_1463,In_2269,In_283);
xor U1464 (N_1464,N_1360,N_1350);
nor U1465 (N_1465,N_692,N_1279);
or U1466 (N_1466,In_1202,In_89);
and U1467 (N_1467,In_2545,N_1178);
xnor U1468 (N_1468,In_1121,N_567);
and U1469 (N_1469,In_704,N_1347);
nor U1470 (N_1470,In_2400,N_1241);
or U1471 (N_1471,N_34,N_1057);
nand U1472 (N_1472,In_208,N_1162);
nand U1473 (N_1473,N_4,In_1450);
and U1474 (N_1474,In_1391,N_21);
nor U1475 (N_1475,N_1341,N_1356);
or U1476 (N_1476,In_2461,In_2801);
xor U1477 (N_1477,In_179,In_83);
and U1478 (N_1478,In_2910,In_582);
nor U1479 (N_1479,N_1264,In_1193);
xnor U1480 (N_1480,N_625,In_1175);
nand U1481 (N_1481,N_1181,In_723);
and U1482 (N_1482,N_755,In_2060);
nand U1483 (N_1483,N_909,In_2883);
nor U1484 (N_1484,In_2458,In_737);
or U1485 (N_1485,In_1559,In_779);
nor U1486 (N_1486,In_103,In_2392);
and U1487 (N_1487,In_1847,In_989);
nor U1488 (N_1488,In_791,N_1122);
xnor U1489 (N_1489,In_232,In_845);
and U1490 (N_1490,N_731,In_1374);
or U1491 (N_1491,N_1090,N_1272);
and U1492 (N_1492,In_2444,In_171);
nor U1493 (N_1493,In_1114,In_2484);
xor U1494 (N_1494,N_1211,N_1029);
xor U1495 (N_1495,In_974,N_175);
nor U1496 (N_1496,In_1055,In_2774);
xor U1497 (N_1497,N_863,In_2707);
nor U1498 (N_1498,N_1131,In_2375);
or U1499 (N_1499,In_1734,N_1100);
nand U1500 (N_1500,In_432,In_618);
and U1501 (N_1501,N_1199,N_1300);
or U1502 (N_1502,In_1132,N_620);
and U1503 (N_1503,N_1235,N_1172);
nor U1504 (N_1504,N_209,N_1189);
or U1505 (N_1505,In_1416,In_1065);
nor U1506 (N_1506,N_1315,N_572);
nand U1507 (N_1507,N_803,In_1332);
and U1508 (N_1508,In_1669,N_1075);
nor U1509 (N_1509,N_1308,In_361);
or U1510 (N_1510,N_394,N_1228);
nor U1511 (N_1511,N_285,N_519);
or U1512 (N_1512,In_813,N_1301);
xor U1513 (N_1513,In_2567,In_2450);
xnor U1514 (N_1514,N_831,N_210);
or U1515 (N_1515,N_35,N_1355);
nand U1516 (N_1516,In_1421,In_174);
nor U1517 (N_1517,In_1336,N_813);
xor U1518 (N_1518,N_706,In_1295);
nand U1519 (N_1519,N_373,In_733);
nor U1520 (N_1520,N_545,In_206);
or U1521 (N_1521,In_1420,N_1210);
xor U1522 (N_1522,N_276,In_2575);
xor U1523 (N_1523,In_2001,N_1018);
nor U1524 (N_1524,N_875,N_261);
or U1525 (N_1525,N_1087,N_1302);
nand U1526 (N_1526,N_631,N_1022);
nor U1527 (N_1527,N_152,N_290);
nand U1528 (N_1528,N_1332,N_1265);
nand U1529 (N_1529,N_881,In_524);
and U1530 (N_1530,In_1981,N_1205);
or U1531 (N_1531,N_1002,N_94);
nor U1532 (N_1532,In_2970,In_1539);
xnor U1533 (N_1533,In_1903,In_384);
nor U1534 (N_1534,N_1392,N_1102);
nand U1535 (N_1535,In_2956,In_1201);
or U1536 (N_1536,In_2614,N_150);
nor U1537 (N_1537,N_1261,In_1610);
xnor U1538 (N_1538,N_854,In_1427);
or U1539 (N_1539,In_835,N_346);
nand U1540 (N_1540,In_2287,In_1545);
nor U1541 (N_1541,In_2223,N_693);
or U1542 (N_1542,In_764,In_1459);
nand U1543 (N_1543,In_1950,In_1932);
and U1544 (N_1544,N_449,In_1713);
and U1545 (N_1545,N_888,In_927);
and U1546 (N_1546,N_1375,In_945);
nor U1547 (N_1547,In_437,In_1270);
nand U1548 (N_1548,N_1290,In_756);
nor U1549 (N_1549,N_214,In_2877);
nor U1550 (N_1550,In_1904,In_627);
xnor U1551 (N_1551,In_667,N_979);
nand U1552 (N_1552,N_136,N_808);
or U1553 (N_1553,In_300,N_658);
xnor U1554 (N_1554,In_1292,In_858);
xnor U1555 (N_1555,N_1165,In_695);
or U1556 (N_1556,N_1348,N_614);
nor U1557 (N_1557,N_954,In_1432);
and U1558 (N_1558,N_352,In_519);
nand U1559 (N_1559,N_751,In_2225);
nor U1560 (N_1560,N_106,In_1379);
nor U1561 (N_1561,N_396,In_1690);
and U1562 (N_1562,N_301,In_2255);
nor U1563 (N_1563,In_1818,N_1255);
nor U1564 (N_1564,N_174,In_1996);
nand U1565 (N_1565,In_1642,N_1368);
or U1566 (N_1566,N_1358,In_1817);
nor U1567 (N_1567,N_608,In_815);
or U1568 (N_1568,N_840,N_1008);
and U1569 (N_1569,In_1268,In_1780);
or U1570 (N_1570,In_683,In_2460);
or U1571 (N_1571,N_970,N_707);
and U1572 (N_1572,N_317,In_2061);
nor U1573 (N_1573,In_770,N_1013);
nand U1574 (N_1574,In_1882,In_1407);
or U1575 (N_1575,N_1336,N_829);
nand U1576 (N_1576,In_2343,In_161);
or U1577 (N_1577,N_603,In_2669);
nor U1578 (N_1578,In_2722,N_1110);
nand U1579 (N_1579,In_1732,In_1247);
xnor U1580 (N_1580,In_1916,N_1340);
nor U1581 (N_1581,In_1812,In_1119);
nor U1582 (N_1582,N_1316,In_2637);
and U1583 (N_1583,N_817,In_562);
or U1584 (N_1584,In_345,N_95);
and U1585 (N_1585,In_397,N_1047);
nor U1586 (N_1586,N_395,N_1159);
or U1587 (N_1587,In_926,N_923);
and U1588 (N_1588,In_2173,In_64);
and U1589 (N_1589,In_2362,N_1224);
and U1590 (N_1590,N_673,In_725);
or U1591 (N_1591,N_616,N_581);
and U1592 (N_1592,N_542,N_564);
and U1593 (N_1593,In_2537,In_1906);
and U1594 (N_1594,N_771,N_741);
and U1595 (N_1595,N_1026,In_1716);
nand U1596 (N_1596,N_1396,N_1240);
or U1597 (N_1597,In_1203,In_1544);
xor U1598 (N_1598,N_287,In_2872);
nand U1599 (N_1599,In_2895,In_2401);
or U1600 (N_1600,In_2261,N_1448);
nand U1601 (N_1601,In_2236,N_228);
or U1602 (N_1602,N_1044,In_2717);
and U1603 (N_1603,In_1303,In_595);
or U1604 (N_1604,In_840,N_1327);
nand U1605 (N_1605,N_1197,N_1105);
nor U1606 (N_1606,In_654,N_1591);
nor U1607 (N_1607,N_1142,In_2232);
or U1608 (N_1608,In_2823,In_2457);
xor U1609 (N_1609,N_418,N_1145);
and U1610 (N_1610,N_1492,N_1527);
and U1611 (N_1611,In_1707,In_2162);
or U1612 (N_1612,In_1917,In_2258);
nor U1613 (N_1613,N_998,N_1596);
nand U1614 (N_1614,In_1931,In_1462);
and U1615 (N_1615,N_220,In_1919);
nor U1616 (N_1616,In_2304,In_2708);
or U1617 (N_1617,N_1536,In_320);
nor U1618 (N_1618,N_548,N_1137);
nand U1619 (N_1619,N_883,In_402);
and U1620 (N_1620,N_1427,N_327);
or U1621 (N_1621,N_1038,N_1313);
xor U1622 (N_1622,In_2763,N_1291);
and U1623 (N_1623,N_1411,N_185);
nor U1624 (N_1624,In_1725,N_864);
nand U1625 (N_1625,N_1225,In_1452);
and U1626 (N_1626,N_112,N_782);
nand U1627 (N_1627,N_1160,In_2348);
nor U1628 (N_1628,N_828,In_1760);
nor U1629 (N_1629,In_1460,N_566);
xor U1630 (N_1630,N_1385,N_916);
and U1631 (N_1631,N_1397,In_2595);
nand U1632 (N_1632,In_2428,In_2748);
or U1633 (N_1633,N_597,N_1462);
xnor U1634 (N_1634,N_960,N_1222);
xor U1635 (N_1635,N_447,N_412);
xor U1636 (N_1636,In_825,In_985);
nor U1637 (N_1637,N_818,N_1449);
and U1638 (N_1638,In_113,In_1758);
or U1639 (N_1639,N_985,N_1345);
and U1640 (N_1640,In_1019,N_811);
nor U1641 (N_1641,N_912,N_1060);
nand U1642 (N_1642,In_731,N_1412);
or U1643 (N_1643,In_851,N_911);
and U1644 (N_1644,N_342,N_1213);
nand U1645 (N_1645,N_1234,N_1231);
xor U1646 (N_1646,N_1594,N_927);
nor U1647 (N_1647,N_972,In_2229);
nor U1648 (N_1648,In_2293,N_1278);
nand U1649 (N_1649,In_352,In_1098);
nand U1650 (N_1650,In_2700,N_1439);
nand U1651 (N_1651,In_1285,In_289);
and U1652 (N_1652,In_1058,N_562);
or U1653 (N_1653,N_1410,N_770);
xnor U1654 (N_1654,N_872,In_2239);
or U1655 (N_1655,N_399,N_1542);
nor U1656 (N_1656,In_1505,In_1094);
and U1657 (N_1657,In_2919,N_43);
and U1658 (N_1658,N_703,N_1074);
or U1659 (N_1659,In_1762,N_980);
nand U1660 (N_1660,N_1303,In_669);
nand U1661 (N_1661,In_2391,N_1578);
nor U1662 (N_1662,In_652,In_2942);
xnor U1663 (N_1663,N_1115,N_1333);
nand U1664 (N_1664,N_1266,N_930);
nand U1665 (N_1665,N_1139,In_2653);
or U1666 (N_1666,In_343,N_732);
nand U1667 (N_1667,N_790,In_1915);
and U1668 (N_1668,In_2568,In_2888);
or U1669 (N_1669,N_1500,N_1366);
or U1670 (N_1670,In_209,In_1013);
nor U1671 (N_1671,In_2732,In_1602);
and U1672 (N_1672,N_1236,N_1035);
nand U1673 (N_1673,N_1476,N_1390);
and U1674 (N_1674,N_113,In_541);
or U1675 (N_1675,N_973,N_451);
or U1676 (N_1676,In_1076,In_153);
xnor U1677 (N_1677,N_1369,In_313);
xnor U1678 (N_1678,N_948,N_861);
nand U1679 (N_1679,In_1784,N_1050);
and U1680 (N_1680,In_2199,N_1465);
nand U1681 (N_1681,N_56,N_1560);
and U1682 (N_1682,N_619,N_842);
xnor U1683 (N_1683,In_192,In_2135);
xnor U1684 (N_1684,In_1033,N_1194);
nor U1685 (N_1685,In_2815,N_339);
or U1686 (N_1686,In_1,In_2283);
and U1687 (N_1687,N_1471,N_1293);
and U1688 (N_1688,In_549,N_1157);
nand U1689 (N_1689,N_1114,In_2235);
nor U1690 (N_1690,N_1138,N_601);
and U1691 (N_1691,In_856,N_1400);
nand U1692 (N_1692,N_938,In_1492);
and U1693 (N_1693,N_1258,N_1311);
or U1694 (N_1694,In_1107,N_1508);
nor U1695 (N_1695,N_1324,N_1503);
xor U1696 (N_1696,N_708,In_2280);
and U1697 (N_1697,N_1561,In_1252);
xor U1698 (N_1698,N_1505,N_139);
and U1699 (N_1699,N_1227,N_1454);
and U1700 (N_1700,In_490,In_1914);
xor U1701 (N_1701,N_1096,N_208);
xnor U1702 (N_1702,N_933,In_9);
nand U1703 (N_1703,In_2480,N_93);
and U1704 (N_1704,N_1023,In_2257);
nor U1705 (N_1705,In_99,N_1021);
nand U1706 (N_1706,In_2580,In_1464);
nor U1707 (N_1707,In_712,In_929);
or U1708 (N_1708,N_1401,In_296);
xnor U1709 (N_1709,In_1884,N_1488);
or U1710 (N_1710,N_1472,N_1245);
xnor U1711 (N_1711,N_1028,N_718);
and U1712 (N_1712,N_908,N_1009);
or U1713 (N_1713,N_200,N_897);
xnor U1714 (N_1714,In_450,N_1305);
nand U1715 (N_1715,In_200,N_1532);
nand U1716 (N_1716,N_801,N_1377);
or U1717 (N_1717,N_641,N_1254);
and U1718 (N_1718,In_1717,In_607);
nor U1719 (N_1719,In_2332,In_379);
xnor U1720 (N_1720,In_315,In_824);
xor U1721 (N_1721,N_1475,N_1595);
and U1722 (N_1722,N_1260,N_221);
and U1723 (N_1723,In_802,N_110);
xor U1724 (N_1724,N_1442,In_982);
nor U1725 (N_1725,N_1534,N_1351);
and U1726 (N_1726,N_952,In_711);
and U1727 (N_1727,In_1826,N_1509);
nand U1728 (N_1728,N_256,N_130);
nor U1729 (N_1729,N_1419,N_1513);
nor U1730 (N_1730,In_852,N_750);
nand U1731 (N_1731,N_443,N_1268);
xor U1732 (N_1732,In_374,In_1072);
nand U1733 (N_1733,In_1860,N_1446);
nand U1734 (N_1734,In_947,N_1175);
nand U1735 (N_1735,N_1409,In_1635);
and U1736 (N_1736,N_698,N_964);
nor U1737 (N_1737,N_724,In_1080);
nor U1738 (N_1738,N_1335,N_1597);
nor U1739 (N_1739,N_1512,N_1277);
or U1740 (N_1740,N_1426,N_1323);
or U1741 (N_1741,N_1510,In_1405);
or U1742 (N_1742,In_891,In_1157);
nor U1743 (N_1743,N_1119,In_1767);
or U1744 (N_1744,N_1477,N_1421);
nand U1745 (N_1745,N_1237,In_1777);
nor U1746 (N_1746,In_2032,N_1402);
or U1747 (N_1747,In_433,In_1210);
nor U1748 (N_1748,In_1874,N_928);
and U1749 (N_1749,N_1338,N_1599);
xnor U1750 (N_1750,In_95,In_2613);
and U1751 (N_1751,In_2087,N_1206);
or U1752 (N_1752,N_272,In_2468);
nor U1753 (N_1753,In_1500,In_2932);
xor U1754 (N_1754,In_601,N_424);
or U1755 (N_1755,N_1541,In_2576);
nand U1756 (N_1756,In_54,N_1429);
or U1757 (N_1757,N_1422,N_1081);
and U1758 (N_1758,N_1339,In_2013);
nor U1759 (N_1759,In_2889,In_250);
xor U1760 (N_1760,N_1574,N_1528);
nor U1761 (N_1761,N_326,In_1112);
nor U1762 (N_1762,N_432,In_2544);
and U1763 (N_1763,In_2429,N_1453);
or U1764 (N_1764,N_1109,N_1056);
or U1765 (N_1765,N_345,In_1009);
and U1766 (N_1766,N_800,In_1371);
xnor U1767 (N_1767,In_1397,N_1581);
xnor U1768 (N_1768,In_77,In_1566);
nand U1769 (N_1769,In_162,In_2147);
and U1770 (N_1770,In_1220,N_1295);
nand U1771 (N_1771,N_1383,N_319);
nand U1772 (N_1772,N_390,In_229);
xnor U1773 (N_1773,N_1147,N_463);
nand U1774 (N_1774,N_1073,In_1160);
or U1775 (N_1775,In_1528,N_1221);
xnor U1776 (N_1776,N_1059,N_1151);
and U1777 (N_1777,In_195,N_1365);
xor U1778 (N_1778,N_1118,N_855);
xor U1779 (N_1779,N_1575,In_2207);
xor U1780 (N_1780,N_1250,N_1470);
nand U1781 (N_1781,In_1503,N_853);
nor U1782 (N_1782,N_267,In_931);
or U1783 (N_1783,N_337,N_1036);
xnor U1784 (N_1784,N_134,N_1485);
xor U1785 (N_1785,N_1322,N_33);
and U1786 (N_1786,In_144,In_918);
xnor U1787 (N_1787,In_2792,N_1156);
and U1788 (N_1788,In_2085,In_1898);
xor U1789 (N_1789,N_1098,N_163);
or U1790 (N_1790,N_1573,In_847);
nand U1791 (N_1791,In_2673,In_2999);
and U1792 (N_1792,N_768,N_1522);
nand U1793 (N_1793,N_7,N_1025);
nand U1794 (N_1794,N_1447,N_502);
and U1795 (N_1795,N_1433,In_2813);
and U1796 (N_1796,In_417,N_1275);
nor U1797 (N_1797,N_870,In_48);
nor U1798 (N_1798,N_1526,In_1859);
nor U1799 (N_1799,N_1095,In_1475);
nor U1800 (N_1800,N_1781,In_2272);
or U1801 (N_1801,N_1354,In_2264);
nor U1802 (N_1802,In_198,In_2124);
and U1803 (N_1803,N_1379,N_1588);
nand U1804 (N_1804,In_1362,In_2716);
xor U1805 (N_1805,In_1328,N_1101);
and U1806 (N_1806,In_393,N_1403);
nor U1807 (N_1807,In_2731,N_1668);
xnor U1808 (N_1808,In_1056,N_1603);
and U1809 (N_1809,N_1598,N_745);
nand U1810 (N_1810,In_2121,N_1031);
or U1811 (N_1811,In_211,N_1012);
or U1812 (N_1812,N_1207,N_1220);
or U1813 (N_1813,In_1046,In_2678);
xor U1814 (N_1814,N_704,N_205);
and U1815 (N_1815,N_1661,N_1686);
and U1816 (N_1816,N_1757,In_1805);
or U1817 (N_1817,N_1604,N_767);
and U1818 (N_1818,N_652,In_23);
xor U1819 (N_1819,In_685,N_1762);
or U1820 (N_1820,N_370,In_321);
or U1821 (N_1821,N_1041,In_877);
or U1822 (N_1822,In_331,In_817);
nand U1823 (N_1823,N_1558,N_1337);
or U1824 (N_1824,N_852,N_1705);
and U1825 (N_1825,N_426,N_945);
nor U1826 (N_1826,In_2702,N_1787);
xnor U1827 (N_1827,N_1247,N_366);
nor U1828 (N_1828,N_1299,N_1128);
xor U1829 (N_1829,In_560,N_105);
nand U1830 (N_1830,In_1955,N_1378);
xor U1831 (N_1831,In_489,N_1718);
nand U1832 (N_1832,N_1744,N_1473);
xnor U1833 (N_1833,N_944,N_580);
xnor U1834 (N_1834,In_415,In_295);
and U1835 (N_1835,N_1784,N_677);
nand U1836 (N_1836,N_1380,N_60);
nand U1837 (N_1837,N_1136,In_125);
nand U1838 (N_1838,N_1144,N_1715);
nor U1839 (N_1839,N_1707,In_2878);
and U1840 (N_1840,N_1782,N_694);
and U1841 (N_1841,N_1329,N_251);
or U1842 (N_1842,In_1695,N_659);
xnor U1843 (N_1843,N_1203,N_1215);
xor U1844 (N_1844,N_413,N_1474);
or U1845 (N_1845,In_298,N_835);
or U1846 (N_1846,In_1016,N_1212);
or U1847 (N_1847,N_737,N_1551);
nand U1848 (N_1848,N_635,In_1772);
xnor U1849 (N_1849,N_1629,N_824);
nor U1850 (N_1850,N_1459,In_1070);
or U1851 (N_1851,N_1662,In_80);
nand U1852 (N_1852,N_1698,N_1789);
nand U1853 (N_1853,N_1732,In_408);
nor U1854 (N_1854,N_1589,N_924);
nor U1855 (N_1855,N_1719,N_1294);
xnor U1856 (N_1856,In_279,N_1743);
nand U1857 (N_1857,N_848,In_995);
nand U1858 (N_1858,N_1506,N_1014);
nor U1859 (N_1859,In_1490,N_1367);
or U1860 (N_1860,N_1330,In_46);
and U1861 (N_1861,N_1700,N_1486);
xor U1862 (N_1862,N_1667,In_2049);
and U1863 (N_1863,N_837,In_792);
or U1864 (N_1864,N_1775,N_1774);
nor U1865 (N_1865,In_306,N_1625);
nor U1866 (N_1866,N_16,In_1356);
xor U1867 (N_1867,In_2250,N_1430);
and U1868 (N_1868,N_951,In_2847);
and U1869 (N_1869,In_85,In_344);
nand U1870 (N_1870,N_1113,N_1673);
xnor U1871 (N_1871,N_830,In_893);
nand U1872 (N_1872,N_1617,In_1849);
nor U1873 (N_1873,In_1574,N_1326);
nand U1874 (N_1874,N_1216,N_929);
nor U1875 (N_1875,N_1564,N_1692);
nand U1876 (N_1876,In_946,N_491);
nand U1877 (N_1877,N_1773,In_2402);
xnor U1878 (N_1878,N_845,N_1671);
nor U1879 (N_1879,In_2051,In_684);
xnor U1880 (N_1880,N_1441,N_1434);
nor U1881 (N_1881,N_330,In_98);
xnor U1882 (N_1882,In_1314,N_1218);
or U1883 (N_1883,N_1576,N_1739);
xnor U1884 (N_1884,N_1404,In_2969);
nor U1885 (N_1885,N_1792,In_1024);
xnor U1886 (N_1886,In_1844,N_1543);
nor U1887 (N_1887,In_134,N_1610);
xor U1888 (N_1888,N_1628,In_2861);
nor U1889 (N_1889,N_1763,N_1734);
nand U1890 (N_1890,In_1363,In_2832);
xnor U1891 (N_1891,N_1793,In_1140);
xor U1892 (N_1892,N_1043,N_1683);
or U1893 (N_1893,In_412,N_1417);
xor U1894 (N_1894,N_1711,N_1554);
or U1895 (N_1895,N_1529,In_1647);
or U1896 (N_1896,In_750,N_1582);
nor U1897 (N_1897,In_52,In_1816);
xor U1898 (N_1898,In_2775,N_882);
xnor U1899 (N_1899,N_1777,N_1498);
nand U1900 (N_1900,N_528,N_1478);
and U1901 (N_1901,N_779,N_1583);
xnor U1902 (N_1902,N_1641,In_2624);
or U1903 (N_1903,N_1452,N_605);
and U1904 (N_1904,In_1633,In_2309);
and U1905 (N_1905,In_2284,In_1850);
and U1906 (N_1906,In_425,N_1693);
xnor U1907 (N_1907,N_1399,In_392);
nor U1908 (N_1908,N_1571,In_72);
nor U1909 (N_1909,N_73,In_1467);
nor U1910 (N_1910,N_1103,In_2807);
nor U1911 (N_1911,N_1461,N_1374);
nand U1912 (N_1912,N_1618,N_901);
nand U1913 (N_1913,In_1593,N_1173);
nor U1914 (N_1914,N_1405,N_1443);
nand U1915 (N_1915,N_1394,In_1409);
nand U1916 (N_1916,N_1524,N_1201);
and U1917 (N_1917,N_1229,In_1166);
xnor U1918 (N_1918,N_1209,N_660);
xor U1919 (N_1919,In_36,N_1325);
nand U1920 (N_1920,N_1507,N_1116);
and U1921 (N_1921,N_1450,N_1202);
and U1922 (N_1922,N_1758,N_1494);
nand U1923 (N_1923,N_286,N_1310);
and U1924 (N_1924,In_78,In_120);
and U1925 (N_1925,In_488,In_1129);
nand U1926 (N_1926,In_58,In_605);
or U1927 (N_1927,N_663,N_1540);
and U1928 (N_1928,N_1149,In_2656);
nor U1929 (N_1929,N_777,In_1433);
and U1930 (N_1930,In_514,N_166);
and U1931 (N_1931,In_2937,In_1556);
xnor U1932 (N_1932,In_2198,In_2950);
or U1933 (N_1933,N_1602,N_165);
xnor U1934 (N_1934,N_1687,N_140);
and U1935 (N_1935,N_1353,N_1737);
nor U1936 (N_1936,N_974,N_1183);
or U1937 (N_1937,N_792,In_1455);
nor U1938 (N_1938,In_341,In_1508);
and U1939 (N_1939,In_1650,N_1238);
or U1940 (N_1940,N_293,N_1720);
or U1941 (N_1941,N_656,In_853);
or U1942 (N_1942,N_1463,N_1735);
xor U1943 (N_1943,In_2089,N_1730);
and U1944 (N_1944,N_1694,N_733);
xor U1945 (N_1945,N_1428,N_1062);
nor U1946 (N_1946,In_1293,N_1217);
or U1947 (N_1947,N_1656,N_552);
and U1948 (N_1948,In_2,N_1587);
or U1949 (N_1949,In_1305,N_1164);
or U1950 (N_1950,N_1093,N_1559);
nor U1951 (N_1951,In_1245,In_2739);
nand U1952 (N_1952,N_738,In_1646);
or U1953 (N_1953,N_1163,N_1660);
nor U1954 (N_1954,In_2415,N_624);
xnor U1955 (N_1955,In_2092,N_1549);
and U1956 (N_1956,In_913,N_487);
nor U1957 (N_1957,N_1055,In_916);
xor U1958 (N_1958,N_1232,In_626);
nor U1959 (N_1959,In_873,N_806);
xor U1960 (N_1960,N_862,In_2994);
nand U1961 (N_1961,N_323,N_1755);
xnor U1962 (N_1962,N_1501,N_1645);
or U1963 (N_1963,N_1516,In_1856);
or U1964 (N_1964,N_147,In_1952);
and U1965 (N_1965,In_1139,In_1733);
and U1966 (N_1966,In_2529,In_1924);
or U1967 (N_1967,In_1426,In_1022);
xor U1968 (N_1968,N_1682,N_571);
xnor U1969 (N_1969,N_1752,N_516);
xnor U1970 (N_1970,N_477,N_554);
nor U1971 (N_1971,In_979,N_1553);
nand U1972 (N_1972,N_1121,In_2662);
and U1973 (N_1973,In_2698,In_810);
or U1974 (N_1974,In_2366,N_1714);
and U1975 (N_1975,In_993,N_1727);
nand U1976 (N_1976,N_1630,N_1635);
nand U1977 (N_1977,N_84,N_1709);
and U1978 (N_1978,N_213,In_2533);
xnor U1979 (N_1979,In_1930,N_2);
nor U1980 (N_1980,N_1246,In_2552);
and U1981 (N_1981,In_326,In_456);
xnor U1982 (N_1982,N_505,N_1626);
xor U1983 (N_1983,N_1381,N_789);
nand U1984 (N_1984,N_1767,N_1633);
and U1985 (N_1985,In_1889,In_1124);
nor U1986 (N_1986,In_1701,In_1979);
nand U1987 (N_1987,In_2288,N_1712);
and U1988 (N_1988,N_299,N_1608);
nor U1989 (N_1989,In_2358,N_1489);
nand U1990 (N_1990,N_376,In_2433);
xnor U1991 (N_1991,N_1651,N_1642);
xor U1992 (N_1992,In_1192,In_1846);
or U1993 (N_1993,In_1620,N_1314);
xnor U1994 (N_1994,In_1366,In_2685);
nand U1995 (N_1995,N_1391,In_389);
and U1996 (N_1996,N_766,In_2513);
or U1997 (N_1997,In_580,In_2406);
or U1998 (N_1998,In_431,In_701);
xnor U1999 (N_1999,In_1798,N_558);
nand U2000 (N_2000,N_987,N_1894);
and U2001 (N_2001,In_1639,N_1580);
nand U2002 (N_2002,N_1780,In_1091);
nand U2003 (N_2003,N_1825,N_266);
xor U2004 (N_2004,N_643,N_1796);
xor U2005 (N_2005,N_1824,N_1616);
nor U2006 (N_2006,N_1425,N_1546);
nand U2007 (N_2007,N_1286,In_2749);
xnor U2008 (N_2008,N_1799,In_2414);
or U2009 (N_2009,In_173,N_1912);
and U2010 (N_2010,N_1960,In_2646);
nand U2011 (N_2011,N_1949,N_9);
nand U2012 (N_2012,N_1933,In_1861);
nor U2013 (N_2013,In_349,In_1324);
and U2014 (N_2014,In_677,N_1768);
nor U2015 (N_2015,N_1893,N_600);
and U2016 (N_2016,N_630,N_961);
xnor U2017 (N_2017,N_690,N_994);
nand U2018 (N_2018,N_546,N_1991);
or U2019 (N_2019,N_1808,N_1954);
nand U2020 (N_2020,N_1904,N_1779);
xor U2021 (N_2021,In_778,In_1600);
xnor U2022 (N_2022,N_1511,N_1871);
xor U2023 (N_2023,N_1208,N_1876);
nor U2024 (N_2024,N_1873,In_2105);
xnor U2025 (N_2025,N_1000,In_1310);
xor U2026 (N_2026,N_1071,N_483);
xor U2027 (N_2027,N_1230,In_1154);
nand U2028 (N_2028,N_1849,N_1487);
xor U2029 (N_2029,In_1279,N_1416);
nor U2030 (N_2030,N_1514,N_61);
nor U2031 (N_2031,N_856,N_599);
xnor U2032 (N_2032,N_1898,N_627);
nor U2033 (N_2033,N_1842,N_1148);
and U2034 (N_2034,N_1803,N_1717);
xnor U2035 (N_2035,N_1841,N_1445);
nor U2036 (N_2036,N_1931,N_1655);
xnor U2037 (N_2037,N_1708,In_118);
xor U2038 (N_2038,N_1288,In_1337);
xnor U2039 (N_2039,In_2627,N_1751);
nand U2040 (N_2040,N_207,N_1080);
xor U2041 (N_2041,In_263,N_1943);
or U2042 (N_2042,N_439,N_1847);
nor U2043 (N_2043,In_1830,N_1962);
nor U2044 (N_2044,N_1866,N_1620);
xnor U2045 (N_2045,N_1525,In_2607);
nor U2046 (N_2046,N_1920,In_1354);
nor U2047 (N_2047,N_1814,N_1815);
or U2048 (N_2048,In_574,N_1716);
xnor U2049 (N_2049,N_1568,N_1045);
and U2050 (N_2050,N_1868,N_815);
and U2051 (N_2051,N_20,In_1123);
xnor U2052 (N_2052,In_1751,N_1967);
nand U2053 (N_2053,In_400,N_1827);
nor U2054 (N_2054,N_1051,In_811);
xor U2055 (N_2055,In_504,In_1403);
or U2056 (N_2056,N_1638,N_1304);
and U2057 (N_2057,In_668,N_1233);
nor U2058 (N_2058,In_1396,In_795);
xor U2059 (N_2059,In_1851,N_1674);
or U2060 (N_2060,In_898,In_890);
and U2061 (N_2061,N_1533,N_1654);
or U2062 (N_2062,N_1312,N_847);
xor U2063 (N_2063,N_1468,N_1243);
nand U2064 (N_2064,N_1809,N_1244);
and U2065 (N_2065,N_1538,N_1831);
nor U2066 (N_2066,In_172,N_1986);
xor U2067 (N_2067,N_1863,N_1908);
nand U2068 (N_2068,In_366,N_231);
and U2069 (N_2069,N_438,N_1653);
nor U2070 (N_2070,In_905,N_1794);
and U2071 (N_2071,N_819,N_536);
and U2072 (N_2072,N_1676,N_1359);
and U2073 (N_2073,N_904,N_1481);
or U2074 (N_2074,In_2022,N_328);
or U2075 (N_2075,In_1089,N_1903);
nor U2076 (N_2076,N_1859,N_1483);
or U2077 (N_2077,N_1065,N_1993);
or U2078 (N_2078,N_1890,N_1049);
and U2079 (N_2079,N_1891,N_1451);
nor U2080 (N_2080,N_1519,In_180);
or U2081 (N_2081,N_1948,N_710);
and U2082 (N_2082,N_1435,N_1318);
nor U2083 (N_2083,In_839,N_1566);
or U2084 (N_2084,N_1922,N_1407);
nand U2085 (N_2085,N_1970,N_1609);
and U2086 (N_2086,N_1907,In_1797);
nor U2087 (N_2087,In_1596,N_914);
and U2088 (N_2088,N_1317,N_1945);
nor U2089 (N_2089,N_1460,N_1458);
and U2090 (N_2090,N_1984,N_1259);
nor U2091 (N_2091,N_494,N_1406);
or U2092 (N_2092,N_230,In_2466);
and U2093 (N_2093,N_1444,N_1106);
nor U2094 (N_2094,In_2451,In_1063);
nor U2095 (N_2095,N_1880,N_1248);
and U2096 (N_2096,In_1778,In_1499);
or U2097 (N_2097,N_1703,In_2997);
and U2098 (N_2098,N_1504,N_1627);
and U2099 (N_2099,In_983,In_2870);
and U2100 (N_2100,N_1788,In_569);
nand U2101 (N_2101,In_2171,N_259);
xnor U2102 (N_2102,In_1067,In_895);
xnor U2103 (N_2103,In_1820,In_2879);
nand U2104 (N_2104,N_1665,N_802);
nand U2105 (N_2105,N_1897,In_1150);
xnor U2106 (N_2106,N_1362,In_1714);
and U2107 (N_2107,N_1436,N_440);
xnor U2108 (N_2108,N_1964,N_1756);
or U2109 (N_2109,N_1584,In_1254);
xor U2110 (N_2110,In_131,N_1909);
or U2111 (N_2111,N_1761,N_748);
nor U2112 (N_2112,N_198,N_859);
and U2113 (N_2113,N_1969,N_1550);
xnor U2114 (N_2114,N_1083,In_2048);
or U2115 (N_2115,In_2860,N_717);
and U2116 (N_2116,In_340,In_828);
nor U2117 (N_2117,N_1681,In_282);
or U2118 (N_2118,N_1974,In_2703);
nor U2119 (N_2119,N_1518,N_340);
or U2120 (N_2120,In_2498,N_760);
nand U2121 (N_2121,N_936,In_1764);
and U2122 (N_2122,N_1760,N_1806);
nor U2123 (N_2123,In_1953,In_2896);
nor U2124 (N_2124,N_1611,In_536);
nor U2125 (N_2125,N_1239,In_2990);
or U2126 (N_2126,N_1988,In_1564);
or U2127 (N_2127,In_2088,N_1996);
or U2128 (N_2128,N_1046,N_967);
or U2129 (N_2129,N_959,In_2492);
xor U2130 (N_2130,N_1331,N_1614);
or U2131 (N_2131,N_1223,N_568);
nand U2132 (N_2132,N_1856,In_2532);
nand U2133 (N_2133,N_1778,N_1992);
and U2134 (N_2134,N_1678,In_1329);
nor U2135 (N_2135,N_1192,N_171);
nand U2136 (N_2136,N_1371,In_1573);
nor U2137 (N_2137,In_1037,N_1357);
nor U2138 (N_2138,N_1352,In_222);
and U2139 (N_2139,N_1600,In_2308);
or U2140 (N_2140,In_686,N_1689);
xnor U2141 (N_2141,N_1414,N_1845);
and U2142 (N_2142,N_1586,N_1069);
xnor U2143 (N_2143,N_1005,N_170);
and U2144 (N_2144,N_1177,N_1328);
and U2145 (N_2145,N_1196,N_177);
xnor U2146 (N_2146,N_1830,N_1952);
xor U2147 (N_2147,N_1226,N_791);
xnor U2148 (N_2148,N_1918,N_1606);
xor U2149 (N_2149,N_1819,In_1813);
and U2150 (N_2150,N_19,N_1998);
xor U2151 (N_2151,In_1576,In_1186);
and U2152 (N_2152,N_1469,N_1697);
xor U2153 (N_2153,N_1740,N_1914);
xor U2154 (N_2154,In_1968,N_664);
and U2155 (N_2155,N_1921,In_798);
nand U2156 (N_2156,N_1273,In_1218);
xnor U2157 (N_2157,N_857,N_1710);
and U2158 (N_2158,N_1530,In_116);
or U2159 (N_2159,N_1965,In_126);
xnor U2160 (N_2160,N_1886,N_1895);
nor U2161 (N_2161,N_1285,In_775);
or U2162 (N_2162,N_1143,In_2535);
nor U2163 (N_2163,N_1040,N_716);
and U2164 (N_2164,N_1408,N_1823);
and U2165 (N_2165,N_1813,N_683);
xor U2166 (N_2166,N_1523,N_1946);
and U2167 (N_2167,N_1741,N_1980);
or U2168 (N_2168,N_753,In_757);
or U2169 (N_2169,In_1886,In_1242);
xor U2170 (N_2170,N_1482,N_1818);
or U2171 (N_2171,N_1464,N_1632);
nand U2172 (N_2172,N_156,N_254);
and U2173 (N_2173,N_827,In_765);
nor U2174 (N_2174,N_1099,In_2292);
nor U2175 (N_2175,N_1791,N_1896);
xnor U2176 (N_2176,N_1413,N_1545);
or U2177 (N_2177,In_546,N_1748);
xnor U2178 (N_2178,N_1639,N_211);
nor U2179 (N_2179,N_1702,N_1721);
xor U2180 (N_2180,N_1479,N_1747);
nand U2181 (N_2181,N_1723,N_1963);
and U2182 (N_2182,N_1146,In_2244);
xor U2183 (N_2183,N_1601,In_90);
and U2184 (N_2184,In_2780,N_1930);
or U2185 (N_2185,N_1669,N_1829);
xor U2186 (N_2186,N_1496,N_1132);
nor U2187 (N_2187,In_2190,N_1826);
or U2188 (N_2188,N_1592,N_898);
and U2189 (N_2189,N_1537,N_939);
nand U2190 (N_2190,In_203,N_1696);
nand U2191 (N_2191,In_228,N_1670);
nor U2192 (N_2192,In_1883,N_1605);
nand U2193 (N_2193,N_132,In_1364);
or U2194 (N_2194,N_403,N_17);
nand U2195 (N_2195,N_1423,N_1934);
or U2196 (N_2196,N_1704,N_1389);
nand U2197 (N_2197,N_18,N_1916);
nand U2198 (N_2198,N_894,N_539);
nor U2199 (N_2199,N_504,N_354);
xor U2200 (N_2200,N_2171,In_193);
and U2201 (N_2201,N_1306,N_2122);
nand U2202 (N_2202,N_2082,N_2129);
nor U2203 (N_2203,N_1517,N_515);
and U2204 (N_2204,N_1307,N_1925);
and U2205 (N_2205,N_1877,N_2149);
nor U2206 (N_2206,N_1274,In_1301);
or U2207 (N_2207,In_2408,N_1997);
nor U2208 (N_2208,N_119,N_1800);
xnor U2209 (N_2209,N_2081,N_1499);
nand U2210 (N_2210,In_1002,N_2127);
or U2211 (N_2211,N_1844,In_181);
nand U2212 (N_2212,N_893,N_1664);
nor U2213 (N_2213,N_583,In_2975);
and U2214 (N_2214,N_1875,N_167);
xnor U2215 (N_2215,N_1999,N_1728);
xor U2216 (N_2216,In_1087,N_917);
nand U2217 (N_2217,N_2118,N_946);
nor U2218 (N_2218,N_2160,N_1759);
xnor U2219 (N_2219,N_270,N_1706);
nand U2220 (N_2220,N_2047,N_1861);
xnor U2221 (N_2221,N_1905,N_950);
nand U2222 (N_2222,In_662,In_2154);
and U2223 (N_2223,N_1885,N_1764);
nand U2224 (N_2224,N_2092,N_1919);
nand U2225 (N_2225,N_1746,N_190);
xnor U2226 (N_2226,N_1901,N_1738);
nor U2227 (N_2227,N_646,N_1786);
nor U2228 (N_2228,N_2067,N_1010);
or U2229 (N_2229,N_816,N_1820);
nand U2230 (N_2230,N_1902,N_2005);
xor U2231 (N_2231,In_2789,N_388);
nor U2232 (N_2232,N_2046,In_1069);
xor U2233 (N_2233,In_327,In_2431);
xnor U2234 (N_2234,N_2099,In_997);
xor U2235 (N_2235,N_2153,N_2146);
and U2236 (N_2236,N_2140,N_1619);
and U2237 (N_2237,N_1376,N_2192);
nor U2238 (N_2238,In_442,In_2417);
or U2239 (N_2239,N_2090,N_353);
nand U2240 (N_2240,In_2666,In_1377);
and U2241 (N_2241,N_2057,N_1972);
xor U2242 (N_2242,In_2844,N_1287);
nand U2243 (N_2243,In_1200,In_1660);
or U2244 (N_2244,N_1940,N_1438);
or U2245 (N_2245,N_1562,N_1652);
nor U2246 (N_2246,In_752,N_1607);
nor U2247 (N_2247,N_1643,In_419);
and U2248 (N_2248,In_896,N_374);
nor U2249 (N_2249,In_1512,In_2713);
nand U2250 (N_2250,In_2686,In_1507);
xor U2251 (N_2251,N_2063,N_2107);
nor U2252 (N_2252,N_1042,N_2064);
or U2253 (N_2253,N_1418,N_1015);
nor U2254 (N_2254,N_2143,In_2599);
xnor U2255 (N_2255,N_579,N_1733);
and U2256 (N_2256,In_427,N_1966);
or U2257 (N_2257,In_1769,In_1081);
xor U2258 (N_2258,N_2056,N_1167);
or U2259 (N_2259,N_2075,N_1535);
nor U2260 (N_2260,N_428,In_240);
and U2261 (N_2261,N_714,N_1804);
and U2262 (N_2262,N_510,N_1944);
nor U2263 (N_2263,N_1296,In_1516);
nand U2264 (N_2264,N_441,N_1384);
nand U2265 (N_2265,N_1882,N_90);
nor U2266 (N_2266,N_145,In_1614);
nor U2267 (N_2267,N_1493,N_1958);
xor U2268 (N_2268,N_1219,N_1797);
nand U2269 (N_2269,N_1491,N_1811);
or U2270 (N_2270,N_2022,In_1912);
nor U2271 (N_2271,N_2108,N_1649);
and U2272 (N_2272,In_1099,N_1349);
xnor U2273 (N_2273,N_238,In_724);
or U2274 (N_2274,N_1855,N_1843);
xnor U2275 (N_2275,N_1415,In_215);
xnor U2276 (N_2276,N_647,N_1749);
nor U2277 (N_2277,In_642,In_2623);
nand U2278 (N_2278,N_187,In_2534);
xor U2279 (N_2279,In_2558,N_1297);
xor U2280 (N_2280,N_1729,In_382);
xor U2281 (N_2281,N_2078,N_1292);
or U2282 (N_2282,N_1981,N_1016);
nor U2283 (N_2283,N_1657,N_381);
and U2284 (N_2284,N_2117,N_1978);
nor U2285 (N_2285,In_2035,N_360);
nand U2286 (N_2286,N_2166,N_2130);
xnor U2287 (N_2287,N_1975,N_1020);
and U2288 (N_2288,N_886,N_1253);
nand U2289 (N_2289,In_592,N_1659);
or U2290 (N_2290,N_1457,In_1603);
and U2291 (N_2291,In_274,N_1198);
or U2292 (N_2292,N_1858,N_1440);
nor U2293 (N_2293,N_1857,N_2037);
or U2294 (N_2294,N_1929,N_1713);
and U2295 (N_2295,N_2165,N_2032);
and U2296 (N_2296,N_1913,N_1783);
and U2297 (N_2297,N_517,N_265);
and U2298 (N_2298,In_160,N_1691);
nand U2299 (N_2299,N_667,N_2004);
nand U2300 (N_2300,N_1612,N_1865);
or U2301 (N_2301,N_1801,N_1520);
nand U2302 (N_2302,N_1973,N_1342);
nor U2303 (N_2303,N_1953,In_1406);
nor U2304 (N_2304,N_699,N_925);
nand U2305 (N_2305,In_2295,N_1807);
nor U2306 (N_2306,N_2189,N_2065);
and U2307 (N_2307,N_99,N_1977);
nor U2308 (N_2308,N_1917,In_2675);
or U2309 (N_2309,N_1679,N_879);
nand U2310 (N_2310,N_1182,N_1947);
and U2311 (N_2311,N_1812,N_1393);
or U2312 (N_2312,N_843,In_803);
nand U2313 (N_2313,N_1431,N_2196);
nand U2314 (N_2314,In_1514,N_2158);
xnor U2315 (N_2315,N_1282,In_1250);
and U2316 (N_2316,N_1848,N_743);
nor U2317 (N_2317,In_2043,N_637);
nand U2318 (N_2318,N_1846,In_2777);
nor U2319 (N_2319,N_1565,N_1750);
xor U2320 (N_2320,N_1795,N_2105);
or U2321 (N_2321,N_1502,N_2188);
nand U2322 (N_2322,N_189,In_252);
and U2323 (N_2323,N_1135,In_1308);
or U2324 (N_2324,N_700,N_1490);
and U2325 (N_2325,N_2042,In_1766);
and U2326 (N_2326,N_2058,N_124);
and U2327 (N_2327,N_1017,N_712);
xor U2328 (N_2328,N_2169,N_2168);
nor U2329 (N_2329,N_1906,N_1852);
xor U2330 (N_2330,N_1979,N_1911);
and U2331 (N_2331,In_762,N_472);
nand U2332 (N_2332,N_1613,N_1985);
nand U2333 (N_2333,N_2123,In_1692);
and U2334 (N_2334,N_2002,N_1467);
xor U2335 (N_2335,N_1420,N_2110);
nor U2336 (N_2336,N_895,N_2030);
nor U2337 (N_2337,N_1928,N_1822);
or U2338 (N_2338,N_906,N_2186);
or U2339 (N_2339,N_1544,N_2020);
nand U2340 (N_2340,N_2154,N_2155);
or U2341 (N_2341,N_1910,N_1899);
and U2342 (N_2342,N_1770,N_2128);
nor U2343 (N_2343,In_1678,N_1976);
xor U2344 (N_2344,N_965,N_1878);
nor U2345 (N_2345,N_1364,N_2085);
xor U2346 (N_2346,N_1585,N_2013);
or U2347 (N_2347,In_2812,N_666);
or U2348 (N_2348,N_1888,In_1977);
and U2349 (N_2349,N_1456,N_665);
and U2350 (N_2350,N_2163,In_2475);
nand U2351 (N_2351,In_1983,N_2103);
xor U2352 (N_2352,N_1990,N_1570);
nor U2353 (N_2353,N_1754,N_1280);
nand U2354 (N_2354,In_2886,N_2026);
or U2355 (N_2355,N_1989,N_2170);
nand U2356 (N_2356,N_1593,N_822);
nor U2357 (N_2357,N_812,N_1432);
xnor U2358 (N_2358,N_1834,N_484);
or U2359 (N_2359,In_2230,N_648);
and U2360 (N_2360,N_2080,N_1982);
nor U2361 (N_2361,N_2124,N_2014);
xnor U2362 (N_2362,N_169,N_2157);
nor U2363 (N_2363,N_2071,N_2087);
xnor U2364 (N_2364,In_1261,In_928);
nand U2365 (N_2365,N_1688,In_1551);
nand U2366 (N_2366,N_1176,In_260);
and U2367 (N_2367,In_531,N_1108);
nand U2368 (N_2368,N_887,N_1776);
nand U2369 (N_2369,N_2138,N_2074);
nand U2370 (N_2370,N_949,N_2016);
xnor U2371 (N_2371,N_1881,N_1150);
and U2372 (N_2372,N_2008,N_1590);
or U2373 (N_2373,In_2820,N_2133);
or U2374 (N_2374,In_45,N_1171);
and U2375 (N_2375,N_1959,N_1838);
nand U2376 (N_2376,N_867,N_2001);
or U2377 (N_2377,N_2035,In_826);
or U2378 (N_2378,N_1092,N_2076);
nor U2379 (N_2379,N_1941,N_1169);
or U2380 (N_2380,N_2176,N_2187);
or U2381 (N_2381,N_1950,N_1851);
and U2382 (N_2382,N_1242,N_1701);
and U2383 (N_2383,N_2006,N_1007);
or U2384 (N_2384,N_2197,N_2152);
and U2385 (N_2385,In_467,N_8);
xor U2386 (N_2386,N_1424,N_1398);
xor U2387 (N_2387,N_1388,N_1862);
or U2388 (N_2388,N_2073,N_1772);
nor U2389 (N_2389,N_2164,N_1539);
or U2390 (N_2390,N_1987,N_2019);
nor U2391 (N_2391,In_84,In_2522);
and U2392 (N_2392,N_1321,N_1027);
and U2393 (N_2393,N_2151,N_468);
and U2394 (N_2394,N_2120,N_1810);
nor U2395 (N_2395,N_2173,N_1556);
or U2396 (N_2396,N_1833,N_1785);
xnor U2397 (N_2397,N_1577,N_2034);
and U2398 (N_2398,N_2000,N_2141);
nand U2399 (N_2399,In_739,In_2120);
and U2400 (N_2400,N_2324,N_2094);
nand U2401 (N_2401,N_2237,N_2320);
xnor U2402 (N_2402,N_1658,In_509);
nor U2403 (N_2403,N_1548,N_2131);
and U2404 (N_2404,N_1690,N_2070);
nor U2405 (N_2405,N_1961,N_1725);
xor U2406 (N_2406,N_1790,N_2308);
or U2407 (N_2407,N_2280,In_15);
xnor U2408 (N_2408,N_2338,N_2093);
xor U2409 (N_2409,N_2359,N_2397);
xor U2410 (N_2410,N_2248,N_415);
or U2411 (N_2411,N_2319,N_2274);
nor U2412 (N_2412,In_1632,N_2309);
nor U2413 (N_2413,N_2242,In_1575);
nand U2414 (N_2414,In_2139,N_448);
xor U2415 (N_2415,N_2373,In_2016);
and U2416 (N_2416,N_2353,N_2114);
nand U2417 (N_2417,In_470,In_50);
and U2418 (N_2418,N_2253,In_678);
xor U2419 (N_2419,N_2315,In_969);
xnor U2420 (N_2420,N_2207,N_2177);
nor U2421 (N_2421,N_2256,N_1935);
and U2422 (N_2422,N_2021,N_2159);
xnor U2423 (N_2423,N_2181,N_2335);
xor U2424 (N_2424,N_2111,In_659);
xor U2425 (N_2425,N_2246,N_1872);
and U2426 (N_2426,N_2330,In_1876);
and U2427 (N_2427,In_1540,N_1860);
nand U2428 (N_2428,N_1995,N_1769);
and U2429 (N_2429,N_2224,N_1923);
xnor U2430 (N_2430,N_2003,N_2331);
xor U2431 (N_2431,In_1858,N_2368);
nand U2432 (N_2432,N_1736,N_2293);
or U2433 (N_2433,N_2066,In_1923);
nand U2434 (N_2434,N_2091,N_2378);
xor U2435 (N_2435,N_1624,N_1869);
nor U2436 (N_2436,N_1724,N_2316);
nand U2437 (N_2437,N_823,In_1185);
nor U2438 (N_2438,N_2211,N_1001);
and U2439 (N_2439,In_365,N_2268);
or U2440 (N_2440,N_2348,N_1936);
nor U2441 (N_2441,N_2312,N_2282);
and U2442 (N_2442,N_2184,N_2244);
and U2443 (N_2443,N_2250,N_2264);
xnor U2444 (N_2444,N_2277,N_2134);
xor U2445 (N_2445,N_2347,N_2278);
and U2446 (N_2446,N_2364,N_2251);
xor U2447 (N_2447,N_1555,N_1091);
or U2448 (N_2448,N_2015,N_1850);
or U2449 (N_2449,N_421,N_2018);
nand U2450 (N_2450,N_1640,In_1052);
xor U2451 (N_2451,N_2208,In_3);
and U2452 (N_2452,N_2052,N_1837);
nand U2453 (N_2453,N_2300,In_117);
xnor U2454 (N_2454,N_1765,N_1547);
nand U2455 (N_2455,N_2322,N_2394);
xnor U2456 (N_2456,N_2135,N_2298);
xnor U2457 (N_2457,N_2150,N_2027);
nor U2458 (N_2458,N_2213,In_2186);
or U2459 (N_2459,N_1892,N_2255);
xnor U2460 (N_2460,N_2317,N_1887);
xor U2461 (N_2461,N_2132,N_2191);
nor U2462 (N_2462,N_678,N_2262);
or U2463 (N_2463,In_1479,In_59);
and U2464 (N_2464,N_1263,N_1276);
and U2465 (N_2465,In_2572,In_1173);
and U2466 (N_2466,In_2067,N_1117);
nand U2467 (N_2467,N_2381,In_2841);
or U2468 (N_2468,N_2229,N_1684);
and U2469 (N_2469,N_1070,N_2265);
and U2470 (N_2470,N_2043,In_499);
nand U2471 (N_2471,N_2367,N_2147);
xor U2472 (N_2472,In_2443,N_1480);
or U2473 (N_2473,N_2356,N_2334);
xnor U2474 (N_2474,N_2222,N_1951);
xnor U2475 (N_2475,N_2179,N_2206);
or U2476 (N_2476,N_832,N_2339);
or U2477 (N_2477,N_2097,N_2398);
xor U2478 (N_2478,N_2238,N_2031);
nor U2479 (N_2479,N_992,N_2346);
and U2480 (N_2480,N_2311,N_1938);
and U2481 (N_2481,N_1271,N_1284);
or U2482 (N_2482,N_968,N_1663);
or U2483 (N_2483,N_2217,In_1209);
xor U2484 (N_2484,N_2365,N_1521);
nor U2485 (N_2485,N_2011,N_2290);
or U2486 (N_2486,In_2398,N_2272);
nand U2487 (N_2487,N_1968,N_2261);
nand U2488 (N_2488,N_2012,N_2288);
xnor U2489 (N_2489,N_1955,N_1373);
and U2490 (N_2490,N_2360,N_1497);
nand U2491 (N_2491,N_2198,N_1883);
nand U2492 (N_2492,In_558,N_2307);
nand U2493 (N_2493,N_2025,N_2040);
xnor U2494 (N_2494,N_1816,N_2369);
or U2495 (N_2495,N_2327,N_2104);
or U2496 (N_2496,N_2193,N_305);
or U2497 (N_2497,N_2247,N_2390);
and U2498 (N_2498,N_2286,N_2024);
nor U2499 (N_2499,N_1864,N_1204);
nand U2500 (N_2500,N_2287,N_2321);
xor U2501 (N_2501,N_2361,N_1853);
and U2502 (N_2502,N_2194,N_2098);
nand U2503 (N_2503,N_2266,N_2382);
and U2504 (N_2504,N_2343,N_1805);
nand U2505 (N_2505,N_1621,N_1884);
xor U2506 (N_2506,N_1623,N_1937);
nand U2507 (N_2507,N_1484,N_389);
nand U2508 (N_2508,N_2054,In_92);
or U2509 (N_2509,N_1154,N_2337);
or U2510 (N_2510,N_2041,N_1646);
or U2511 (N_2511,N_1870,N_662);
or U2512 (N_2512,N_243,N_1821);
nor U2513 (N_2513,In_2493,N_2345);
and U2514 (N_2514,N_1320,N_1854);
nand U2515 (N_2515,N_2017,In_2123);
xnor U2516 (N_2516,N_1766,N_2121);
xor U2517 (N_2517,N_2119,In_1084);
nor U2518 (N_2518,N_1179,N_2212);
nand U2519 (N_2519,N_2178,N_2254);
nand U2520 (N_2520,In_109,N_2236);
or U2521 (N_2521,N_2045,N_2281);
and U2522 (N_2522,In_237,N_2396);
and U2523 (N_2523,N_2295,In_199);
or U2524 (N_2524,In_1325,N_2318);
nor U2525 (N_2525,N_1699,N_2372);
nor U2526 (N_2526,N_2350,In_312);
nand U2527 (N_2527,In_2989,N_2175);
nor U2528 (N_2528,N_1631,N_2084);
and U2529 (N_2529,N_1572,N_31);
xor U2530 (N_2530,N_1563,N_2285);
and U2531 (N_2531,In_259,In_1287);
nor U2532 (N_2532,N_769,N_2358);
nand U2533 (N_2533,N_1636,N_2328);
or U2534 (N_2534,N_2245,N_2340);
or U2535 (N_2535,N_2276,N_2028);
or U2536 (N_2536,N_2374,N_2326);
and U2537 (N_2537,N_2039,In_2536);
nor U2538 (N_2538,N_1926,In_2111);
or U2539 (N_2539,N_2297,N_2383);
xor U2540 (N_2540,N_2259,N_2332);
xnor U2541 (N_2541,N_999,In_545);
and U2542 (N_2542,N_701,N_1971);
nor U2543 (N_2543,N_2271,N_1515);
and U2544 (N_2544,In_483,In_2008);
xnor U2545 (N_2545,N_1019,N_102);
and U2546 (N_2546,N_2239,N_2226);
xor U2547 (N_2547,N_2235,N_2180);
nand U2548 (N_2548,In_655,N_1455);
nor U2549 (N_2549,N_2200,N_1648);
nor U2550 (N_2550,N_1053,N_2007);
and U2551 (N_2551,N_2392,N_2139);
nor U2552 (N_2552,N_1879,N_2258);
or U2553 (N_2553,N_362,N_1186);
and U2554 (N_2554,N_2341,N_1078);
nand U2555 (N_2555,N_2391,N_1695);
or U2556 (N_2556,In_2122,N_2162);
or U2557 (N_2557,N_2257,N_2233);
xnor U2558 (N_2558,N_531,N_1835);
nor U2559 (N_2559,N_1281,In_1637);
nor U2560 (N_2560,N_1900,N_2029);
nor U2561 (N_2561,N_2303,N_1077);
nor U2562 (N_2562,N_2049,N_2095);
and U2563 (N_2563,N_2215,N_2363);
and U2564 (N_2564,N_2314,N_2137);
xnor U2565 (N_2565,N_2249,N_2112);
and U2566 (N_2566,N_1395,In_865);
or U2567 (N_2567,In_2929,N_2174);
and U2568 (N_2568,N_1828,N_2161);
and U2569 (N_2569,N_2227,N_2267);
nand U2570 (N_2570,N_1745,N_2379);
nor U2571 (N_2571,N_52,N_1094);
and U2572 (N_2572,In_776,N_1983);
and U2573 (N_2573,N_2296,In_801);
xor U2574 (N_2574,N_1753,In_414);
and U2575 (N_2575,N_2223,N_2106);
xnor U2576 (N_2576,N_1637,N_2096);
or U2577 (N_2577,N_1567,N_2089);
nor U2578 (N_2578,N_1771,In_2834);
nand U2579 (N_2579,In_1378,N_2385);
nor U2580 (N_2580,N_2355,N_612);
nand U2581 (N_2581,N_2216,N_1726);
nand U2582 (N_2582,N_1650,N_2010);
nand U2583 (N_2583,N_1839,N_2323);
and U2584 (N_2584,N_2386,N_2172);
or U2585 (N_2585,N_2275,N_2384);
and U2586 (N_2586,In_2918,N_1193);
xnor U2587 (N_2587,N_2228,N_2023);
nor U2588 (N_2588,N_2061,N_2086);
or U2589 (N_2589,N_2260,N_2305);
nand U2590 (N_2590,N_2395,In_1294);
nand U2591 (N_2591,N_1915,N_2209);
or U2592 (N_2592,N_2375,N_2393);
or U2593 (N_2593,In_2347,N_640);
or U2594 (N_2594,In_1537,N_2126);
or U2595 (N_2595,N_1957,N_1289);
or U2596 (N_2596,N_2232,N_2352);
or U2597 (N_2597,N_1677,N_2148);
nor U2598 (N_2598,N_2389,N_1832);
xor U2599 (N_2599,N_2357,N_2231);
xor U2600 (N_2600,N_2518,N_2511);
and U2601 (N_2601,N_2273,N_2473);
xor U2602 (N_2602,N_2493,N_2060);
and U2603 (N_2603,N_2575,N_2451);
xor U2604 (N_2604,N_2519,N_2490);
and U2605 (N_2605,N_2144,N_2513);
and U2606 (N_2606,N_2547,N_2520);
nor U2607 (N_2607,N_2533,N_2136);
nor U2608 (N_2608,In_204,N_2366);
and U2609 (N_2609,N_1495,N_2221);
and U2610 (N_2610,N_2289,In_1719);
and U2611 (N_2611,N_2294,N_2342);
xor U2612 (N_2612,N_2036,N_2203);
xnor U2613 (N_2613,N_2292,N_2304);
nand U2614 (N_2614,N_1742,N_2582);
xor U2615 (N_2615,N_2469,N_2439);
nor U2616 (N_2616,N_2263,In_1535);
or U2617 (N_2617,N_2464,N_2500);
nand U2618 (N_2618,N_1531,N_2474);
nor U2619 (N_2619,N_2413,N_2580);
and U2620 (N_2620,N_2313,N_2387);
nand U2621 (N_2621,N_2291,N_2587);
and U2622 (N_2622,N_1052,In_806);
nand U2623 (N_2623,N_2408,N_1932);
and U2624 (N_2624,N_1133,In_1649);
or U2625 (N_2625,N_877,N_2479);
nand U2626 (N_2626,N_2492,N_2512);
nor U2627 (N_2627,In_2090,N_796);
and U2628 (N_2628,N_1672,N_2578);
and U2629 (N_2629,N_1569,N_2156);
or U2630 (N_2630,N_1309,N_1262);
or U2631 (N_2631,In_1353,N_1647);
or U2632 (N_2632,N_2594,N_1924);
xnor U2633 (N_2633,N_2584,N_1956);
nand U2634 (N_2634,N_2586,N_844);
xor U2635 (N_2635,N_2301,In_2145);
or U2636 (N_2636,N_2471,N_2557);
nand U2637 (N_2637,N_2426,N_2489);
nor U2638 (N_2638,N_2424,N_2284);
or U2639 (N_2639,In_10,N_880);
nand U2640 (N_2640,N_2545,N_1387);
and U2641 (N_2641,N_2475,N_891);
nor U2642 (N_2642,N_2195,N_1269);
xor U2643 (N_2643,N_2351,N_2581);
or U2644 (N_2644,In_314,N_2544);
and U2645 (N_2645,N_2420,N_2048);
or U2646 (N_2646,N_2399,In_2265);
nor U2647 (N_2647,N_2409,N_2199);
nand U2648 (N_2648,N_2333,N_2531);
nor U2649 (N_2649,N_1127,N_2401);
nand U2650 (N_2650,N_986,N_2218);
xnor U2651 (N_2651,N_2062,N_2411);
or U2652 (N_2652,N_1361,N_2537);
and U2653 (N_2653,N_2536,N_2243);
nor U2654 (N_2654,N_2507,N_2491);
and U2655 (N_2655,N_618,N_2525);
nor U2656 (N_2656,N_2468,N_2552);
or U2657 (N_2657,N_2567,N_2461);
and U2658 (N_2658,N_2302,N_2463);
and U2659 (N_2659,N_2418,In_972);
nand U2660 (N_2660,N_2433,N_2402);
and U2661 (N_2661,N_2053,N_2466);
or U2662 (N_2662,N_2457,N_2038);
or U2663 (N_2663,N_2502,In_2478);
or U2664 (N_2664,N_2412,In_2520);
nor U2665 (N_2665,N_2102,N_2495);
xnor U2666 (N_2666,N_2577,N_2240);
or U2667 (N_2667,N_2079,N_2458);
nand U2668 (N_2668,N_2444,N_2508);
nor U2669 (N_2669,N_2100,N_2428);
and U2670 (N_2670,N_2561,N_2182);
or U2671 (N_2671,N_2516,In_1010);
and U2672 (N_2672,N_2183,N_2450);
or U2673 (N_2673,In_1711,N_2551);
nand U2674 (N_2674,N_1927,N_2535);
nor U2675 (N_2675,In_911,N_2325);
and U2676 (N_2676,N_2569,N_851);
and U2677 (N_2677,N_2050,In_735);
and U2678 (N_2678,N_2515,N_1267);
nor U2679 (N_2679,N_369,N_2344);
nor U2680 (N_2680,N_2540,N_940);
and U2681 (N_2681,N_2509,N_2310);
nor U2682 (N_2682,N_2599,N_2438);
or U2683 (N_2683,N_2455,N_1666);
or U2684 (N_2684,N_2480,N_2055);
and U2685 (N_2685,N_1466,N_2269);
xnor U2686 (N_2686,N_2534,N_1722);
nor U2687 (N_2687,N_2579,In_2772);
and U2688 (N_2688,N_2219,N_2230);
nand U2689 (N_2689,N_2592,N_2478);
nand U2690 (N_2690,N_2205,N_2470);
nand U2691 (N_2691,N_2432,N_2554);
xnor U2692 (N_2692,N_2564,N_2101);
nor U2693 (N_2693,N_2538,In_2057);
nand U2694 (N_2694,N_2596,N_1067);
and U2695 (N_2695,N_2483,N_2069);
or U2696 (N_2696,N_2530,N_2306);
nor U2697 (N_2697,N_1372,N_2068);
or U2698 (N_2698,N_1346,N_2454);
nand U2699 (N_2699,N_2528,N_2431);
nor U2700 (N_2700,N_2499,N_2279);
and U2701 (N_2701,In_1819,N_2403);
nor U2702 (N_2702,N_2459,N_2562);
nand U2703 (N_2703,N_2430,N_2484);
or U2704 (N_2704,N_2407,N_2145);
and U2705 (N_2705,N_2427,N_2494);
or U2706 (N_2706,N_2595,N_1802);
nor U2707 (N_2707,N_2472,N_2546);
and U2708 (N_2708,N_2568,N_2498);
nor U2709 (N_2709,N_2589,N_2497);
xor U2710 (N_2710,N_2446,N_2416);
nand U2711 (N_2711,N_1994,N_2113);
xor U2712 (N_2712,N_2548,N_2588);
or U2713 (N_2713,N_488,N_2510);
nor U2714 (N_2714,N_759,N_2434);
nor U2715 (N_2715,N_2425,N_1675);
nor U2716 (N_2716,N_2414,N_1622);
nor U2717 (N_2717,N_2436,N_2467);
nand U2718 (N_2718,N_2116,In_2980);
or U2719 (N_2719,N_2524,N_2190);
and U2720 (N_2720,N_2443,N_2329);
or U2721 (N_2721,N_2437,N_2210);
nand U2722 (N_2722,N_2558,N_1685);
nor U2723 (N_2723,N_2563,N_2591);
xnor U2724 (N_2724,N_1874,N_2142);
or U2725 (N_2725,In_1236,N_2541);
nor U2726 (N_2726,N_2435,N_2241);
nor U2727 (N_2727,N_2550,N_2593);
xnor U2728 (N_2728,N_2456,N_2448);
xor U2729 (N_2729,N_2072,In_2655);
nand U2730 (N_2730,N_2532,N_2503);
nand U2731 (N_2731,N_2370,N_1634);
and U2732 (N_2732,N_2477,N_2585);
and U2733 (N_2733,N_1615,N_2522);
or U2734 (N_2734,N_2501,N_2009);
nor U2735 (N_2735,N_2201,N_2299);
xnor U2736 (N_2736,N_2204,N_2573);
and U2737 (N_2737,N_2421,In_1599);
and U2738 (N_2738,In_2328,N_2380);
nand U2739 (N_2739,N_423,In_293);
nand U2740 (N_2740,N_2252,N_2440);
nand U2741 (N_2741,N_2044,N_2417);
nand U2742 (N_2742,N_2583,N_2559);
and U2743 (N_2743,N_2571,N_2423);
nand U2744 (N_2744,N_2542,N_2590);
nand U2745 (N_2745,N_2543,N_2234);
nor U2746 (N_2746,N_836,N_2400);
nand U2747 (N_2747,N_1552,N_2539);
and U2748 (N_2748,N_1437,N_2462);
and U2749 (N_2749,N_2376,N_2476);
nor U2750 (N_2750,N_2460,N_1867);
nor U2751 (N_2751,N_2496,N_2505);
nor U2752 (N_2752,N_2371,N_2033);
xor U2753 (N_2753,In_2161,N_2574);
xnor U2754 (N_2754,N_966,N_2449);
nand U2755 (N_2755,N_2517,N_1298);
nor U2756 (N_2756,N_2565,N_1836);
xnor U2757 (N_2757,N_2485,N_2214);
xor U2758 (N_2758,N_2405,N_2506);
nor U2759 (N_2759,N_2465,N_1680);
nor U2760 (N_2760,N_2526,N_2225);
nor U2761 (N_2761,N_2125,N_2442);
nand U2762 (N_2762,N_2487,N_2453);
or U2763 (N_2763,N_2598,N_2441);
or U2764 (N_2764,N_1644,N_1579);
or U2765 (N_2765,N_2597,N_2422);
and U2766 (N_2766,In_2947,N_2521);
or U2767 (N_2767,N_2452,N_2202);
nor U2768 (N_2768,N_2336,N_2077);
or U2769 (N_2769,N_2404,N_781);
or U2770 (N_2770,N_2566,N_2576);
and U2771 (N_2771,N_2482,N_2283);
nand U2772 (N_2772,N_2354,N_2059);
or U2773 (N_2773,N_2109,N_2549);
nor U2774 (N_2774,N_2167,N_2419);
nand U2775 (N_2775,N_2115,N_1817);
nand U2776 (N_2776,N_2445,N_465);
or U2777 (N_2777,N_2051,N_2088);
nor U2778 (N_2778,N_2377,N_2488);
xnor U2779 (N_2779,N_1798,N_2570);
nor U2780 (N_2780,N_2429,N_2220);
nand U2781 (N_2781,N_1939,N_1889);
nand U2782 (N_2782,N_2362,N_2553);
nand U2783 (N_2783,N_2556,N_807);
xnor U2784 (N_2784,N_1104,N_2560);
or U2785 (N_2785,N_2529,N_2527);
nand U2786 (N_2786,N_2523,N_2185);
nand U2787 (N_2787,N_2083,N_2486);
and U2788 (N_2788,N_2481,N_1003);
and U2789 (N_2789,N_2270,N_1557);
and U2790 (N_2790,In_632,N_2388);
nand U2791 (N_2791,N_2415,N_2410);
and U2792 (N_2792,N_1942,N_2349);
or U2793 (N_2793,In_1684,N_2572);
nor U2794 (N_2794,N_1731,N_2447);
xor U2795 (N_2795,In_1651,N_2514);
nand U2796 (N_2796,N_2504,N_108);
and U2797 (N_2797,In_1212,In_8);
xnor U2798 (N_2798,N_1840,N_2555);
and U2799 (N_2799,N_2406,N_143);
nand U2800 (N_2800,N_2703,N_2789);
and U2801 (N_2801,N_2690,N_2606);
nand U2802 (N_2802,N_2769,N_2711);
nor U2803 (N_2803,N_2615,N_2735);
nor U2804 (N_2804,N_2607,N_2748);
and U2805 (N_2805,N_2698,N_2635);
or U2806 (N_2806,N_2609,N_2772);
or U2807 (N_2807,N_2693,N_2740);
or U2808 (N_2808,N_2654,N_2670);
or U2809 (N_2809,N_2619,N_2684);
or U2810 (N_2810,N_2734,N_2617);
nand U2811 (N_2811,N_2702,N_2603);
xor U2812 (N_2812,N_2645,N_2666);
nand U2813 (N_2813,N_2750,N_2785);
nand U2814 (N_2814,N_2637,N_2731);
or U2815 (N_2815,N_2792,N_2732);
nand U2816 (N_2816,N_2741,N_2714);
xor U2817 (N_2817,N_2691,N_2697);
nand U2818 (N_2818,N_2737,N_2701);
and U2819 (N_2819,N_2745,N_2794);
or U2820 (N_2820,N_2762,N_2608);
or U2821 (N_2821,N_2664,N_2708);
nand U2822 (N_2822,N_2719,N_2689);
xnor U2823 (N_2823,N_2612,N_2793);
xor U2824 (N_2824,N_2626,N_2660);
nand U2825 (N_2825,N_2787,N_2685);
nand U2826 (N_2826,N_2622,N_2754);
xor U2827 (N_2827,N_2797,N_2720);
nand U2828 (N_2828,N_2791,N_2677);
and U2829 (N_2829,N_2669,N_2623);
and U2830 (N_2830,N_2651,N_2705);
nand U2831 (N_2831,N_2774,N_2781);
xor U2832 (N_2832,N_2766,N_2646);
and U2833 (N_2833,N_2667,N_2620);
nand U2834 (N_2834,N_2674,N_2710);
or U2835 (N_2835,N_2699,N_2728);
nand U2836 (N_2836,N_2724,N_2632);
and U2837 (N_2837,N_2770,N_2717);
and U2838 (N_2838,N_2638,N_2752);
nor U2839 (N_2839,N_2618,N_2768);
nor U2840 (N_2840,N_2780,N_2727);
xnor U2841 (N_2841,N_2647,N_2747);
or U2842 (N_2842,N_2629,N_2678);
nor U2843 (N_2843,N_2663,N_2650);
xor U2844 (N_2844,N_2653,N_2763);
and U2845 (N_2845,N_2640,N_2739);
nand U2846 (N_2846,N_2634,N_2605);
nand U2847 (N_2847,N_2729,N_2744);
or U2848 (N_2848,N_2743,N_2649);
nor U2849 (N_2849,N_2773,N_2671);
nor U2850 (N_2850,N_2628,N_2659);
xnor U2851 (N_2851,N_2662,N_2784);
nor U2852 (N_2852,N_2798,N_2604);
or U2853 (N_2853,N_2633,N_2786);
nand U2854 (N_2854,N_2704,N_2709);
xnor U2855 (N_2855,N_2627,N_2776);
xor U2856 (N_2856,N_2624,N_2679);
and U2857 (N_2857,N_2656,N_2713);
nor U2858 (N_2858,N_2601,N_2742);
xnor U2859 (N_2859,N_2783,N_2707);
xor U2860 (N_2860,N_2652,N_2673);
nor U2861 (N_2861,N_2777,N_2755);
and U2862 (N_2862,N_2648,N_2665);
and U2863 (N_2863,N_2778,N_2782);
nand U2864 (N_2864,N_2779,N_2644);
and U2865 (N_2865,N_2641,N_2700);
nand U2866 (N_2866,N_2759,N_2643);
or U2867 (N_2867,N_2733,N_2799);
and U2868 (N_2868,N_2716,N_2655);
or U2869 (N_2869,N_2736,N_2625);
and U2870 (N_2870,N_2753,N_2682);
nand U2871 (N_2871,N_2694,N_2757);
nor U2872 (N_2872,N_2611,N_2630);
and U2873 (N_2873,N_2761,N_2692);
or U2874 (N_2874,N_2760,N_2738);
xor U2875 (N_2875,N_2765,N_2746);
nand U2876 (N_2876,N_2613,N_2642);
xnor U2877 (N_2877,N_2658,N_2614);
xnor U2878 (N_2878,N_2657,N_2771);
nand U2879 (N_2879,N_2764,N_2621);
nor U2880 (N_2880,N_2730,N_2796);
nor U2881 (N_2881,N_2706,N_2726);
or U2882 (N_2882,N_2775,N_2672);
and U2883 (N_2883,N_2767,N_2668);
and U2884 (N_2884,N_2758,N_2602);
nand U2885 (N_2885,N_2790,N_2751);
nor U2886 (N_2886,N_2610,N_2695);
or U2887 (N_2887,N_2749,N_2676);
or U2888 (N_2888,N_2681,N_2723);
nor U2889 (N_2889,N_2639,N_2718);
and U2890 (N_2890,N_2756,N_2683);
nand U2891 (N_2891,N_2688,N_2616);
nor U2892 (N_2892,N_2636,N_2680);
xnor U2893 (N_2893,N_2675,N_2686);
and U2894 (N_2894,N_2600,N_2687);
nor U2895 (N_2895,N_2795,N_2715);
xnor U2896 (N_2896,N_2788,N_2721);
or U2897 (N_2897,N_2725,N_2696);
xnor U2898 (N_2898,N_2712,N_2722);
and U2899 (N_2899,N_2661,N_2631);
and U2900 (N_2900,N_2712,N_2717);
nor U2901 (N_2901,N_2638,N_2758);
and U2902 (N_2902,N_2780,N_2732);
nand U2903 (N_2903,N_2736,N_2689);
nor U2904 (N_2904,N_2709,N_2635);
or U2905 (N_2905,N_2646,N_2685);
and U2906 (N_2906,N_2789,N_2602);
or U2907 (N_2907,N_2768,N_2780);
or U2908 (N_2908,N_2662,N_2701);
xor U2909 (N_2909,N_2621,N_2627);
nand U2910 (N_2910,N_2731,N_2724);
xor U2911 (N_2911,N_2712,N_2638);
or U2912 (N_2912,N_2767,N_2789);
or U2913 (N_2913,N_2705,N_2634);
nand U2914 (N_2914,N_2750,N_2790);
nand U2915 (N_2915,N_2621,N_2607);
and U2916 (N_2916,N_2628,N_2776);
and U2917 (N_2917,N_2694,N_2725);
or U2918 (N_2918,N_2689,N_2741);
nand U2919 (N_2919,N_2741,N_2729);
or U2920 (N_2920,N_2789,N_2628);
xnor U2921 (N_2921,N_2652,N_2789);
nor U2922 (N_2922,N_2605,N_2639);
or U2923 (N_2923,N_2777,N_2641);
and U2924 (N_2924,N_2633,N_2611);
or U2925 (N_2925,N_2668,N_2663);
and U2926 (N_2926,N_2775,N_2667);
nor U2927 (N_2927,N_2685,N_2698);
and U2928 (N_2928,N_2676,N_2721);
nand U2929 (N_2929,N_2767,N_2701);
nor U2930 (N_2930,N_2769,N_2641);
nand U2931 (N_2931,N_2786,N_2642);
or U2932 (N_2932,N_2774,N_2777);
nand U2933 (N_2933,N_2731,N_2783);
nor U2934 (N_2934,N_2745,N_2702);
and U2935 (N_2935,N_2797,N_2765);
xnor U2936 (N_2936,N_2765,N_2789);
nand U2937 (N_2937,N_2685,N_2740);
xnor U2938 (N_2938,N_2628,N_2752);
nand U2939 (N_2939,N_2661,N_2710);
and U2940 (N_2940,N_2648,N_2779);
and U2941 (N_2941,N_2685,N_2619);
xnor U2942 (N_2942,N_2798,N_2600);
nor U2943 (N_2943,N_2684,N_2643);
or U2944 (N_2944,N_2619,N_2707);
nor U2945 (N_2945,N_2760,N_2727);
nor U2946 (N_2946,N_2701,N_2707);
xor U2947 (N_2947,N_2601,N_2785);
xor U2948 (N_2948,N_2696,N_2657);
nor U2949 (N_2949,N_2768,N_2737);
xor U2950 (N_2950,N_2640,N_2782);
or U2951 (N_2951,N_2634,N_2767);
and U2952 (N_2952,N_2712,N_2744);
or U2953 (N_2953,N_2692,N_2771);
nand U2954 (N_2954,N_2725,N_2722);
nand U2955 (N_2955,N_2624,N_2758);
xor U2956 (N_2956,N_2608,N_2781);
or U2957 (N_2957,N_2717,N_2707);
or U2958 (N_2958,N_2795,N_2628);
and U2959 (N_2959,N_2711,N_2795);
nor U2960 (N_2960,N_2741,N_2671);
nand U2961 (N_2961,N_2737,N_2624);
and U2962 (N_2962,N_2625,N_2710);
and U2963 (N_2963,N_2751,N_2730);
nand U2964 (N_2964,N_2622,N_2720);
or U2965 (N_2965,N_2620,N_2668);
nor U2966 (N_2966,N_2780,N_2609);
xnor U2967 (N_2967,N_2750,N_2694);
or U2968 (N_2968,N_2761,N_2625);
and U2969 (N_2969,N_2789,N_2630);
nor U2970 (N_2970,N_2734,N_2783);
xnor U2971 (N_2971,N_2732,N_2639);
xor U2972 (N_2972,N_2631,N_2776);
nor U2973 (N_2973,N_2627,N_2602);
and U2974 (N_2974,N_2634,N_2784);
nor U2975 (N_2975,N_2744,N_2732);
nand U2976 (N_2976,N_2670,N_2638);
xnor U2977 (N_2977,N_2699,N_2620);
nor U2978 (N_2978,N_2652,N_2798);
or U2979 (N_2979,N_2781,N_2613);
xor U2980 (N_2980,N_2726,N_2668);
nand U2981 (N_2981,N_2665,N_2608);
nor U2982 (N_2982,N_2659,N_2649);
and U2983 (N_2983,N_2697,N_2763);
nor U2984 (N_2984,N_2646,N_2670);
and U2985 (N_2985,N_2796,N_2649);
nor U2986 (N_2986,N_2730,N_2677);
nand U2987 (N_2987,N_2712,N_2631);
and U2988 (N_2988,N_2621,N_2788);
and U2989 (N_2989,N_2683,N_2676);
or U2990 (N_2990,N_2651,N_2775);
or U2991 (N_2991,N_2705,N_2633);
nand U2992 (N_2992,N_2698,N_2792);
xor U2993 (N_2993,N_2635,N_2771);
and U2994 (N_2994,N_2688,N_2668);
and U2995 (N_2995,N_2683,N_2700);
or U2996 (N_2996,N_2792,N_2753);
xnor U2997 (N_2997,N_2626,N_2787);
and U2998 (N_2998,N_2742,N_2677);
nand U2999 (N_2999,N_2619,N_2754);
xnor U3000 (N_3000,N_2933,N_2942);
and U3001 (N_3001,N_2990,N_2910);
nor U3002 (N_3002,N_2987,N_2943);
nand U3003 (N_3003,N_2883,N_2863);
and U3004 (N_3004,N_2868,N_2970);
nor U3005 (N_3005,N_2825,N_2823);
nor U3006 (N_3006,N_2866,N_2912);
xor U3007 (N_3007,N_2814,N_2929);
and U3008 (N_3008,N_2934,N_2859);
and U3009 (N_3009,N_2837,N_2909);
or U3010 (N_3010,N_2851,N_2955);
or U3011 (N_3011,N_2925,N_2928);
nor U3012 (N_3012,N_2892,N_2827);
or U3013 (N_3013,N_2980,N_2979);
xor U3014 (N_3014,N_2963,N_2958);
xor U3015 (N_3015,N_2961,N_2875);
and U3016 (N_3016,N_2874,N_2916);
xor U3017 (N_3017,N_2893,N_2903);
xor U3018 (N_3018,N_2962,N_2890);
nor U3019 (N_3019,N_2832,N_2895);
nor U3020 (N_3020,N_2836,N_2994);
xor U3021 (N_3021,N_2948,N_2968);
xnor U3022 (N_3022,N_2996,N_2927);
and U3023 (N_3023,N_2959,N_2969);
xor U3024 (N_3024,N_2905,N_2804);
or U3025 (N_3025,N_2867,N_2820);
or U3026 (N_3026,N_2973,N_2880);
and U3027 (N_3027,N_2860,N_2900);
xnor U3028 (N_3028,N_2841,N_2908);
and U3029 (N_3029,N_2992,N_2865);
nand U3030 (N_3030,N_2915,N_2989);
nor U3031 (N_3031,N_2940,N_2956);
or U3032 (N_3032,N_2998,N_2920);
or U3033 (N_3033,N_2878,N_2977);
nand U3034 (N_3034,N_2843,N_2966);
xor U3035 (N_3035,N_2848,N_2995);
and U3036 (N_3036,N_2824,N_2826);
nor U3037 (N_3037,N_2862,N_2801);
nand U3038 (N_3038,N_2864,N_2967);
xnor U3039 (N_3039,N_2924,N_2870);
and U3040 (N_3040,N_2815,N_2991);
xnor U3041 (N_3041,N_2816,N_2853);
nor U3042 (N_3042,N_2930,N_2803);
xor U3043 (N_3043,N_2918,N_2896);
xnor U3044 (N_3044,N_2986,N_2839);
or U3045 (N_3045,N_2904,N_2984);
and U3046 (N_3046,N_2831,N_2951);
or U3047 (N_3047,N_2964,N_2894);
xnor U3048 (N_3048,N_2953,N_2976);
and U3049 (N_3049,N_2871,N_2949);
xor U3050 (N_3050,N_2957,N_2960);
nand U3051 (N_3051,N_2861,N_2842);
nand U3052 (N_3052,N_2885,N_2919);
or U3053 (N_3053,N_2985,N_2844);
and U3054 (N_3054,N_2931,N_2811);
and U3055 (N_3055,N_2952,N_2906);
and U3056 (N_3056,N_2809,N_2902);
nand U3057 (N_3057,N_2800,N_2805);
xnor U3058 (N_3058,N_2965,N_2850);
or U3059 (N_3059,N_2838,N_2852);
nor U3060 (N_3060,N_2829,N_2954);
and U3061 (N_3061,N_2899,N_2849);
and U3062 (N_3062,N_2822,N_2802);
xor U3063 (N_3063,N_2869,N_2999);
xor U3064 (N_3064,N_2944,N_2819);
nor U3065 (N_3065,N_2974,N_2898);
nor U3066 (N_3066,N_2807,N_2887);
and U3067 (N_3067,N_2840,N_2886);
nand U3068 (N_3068,N_2945,N_2858);
xnor U3069 (N_3069,N_2972,N_2813);
nand U3070 (N_3070,N_2856,N_2854);
or U3071 (N_3071,N_2971,N_2941);
xnor U3072 (N_3072,N_2810,N_2935);
nand U3073 (N_3073,N_2917,N_2932);
xnor U3074 (N_3074,N_2938,N_2879);
nor U3075 (N_3075,N_2975,N_2926);
xor U3076 (N_3076,N_2907,N_2812);
nand U3077 (N_3077,N_2857,N_2821);
and U3078 (N_3078,N_2947,N_2946);
and U3079 (N_3079,N_2806,N_2888);
and U3080 (N_3080,N_2818,N_2921);
and U3081 (N_3081,N_2847,N_2983);
and U3082 (N_3082,N_2897,N_2877);
and U3083 (N_3083,N_2993,N_2884);
xnor U3084 (N_3084,N_2872,N_2876);
or U3085 (N_3085,N_2846,N_2923);
nor U3086 (N_3086,N_2914,N_2913);
and U3087 (N_3087,N_2828,N_2808);
and U3088 (N_3088,N_2845,N_2982);
xor U3089 (N_3089,N_2922,N_2833);
nand U3090 (N_3090,N_2981,N_2891);
nand U3091 (N_3091,N_2835,N_2936);
nand U3092 (N_3092,N_2939,N_2855);
nand U3093 (N_3093,N_2901,N_2882);
and U3094 (N_3094,N_2889,N_2937);
and U3095 (N_3095,N_2834,N_2881);
nand U3096 (N_3096,N_2830,N_2950);
nor U3097 (N_3097,N_2911,N_2988);
and U3098 (N_3098,N_2978,N_2817);
nand U3099 (N_3099,N_2997,N_2873);
nor U3100 (N_3100,N_2816,N_2917);
nand U3101 (N_3101,N_2954,N_2804);
xor U3102 (N_3102,N_2962,N_2913);
nand U3103 (N_3103,N_2841,N_2899);
and U3104 (N_3104,N_2928,N_2823);
xor U3105 (N_3105,N_2913,N_2924);
nor U3106 (N_3106,N_2968,N_2842);
nand U3107 (N_3107,N_2841,N_2907);
xnor U3108 (N_3108,N_2819,N_2805);
or U3109 (N_3109,N_2899,N_2813);
or U3110 (N_3110,N_2896,N_2885);
or U3111 (N_3111,N_2948,N_2936);
nor U3112 (N_3112,N_2802,N_2830);
and U3113 (N_3113,N_2948,N_2875);
xor U3114 (N_3114,N_2875,N_2942);
and U3115 (N_3115,N_2809,N_2873);
and U3116 (N_3116,N_2883,N_2952);
or U3117 (N_3117,N_2917,N_2998);
or U3118 (N_3118,N_2924,N_2838);
nand U3119 (N_3119,N_2856,N_2890);
or U3120 (N_3120,N_2825,N_2835);
and U3121 (N_3121,N_2834,N_2827);
and U3122 (N_3122,N_2932,N_2939);
nand U3123 (N_3123,N_2873,N_2941);
nand U3124 (N_3124,N_2879,N_2911);
xnor U3125 (N_3125,N_2950,N_2957);
xor U3126 (N_3126,N_2897,N_2905);
nor U3127 (N_3127,N_2892,N_2839);
and U3128 (N_3128,N_2845,N_2873);
xor U3129 (N_3129,N_2927,N_2919);
nor U3130 (N_3130,N_2824,N_2965);
or U3131 (N_3131,N_2992,N_2826);
and U3132 (N_3132,N_2835,N_2805);
nand U3133 (N_3133,N_2995,N_2874);
or U3134 (N_3134,N_2918,N_2841);
nor U3135 (N_3135,N_2998,N_2827);
and U3136 (N_3136,N_2847,N_2867);
nand U3137 (N_3137,N_2842,N_2927);
or U3138 (N_3138,N_2859,N_2872);
xnor U3139 (N_3139,N_2847,N_2903);
xor U3140 (N_3140,N_2971,N_2873);
or U3141 (N_3141,N_2847,N_2932);
or U3142 (N_3142,N_2971,N_2952);
nor U3143 (N_3143,N_2916,N_2912);
nand U3144 (N_3144,N_2818,N_2815);
or U3145 (N_3145,N_2917,N_2985);
nor U3146 (N_3146,N_2912,N_2856);
or U3147 (N_3147,N_2936,N_2864);
nand U3148 (N_3148,N_2837,N_2984);
nor U3149 (N_3149,N_2893,N_2899);
or U3150 (N_3150,N_2924,N_2971);
nor U3151 (N_3151,N_2956,N_2816);
or U3152 (N_3152,N_2804,N_2927);
xor U3153 (N_3153,N_2890,N_2880);
or U3154 (N_3154,N_2952,N_2872);
or U3155 (N_3155,N_2837,N_2930);
and U3156 (N_3156,N_2961,N_2923);
xor U3157 (N_3157,N_2921,N_2836);
nor U3158 (N_3158,N_2806,N_2878);
or U3159 (N_3159,N_2934,N_2972);
xor U3160 (N_3160,N_2979,N_2801);
nand U3161 (N_3161,N_2908,N_2914);
nand U3162 (N_3162,N_2981,N_2820);
nand U3163 (N_3163,N_2834,N_2801);
or U3164 (N_3164,N_2944,N_2897);
nand U3165 (N_3165,N_2977,N_2822);
xnor U3166 (N_3166,N_2812,N_2800);
nand U3167 (N_3167,N_2922,N_2812);
or U3168 (N_3168,N_2966,N_2893);
nor U3169 (N_3169,N_2932,N_2849);
or U3170 (N_3170,N_2825,N_2962);
xnor U3171 (N_3171,N_2801,N_2828);
xor U3172 (N_3172,N_2883,N_2892);
or U3173 (N_3173,N_2919,N_2944);
and U3174 (N_3174,N_2879,N_2813);
or U3175 (N_3175,N_2875,N_2833);
nand U3176 (N_3176,N_2844,N_2832);
nor U3177 (N_3177,N_2836,N_2995);
nor U3178 (N_3178,N_2940,N_2911);
and U3179 (N_3179,N_2897,N_2850);
nor U3180 (N_3180,N_2845,N_2975);
and U3181 (N_3181,N_2826,N_2888);
nor U3182 (N_3182,N_2969,N_2920);
and U3183 (N_3183,N_2998,N_2923);
and U3184 (N_3184,N_2831,N_2976);
nand U3185 (N_3185,N_2907,N_2837);
or U3186 (N_3186,N_2951,N_2833);
nor U3187 (N_3187,N_2933,N_2856);
xor U3188 (N_3188,N_2889,N_2913);
and U3189 (N_3189,N_2973,N_2897);
nor U3190 (N_3190,N_2940,N_2986);
xor U3191 (N_3191,N_2847,N_2937);
nor U3192 (N_3192,N_2986,N_2917);
nor U3193 (N_3193,N_2867,N_2941);
and U3194 (N_3194,N_2872,N_2927);
and U3195 (N_3195,N_2856,N_2905);
xor U3196 (N_3196,N_2886,N_2975);
nor U3197 (N_3197,N_2926,N_2981);
and U3198 (N_3198,N_2977,N_2981);
xnor U3199 (N_3199,N_2901,N_2957);
nand U3200 (N_3200,N_3178,N_3173);
nor U3201 (N_3201,N_3167,N_3080);
nor U3202 (N_3202,N_3076,N_3131);
xor U3203 (N_3203,N_3175,N_3078);
nor U3204 (N_3204,N_3084,N_3026);
nor U3205 (N_3205,N_3031,N_3169);
xor U3206 (N_3206,N_3109,N_3138);
and U3207 (N_3207,N_3064,N_3044);
and U3208 (N_3208,N_3099,N_3139);
or U3209 (N_3209,N_3194,N_3004);
nor U3210 (N_3210,N_3006,N_3079);
nand U3211 (N_3211,N_3196,N_3003);
and U3212 (N_3212,N_3186,N_3033);
nand U3213 (N_3213,N_3012,N_3085);
xor U3214 (N_3214,N_3089,N_3171);
and U3215 (N_3215,N_3111,N_3100);
nand U3216 (N_3216,N_3071,N_3093);
nor U3217 (N_3217,N_3114,N_3025);
nor U3218 (N_3218,N_3094,N_3176);
and U3219 (N_3219,N_3145,N_3018);
and U3220 (N_3220,N_3082,N_3120);
xor U3221 (N_3221,N_3068,N_3188);
and U3222 (N_3222,N_3198,N_3141);
and U3223 (N_3223,N_3050,N_3092);
or U3224 (N_3224,N_3001,N_3197);
nor U3225 (N_3225,N_3143,N_3155);
or U3226 (N_3226,N_3177,N_3199);
and U3227 (N_3227,N_3190,N_3115);
or U3228 (N_3228,N_3156,N_3095);
nand U3229 (N_3229,N_3163,N_3191);
or U3230 (N_3230,N_3075,N_3021);
xnor U3231 (N_3231,N_3116,N_3187);
nor U3232 (N_3232,N_3052,N_3067);
or U3233 (N_3233,N_3136,N_3108);
or U3234 (N_3234,N_3192,N_3010);
xnor U3235 (N_3235,N_3154,N_3150);
or U3236 (N_3236,N_3124,N_3106);
and U3237 (N_3237,N_3184,N_3013);
or U3238 (N_3238,N_3066,N_3165);
nor U3239 (N_3239,N_3024,N_3090);
xor U3240 (N_3240,N_3107,N_3158);
or U3241 (N_3241,N_3053,N_3164);
and U3242 (N_3242,N_3129,N_3170);
nor U3243 (N_3243,N_3029,N_3030);
nand U3244 (N_3244,N_3023,N_3000);
and U3245 (N_3245,N_3069,N_3051);
nand U3246 (N_3246,N_3137,N_3047);
nor U3247 (N_3247,N_3179,N_3020);
or U3248 (N_3248,N_3042,N_3022);
nand U3249 (N_3249,N_3102,N_3027);
nand U3250 (N_3250,N_3034,N_3151);
or U3251 (N_3251,N_3162,N_3110);
nand U3252 (N_3252,N_3086,N_3101);
nor U3253 (N_3253,N_3134,N_3038);
xnor U3254 (N_3254,N_3011,N_3081);
nor U3255 (N_3255,N_3103,N_3056);
nor U3256 (N_3256,N_3127,N_3189);
and U3257 (N_3257,N_3148,N_3174);
or U3258 (N_3258,N_3055,N_3161);
xor U3259 (N_3259,N_3077,N_3183);
and U3260 (N_3260,N_3028,N_3009);
xnor U3261 (N_3261,N_3017,N_3125);
nand U3262 (N_3262,N_3104,N_3152);
or U3263 (N_3263,N_3063,N_3065);
nor U3264 (N_3264,N_3181,N_3096);
or U3265 (N_3265,N_3097,N_3153);
or U3266 (N_3266,N_3160,N_3083);
nor U3267 (N_3267,N_3180,N_3149);
xor U3268 (N_3268,N_3126,N_3048);
xnor U3269 (N_3269,N_3135,N_3061);
and U3270 (N_3270,N_3037,N_3032);
nor U3271 (N_3271,N_3117,N_3128);
and U3272 (N_3272,N_3123,N_3087);
nand U3273 (N_3273,N_3122,N_3057);
nand U3274 (N_3274,N_3014,N_3168);
nor U3275 (N_3275,N_3147,N_3062);
and U3276 (N_3276,N_3016,N_3113);
or U3277 (N_3277,N_3088,N_3008);
xor U3278 (N_3278,N_3146,N_3072);
xor U3279 (N_3279,N_3049,N_3121);
nand U3280 (N_3280,N_3144,N_3005);
and U3281 (N_3281,N_3185,N_3074);
nand U3282 (N_3282,N_3058,N_3105);
xor U3283 (N_3283,N_3119,N_3002);
or U3284 (N_3284,N_3036,N_3045);
nand U3285 (N_3285,N_3172,N_3060);
xor U3286 (N_3286,N_3041,N_3073);
nand U3287 (N_3287,N_3007,N_3133);
nand U3288 (N_3288,N_3091,N_3130);
nand U3289 (N_3289,N_3040,N_3015);
and U3290 (N_3290,N_3195,N_3054);
xor U3291 (N_3291,N_3157,N_3159);
xor U3292 (N_3292,N_3046,N_3142);
nor U3293 (N_3293,N_3059,N_3035);
nand U3294 (N_3294,N_3118,N_3070);
nand U3295 (N_3295,N_3039,N_3019);
or U3296 (N_3296,N_3182,N_3166);
or U3297 (N_3297,N_3112,N_3140);
nand U3298 (N_3298,N_3132,N_3193);
xor U3299 (N_3299,N_3098,N_3043);
and U3300 (N_3300,N_3089,N_3136);
nor U3301 (N_3301,N_3141,N_3059);
nand U3302 (N_3302,N_3170,N_3134);
nor U3303 (N_3303,N_3142,N_3117);
and U3304 (N_3304,N_3047,N_3050);
or U3305 (N_3305,N_3056,N_3110);
nor U3306 (N_3306,N_3007,N_3067);
and U3307 (N_3307,N_3134,N_3071);
xnor U3308 (N_3308,N_3116,N_3097);
and U3309 (N_3309,N_3100,N_3092);
xor U3310 (N_3310,N_3199,N_3044);
nand U3311 (N_3311,N_3153,N_3005);
or U3312 (N_3312,N_3078,N_3013);
and U3313 (N_3313,N_3056,N_3163);
nand U3314 (N_3314,N_3174,N_3027);
xnor U3315 (N_3315,N_3129,N_3191);
and U3316 (N_3316,N_3088,N_3104);
or U3317 (N_3317,N_3097,N_3105);
or U3318 (N_3318,N_3095,N_3059);
and U3319 (N_3319,N_3095,N_3174);
nand U3320 (N_3320,N_3111,N_3133);
or U3321 (N_3321,N_3009,N_3193);
xor U3322 (N_3322,N_3038,N_3118);
nor U3323 (N_3323,N_3101,N_3053);
and U3324 (N_3324,N_3181,N_3098);
nand U3325 (N_3325,N_3193,N_3052);
and U3326 (N_3326,N_3003,N_3102);
or U3327 (N_3327,N_3027,N_3157);
and U3328 (N_3328,N_3019,N_3147);
or U3329 (N_3329,N_3183,N_3138);
and U3330 (N_3330,N_3039,N_3103);
nor U3331 (N_3331,N_3022,N_3191);
nand U3332 (N_3332,N_3113,N_3036);
nor U3333 (N_3333,N_3142,N_3126);
xor U3334 (N_3334,N_3087,N_3097);
nand U3335 (N_3335,N_3141,N_3019);
or U3336 (N_3336,N_3047,N_3101);
nor U3337 (N_3337,N_3052,N_3155);
and U3338 (N_3338,N_3162,N_3172);
nand U3339 (N_3339,N_3092,N_3080);
xor U3340 (N_3340,N_3166,N_3176);
or U3341 (N_3341,N_3146,N_3119);
or U3342 (N_3342,N_3047,N_3078);
and U3343 (N_3343,N_3073,N_3001);
or U3344 (N_3344,N_3123,N_3014);
nand U3345 (N_3345,N_3159,N_3148);
nand U3346 (N_3346,N_3044,N_3045);
and U3347 (N_3347,N_3157,N_3026);
and U3348 (N_3348,N_3151,N_3051);
nor U3349 (N_3349,N_3077,N_3055);
xor U3350 (N_3350,N_3169,N_3165);
and U3351 (N_3351,N_3178,N_3174);
or U3352 (N_3352,N_3183,N_3042);
and U3353 (N_3353,N_3148,N_3086);
nor U3354 (N_3354,N_3152,N_3139);
and U3355 (N_3355,N_3199,N_3119);
nand U3356 (N_3356,N_3152,N_3032);
xnor U3357 (N_3357,N_3000,N_3158);
nor U3358 (N_3358,N_3141,N_3018);
xor U3359 (N_3359,N_3082,N_3038);
or U3360 (N_3360,N_3058,N_3160);
or U3361 (N_3361,N_3128,N_3143);
or U3362 (N_3362,N_3046,N_3113);
or U3363 (N_3363,N_3045,N_3157);
and U3364 (N_3364,N_3182,N_3163);
xnor U3365 (N_3365,N_3168,N_3130);
nand U3366 (N_3366,N_3038,N_3025);
or U3367 (N_3367,N_3164,N_3153);
nand U3368 (N_3368,N_3157,N_3142);
nand U3369 (N_3369,N_3109,N_3143);
nand U3370 (N_3370,N_3034,N_3038);
nand U3371 (N_3371,N_3155,N_3164);
or U3372 (N_3372,N_3151,N_3183);
nand U3373 (N_3373,N_3182,N_3125);
and U3374 (N_3374,N_3037,N_3117);
and U3375 (N_3375,N_3149,N_3080);
nand U3376 (N_3376,N_3123,N_3198);
nand U3377 (N_3377,N_3155,N_3158);
nand U3378 (N_3378,N_3051,N_3045);
nand U3379 (N_3379,N_3030,N_3172);
xor U3380 (N_3380,N_3189,N_3001);
or U3381 (N_3381,N_3005,N_3078);
or U3382 (N_3382,N_3056,N_3067);
nand U3383 (N_3383,N_3087,N_3045);
or U3384 (N_3384,N_3041,N_3037);
nand U3385 (N_3385,N_3058,N_3116);
or U3386 (N_3386,N_3039,N_3085);
nor U3387 (N_3387,N_3023,N_3137);
nand U3388 (N_3388,N_3137,N_3028);
xnor U3389 (N_3389,N_3039,N_3199);
nand U3390 (N_3390,N_3172,N_3165);
xnor U3391 (N_3391,N_3129,N_3134);
nor U3392 (N_3392,N_3137,N_3084);
nor U3393 (N_3393,N_3024,N_3017);
and U3394 (N_3394,N_3148,N_3031);
xnor U3395 (N_3395,N_3158,N_3109);
or U3396 (N_3396,N_3037,N_3153);
xnor U3397 (N_3397,N_3198,N_3021);
or U3398 (N_3398,N_3108,N_3086);
nor U3399 (N_3399,N_3014,N_3054);
or U3400 (N_3400,N_3366,N_3392);
or U3401 (N_3401,N_3310,N_3381);
or U3402 (N_3402,N_3210,N_3208);
xnor U3403 (N_3403,N_3351,N_3204);
xor U3404 (N_3404,N_3397,N_3279);
or U3405 (N_3405,N_3211,N_3395);
nand U3406 (N_3406,N_3382,N_3336);
nor U3407 (N_3407,N_3353,N_3333);
xnor U3408 (N_3408,N_3317,N_3268);
nor U3409 (N_3409,N_3322,N_3232);
xor U3410 (N_3410,N_3393,N_3378);
nor U3411 (N_3411,N_3386,N_3238);
nand U3412 (N_3412,N_3389,N_3315);
nor U3413 (N_3413,N_3359,N_3229);
and U3414 (N_3414,N_3228,N_3251);
and U3415 (N_3415,N_3246,N_3379);
nor U3416 (N_3416,N_3242,N_3349);
and U3417 (N_3417,N_3244,N_3354);
or U3418 (N_3418,N_3266,N_3258);
nand U3419 (N_3419,N_3295,N_3287);
or U3420 (N_3420,N_3285,N_3290);
and U3421 (N_3421,N_3280,N_3203);
xor U3422 (N_3422,N_3223,N_3339);
xor U3423 (N_3423,N_3355,N_3236);
nand U3424 (N_3424,N_3293,N_3248);
nand U3425 (N_3425,N_3252,N_3342);
xor U3426 (N_3426,N_3256,N_3284);
nor U3427 (N_3427,N_3220,N_3292);
and U3428 (N_3428,N_3318,N_3249);
nor U3429 (N_3429,N_3334,N_3347);
nor U3430 (N_3430,N_3344,N_3301);
or U3431 (N_3431,N_3328,N_3300);
nor U3432 (N_3432,N_3222,N_3320);
and U3433 (N_3433,N_3274,N_3371);
or U3434 (N_3434,N_3216,N_3313);
xnor U3435 (N_3435,N_3350,N_3373);
xnor U3436 (N_3436,N_3296,N_3370);
xor U3437 (N_3437,N_3218,N_3281);
and U3438 (N_3438,N_3270,N_3376);
xor U3439 (N_3439,N_3213,N_3399);
or U3440 (N_3440,N_3321,N_3235);
nand U3441 (N_3441,N_3352,N_3231);
and U3442 (N_3442,N_3230,N_3253);
nor U3443 (N_3443,N_3233,N_3247);
and U3444 (N_3444,N_3234,N_3390);
and U3445 (N_3445,N_3269,N_3341);
nand U3446 (N_3446,N_3338,N_3363);
nand U3447 (N_3447,N_3312,N_3329);
nand U3448 (N_3448,N_3225,N_3245);
nand U3449 (N_3449,N_3297,N_3276);
xnor U3450 (N_3450,N_3314,N_3388);
xor U3451 (N_3451,N_3375,N_3367);
nor U3452 (N_3452,N_3387,N_3306);
nand U3453 (N_3453,N_3205,N_3298);
nand U3454 (N_3454,N_3374,N_3267);
nor U3455 (N_3455,N_3364,N_3377);
nand U3456 (N_3456,N_3368,N_3391);
nand U3457 (N_3457,N_3277,N_3286);
or U3458 (N_3458,N_3271,N_3291);
and U3459 (N_3459,N_3326,N_3308);
nor U3460 (N_3460,N_3332,N_3224);
or U3461 (N_3461,N_3282,N_3250);
and U3462 (N_3462,N_3275,N_3207);
nor U3463 (N_3463,N_3324,N_3360);
nor U3464 (N_3464,N_3331,N_3396);
or U3465 (N_3465,N_3335,N_3265);
nand U3466 (N_3466,N_3383,N_3263);
or U3467 (N_3467,N_3262,N_3219);
and U3468 (N_3468,N_3254,N_3358);
and U3469 (N_3469,N_3200,N_3348);
xor U3470 (N_3470,N_3257,N_3302);
nand U3471 (N_3471,N_3209,N_3201);
xor U3472 (N_3472,N_3304,N_3398);
xnor U3473 (N_3473,N_3227,N_3202);
or U3474 (N_3474,N_3340,N_3259);
nor U3475 (N_3475,N_3307,N_3361);
xnor U3476 (N_3476,N_3316,N_3243);
or U3477 (N_3477,N_3206,N_3319);
and U3478 (N_3478,N_3380,N_3372);
nand U3479 (N_3479,N_3240,N_3264);
or U3480 (N_3480,N_3356,N_3260);
nand U3481 (N_3481,N_3294,N_3214);
and U3482 (N_3482,N_3309,N_3384);
or U3483 (N_3483,N_3385,N_3369);
nand U3484 (N_3484,N_3299,N_3261);
or U3485 (N_3485,N_3325,N_3272);
xnor U3486 (N_3486,N_3283,N_3221);
xor U3487 (N_3487,N_3289,N_3255);
nand U3488 (N_3488,N_3226,N_3394);
nor U3489 (N_3489,N_3337,N_3362);
nand U3490 (N_3490,N_3330,N_3212);
and U3491 (N_3491,N_3311,N_3239);
nor U3492 (N_3492,N_3357,N_3343);
xnor U3493 (N_3493,N_3215,N_3273);
nor U3494 (N_3494,N_3237,N_3323);
nor U3495 (N_3495,N_3365,N_3241);
xor U3496 (N_3496,N_3303,N_3327);
nand U3497 (N_3497,N_3288,N_3278);
or U3498 (N_3498,N_3346,N_3345);
nor U3499 (N_3499,N_3305,N_3217);
or U3500 (N_3500,N_3227,N_3263);
or U3501 (N_3501,N_3283,N_3241);
nand U3502 (N_3502,N_3229,N_3382);
nand U3503 (N_3503,N_3311,N_3220);
nand U3504 (N_3504,N_3245,N_3398);
and U3505 (N_3505,N_3279,N_3257);
and U3506 (N_3506,N_3310,N_3261);
or U3507 (N_3507,N_3213,N_3355);
and U3508 (N_3508,N_3273,N_3240);
or U3509 (N_3509,N_3241,N_3274);
and U3510 (N_3510,N_3381,N_3332);
nor U3511 (N_3511,N_3217,N_3301);
nand U3512 (N_3512,N_3294,N_3398);
or U3513 (N_3513,N_3392,N_3290);
nor U3514 (N_3514,N_3234,N_3321);
xnor U3515 (N_3515,N_3248,N_3345);
nor U3516 (N_3516,N_3308,N_3284);
nand U3517 (N_3517,N_3385,N_3371);
xor U3518 (N_3518,N_3329,N_3202);
or U3519 (N_3519,N_3238,N_3382);
nand U3520 (N_3520,N_3370,N_3391);
nor U3521 (N_3521,N_3368,N_3252);
nor U3522 (N_3522,N_3253,N_3239);
nor U3523 (N_3523,N_3365,N_3232);
or U3524 (N_3524,N_3290,N_3390);
nand U3525 (N_3525,N_3219,N_3363);
nand U3526 (N_3526,N_3336,N_3298);
nor U3527 (N_3527,N_3281,N_3313);
nor U3528 (N_3528,N_3249,N_3262);
nand U3529 (N_3529,N_3307,N_3212);
nor U3530 (N_3530,N_3236,N_3237);
xnor U3531 (N_3531,N_3333,N_3321);
nand U3532 (N_3532,N_3205,N_3206);
and U3533 (N_3533,N_3390,N_3302);
and U3534 (N_3534,N_3347,N_3204);
xor U3535 (N_3535,N_3380,N_3303);
nand U3536 (N_3536,N_3294,N_3237);
and U3537 (N_3537,N_3239,N_3308);
nor U3538 (N_3538,N_3263,N_3257);
xor U3539 (N_3539,N_3288,N_3222);
nor U3540 (N_3540,N_3285,N_3388);
xnor U3541 (N_3541,N_3307,N_3325);
nand U3542 (N_3542,N_3353,N_3393);
xnor U3543 (N_3543,N_3254,N_3208);
xor U3544 (N_3544,N_3296,N_3304);
nand U3545 (N_3545,N_3342,N_3318);
nor U3546 (N_3546,N_3361,N_3283);
and U3547 (N_3547,N_3286,N_3377);
xor U3548 (N_3548,N_3347,N_3310);
and U3549 (N_3549,N_3330,N_3210);
or U3550 (N_3550,N_3280,N_3219);
xnor U3551 (N_3551,N_3334,N_3289);
and U3552 (N_3552,N_3326,N_3255);
xnor U3553 (N_3553,N_3212,N_3292);
nor U3554 (N_3554,N_3394,N_3231);
xor U3555 (N_3555,N_3255,N_3263);
nor U3556 (N_3556,N_3351,N_3254);
or U3557 (N_3557,N_3330,N_3302);
nand U3558 (N_3558,N_3330,N_3312);
or U3559 (N_3559,N_3224,N_3313);
and U3560 (N_3560,N_3357,N_3261);
or U3561 (N_3561,N_3302,N_3254);
nand U3562 (N_3562,N_3394,N_3205);
xnor U3563 (N_3563,N_3379,N_3311);
nor U3564 (N_3564,N_3252,N_3251);
nand U3565 (N_3565,N_3275,N_3237);
or U3566 (N_3566,N_3289,N_3312);
xor U3567 (N_3567,N_3368,N_3369);
nand U3568 (N_3568,N_3274,N_3305);
or U3569 (N_3569,N_3294,N_3303);
or U3570 (N_3570,N_3343,N_3358);
xnor U3571 (N_3571,N_3383,N_3390);
xnor U3572 (N_3572,N_3388,N_3384);
xnor U3573 (N_3573,N_3373,N_3243);
or U3574 (N_3574,N_3325,N_3314);
and U3575 (N_3575,N_3206,N_3296);
and U3576 (N_3576,N_3396,N_3362);
or U3577 (N_3577,N_3371,N_3340);
and U3578 (N_3578,N_3394,N_3285);
xnor U3579 (N_3579,N_3323,N_3360);
or U3580 (N_3580,N_3379,N_3269);
and U3581 (N_3581,N_3220,N_3260);
xor U3582 (N_3582,N_3321,N_3209);
and U3583 (N_3583,N_3246,N_3271);
xor U3584 (N_3584,N_3380,N_3273);
and U3585 (N_3585,N_3319,N_3268);
xor U3586 (N_3586,N_3272,N_3356);
nor U3587 (N_3587,N_3230,N_3342);
nand U3588 (N_3588,N_3250,N_3388);
nand U3589 (N_3589,N_3306,N_3390);
nand U3590 (N_3590,N_3392,N_3237);
or U3591 (N_3591,N_3341,N_3205);
xnor U3592 (N_3592,N_3236,N_3394);
or U3593 (N_3593,N_3347,N_3284);
nand U3594 (N_3594,N_3328,N_3204);
nor U3595 (N_3595,N_3326,N_3279);
and U3596 (N_3596,N_3383,N_3299);
nand U3597 (N_3597,N_3274,N_3279);
nand U3598 (N_3598,N_3265,N_3396);
and U3599 (N_3599,N_3318,N_3361);
and U3600 (N_3600,N_3538,N_3451);
or U3601 (N_3601,N_3432,N_3569);
nor U3602 (N_3602,N_3426,N_3549);
nand U3603 (N_3603,N_3449,N_3407);
and U3604 (N_3604,N_3579,N_3425);
xor U3605 (N_3605,N_3502,N_3563);
or U3606 (N_3606,N_3543,N_3535);
or U3607 (N_3607,N_3442,N_3592);
nand U3608 (N_3608,N_3486,N_3530);
nand U3609 (N_3609,N_3534,N_3459);
nand U3610 (N_3610,N_3420,N_3401);
nand U3611 (N_3611,N_3562,N_3533);
nor U3612 (N_3612,N_3469,N_3542);
and U3613 (N_3613,N_3552,N_3590);
xnor U3614 (N_3614,N_3404,N_3496);
nand U3615 (N_3615,N_3561,N_3595);
and U3616 (N_3616,N_3421,N_3585);
xnor U3617 (N_3617,N_3591,N_3488);
nor U3618 (N_3618,N_3566,N_3540);
nand U3619 (N_3619,N_3487,N_3443);
nand U3620 (N_3620,N_3429,N_3567);
nor U3621 (N_3621,N_3597,N_3531);
nor U3622 (N_3622,N_3501,N_3415);
and U3623 (N_3623,N_3500,N_3507);
nor U3624 (N_3624,N_3524,N_3472);
xor U3625 (N_3625,N_3571,N_3482);
and U3626 (N_3626,N_3453,N_3427);
or U3627 (N_3627,N_3445,N_3495);
nand U3628 (N_3628,N_3550,N_3458);
and U3629 (N_3629,N_3478,N_3479);
xor U3630 (N_3630,N_3525,N_3438);
and U3631 (N_3631,N_3460,N_3412);
nor U3632 (N_3632,N_3466,N_3548);
or U3633 (N_3633,N_3435,N_3536);
nand U3634 (N_3634,N_3439,N_3411);
nand U3635 (N_3635,N_3428,N_3514);
nand U3636 (N_3636,N_3532,N_3450);
nand U3637 (N_3637,N_3494,N_3511);
nand U3638 (N_3638,N_3584,N_3546);
xor U3639 (N_3639,N_3462,N_3456);
nor U3640 (N_3640,N_3491,N_3572);
nor U3641 (N_3641,N_3512,N_3498);
nand U3642 (N_3642,N_3518,N_3454);
nor U3643 (N_3643,N_3430,N_3422);
and U3644 (N_3644,N_3523,N_3473);
and U3645 (N_3645,N_3434,N_3544);
and U3646 (N_3646,N_3489,N_3527);
and U3647 (N_3647,N_3416,N_3461);
nor U3648 (N_3648,N_3481,N_3475);
or U3649 (N_3649,N_3526,N_3519);
xor U3650 (N_3650,N_3455,N_3499);
xor U3651 (N_3651,N_3589,N_3485);
and U3652 (N_3652,N_3587,N_3557);
and U3653 (N_3653,N_3483,N_3441);
xor U3654 (N_3654,N_3529,N_3594);
or U3655 (N_3655,N_3477,N_3419);
xor U3656 (N_3656,N_3431,N_3560);
and U3657 (N_3657,N_3586,N_3505);
xnor U3658 (N_3658,N_3446,N_3463);
nor U3659 (N_3659,N_3440,N_3577);
and U3660 (N_3660,N_3554,N_3464);
xnor U3661 (N_3661,N_3433,N_3410);
nor U3662 (N_3662,N_3509,N_3582);
nor U3663 (N_3663,N_3539,N_3490);
and U3664 (N_3664,N_3564,N_3403);
nand U3665 (N_3665,N_3413,N_3555);
or U3666 (N_3666,N_3553,N_3418);
and U3667 (N_3667,N_3470,N_3405);
nand U3668 (N_3668,N_3468,N_3508);
nor U3669 (N_3669,N_3574,N_3402);
and U3670 (N_3670,N_3575,N_3520);
nand U3671 (N_3671,N_3510,N_3424);
and U3672 (N_3672,N_3598,N_3408);
xnor U3673 (N_3673,N_3559,N_3522);
xor U3674 (N_3674,N_3588,N_3581);
nor U3675 (N_3675,N_3580,N_3506);
nand U3676 (N_3676,N_3596,N_3493);
xor U3677 (N_3677,N_3578,N_3537);
xor U3678 (N_3678,N_3504,N_3516);
and U3679 (N_3679,N_3568,N_3573);
nor U3680 (N_3680,N_3558,N_3406);
or U3681 (N_3681,N_3593,N_3476);
nand U3682 (N_3682,N_3503,N_3417);
or U3683 (N_3683,N_3400,N_3556);
nand U3684 (N_3684,N_3576,N_3471);
xor U3685 (N_3685,N_3551,N_3545);
nor U3686 (N_3686,N_3515,N_3423);
nand U3687 (N_3687,N_3465,N_3513);
nand U3688 (N_3688,N_3448,N_3565);
or U3689 (N_3689,N_3447,N_3457);
nor U3690 (N_3690,N_3492,N_3409);
or U3691 (N_3691,N_3480,N_3452);
and U3692 (N_3692,N_3517,N_3528);
nor U3693 (N_3693,N_3521,N_3484);
nand U3694 (N_3694,N_3570,N_3467);
and U3695 (N_3695,N_3547,N_3436);
and U3696 (N_3696,N_3474,N_3414);
nand U3697 (N_3697,N_3497,N_3444);
and U3698 (N_3698,N_3437,N_3583);
xor U3699 (N_3699,N_3541,N_3599);
nor U3700 (N_3700,N_3542,N_3451);
nor U3701 (N_3701,N_3592,N_3484);
and U3702 (N_3702,N_3531,N_3518);
and U3703 (N_3703,N_3459,N_3431);
xnor U3704 (N_3704,N_3451,N_3449);
or U3705 (N_3705,N_3598,N_3438);
and U3706 (N_3706,N_3574,N_3581);
and U3707 (N_3707,N_3538,N_3485);
xor U3708 (N_3708,N_3522,N_3540);
and U3709 (N_3709,N_3497,N_3443);
and U3710 (N_3710,N_3400,N_3585);
and U3711 (N_3711,N_3432,N_3578);
xor U3712 (N_3712,N_3595,N_3494);
nand U3713 (N_3713,N_3525,N_3578);
and U3714 (N_3714,N_3412,N_3503);
or U3715 (N_3715,N_3434,N_3557);
xor U3716 (N_3716,N_3452,N_3423);
xor U3717 (N_3717,N_3542,N_3434);
nand U3718 (N_3718,N_3415,N_3556);
nand U3719 (N_3719,N_3400,N_3479);
nand U3720 (N_3720,N_3434,N_3422);
xor U3721 (N_3721,N_3414,N_3515);
nand U3722 (N_3722,N_3581,N_3528);
or U3723 (N_3723,N_3419,N_3489);
nor U3724 (N_3724,N_3426,N_3571);
nand U3725 (N_3725,N_3470,N_3595);
and U3726 (N_3726,N_3485,N_3519);
nor U3727 (N_3727,N_3483,N_3574);
nand U3728 (N_3728,N_3568,N_3402);
xnor U3729 (N_3729,N_3472,N_3439);
nor U3730 (N_3730,N_3506,N_3473);
xor U3731 (N_3731,N_3580,N_3480);
nand U3732 (N_3732,N_3589,N_3575);
or U3733 (N_3733,N_3590,N_3562);
or U3734 (N_3734,N_3480,N_3559);
and U3735 (N_3735,N_3439,N_3587);
or U3736 (N_3736,N_3498,N_3429);
or U3737 (N_3737,N_3563,N_3448);
nor U3738 (N_3738,N_3494,N_3528);
nand U3739 (N_3739,N_3401,N_3409);
or U3740 (N_3740,N_3574,N_3532);
or U3741 (N_3741,N_3506,N_3460);
nor U3742 (N_3742,N_3509,N_3492);
xor U3743 (N_3743,N_3587,N_3519);
nor U3744 (N_3744,N_3562,N_3473);
and U3745 (N_3745,N_3556,N_3428);
or U3746 (N_3746,N_3527,N_3575);
or U3747 (N_3747,N_3503,N_3546);
or U3748 (N_3748,N_3411,N_3428);
or U3749 (N_3749,N_3530,N_3466);
nor U3750 (N_3750,N_3585,N_3517);
nor U3751 (N_3751,N_3415,N_3487);
and U3752 (N_3752,N_3481,N_3558);
nor U3753 (N_3753,N_3437,N_3406);
nor U3754 (N_3754,N_3559,N_3551);
and U3755 (N_3755,N_3596,N_3579);
or U3756 (N_3756,N_3498,N_3518);
xnor U3757 (N_3757,N_3583,N_3444);
or U3758 (N_3758,N_3570,N_3508);
or U3759 (N_3759,N_3432,N_3517);
nor U3760 (N_3760,N_3545,N_3482);
nor U3761 (N_3761,N_3532,N_3416);
nor U3762 (N_3762,N_3588,N_3554);
or U3763 (N_3763,N_3488,N_3455);
nor U3764 (N_3764,N_3531,N_3460);
or U3765 (N_3765,N_3413,N_3479);
xnor U3766 (N_3766,N_3419,N_3423);
or U3767 (N_3767,N_3561,N_3412);
or U3768 (N_3768,N_3585,N_3563);
and U3769 (N_3769,N_3422,N_3522);
xor U3770 (N_3770,N_3450,N_3481);
nand U3771 (N_3771,N_3539,N_3410);
nand U3772 (N_3772,N_3421,N_3453);
nand U3773 (N_3773,N_3403,N_3561);
or U3774 (N_3774,N_3452,N_3556);
and U3775 (N_3775,N_3403,N_3412);
and U3776 (N_3776,N_3565,N_3526);
xor U3777 (N_3777,N_3431,N_3457);
xor U3778 (N_3778,N_3548,N_3435);
nand U3779 (N_3779,N_3544,N_3588);
or U3780 (N_3780,N_3539,N_3515);
or U3781 (N_3781,N_3463,N_3570);
or U3782 (N_3782,N_3498,N_3487);
or U3783 (N_3783,N_3479,N_3466);
xnor U3784 (N_3784,N_3417,N_3492);
nand U3785 (N_3785,N_3449,N_3402);
nand U3786 (N_3786,N_3436,N_3478);
nor U3787 (N_3787,N_3599,N_3433);
nand U3788 (N_3788,N_3415,N_3545);
and U3789 (N_3789,N_3462,N_3571);
xor U3790 (N_3790,N_3513,N_3516);
and U3791 (N_3791,N_3560,N_3500);
and U3792 (N_3792,N_3415,N_3516);
xor U3793 (N_3793,N_3412,N_3532);
and U3794 (N_3794,N_3527,N_3452);
nand U3795 (N_3795,N_3596,N_3458);
nand U3796 (N_3796,N_3421,N_3580);
nor U3797 (N_3797,N_3561,N_3490);
or U3798 (N_3798,N_3478,N_3532);
and U3799 (N_3799,N_3589,N_3527);
nand U3800 (N_3800,N_3630,N_3759);
nor U3801 (N_3801,N_3605,N_3701);
nand U3802 (N_3802,N_3719,N_3609);
or U3803 (N_3803,N_3787,N_3707);
or U3804 (N_3804,N_3780,N_3722);
xor U3805 (N_3805,N_3673,N_3753);
and U3806 (N_3806,N_3634,N_3694);
or U3807 (N_3807,N_3734,N_3785);
or U3808 (N_3808,N_3705,N_3614);
nor U3809 (N_3809,N_3711,N_3791);
or U3810 (N_3810,N_3714,N_3782);
or U3811 (N_3811,N_3706,N_3740);
nand U3812 (N_3812,N_3619,N_3709);
or U3813 (N_3813,N_3604,N_3655);
xor U3814 (N_3814,N_3646,N_3687);
nor U3815 (N_3815,N_3799,N_3767);
xor U3816 (N_3816,N_3679,N_3750);
or U3817 (N_3817,N_3712,N_3738);
or U3818 (N_3818,N_3650,N_3690);
nand U3819 (N_3819,N_3716,N_3657);
xor U3820 (N_3820,N_3798,N_3635);
nand U3821 (N_3821,N_3676,N_3731);
nand U3822 (N_3822,N_3662,N_3652);
or U3823 (N_3823,N_3645,N_3729);
nor U3824 (N_3824,N_3728,N_3717);
and U3825 (N_3825,N_3675,N_3770);
nor U3826 (N_3826,N_3772,N_3749);
nand U3827 (N_3827,N_3744,N_3765);
nor U3828 (N_3828,N_3625,N_3684);
and U3829 (N_3829,N_3617,N_3653);
or U3830 (N_3830,N_3726,N_3794);
xnor U3831 (N_3831,N_3797,N_3760);
xor U3832 (N_3832,N_3697,N_3761);
nor U3833 (N_3833,N_3695,N_3627);
nor U3834 (N_3834,N_3763,N_3677);
nand U3835 (N_3835,N_3668,N_3642);
nor U3836 (N_3836,N_3660,N_3764);
nand U3837 (N_3837,N_3735,N_3688);
nand U3838 (N_3838,N_3793,N_3727);
and U3839 (N_3839,N_3643,N_3710);
or U3840 (N_3840,N_3628,N_3626);
xor U3841 (N_3841,N_3664,N_3757);
and U3842 (N_3842,N_3631,N_3752);
and U3843 (N_3843,N_3689,N_3732);
and U3844 (N_3844,N_3699,N_3641);
xnor U3845 (N_3845,N_3755,N_3708);
nand U3846 (N_3846,N_3762,N_3723);
nor U3847 (N_3847,N_3746,N_3777);
or U3848 (N_3848,N_3637,N_3665);
and U3849 (N_3849,N_3640,N_3651);
xnor U3850 (N_3850,N_3685,N_3747);
or U3851 (N_3851,N_3788,N_3769);
xnor U3852 (N_3852,N_3779,N_3766);
xnor U3853 (N_3853,N_3667,N_3721);
nor U3854 (N_3854,N_3683,N_3629);
and U3855 (N_3855,N_3718,N_3774);
xnor U3856 (N_3856,N_3666,N_3636);
xnor U3857 (N_3857,N_3678,N_3790);
nand U3858 (N_3858,N_3648,N_3622);
nor U3859 (N_3859,N_3702,N_3670);
nor U3860 (N_3860,N_3671,N_3700);
and U3861 (N_3861,N_3692,N_3743);
and U3862 (N_3862,N_3783,N_3720);
nand U3863 (N_3863,N_3616,N_3672);
nor U3864 (N_3864,N_3748,N_3610);
and U3865 (N_3865,N_3795,N_3758);
nor U3866 (N_3866,N_3620,N_3644);
and U3867 (N_3867,N_3775,N_3613);
nor U3868 (N_3868,N_3773,N_3789);
or U3869 (N_3869,N_3786,N_3698);
and U3870 (N_3870,N_3618,N_3715);
nor U3871 (N_3871,N_3612,N_3600);
nor U3872 (N_3872,N_3658,N_3686);
nand U3873 (N_3873,N_3754,N_3781);
xnor U3874 (N_3874,N_3725,N_3654);
nand U3875 (N_3875,N_3776,N_3661);
nor U3876 (N_3876,N_3792,N_3739);
or U3877 (N_3877,N_3649,N_3611);
nand U3878 (N_3878,N_3768,N_3771);
nor U3879 (N_3879,N_3601,N_3669);
or U3880 (N_3880,N_3713,N_3615);
and U3881 (N_3881,N_3736,N_3733);
xnor U3882 (N_3882,N_3742,N_3638);
and U3883 (N_3883,N_3663,N_3607);
or U3884 (N_3884,N_3778,N_3730);
xor U3885 (N_3885,N_3756,N_3696);
and U3886 (N_3886,N_3693,N_3632);
nor U3887 (N_3887,N_3674,N_3703);
nand U3888 (N_3888,N_3659,N_3784);
nor U3889 (N_3889,N_3602,N_3681);
and U3890 (N_3890,N_3737,N_3796);
or U3891 (N_3891,N_3724,N_3603);
or U3892 (N_3892,N_3639,N_3633);
xnor U3893 (N_3893,N_3751,N_3647);
nor U3894 (N_3894,N_3621,N_3623);
nor U3895 (N_3895,N_3682,N_3608);
nor U3896 (N_3896,N_3704,N_3745);
xor U3897 (N_3897,N_3624,N_3656);
nor U3898 (N_3898,N_3606,N_3741);
and U3899 (N_3899,N_3680,N_3691);
and U3900 (N_3900,N_3623,N_3692);
nor U3901 (N_3901,N_3701,N_3792);
nor U3902 (N_3902,N_3603,N_3670);
xor U3903 (N_3903,N_3616,N_3705);
nor U3904 (N_3904,N_3726,N_3602);
nor U3905 (N_3905,N_3795,N_3775);
xor U3906 (N_3906,N_3632,N_3622);
xnor U3907 (N_3907,N_3618,N_3606);
xnor U3908 (N_3908,N_3630,N_3750);
and U3909 (N_3909,N_3731,N_3624);
and U3910 (N_3910,N_3688,N_3696);
nor U3911 (N_3911,N_3799,N_3688);
nor U3912 (N_3912,N_3656,N_3737);
and U3913 (N_3913,N_3656,N_3761);
nand U3914 (N_3914,N_3772,N_3764);
or U3915 (N_3915,N_3649,N_3740);
and U3916 (N_3916,N_3722,N_3775);
and U3917 (N_3917,N_3725,N_3644);
nand U3918 (N_3918,N_3762,N_3616);
xor U3919 (N_3919,N_3674,N_3624);
or U3920 (N_3920,N_3634,N_3758);
xnor U3921 (N_3921,N_3688,N_3654);
xnor U3922 (N_3922,N_3781,N_3714);
and U3923 (N_3923,N_3669,N_3699);
nor U3924 (N_3924,N_3799,N_3697);
nor U3925 (N_3925,N_3606,N_3651);
nor U3926 (N_3926,N_3746,N_3710);
nor U3927 (N_3927,N_3630,N_3730);
nor U3928 (N_3928,N_3715,N_3718);
xnor U3929 (N_3929,N_3753,N_3706);
and U3930 (N_3930,N_3740,N_3748);
nand U3931 (N_3931,N_3665,N_3722);
and U3932 (N_3932,N_3732,N_3662);
nor U3933 (N_3933,N_3759,N_3799);
or U3934 (N_3934,N_3798,N_3779);
nor U3935 (N_3935,N_3625,N_3680);
nor U3936 (N_3936,N_3713,N_3778);
or U3937 (N_3937,N_3635,N_3782);
and U3938 (N_3938,N_3776,N_3610);
or U3939 (N_3939,N_3677,N_3704);
nand U3940 (N_3940,N_3780,N_3726);
nor U3941 (N_3941,N_3773,N_3628);
and U3942 (N_3942,N_3603,N_3651);
or U3943 (N_3943,N_3758,N_3717);
nand U3944 (N_3944,N_3787,N_3725);
or U3945 (N_3945,N_3744,N_3700);
or U3946 (N_3946,N_3710,N_3632);
and U3947 (N_3947,N_3654,N_3746);
and U3948 (N_3948,N_3605,N_3671);
nand U3949 (N_3949,N_3634,N_3612);
and U3950 (N_3950,N_3605,N_3729);
xor U3951 (N_3951,N_3749,N_3780);
xnor U3952 (N_3952,N_3642,N_3760);
nand U3953 (N_3953,N_3623,N_3735);
nand U3954 (N_3954,N_3617,N_3630);
nand U3955 (N_3955,N_3655,N_3631);
nand U3956 (N_3956,N_3722,N_3668);
and U3957 (N_3957,N_3781,N_3641);
nand U3958 (N_3958,N_3798,N_3668);
xnor U3959 (N_3959,N_3603,N_3689);
nand U3960 (N_3960,N_3702,N_3602);
nor U3961 (N_3961,N_3734,N_3689);
nor U3962 (N_3962,N_3698,N_3705);
xnor U3963 (N_3963,N_3632,N_3793);
xnor U3964 (N_3964,N_3717,N_3790);
xnor U3965 (N_3965,N_3667,N_3654);
xor U3966 (N_3966,N_3732,N_3770);
or U3967 (N_3967,N_3699,N_3773);
nand U3968 (N_3968,N_3783,N_3727);
nor U3969 (N_3969,N_3790,N_3793);
and U3970 (N_3970,N_3602,N_3712);
or U3971 (N_3971,N_3726,N_3768);
nand U3972 (N_3972,N_3702,N_3611);
and U3973 (N_3973,N_3635,N_3793);
or U3974 (N_3974,N_3605,N_3608);
or U3975 (N_3975,N_3677,N_3788);
and U3976 (N_3976,N_3722,N_3756);
or U3977 (N_3977,N_3705,N_3730);
nor U3978 (N_3978,N_3620,N_3735);
nor U3979 (N_3979,N_3795,N_3756);
nor U3980 (N_3980,N_3608,N_3767);
and U3981 (N_3981,N_3718,N_3708);
and U3982 (N_3982,N_3639,N_3733);
and U3983 (N_3983,N_3782,N_3709);
and U3984 (N_3984,N_3766,N_3661);
xor U3985 (N_3985,N_3603,N_3778);
nor U3986 (N_3986,N_3685,N_3789);
xnor U3987 (N_3987,N_3709,N_3665);
and U3988 (N_3988,N_3734,N_3799);
or U3989 (N_3989,N_3749,N_3750);
and U3990 (N_3990,N_3732,N_3787);
nor U3991 (N_3991,N_3612,N_3726);
xor U3992 (N_3992,N_3721,N_3712);
nor U3993 (N_3993,N_3674,N_3713);
or U3994 (N_3994,N_3765,N_3779);
nand U3995 (N_3995,N_3757,N_3684);
or U3996 (N_3996,N_3738,N_3732);
and U3997 (N_3997,N_3643,N_3777);
or U3998 (N_3998,N_3699,N_3759);
nand U3999 (N_3999,N_3651,N_3612);
nand U4000 (N_4000,N_3999,N_3809);
or U4001 (N_4001,N_3909,N_3963);
or U4002 (N_4002,N_3967,N_3848);
and U4003 (N_4003,N_3878,N_3859);
nand U4004 (N_4004,N_3853,N_3997);
nor U4005 (N_4005,N_3815,N_3883);
nor U4006 (N_4006,N_3956,N_3846);
nor U4007 (N_4007,N_3960,N_3904);
nor U4008 (N_4008,N_3869,N_3905);
nand U4009 (N_4009,N_3913,N_3924);
xor U4010 (N_4010,N_3941,N_3868);
nor U4011 (N_4011,N_3840,N_3977);
nor U4012 (N_4012,N_3887,N_3919);
nor U4013 (N_4013,N_3986,N_3979);
or U4014 (N_4014,N_3929,N_3942);
xor U4015 (N_4015,N_3871,N_3945);
or U4016 (N_4016,N_3981,N_3816);
or U4017 (N_4017,N_3818,N_3961);
nand U4018 (N_4018,N_3896,N_3988);
or U4019 (N_4019,N_3861,N_3824);
and U4020 (N_4020,N_3899,N_3827);
nand U4021 (N_4021,N_3870,N_3922);
xor U4022 (N_4022,N_3849,N_3806);
nand U4023 (N_4023,N_3978,N_3838);
or U4024 (N_4024,N_3923,N_3921);
xnor U4025 (N_4025,N_3947,N_3959);
xor U4026 (N_4026,N_3857,N_3898);
or U4027 (N_4027,N_3886,N_3937);
nand U4028 (N_4028,N_3835,N_3845);
nor U4029 (N_4029,N_3987,N_3800);
nor U4030 (N_4030,N_3889,N_3933);
or U4031 (N_4031,N_3864,N_3990);
nand U4032 (N_4032,N_3844,N_3943);
or U4033 (N_4033,N_3952,N_3865);
or U4034 (N_4034,N_3917,N_3993);
xnor U4035 (N_4035,N_3811,N_3821);
and U4036 (N_4036,N_3877,N_3953);
xor U4037 (N_4037,N_3955,N_3931);
or U4038 (N_4038,N_3927,N_3957);
xor U4039 (N_4039,N_3936,N_3969);
nor U4040 (N_4040,N_3879,N_3810);
nor U4041 (N_4041,N_3822,N_3949);
nand U4042 (N_4042,N_3855,N_3801);
or U4043 (N_4043,N_3926,N_3973);
xnor U4044 (N_4044,N_3964,N_3894);
or U4045 (N_4045,N_3895,N_3841);
xnor U4046 (N_4046,N_3954,N_3884);
nand U4047 (N_4047,N_3902,N_3828);
xor U4048 (N_4048,N_3836,N_3880);
and U4049 (N_4049,N_3834,N_3950);
nor U4050 (N_4050,N_3854,N_3995);
nor U4051 (N_4051,N_3819,N_3803);
and U4052 (N_4052,N_3860,N_3866);
nor U4053 (N_4053,N_3812,N_3872);
and U4054 (N_4054,N_3901,N_3984);
xnor U4055 (N_4055,N_3968,N_3831);
nand U4056 (N_4056,N_3826,N_3925);
xor U4057 (N_4057,N_3888,N_3862);
nor U4058 (N_4058,N_3948,N_3802);
or U4059 (N_4059,N_3971,N_3992);
nand U4060 (N_4060,N_3873,N_3946);
or U4061 (N_4061,N_3980,N_3970);
nor U4062 (N_4062,N_3874,N_3972);
nor U4063 (N_4063,N_3885,N_3911);
nand U4064 (N_4064,N_3897,N_3983);
nand U4065 (N_4065,N_3890,N_3918);
or U4066 (N_4066,N_3991,N_3938);
nor U4067 (N_4067,N_3935,N_3998);
nor U4068 (N_4068,N_3996,N_3944);
xor U4069 (N_4069,N_3814,N_3876);
xor U4070 (N_4070,N_3843,N_3832);
nor U4071 (N_4071,N_3804,N_3934);
nand U4072 (N_4072,N_3856,N_3908);
nor U4073 (N_4073,N_3975,N_3820);
and U4074 (N_4074,N_3842,N_3867);
nor U4075 (N_4075,N_3893,N_3976);
or U4076 (N_4076,N_3858,N_3966);
nor U4077 (N_4077,N_3982,N_3850);
nor U4078 (N_4078,N_3863,N_3823);
nand U4079 (N_4079,N_3833,N_3951);
and U4080 (N_4080,N_3875,N_3965);
nand U4081 (N_4081,N_3881,N_3932);
and U4082 (N_4082,N_3906,N_3910);
nand U4083 (N_4083,N_3807,N_3962);
nand U4084 (N_4084,N_3985,N_3808);
nor U4085 (N_4085,N_3830,N_3851);
and U4086 (N_4086,N_3891,N_3837);
nand U4087 (N_4087,N_3892,N_3916);
nor U4088 (N_4088,N_3914,N_3930);
xor U4089 (N_4089,N_3847,N_3817);
nor U4090 (N_4090,N_3928,N_3825);
or U4091 (N_4091,N_3852,N_3829);
and U4092 (N_4092,N_3839,N_3920);
or U4093 (N_4093,N_3939,N_3813);
and U4094 (N_4094,N_3912,N_3989);
xnor U4095 (N_4095,N_3994,N_3900);
and U4096 (N_4096,N_3903,N_3805);
or U4097 (N_4097,N_3974,N_3907);
xnor U4098 (N_4098,N_3882,N_3915);
nand U4099 (N_4099,N_3940,N_3958);
and U4100 (N_4100,N_3822,N_3870);
nand U4101 (N_4101,N_3952,N_3923);
nor U4102 (N_4102,N_3889,N_3977);
nand U4103 (N_4103,N_3957,N_3899);
and U4104 (N_4104,N_3855,N_3911);
and U4105 (N_4105,N_3835,N_3876);
xor U4106 (N_4106,N_3828,N_3944);
and U4107 (N_4107,N_3825,N_3834);
nor U4108 (N_4108,N_3922,N_3903);
nor U4109 (N_4109,N_3888,N_3884);
nand U4110 (N_4110,N_3939,N_3891);
xnor U4111 (N_4111,N_3889,N_3966);
nor U4112 (N_4112,N_3947,N_3885);
and U4113 (N_4113,N_3992,N_3893);
nor U4114 (N_4114,N_3850,N_3978);
nor U4115 (N_4115,N_3845,N_3818);
nand U4116 (N_4116,N_3804,N_3887);
nor U4117 (N_4117,N_3803,N_3809);
and U4118 (N_4118,N_3887,N_3935);
or U4119 (N_4119,N_3816,N_3889);
nor U4120 (N_4120,N_3997,N_3887);
nand U4121 (N_4121,N_3860,N_3885);
and U4122 (N_4122,N_3922,N_3900);
nor U4123 (N_4123,N_3913,N_3942);
or U4124 (N_4124,N_3828,N_3886);
xnor U4125 (N_4125,N_3887,N_3811);
and U4126 (N_4126,N_3872,N_3996);
xnor U4127 (N_4127,N_3982,N_3861);
and U4128 (N_4128,N_3913,N_3803);
nor U4129 (N_4129,N_3827,N_3923);
nand U4130 (N_4130,N_3869,N_3808);
nor U4131 (N_4131,N_3855,N_3937);
and U4132 (N_4132,N_3829,N_3837);
nand U4133 (N_4133,N_3892,N_3893);
and U4134 (N_4134,N_3830,N_3936);
nand U4135 (N_4135,N_3981,N_3996);
and U4136 (N_4136,N_3849,N_3891);
and U4137 (N_4137,N_3840,N_3994);
nand U4138 (N_4138,N_3973,N_3894);
and U4139 (N_4139,N_3917,N_3912);
or U4140 (N_4140,N_3867,N_3853);
nor U4141 (N_4141,N_3908,N_3948);
nor U4142 (N_4142,N_3817,N_3914);
xnor U4143 (N_4143,N_3975,N_3876);
or U4144 (N_4144,N_3902,N_3903);
nand U4145 (N_4145,N_3870,N_3982);
nand U4146 (N_4146,N_3861,N_3912);
and U4147 (N_4147,N_3966,N_3927);
xor U4148 (N_4148,N_3833,N_3941);
and U4149 (N_4149,N_3877,N_3952);
and U4150 (N_4150,N_3962,N_3853);
and U4151 (N_4151,N_3900,N_3995);
xor U4152 (N_4152,N_3853,N_3922);
nor U4153 (N_4153,N_3964,N_3921);
nor U4154 (N_4154,N_3808,N_3966);
or U4155 (N_4155,N_3846,N_3831);
or U4156 (N_4156,N_3992,N_3833);
and U4157 (N_4157,N_3913,N_3963);
xor U4158 (N_4158,N_3817,N_3974);
and U4159 (N_4159,N_3906,N_3884);
nand U4160 (N_4160,N_3844,N_3924);
and U4161 (N_4161,N_3942,N_3921);
xor U4162 (N_4162,N_3853,N_3924);
nand U4163 (N_4163,N_3891,N_3812);
nor U4164 (N_4164,N_3920,N_3913);
and U4165 (N_4165,N_3879,N_3921);
nand U4166 (N_4166,N_3880,N_3837);
or U4167 (N_4167,N_3920,N_3909);
nand U4168 (N_4168,N_3939,N_3833);
nand U4169 (N_4169,N_3934,N_3855);
nor U4170 (N_4170,N_3805,N_3987);
xnor U4171 (N_4171,N_3964,N_3906);
or U4172 (N_4172,N_3844,N_3931);
xnor U4173 (N_4173,N_3812,N_3818);
nor U4174 (N_4174,N_3969,N_3811);
nor U4175 (N_4175,N_3821,N_3882);
xor U4176 (N_4176,N_3801,N_3813);
xor U4177 (N_4177,N_3866,N_3915);
and U4178 (N_4178,N_3838,N_3996);
and U4179 (N_4179,N_3933,N_3944);
nand U4180 (N_4180,N_3971,N_3887);
nor U4181 (N_4181,N_3947,N_3913);
nor U4182 (N_4182,N_3865,N_3878);
or U4183 (N_4183,N_3892,N_3811);
or U4184 (N_4184,N_3801,N_3870);
nor U4185 (N_4185,N_3819,N_3993);
and U4186 (N_4186,N_3881,N_3974);
or U4187 (N_4187,N_3847,N_3904);
and U4188 (N_4188,N_3807,N_3936);
or U4189 (N_4189,N_3851,N_3952);
and U4190 (N_4190,N_3870,N_3837);
and U4191 (N_4191,N_3842,N_3884);
or U4192 (N_4192,N_3833,N_3817);
nor U4193 (N_4193,N_3933,N_3931);
or U4194 (N_4194,N_3929,N_3955);
nor U4195 (N_4195,N_3920,N_3896);
and U4196 (N_4196,N_3841,N_3902);
nor U4197 (N_4197,N_3849,N_3853);
xnor U4198 (N_4198,N_3970,N_3948);
or U4199 (N_4199,N_3931,N_3800);
nand U4200 (N_4200,N_4098,N_4023);
or U4201 (N_4201,N_4179,N_4134);
xnor U4202 (N_4202,N_4072,N_4198);
xnor U4203 (N_4203,N_4103,N_4114);
nor U4204 (N_4204,N_4142,N_4094);
nand U4205 (N_4205,N_4025,N_4045);
nor U4206 (N_4206,N_4050,N_4054);
xnor U4207 (N_4207,N_4136,N_4085);
nand U4208 (N_4208,N_4150,N_4010);
nand U4209 (N_4209,N_4173,N_4194);
or U4210 (N_4210,N_4124,N_4182);
and U4211 (N_4211,N_4158,N_4063);
xor U4212 (N_4212,N_4138,N_4057);
and U4213 (N_4213,N_4119,N_4191);
and U4214 (N_4214,N_4160,N_4051);
and U4215 (N_4215,N_4026,N_4192);
xnor U4216 (N_4216,N_4177,N_4180);
nand U4217 (N_4217,N_4126,N_4049);
nand U4218 (N_4218,N_4017,N_4147);
nand U4219 (N_4219,N_4083,N_4011);
nor U4220 (N_4220,N_4110,N_4084);
xnor U4221 (N_4221,N_4047,N_4044);
xor U4222 (N_4222,N_4022,N_4125);
nand U4223 (N_4223,N_4118,N_4028);
nor U4224 (N_4224,N_4154,N_4193);
nand U4225 (N_4225,N_4165,N_4184);
nor U4226 (N_4226,N_4031,N_4055);
nand U4227 (N_4227,N_4133,N_4037);
nand U4228 (N_4228,N_4157,N_4066);
xor U4229 (N_4229,N_4162,N_4129);
nand U4230 (N_4230,N_4121,N_4078);
or U4231 (N_4231,N_4088,N_4117);
nor U4232 (N_4232,N_4164,N_4016);
nor U4233 (N_4233,N_4123,N_4032);
nor U4234 (N_4234,N_4056,N_4145);
and U4235 (N_4235,N_4067,N_4082);
and U4236 (N_4236,N_4181,N_4012);
xnor U4237 (N_4237,N_4062,N_4195);
and U4238 (N_4238,N_4073,N_4090);
or U4239 (N_4239,N_4113,N_4116);
nor U4240 (N_4240,N_4105,N_4009);
nor U4241 (N_4241,N_4015,N_4036);
nand U4242 (N_4242,N_4167,N_4199);
or U4243 (N_4243,N_4058,N_4183);
nand U4244 (N_4244,N_4178,N_4127);
nor U4245 (N_4245,N_4153,N_4076);
or U4246 (N_4246,N_4106,N_4091);
nor U4247 (N_4247,N_4020,N_4108);
nand U4248 (N_4248,N_4107,N_4149);
nor U4249 (N_4249,N_4087,N_4131);
nand U4250 (N_4250,N_4111,N_4139);
xnor U4251 (N_4251,N_4143,N_4069);
nor U4252 (N_4252,N_4135,N_4163);
nor U4253 (N_4253,N_4052,N_4074);
nor U4254 (N_4254,N_4075,N_4166);
or U4255 (N_4255,N_4122,N_4109);
and U4256 (N_4256,N_4034,N_4132);
or U4257 (N_4257,N_4140,N_4099);
or U4258 (N_4258,N_4030,N_4169);
nand U4259 (N_4259,N_4128,N_4000);
nor U4260 (N_4260,N_4024,N_4080);
nand U4261 (N_4261,N_4019,N_4004);
and U4262 (N_4262,N_4185,N_4120);
nor U4263 (N_4263,N_4048,N_4071);
xnor U4264 (N_4264,N_4092,N_4104);
nor U4265 (N_4265,N_4041,N_4176);
or U4266 (N_4266,N_4159,N_4081);
and U4267 (N_4267,N_4102,N_4151);
nor U4268 (N_4268,N_4046,N_4170);
xnor U4269 (N_4269,N_4040,N_4130);
or U4270 (N_4270,N_4137,N_4175);
nand U4271 (N_4271,N_4141,N_4059);
or U4272 (N_4272,N_4171,N_4156);
xor U4273 (N_4273,N_4053,N_4027);
xor U4274 (N_4274,N_4039,N_4172);
nand U4275 (N_4275,N_4033,N_4003);
nand U4276 (N_4276,N_4196,N_4068);
or U4277 (N_4277,N_4144,N_4079);
xnor U4278 (N_4278,N_4021,N_4043);
nor U4279 (N_4279,N_4014,N_4064);
and U4280 (N_4280,N_4190,N_4008);
and U4281 (N_4281,N_4065,N_4174);
nand U4282 (N_4282,N_4005,N_4013);
and U4283 (N_4283,N_4096,N_4152);
and U4284 (N_4284,N_4060,N_4115);
and U4285 (N_4285,N_4086,N_4168);
xor U4286 (N_4286,N_4188,N_4018);
nand U4287 (N_4287,N_4038,N_4101);
or U4288 (N_4288,N_4029,N_4148);
nor U4289 (N_4289,N_4006,N_4095);
nand U4290 (N_4290,N_4197,N_4189);
or U4291 (N_4291,N_4093,N_4077);
nor U4292 (N_4292,N_4042,N_4146);
nand U4293 (N_4293,N_4061,N_4186);
nand U4294 (N_4294,N_4007,N_4089);
xnor U4295 (N_4295,N_4097,N_4001);
nand U4296 (N_4296,N_4070,N_4100);
nor U4297 (N_4297,N_4035,N_4112);
or U4298 (N_4298,N_4002,N_4155);
or U4299 (N_4299,N_4161,N_4187);
nor U4300 (N_4300,N_4069,N_4141);
and U4301 (N_4301,N_4163,N_4038);
xnor U4302 (N_4302,N_4105,N_4168);
nand U4303 (N_4303,N_4108,N_4167);
or U4304 (N_4304,N_4104,N_4061);
nand U4305 (N_4305,N_4088,N_4145);
nand U4306 (N_4306,N_4188,N_4196);
and U4307 (N_4307,N_4052,N_4170);
nand U4308 (N_4308,N_4155,N_4145);
and U4309 (N_4309,N_4157,N_4046);
or U4310 (N_4310,N_4081,N_4143);
or U4311 (N_4311,N_4186,N_4058);
nand U4312 (N_4312,N_4186,N_4090);
nor U4313 (N_4313,N_4175,N_4000);
nor U4314 (N_4314,N_4175,N_4120);
nand U4315 (N_4315,N_4110,N_4180);
nor U4316 (N_4316,N_4041,N_4097);
nand U4317 (N_4317,N_4067,N_4126);
or U4318 (N_4318,N_4037,N_4023);
and U4319 (N_4319,N_4160,N_4115);
nor U4320 (N_4320,N_4147,N_4189);
nand U4321 (N_4321,N_4021,N_4061);
xor U4322 (N_4322,N_4098,N_4142);
or U4323 (N_4323,N_4072,N_4112);
xnor U4324 (N_4324,N_4087,N_4151);
or U4325 (N_4325,N_4196,N_4164);
and U4326 (N_4326,N_4197,N_4016);
and U4327 (N_4327,N_4067,N_4006);
nand U4328 (N_4328,N_4180,N_4127);
or U4329 (N_4329,N_4183,N_4162);
and U4330 (N_4330,N_4047,N_4021);
and U4331 (N_4331,N_4069,N_4082);
xor U4332 (N_4332,N_4020,N_4054);
or U4333 (N_4333,N_4105,N_4070);
or U4334 (N_4334,N_4132,N_4139);
xor U4335 (N_4335,N_4060,N_4095);
or U4336 (N_4336,N_4192,N_4055);
xnor U4337 (N_4337,N_4100,N_4002);
xor U4338 (N_4338,N_4047,N_4197);
nand U4339 (N_4339,N_4168,N_4127);
xor U4340 (N_4340,N_4064,N_4180);
xor U4341 (N_4341,N_4038,N_4164);
nor U4342 (N_4342,N_4075,N_4047);
or U4343 (N_4343,N_4127,N_4090);
xnor U4344 (N_4344,N_4058,N_4075);
nor U4345 (N_4345,N_4007,N_4030);
or U4346 (N_4346,N_4037,N_4087);
xor U4347 (N_4347,N_4036,N_4025);
nor U4348 (N_4348,N_4055,N_4145);
nor U4349 (N_4349,N_4003,N_4008);
and U4350 (N_4350,N_4170,N_4068);
or U4351 (N_4351,N_4135,N_4043);
nor U4352 (N_4352,N_4114,N_4096);
nand U4353 (N_4353,N_4067,N_4083);
nor U4354 (N_4354,N_4100,N_4114);
nor U4355 (N_4355,N_4181,N_4077);
xor U4356 (N_4356,N_4019,N_4044);
nor U4357 (N_4357,N_4008,N_4076);
nor U4358 (N_4358,N_4040,N_4077);
or U4359 (N_4359,N_4098,N_4017);
or U4360 (N_4360,N_4109,N_4153);
xor U4361 (N_4361,N_4115,N_4168);
xnor U4362 (N_4362,N_4093,N_4080);
nor U4363 (N_4363,N_4146,N_4077);
or U4364 (N_4364,N_4073,N_4153);
nor U4365 (N_4365,N_4120,N_4164);
and U4366 (N_4366,N_4103,N_4176);
and U4367 (N_4367,N_4193,N_4047);
xor U4368 (N_4368,N_4192,N_4132);
xor U4369 (N_4369,N_4079,N_4193);
xnor U4370 (N_4370,N_4114,N_4147);
nor U4371 (N_4371,N_4187,N_4079);
nor U4372 (N_4372,N_4040,N_4148);
nand U4373 (N_4373,N_4125,N_4067);
nand U4374 (N_4374,N_4078,N_4061);
nor U4375 (N_4375,N_4048,N_4172);
xor U4376 (N_4376,N_4021,N_4092);
and U4377 (N_4377,N_4082,N_4073);
and U4378 (N_4378,N_4195,N_4098);
and U4379 (N_4379,N_4104,N_4127);
xnor U4380 (N_4380,N_4025,N_4181);
or U4381 (N_4381,N_4169,N_4158);
nor U4382 (N_4382,N_4176,N_4096);
nor U4383 (N_4383,N_4177,N_4054);
nand U4384 (N_4384,N_4107,N_4106);
nor U4385 (N_4385,N_4101,N_4152);
nor U4386 (N_4386,N_4140,N_4060);
xnor U4387 (N_4387,N_4168,N_4000);
or U4388 (N_4388,N_4102,N_4148);
and U4389 (N_4389,N_4152,N_4005);
nor U4390 (N_4390,N_4019,N_4076);
nand U4391 (N_4391,N_4047,N_4174);
or U4392 (N_4392,N_4009,N_4178);
xnor U4393 (N_4393,N_4011,N_4187);
nor U4394 (N_4394,N_4141,N_4177);
and U4395 (N_4395,N_4039,N_4146);
or U4396 (N_4396,N_4027,N_4040);
and U4397 (N_4397,N_4174,N_4186);
nand U4398 (N_4398,N_4176,N_4134);
nand U4399 (N_4399,N_4103,N_4172);
nor U4400 (N_4400,N_4384,N_4219);
or U4401 (N_4401,N_4261,N_4287);
or U4402 (N_4402,N_4388,N_4211);
nand U4403 (N_4403,N_4315,N_4340);
and U4404 (N_4404,N_4216,N_4396);
nor U4405 (N_4405,N_4209,N_4299);
xnor U4406 (N_4406,N_4372,N_4231);
and U4407 (N_4407,N_4376,N_4297);
xnor U4408 (N_4408,N_4381,N_4205);
nor U4409 (N_4409,N_4243,N_4227);
xnor U4410 (N_4410,N_4223,N_4336);
nor U4411 (N_4411,N_4329,N_4339);
xor U4412 (N_4412,N_4397,N_4322);
nor U4413 (N_4413,N_4343,N_4309);
and U4414 (N_4414,N_4253,N_4303);
or U4415 (N_4415,N_4352,N_4356);
xnor U4416 (N_4416,N_4290,N_4200);
nor U4417 (N_4417,N_4282,N_4232);
xnor U4418 (N_4418,N_4236,N_4327);
and U4419 (N_4419,N_4267,N_4370);
or U4420 (N_4420,N_4260,N_4398);
and U4421 (N_4421,N_4353,N_4344);
or U4422 (N_4422,N_4271,N_4318);
nor U4423 (N_4423,N_4366,N_4312);
or U4424 (N_4424,N_4331,N_4338);
nand U4425 (N_4425,N_4269,N_4291);
xnor U4426 (N_4426,N_4240,N_4298);
xor U4427 (N_4427,N_4214,N_4319);
nor U4428 (N_4428,N_4255,N_4239);
or U4429 (N_4429,N_4272,N_4302);
and U4430 (N_4430,N_4257,N_4306);
nand U4431 (N_4431,N_4391,N_4389);
and U4432 (N_4432,N_4235,N_4333);
and U4433 (N_4433,N_4348,N_4277);
xnor U4434 (N_4434,N_4278,N_4207);
xor U4435 (N_4435,N_4358,N_4259);
xor U4436 (N_4436,N_4347,N_4226);
and U4437 (N_4437,N_4307,N_4364);
or U4438 (N_4438,N_4201,N_4374);
nor U4439 (N_4439,N_4222,N_4279);
or U4440 (N_4440,N_4203,N_4301);
nor U4441 (N_4441,N_4317,N_4304);
and U4442 (N_4442,N_4218,N_4220);
and U4443 (N_4443,N_4288,N_4320);
xnor U4444 (N_4444,N_4354,N_4264);
nand U4445 (N_4445,N_4208,N_4215);
nand U4446 (N_4446,N_4258,N_4345);
or U4447 (N_4447,N_4386,N_4385);
nand U4448 (N_4448,N_4308,N_4270);
and U4449 (N_4449,N_4300,N_4229);
and U4450 (N_4450,N_4246,N_4275);
nand U4451 (N_4451,N_4276,N_4369);
and U4452 (N_4452,N_4292,N_4286);
nand U4453 (N_4453,N_4359,N_4395);
xnor U4454 (N_4454,N_4332,N_4375);
and U4455 (N_4455,N_4313,N_4305);
and U4456 (N_4456,N_4285,N_4378);
nor U4457 (N_4457,N_4252,N_4233);
nor U4458 (N_4458,N_4314,N_4393);
xnor U4459 (N_4459,N_4265,N_4311);
nand U4460 (N_4460,N_4392,N_4210);
xor U4461 (N_4461,N_4262,N_4373);
nor U4462 (N_4462,N_4365,N_4230);
or U4463 (N_4463,N_4310,N_4251);
or U4464 (N_4464,N_4284,N_4295);
nand U4465 (N_4465,N_4202,N_4249);
xor U4466 (N_4466,N_4296,N_4382);
or U4467 (N_4467,N_4204,N_4399);
nand U4468 (N_4468,N_4245,N_4324);
xor U4469 (N_4469,N_4247,N_4263);
and U4470 (N_4470,N_4293,N_4390);
nor U4471 (N_4471,N_4206,N_4351);
or U4472 (N_4472,N_4273,N_4221);
xnor U4473 (N_4473,N_4256,N_4361);
nor U4474 (N_4474,N_4321,N_4346);
nor U4475 (N_4475,N_4213,N_4377);
nor U4476 (N_4476,N_4250,N_4328);
nand U4477 (N_4477,N_4334,N_4362);
nand U4478 (N_4478,N_4316,N_4238);
and U4479 (N_4479,N_4248,N_4326);
or U4480 (N_4480,N_4212,N_4268);
nand U4481 (N_4481,N_4254,N_4281);
xnor U4482 (N_4482,N_4325,N_4234);
xor U4483 (N_4483,N_4323,N_4283);
xnor U4484 (N_4484,N_4349,N_4350);
xor U4485 (N_4485,N_4357,N_4274);
and U4486 (N_4486,N_4367,N_4394);
nand U4487 (N_4487,N_4241,N_4368);
nand U4488 (N_4488,N_4294,N_4266);
xnor U4489 (N_4489,N_4383,N_4224);
nand U4490 (N_4490,N_4242,N_4341);
nor U4491 (N_4491,N_4228,N_4280);
xnor U4492 (N_4492,N_4342,N_4355);
or U4493 (N_4493,N_4337,N_4379);
and U4494 (N_4494,N_4330,N_4244);
xor U4495 (N_4495,N_4217,N_4289);
nand U4496 (N_4496,N_4335,N_4237);
or U4497 (N_4497,N_4371,N_4225);
nor U4498 (N_4498,N_4387,N_4360);
nor U4499 (N_4499,N_4380,N_4363);
nor U4500 (N_4500,N_4350,N_4360);
and U4501 (N_4501,N_4281,N_4325);
xnor U4502 (N_4502,N_4281,N_4301);
and U4503 (N_4503,N_4369,N_4335);
or U4504 (N_4504,N_4353,N_4308);
or U4505 (N_4505,N_4250,N_4209);
nand U4506 (N_4506,N_4201,N_4379);
nor U4507 (N_4507,N_4278,N_4277);
or U4508 (N_4508,N_4300,N_4369);
or U4509 (N_4509,N_4259,N_4382);
nand U4510 (N_4510,N_4306,N_4260);
or U4511 (N_4511,N_4244,N_4231);
and U4512 (N_4512,N_4222,N_4226);
nor U4513 (N_4513,N_4398,N_4351);
nand U4514 (N_4514,N_4269,N_4217);
nor U4515 (N_4515,N_4383,N_4209);
and U4516 (N_4516,N_4331,N_4278);
xnor U4517 (N_4517,N_4271,N_4309);
nand U4518 (N_4518,N_4211,N_4301);
nand U4519 (N_4519,N_4394,N_4368);
nand U4520 (N_4520,N_4351,N_4332);
nor U4521 (N_4521,N_4201,N_4227);
nand U4522 (N_4522,N_4288,N_4265);
xor U4523 (N_4523,N_4258,N_4230);
nor U4524 (N_4524,N_4390,N_4351);
nand U4525 (N_4525,N_4241,N_4293);
nor U4526 (N_4526,N_4204,N_4263);
xnor U4527 (N_4527,N_4241,N_4304);
and U4528 (N_4528,N_4396,N_4260);
or U4529 (N_4529,N_4349,N_4385);
nand U4530 (N_4530,N_4267,N_4329);
xnor U4531 (N_4531,N_4260,N_4324);
nor U4532 (N_4532,N_4391,N_4211);
xnor U4533 (N_4533,N_4246,N_4258);
nand U4534 (N_4534,N_4266,N_4263);
nor U4535 (N_4535,N_4346,N_4305);
nand U4536 (N_4536,N_4200,N_4364);
or U4537 (N_4537,N_4326,N_4220);
nand U4538 (N_4538,N_4201,N_4231);
and U4539 (N_4539,N_4256,N_4208);
nand U4540 (N_4540,N_4386,N_4397);
nand U4541 (N_4541,N_4228,N_4324);
and U4542 (N_4542,N_4380,N_4234);
nand U4543 (N_4543,N_4235,N_4242);
nor U4544 (N_4544,N_4279,N_4305);
nand U4545 (N_4545,N_4357,N_4285);
nor U4546 (N_4546,N_4205,N_4259);
xor U4547 (N_4547,N_4215,N_4227);
xnor U4548 (N_4548,N_4276,N_4399);
nand U4549 (N_4549,N_4308,N_4278);
or U4550 (N_4550,N_4326,N_4337);
and U4551 (N_4551,N_4270,N_4390);
xnor U4552 (N_4552,N_4250,N_4359);
or U4553 (N_4553,N_4269,N_4349);
or U4554 (N_4554,N_4342,N_4271);
nor U4555 (N_4555,N_4215,N_4377);
nand U4556 (N_4556,N_4340,N_4252);
nor U4557 (N_4557,N_4244,N_4268);
or U4558 (N_4558,N_4287,N_4349);
nor U4559 (N_4559,N_4252,N_4322);
or U4560 (N_4560,N_4283,N_4317);
nand U4561 (N_4561,N_4346,N_4352);
and U4562 (N_4562,N_4238,N_4252);
xor U4563 (N_4563,N_4280,N_4227);
or U4564 (N_4564,N_4376,N_4315);
or U4565 (N_4565,N_4361,N_4340);
or U4566 (N_4566,N_4358,N_4355);
xor U4567 (N_4567,N_4335,N_4298);
nand U4568 (N_4568,N_4307,N_4347);
and U4569 (N_4569,N_4226,N_4374);
nand U4570 (N_4570,N_4373,N_4321);
xor U4571 (N_4571,N_4313,N_4367);
and U4572 (N_4572,N_4264,N_4209);
and U4573 (N_4573,N_4351,N_4361);
and U4574 (N_4574,N_4311,N_4241);
xor U4575 (N_4575,N_4341,N_4322);
nor U4576 (N_4576,N_4234,N_4227);
xor U4577 (N_4577,N_4261,N_4271);
or U4578 (N_4578,N_4309,N_4339);
xor U4579 (N_4579,N_4314,N_4356);
and U4580 (N_4580,N_4255,N_4389);
nor U4581 (N_4581,N_4342,N_4347);
xnor U4582 (N_4582,N_4284,N_4390);
xor U4583 (N_4583,N_4256,N_4236);
nor U4584 (N_4584,N_4339,N_4379);
nand U4585 (N_4585,N_4230,N_4387);
nand U4586 (N_4586,N_4219,N_4243);
and U4587 (N_4587,N_4337,N_4356);
nand U4588 (N_4588,N_4348,N_4385);
or U4589 (N_4589,N_4394,N_4279);
xor U4590 (N_4590,N_4295,N_4301);
nor U4591 (N_4591,N_4385,N_4282);
or U4592 (N_4592,N_4271,N_4354);
and U4593 (N_4593,N_4311,N_4292);
and U4594 (N_4594,N_4320,N_4341);
xor U4595 (N_4595,N_4352,N_4385);
nor U4596 (N_4596,N_4248,N_4328);
and U4597 (N_4597,N_4337,N_4264);
or U4598 (N_4598,N_4304,N_4285);
or U4599 (N_4599,N_4285,N_4324);
or U4600 (N_4600,N_4584,N_4410);
or U4601 (N_4601,N_4466,N_4592);
nand U4602 (N_4602,N_4510,N_4479);
and U4603 (N_4603,N_4418,N_4559);
and U4604 (N_4604,N_4441,N_4414);
or U4605 (N_4605,N_4405,N_4585);
xor U4606 (N_4606,N_4457,N_4459);
xor U4607 (N_4607,N_4516,N_4495);
xnor U4608 (N_4608,N_4534,N_4508);
nor U4609 (N_4609,N_4536,N_4589);
and U4610 (N_4610,N_4499,N_4404);
xnor U4611 (N_4611,N_4489,N_4474);
or U4612 (N_4612,N_4443,N_4408);
xnor U4613 (N_4613,N_4543,N_4452);
or U4614 (N_4614,N_4472,N_4554);
or U4615 (N_4615,N_4402,N_4556);
nand U4616 (N_4616,N_4531,N_4542);
or U4617 (N_4617,N_4519,N_4595);
nor U4618 (N_4618,N_4488,N_4540);
nor U4619 (N_4619,N_4447,N_4500);
or U4620 (N_4620,N_4409,N_4575);
xnor U4621 (N_4621,N_4497,N_4477);
xnor U4622 (N_4622,N_4442,N_4512);
or U4623 (N_4623,N_4415,N_4533);
or U4624 (N_4624,N_4434,N_4552);
and U4625 (N_4625,N_4530,N_4451);
xor U4626 (N_4626,N_4429,N_4563);
xnor U4627 (N_4627,N_4526,N_4566);
nand U4628 (N_4628,N_4453,N_4576);
nand U4629 (N_4629,N_4524,N_4440);
and U4630 (N_4630,N_4427,N_4445);
xnor U4631 (N_4631,N_4511,N_4550);
nand U4632 (N_4632,N_4549,N_4527);
nor U4633 (N_4633,N_4564,N_4528);
and U4634 (N_4634,N_4432,N_4590);
and U4635 (N_4635,N_4560,N_4487);
or U4636 (N_4636,N_4401,N_4450);
and U4637 (N_4637,N_4422,N_4598);
or U4638 (N_4638,N_4503,N_4517);
and U4639 (N_4639,N_4426,N_4596);
and U4640 (N_4640,N_4496,N_4423);
xor U4641 (N_4641,N_4593,N_4523);
xor U4642 (N_4642,N_4514,N_4455);
nand U4643 (N_4643,N_4521,N_4518);
nor U4644 (N_4644,N_4562,N_4412);
xor U4645 (N_4645,N_4492,N_4509);
xnor U4646 (N_4646,N_4544,N_4465);
nand U4647 (N_4647,N_4400,N_4435);
or U4648 (N_4648,N_4532,N_4431);
and U4649 (N_4649,N_4557,N_4491);
nand U4650 (N_4650,N_4444,N_4574);
nand U4651 (N_4651,N_4490,N_4437);
nand U4652 (N_4652,N_4476,N_4506);
nor U4653 (N_4653,N_4541,N_4546);
nor U4654 (N_4654,N_4458,N_4580);
xnor U4655 (N_4655,N_4416,N_4480);
or U4656 (N_4656,N_4498,N_4545);
xor U4657 (N_4657,N_4504,N_4565);
nor U4658 (N_4658,N_4470,N_4473);
xor U4659 (N_4659,N_4425,N_4411);
and U4660 (N_4660,N_4471,N_4483);
xor U4661 (N_4661,N_4421,N_4591);
and U4662 (N_4662,N_4553,N_4529);
nor U4663 (N_4663,N_4581,N_4555);
nand U4664 (N_4664,N_4484,N_4558);
xor U4665 (N_4665,N_4462,N_4403);
and U4666 (N_4666,N_4494,N_4597);
nor U4667 (N_4667,N_4424,N_4569);
nand U4668 (N_4668,N_4573,N_4482);
nor U4669 (N_4669,N_4485,N_4467);
nand U4670 (N_4670,N_4588,N_4433);
nor U4671 (N_4671,N_4561,N_4539);
or U4672 (N_4672,N_4525,N_4428);
and U4673 (N_4673,N_4599,N_4582);
and U4674 (N_4674,N_4478,N_4413);
nand U4675 (N_4675,N_4436,N_4449);
and U4676 (N_4676,N_4448,N_4535);
nor U4677 (N_4677,N_4572,N_4502);
or U4678 (N_4678,N_4481,N_4501);
nand U4679 (N_4679,N_4417,N_4430);
xnor U4680 (N_4680,N_4548,N_4505);
or U4681 (N_4681,N_4570,N_4551);
nor U4682 (N_4682,N_4469,N_4583);
and U4683 (N_4683,N_4464,N_4507);
xnor U4684 (N_4684,N_4438,N_4568);
nand U4685 (N_4685,N_4567,N_4579);
nand U4686 (N_4686,N_4406,N_4493);
and U4687 (N_4687,N_4419,N_4513);
or U4688 (N_4688,N_4486,N_4439);
nand U4689 (N_4689,N_4547,N_4420);
and U4690 (N_4690,N_4461,N_4520);
and U4691 (N_4691,N_4538,N_4522);
and U4692 (N_4692,N_4515,N_4407);
nor U4693 (N_4693,N_4463,N_4577);
nor U4694 (N_4694,N_4456,N_4475);
and U4695 (N_4695,N_4460,N_4594);
nor U4696 (N_4696,N_4446,N_4537);
or U4697 (N_4697,N_4454,N_4586);
xor U4698 (N_4698,N_4571,N_4587);
or U4699 (N_4699,N_4578,N_4468);
nor U4700 (N_4700,N_4442,N_4538);
xor U4701 (N_4701,N_4427,N_4440);
nor U4702 (N_4702,N_4492,N_4595);
and U4703 (N_4703,N_4475,N_4447);
or U4704 (N_4704,N_4528,N_4469);
or U4705 (N_4705,N_4400,N_4520);
or U4706 (N_4706,N_4583,N_4404);
or U4707 (N_4707,N_4530,N_4496);
xnor U4708 (N_4708,N_4446,N_4410);
or U4709 (N_4709,N_4577,N_4439);
nor U4710 (N_4710,N_4551,N_4492);
or U4711 (N_4711,N_4506,N_4442);
or U4712 (N_4712,N_4480,N_4578);
or U4713 (N_4713,N_4417,N_4414);
nand U4714 (N_4714,N_4593,N_4504);
nor U4715 (N_4715,N_4516,N_4494);
or U4716 (N_4716,N_4597,N_4404);
nor U4717 (N_4717,N_4430,N_4565);
xor U4718 (N_4718,N_4556,N_4511);
or U4719 (N_4719,N_4426,N_4571);
xor U4720 (N_4720,N_4409,N_4468);
nand U4721 (N_4721,N_4513,N_4505);
nor U4722 (N_4722,N_4414,N_4420);
nand U4723 (N_4723,N_4434,N_4522);
xor U4724 (N_4724,N_4544,N_4561);
nor U4725 (N_4725,N_4430,N_4547);
nor U4726 (N_4726,N_4507,N_4425);
or U4727 (N_4727,N_4438,N_4559);
and U4728 (N_4728,N_4491,N_4511);
nor U4729 (N_4729,N_4563,N_4517);
nand U4730 (N_4730,N_4482,N_4508);
and U4731 (N_4731,N_4401,N_4508);
or U4732 (N_4732,N_4459,N_4489);
xor U4733 (N_4733,N_4581,N_4560);
xnor U4734 (N_4734,N_4542,N_4535);
and U4735 (N_4735,N_4424,N_4475);
xnor U4736 (N_4736,N_4547,N_4520);
xor U4737 (N_4737,N_4574,N_4430);
or U4738 (N_4738,N_4446,N_4571);
and U4739 (N_4739,N_4404,N_4506);
or U4740 (N_4740,N_4468,N_4540);
or U4741 (N_4741,N_4409,N_4594);
nand U4742 (N_4742,N_4541,N_4524);
or U4743 (N_4743,N_4578,N_4427);
nand U4744 (N_4744,N_4588,N_4569);
nor U4745 (N_4745,N_4533,N_4405);
xnor U4746 (N_4746,N_4541,N_4594);
nor U4747 (N_4747,N_4457,N_4511);
and U4748 (N_4748,N_4526,N_4494);
nand U4749 (N_4749,N_4493,N_4484);
xor U4750 (N_4750,N_4590,N_4585);
and U4751 (N_4751,N_4545,N_4567);
nand U4752 (N_4752,N_4500,N_4468);
or U4753 (N_4753,N_4514,N_4414);
xnor U4754 (N_4754,N_4403,N_4412);
nor U4755 (N_4755,N_4562,N_4420);
xor U4756 (N_4756,N_4412,N_4536);
and U4757 (N_4757,N_4595,N_4407);
nand U4758 (N_4758,N_4542,N_4586);
nor U4759 (N_4759,N_4422,N_4511);
or U4760 (N_4760,N_4519,N_4539);
nor U4761 (N_4761,N_4569,N_4592);
nand U4762 (N_4762,N_4535,N_4451);
nor U4763 (N_4763,N_4461,N_4425);
and U4764 (N_4764,N_4516,N_4508);
nand U4765 (N_4765,N_4478,N_4592);
nand U4766 (N_4766,N_4499,N_4478);
nor U4767 (N_4767,N_4419,N_4434);
xor U4768 (N_4768,N_4551,N_4438);
xor U4769 (N_4769,N_4575,N_4446);
xnor U4770 (N_4770,N_4533,N_4445);
xor U4771 (N_4771,N_4447,N_4508);
or U4772 (N_4772,N_4539,N_4466);
nor U4773 (N_4773,N_4553,N_4490);
and U4774 (N_4774,N_4424,N_4561);
and U4775 (N_4775,N_4517,N_4573);
and U4776 (N_4776,N_4537,N_4405);
and U4777 (N_4777,N_4553,N_4415);
xor U4778 (N_4778,N_4578,N_4474);
nor U4779 (N_4779,N_4593,N_4475);
and U4780 (N_4780,N_4406,N_4592);
nor U4781 (N_4781,N_4506,N_4419);
nand U4782 (N_4782,N_4485,N_4507);
xor U4783 (N_4783,N_4582,N_4508);
nand U4784 (N_4784,N_4445,N_4554);
xor U4785 (N_4785,N_4419,N_4548);
xnor U4786 (N_4786,N_4504,N_4479);
xnor U4787 (N_4787,N_4577,N_4428);
and U4788 (N_4788,N_4491,N_4425);
and U4789 (N_4789,N_4595,N_4542);
nor U4790 (N_4790,N_4417,N_4431);
or U4791 (N_4791,N_4599,N_4532);
nor U4792 (N_4792,N_4531,N_4572);
or U4793 (N_4793,N_4524,N_4599);
or U4794 (N_4794,N_4428,N_4402);
nor U4795 (N_4795,N_4405,N_4579);
nand U4796 (N_4796,N_4404,N_4468);
nor U4797 (N_4797,N_4436,N_4509);
xnor U4798 (N_4798,N_4482,N_4569);
and U4799 (N_4799,N_4449,N_4555);
or U4800 (N_4800,N_4665,N_4611);
xnor U4801 (N_4801,N_4663,N_4798);
nor U4802 (N_4802,N_4741,N_4732);
nand U4803 (N_4803,N_4751,N_4729);
nand U4804 (N_4804,N_4627,N_4637);
nor U4805 (N_4805,N_4670,N_4648);
xor U4806 (N_4806,N_4768,N_4685);
and U4807 (N_4807,N_4767,N_4765);
or U4808 (N_4808,N_4789,N_4695);
and U4809 (N_4809,N_4702,N_4677);
or U4810 (N_4810,N_4701,N_4600);
nand U4811 (N_4811,N_4620,N_4615);
and U4812 (N_4812,N_4649,N_4784);
or U4813 (N_4813,N_4775,N_4779);
nor U4814 (N_4814,N_4740,N_4721);
nor U4815 (N_4815,N_4745,N_4681);
and U4816 (N_4816,N_4763,N_4796);
nor U4817 (N_4817,N_4679,N_4684);
or U4818 (N_4818,N_4749,N_4601);
xor U4819 (N_4819,N_4706,N_4633);
xnor U4820 (N_4820,N_4756,N_4638);
nor U4821 (N_4821,N_4658,N_4748);
xor U4822 (N_4822,N_4641,N_4647);
or U4823 (N_4823,N_4672,N_4696);
nor U4824 (N_4824,N_4755,N_4776);
and U4825 (N_4825,N_4608,N_4698);
nor U4826 (N_4826,N_4709,N_4643);
nand U4827 (N_4827,N_4625,N_4668);
and U4828 (N_4828,N_4712,N_4640);
or U4829 (N_4829,N_4752,N_4703);
and U4830 (N_4830,N_4735,N_4726);
nor U4831 (N_4831,N_4799,N_4780);
xor U4832 (N_4832,N_4682,N_4715);
or U4833 (N_4833,N_4656,N_4705);
xor U4834 (N_4834,N_4666,N_4753);
nor U4835 (N_4835,N_4700,N_4607);
or U4836 (N_4836,N_4609,N_4713);
or U4837 (N_4837,N_4687,N_4739);
nand U4838 (N_4838,N_4619,N_4688);
nand U4839 (N_4839,N_4629,N_4782);
xor U4840 (N_4840,N_4731,N_4602);
xor U4841 (N_4841,N_4714,N_4655);
and U4842 (N_4842,N_4664,N_4686);
or U4843 (N_4843,N_4628,N_4720);
and U4844 (N_4844,N_4635,N_4614);
nor U4845 (N_4845,N_4764,N_4758);
xnor U4846 (N_4846,N_4777,N_4722);
nor U4847 (N_4847,N_4719,N_4630);
nor U4848 (N_4848,N_4654,N_4730);
and U4849 (N_4849,N_4623,N_4787);
nor U4850 (N_4850,N_4744,N_4667);
xor U4851 (N_4851,N_4728,N_4645);
nand U4852 (N_4852,N_4785,N_4636);
or U4853 (N_4853,N_4788,N_4691);
nand U4854 (N_4854,N_4644,N_4725);
or U4855 (N_4855,N_4792,N_4651);
and U4856 (N_4856,N_4708,N_4727);
and U4857 (N_4857,N_4653,N_4738);
or U4858 (N_4858,N_4692,N_4772);
or U4859 (N_4859,N_4761,N_4642);
nor U4860 (N_4860,N_4657,N_4759);
xor U4861 (N_4861,N_4734,N_4716);
or U4862 (N_4862,N_4631,N_4659);
nand U4863 (N_4863,N_4791,N_4786);
nor U4864 (N_4864,N_4757,N_4742);
nand U4865 (N_4865,N_4604,N_4634);
xnor U4866 (N_4866,N_4613,N_4724);
or U4867 (N_4867,N_4718,N_4746);
nand U4868 (N_4868,N_4697,N_4676);
and U4869 (N_4869,N_4610,N_4603);
and U4870 (N_4870,N_4710,N_4773);
or U4871 (N_4871,N_4618,N_4778);
nor U4872 (N_4872,N_4795,N_4671);
nand U4873 (N_4873,N_4673,N_4790);
nor U4874 (N_4874,N_4661,N_4704);
nand U4875 (N_4875,N_4617,N_4605);
and U4876 (N_4876,N_4793,N_4771);
and U4877 (N_4877,N_4639,N_4646);
xor U4878 (N_4878,N_4689,N_4675);
and U4879 (N_4879,N_4683,N_4774);
or U4880 (N_4880,N_4766,N_4769);
and U4881 (N_4881,N_4674,N_4762);
and U4882 (N_4882,N_4626,N_4717);
and U4883 (N_4883,N_4699,N_4612);
xnor U4884 (N_4884,N_4662,N_4606);
xor U4885 (N_4885,N_4750,N_4707);
nand U4886 (N_4886,N_4737,N_4783);
xnor U4887 (N_4887,N_4660,N_4678);
nand U4888 (N_4888,N_4624,N_4743);
and U4889 (N_4889,N_4622,N_4760);
and U4890 (N_4890,N_4680,N_4652);
xnor U4891 (N_4891,N_4797,N_4723);
or U4892 (N_4892,N_4711,N_4650);
xor U4893 (N_4893,N_4616,N_4794);
nor U4894 (N_4894,N_4621,N_4690);
and U4895 (N_4895,N_4693,N_4694);
or U4896 (N_4896,N_4736,N_4770);
nor U4897 (N_4897,N_4747,N_4669);
xor U4898 (N_4898,N_4754,N_4781);
xor U4899 (N_4899,N_4733,N_4632);
nor U4900 (N_4900,N_4662,N_4710);
nor U4901 (N_4901,N_4605,N_4654);
nor U4902 (N_4902,N_4753,N_4775);
or U4903 (N_4903,N_4704,N_4615);
or U4904 (N_4904,N_4613,N_4692);
nor U4905 (N_4905,N_4691,N_4680);
and U4906 (N_4906,N_4788,N_4794);
and U4907 (N_4907,N_4653,N_4715);
and U4908 (N_4908,N_4780,N_4788);
nor U4909 (N_4909,N_4733,N_4615);
xnor U4910 (N_4910,N_4692,N_4686);
nand U4911 (N_4911,N_4685,N_4798);
or U4912 (N_4912,N_4681,N_4601);
nand U4913 (N_4913,N_4789,N_4607);
xnor U4914 (N_4914,N_4686,N_4793);
nand U4915 (N_4915,N_4638,N_4647);
or U4916 (N_4916,N_4779,N_4692);
xnor U4917 (N_4917,N_4644,N_4686);
xor U4918 (N_4918,N_4689,N_4705);
nand U4919 (N_4919,N_4608,N_4691);
and U4920 (N_4920,N_4762,N_4689);
xor U4921 (N_4921,N_4707,N_4666);
nor U4922 (N_4922,N_4665,N_4750);
or U4923 (N_4923,N_4604,N_4775);
nor U4924 (N_4924,N_4710,N_4793);
and U4925 (N_4925,N_4795,N_4712);
xnor U4926 (N_4926,N_4659,N_4695);
nor U4927 (N_4927,N_4692,N_4786);
or U4928 (N_4928,N_4750,N_4658);
xor U4929 (N_4929,N_4783,N_4605);
or U4930 (N_4930,N_4654,N_4677);
and U4931 (N_4931,N_4636,N_4738);
nand U4932 (N_4932,N_4609,N_4765);
nor U4933 (N_4933,N_4667,N_4677);
xor U4934 (N_4934,N_4736,N_4699);
xor U4935 (N_4935,N_4680,N_4778);
nand U4936 (N_4936,N_4680,N_4620);
or U4937 (N_4937,N_4714,N_4683);
or U4938 (N_4938,N_4684,N_4644);
or U4939 (N_4939,N_4724,N_4735);
nand U4940 (N_4940,N_4778,N_4692);
nor U4941 (N_4941,N_4718,N_4661);
or U4942 (N_4942,N_4753,N_4645);
nor U4943 (N_4943,N_4784,N_4712);
xor U4944 (N_4944,N_4789,N_4719);
nor U4945 (N_4945,N_4667,N_4752);
xnor U4946 (N_4946,N_4622,N_4792);
xor U4947 (N_4947,N_4624,N_4784);
or U4948 (N_4948,N_4668,N_4720);
xnor U4949 (N_4949,N_4758,N_4791);
xnor U4950 (N_4950,N_4777,N_4753);
or U4951 (N_4951,N_4643,N_4698);
nand U4952 (N_4952,N_4644,N_4753);
xor U4953 (N_4953,N_4751,N_4690);
nand U4954 (N_4954,N_4752,N_4641);
nor U4955 (N_4955,N_4784,N_4614);
nand U4956 (N_4956,N_4746,N_4790);
or U4957 (N_4957,N_4735,N_4623);
or U4958 (N_4958,N_4749,N_4713);
and U4959 (N_4959,N_4746,N_4645);
and U4960 (N_4960,N_4790,N_4743);
or U4961 (N_4961,N_4711,N_4795);
nor U4962 (N_4962,N_4694,N_4655);
xor U4963 (N_4963,N_4623,N_4783);
nor U4964 (N_4964,N_4680,N_4782);
or U4965 (N_4965,N_4779,N_4622);
and U4966 (N_4966,N_4747,N_4681);
and U4967 (N_4967,N_4746,N_4772);
nor U4968 (N_4968,N_4792,N_4625);
or U4969 (N_4969,N_4645,N_4656);
xor U4970 (N_4970,N_4657,N_4671);
nor U4971 (N_4971,N_4794,N_4700);
or U4972 (N_4972,N_4746,N_4619);
nor U4973 (N_4973,N_4701,N_4767);
xor U4974 (N_4974,N_4781,N_4749);
or U4975 (N_4975,N_4756,N_4671);
nand U4976 (N_4976,N_4679,N_4795);
nand U4977 (N_4977,N_4656,N_4788);
nor U4978 (N_4978,N_4756,N_4743);
nand U4979 (N_4979,N_4762,N_4732);
nand U4980 (N_4980,N_4633,N_4677);
nand U4981 (N_4981,N_4667,N_4670);
xor U4982 (N_4982,N_4661,N_4792);
xor U4983 (N_4983,N_4617,N_4724);
xnor U4984 (N_4984,N_4794,N_4799);
and U4985 (N_4985,N_4797,N_4664);
xor U4986 (N_4986,N_4689,N_4707);
and U4987 (N_4987,N_4663,N_4780);
and U4988 (N_4988,N_4639,N_4626);
and U4989 (N_4989,N_4758,N_4760);
xnor U4990 (N_4990,N_4766,N_4654);
or U4991 (N_4991,N_4762,N_4601);
and U4992 (N_4992,N_4714,N_4766);
xor U4993 (N_4993,N_4664,N_4656);
and U4994 (N_4994,N_4723,N_4644);
and U4995 (N_4995,N_4730,N_4635);
xor U4996 (N_4996,N_4611,N_4694);
and U4997 (N_4997,N_4706,N_4766);
nand U4998 (N_4998,N_4753,N_4707);
nor U4999 (N_4999,N_4733,N_4697);
and U5000 (N_5000,N_4921,N_4910);
or U5001 (N_5001,N_4934,N_4919);
and U5002 (N_5002,N_4927,N_4855);
nor U5003 (N_5003,N_4998,N_4994);
and U5004 (N_5004,N_4899,N_4966);
nand U5005 (N_5005,N_4871,N_4961);
and U5006 (N_5006,N_4814,N_4918);
xor U5007 (N_5007,N_4864,N_4977);
xor U5008 (N_5008,N_4817,N_4876);
xnor U5009 (N_5009,N_4945,N_4852);
nor U5010 (N_5010,N_4965,N_4924);
nor U5011 (N_5011,N_4987,N_4922);
or U5012 (N_5012,N_4898,N_4807);
or U5013 (N_5013,N_4854,N_4951);
nor U5014 (N_5014,N_4949,N_4908);
nand U5015 (N_5015,N_4978,N_4912);
nor U5016 (N_5016,N_4818,N_4816);
nand U5017 (N_5017,N_4835,N_4942);
and U5018 (N_5018,N_4810,N_4941);
xor U5019 (N_5019,N_4888,N_4939);
xor U5020 (N_5020,N_4878,N_4819);
xor U5021 (N_5021,N_4893,N_4901);
nor U5022 (N_5022,N_4986,N_4857);
nor U5023 (N_5023,N_4874,N_4952);
xor U5024 (N_5024,N_4999,N_4859);
nand U5025 (N_5025,N_4851,N_4950);
xor U5026 (N_5026,N_4838,N_4823);
or U5027 (N_5027,N_4970,N_4873);
or U5028 (N_5028,N_4809,N_4868);
and U5029 (N_5029,N_4875,N_4937);
or U5030 (N_5030,N_4828,N_4897);
and U5031 (N_5031,N_4806,N_4825);
nor U5032 (N_5032,N_4991,N_4968);
nor U5033 (N_5033,N_4803,N_4920);
or U5034 (N_5034,N_4836,N_4933);
or U5035 (N_5035,N_4982,N_4971);
xnor U5036 (N_5036,N_4895,N_4954);
nor U5037 (N_5037,N_4929,N_4953);
nand U5038 (N_5038,N_4904,N_4846);
or U5039 (N_5039,N_4869,N_4858);
and U5040 (N_5040,N_4867,N_4957);
or U5041 (N_5041,N_4903,N_4879);
xnor U5042 (N_5042,N_4902,N_4894);
xor U5043 (N_5043,N_4990,N_4975);
or U5044 (N_5044,N_4829,N_4995);
xor U5045 (N_5045,N_4930,N_4989);
nor U5046 (N_5046,N_4905,N_4863);
or U5047 (N_5047,N_4800,N_4860);
nor U5048 (N_5048,N_4805,N_4972);
or U5049 (N_5049,N_4997,N_4808);
nand U5050 (N_5050,N_4946,N_4911);
nand U5051 (N_5051,N_4812,N_4958);
and U5052 (N_5052,N_4947,N_4880);
and U5053 (N_5053,N_4960,N_4843);
nand U5054 (N_5054,N_4913,N_4827);
and U5055 (N_5055,N_4882,N_4955);
xor U5056 (N_5056,N_4931,N_4916);
and U5057 (N_5057,N_4820,N_4821);
xor U5058 (N_5058,N_4847,N_4861);
nand U5059 (N_5059,N_4872,N_4865);
and U5060 (N_5060,N_4962,N_4943);
xnor U5061 (N_5061,N_4884,N_4907);
xnor U5062 (N_5062,N_4974,N_4938);
or U5063 (N_5063,N_4923,N_4906);
and U5064 (N_5064,N_4900,N_4935);
or U5065 (N_5065,N_4956,N_4944);
nand U5066 (N_5066,N_4926,N_4862);
nand U5067 (N_5067,N_4885,N_4849);
and U5068 (N_5068,N_4841,N_4896);
and U5069 (N_5069,N_4985,N_4889);
or U5070 (N_5070,N_4964,N_4840);
and U5071 (N_5071,N_4996,N_4967);
xor U5072 (N_5072,N_4973,N_4881);
or U5073 (N_5073,N_4940,N_4932);
and U5074 (N_5074,N_4815,N_4976);
or U5075 (N_5075,N_4870,N_4984);
or U5076 (N_5076,N_4936,N_4917);
nand U5077 (N_5077,N_4909,N_4981);
or U5078 (N_5078,N_4811,N_4992);
or U5079 (N_5079,N_4833,N_4831);
or U5080 (N_5080,N_4928,N_4988);
and U5081 (N_5081,N_4883,N_4844);
and U5082 (N_5082,N_4813,N_4850);
nor U5083 (N_5083,N_4832,N_4834);
nor U5084 (N_5084,N_4969,N_4822);
and U5085 (N_5085,N_4891,N_4804);
and U5086 (N_5086,N_4842,N_4826);
xor U5087 (N_5087,N_4979,N_4963);
nand U5088 (N_5088,N_4959,N_4824);
and U5089 (N_5089,N_4914,N_4983);
and U5090 (N_5090,N_4925,N_4877);
nor U5091 (N_5091,N_4890,N_4839);
nand U5092 (N_5092,N_4915,N_4892);
or U5093 (N_5093,N_4837,N_4848);
nor U5094 (N_5094,N_4830,N_4856);
and U5095 (N_5095,N_4886,N_4980);
xnor U5096 (N_5096,N_4866,N_4845);
nor U5097 (N_5097,N_4887,N_4853);
nand U5098 (N_5098,N_4802,N_4993);
or U5099 (N_5099,N_4801,N_4948);
or U5100 (N_5100,N_4993,N_4914);
xnor U5101 (N_5101,N_4913,N_4987);
nor U5102 (N_5102,N_4815,N_4954);
or U5103 (N_5103,N_4938,N_4854);
nor U5104 (N_5104,N_4951,N_4835);
nor U5105 (N_5105,N_4832,N_4845);
nand U5106 (N_5106,N_4898,N_4914);
or U5107 (N_5107,N_4972,N_4874);
or U5108 (N_5108,N_4890,N_4842);
or U5109 (N_5109,N_4818,N_4801);
nor U5110 (N_5110,N_4856,N_4887);
xor U5111 (N_5111,N_4852,N_4935);
nor U5112 (N_5112,N_4948,N_4857);
or U5113 (N_5113,N_4826,N_4994);
nand U5114 (N_5114,N_4907,N_4863);
nor U5115 (N_5115,N_4825,N_4954);
xnor U5116 (N_5116,N_4851,N_4810);
xor U5117 (N_5117,N_4889,N_4974);
xor U5118 (N_5118,N_4996,N_4802);
xor U5119 (N_5119,N_4980,N_4842);
xor U5120 (N_5120,N_4835,N_4836);
xnor U5121 (N_5121,N_4903,N_4989);
nor U5122 (N_5122,N_4841,N_4977);
nand U5123 (N_5123,N_4929,N_4825);
nor U5124 (N_5124,N_4979,N_4966);
nor U5125 (N_5125,N_4892,N_4809);
xnor U5126 (N_5126,N_4933,N_4864);
xnor U5127 (N_5127,N_4980,N_4923);
nand U5128 (N_5128,N_4971,N_4837);
and U5129 (N_5129,N_4933,N_4994);
nor U5130 (N_5130,N_4955,N_4906);
xor U5131 (N_5131,N_4979,N_4816);
nand U5132 (N_5132,N_4831,N_4946);
nand U5133 (N_5133,N_4970,N_4909);
nor U5134 (N_5134,N_4861,N_4873);
nor U5135 (N_5135,N_4892,N_4975);
xor U5136 (N_5136,N_4895,N_4917);
nand U5137 (N_5137,N_4861,N_4818);
xnor U5138 (N_5138,N_4919,N_4959);
or U5139 (N_5139,N_4902,N_4805);
and U5140 (N_5140,N_4984,N_4824);
nor U5141 (N_5141,N_4906,N_4838);
xor U5142 (N_5142,N_4886,N_4880);
and U5143 (N_5143,N_4861,N_4903);
xnor U5144 (N_5144,N_4911,N_4992);
nor U5145 (N_5145,N_4834,N_4823);
nor U5146 (N_5146,N_4876,N_4818);
xnor U5147 (N_5147,N_4977,N_4800);
nand U5148 (N_5148,N_4917,N_4905);
xor U5149 (N_5149,N_4961,N_4852);
and U5150 (N_5150,N_4930,N_4993);
or U5151 (N_5151,N_4945,N_4942);
nor U5152 (N_5152,N_4971,N_4827);
and U5153 (N_5153,N_4893,N_4934);
nor U5154 (N_5154,N_4864,N_4986);
nand U5155 (N_5155,N_4861,N_4905);
or U5156 (N_5156,N_4929,N_4893);
and U5157 (N_5157,N_4879,N_4826);
and U5158 (N_5158,N_4872,N_4927);
and U5159 (N_5159,N_4937,N_4879);
nand U5160 (N_5160,N_4936,N_4903);
nand U5161 (N_5161,N_4969,N_4876);
or U5162 (N_5162,N_4804,N_4993);
nor U5163 (N_5163,N_4893,N_4882);
nand U5164 (N_5164,N_4914,N_4916);
or U5165 (N_5165,N_4911,N_4880);
nand U5166 (N_5166,N_4809,N_4874);
and U5167 (N_5167,N_4936,N_4966);
nand U5168 (N_5168,N_4811,N_4889);
nor U5169 (N_5169,N_4948,N_4889);
nor U5170 (N_5170,N_4970,N_4943);
and U5171 (N_5171,N_4807,N_4946);
nor U5172 (N_5172,N_4837,N_4918);
nor U5173 (N_5173,N_4819,N_4820);
and U5174 (N_5174,N_4971,N_4966);
or U5175 (N_5175,N_4812,N_4859);
nor U5176 (N_5176,N_4994,N_4917);
and U5177 (N_5177,N_4853,N_4876);
nor U5178 (N_5178,N_4993,N_4845);
and U5179 (N_5179,N_4863,N_4948);
and U5180 (N_5180,N_4911,N_4974);
nor U5181 (N_5181,N_4971,N_4887);
or U5182 (N_5182,N_4869,N_4801);
and U5183 (N_5183,N_4932,N_4828);
nor U5184 (N_5184,N_4806,N_4807);
nand U5185 (N_5185,N_4901,N_4845);
nand U5186 (N_5186,N_4982,N_4902);
nor U5187 (N_5187,N_4954,N_4830);
or U5188 (N_5188,N_4934,N_4888);
nand U5189 (N_5189,N_4961,N_4805);
xor U5190 (N_5190,N_4906,N_4952);
and U5191 (N_5191,N_4911,N_4978);
nand U5192 (N_5192,N_4931,N_4996);
nand U5193 (N_5193,N_4824,N_4827);
nand U5194 (N_5194,N_4942,N_4915);
nor U5195 (N_5195,N_4997,N_4873);
nor U5196 (N_5196,N_4835,N_4979);
xor U5197 (N_5197,N_4809,N_4968);
or U5198 (N_5198,N_4909,N_4964);
and U5199 (N_5199,N_4965,N_4829);
and U5200 (N_5200,N_5045,N_5057);
and U5201 (N_5201,N_5085,N_5127);
xnor U5202 (N_5202,N_5107,N_5138);
and U5203 (N_5203,N_5088,N_5163);
nand U5204 (N_5204,N_5033,N_5087);
nand U5205 (N_5205,N_5095,N_5185);
nand U5206 (N_5206,N_5183,N_5065);
and U5207 (N_5207,N_5113,N_5132);
nand U5208 (N_5208,N_5039,N_5139);
xnor U5209 (N_5209,N_5090,N_5110);
xnor U5210 (N_5210,N_5082,N_5024);
and U5211 (N_5211,N_5135,N_5008);
or U5212 (N_5212,N_5066,N_5018);
xnor U5213 (N_5213,N_5176,N_5136);
and U5214 (N_5214,N_5188,N_5131);
nand U5215 (N_5215,N_5058,N_5011);
nand U5216 (N_5216,N_5072,N_5195);
nor U5217 (N_5217,N_5111,N_5196);
nand U5218 (N_5218,N_5165,N_5161);
and U5219 (N_5219,N_5180,N_5112);
xnor U5220 (N_5220,N_5137,N_5098);
and U5221 (N_5221,N_5047,N_5105);
or U5222 (N_5222,N_5159,N_5056);
xor U5223 (N_5223,N_5120,N_5145);
nor U5224 (N_5224,N_5099,N_5070);
and U5225 (N_5225,N_5141,N_5108);
nor U5226 (N_5226,N_5148,N_5192);
or U5227 (N_5227,N_5106,N_5022);
or U5228 (N_5228,N_5009,N_5093);
nor U5229 (N_5229,N_5027,N_5020);
nor U5230 (N_5230,N_5186,N_5144);
nand U5231 (N_5231,N_5103,N_5094);
or U5232 (N_5232,N_5063,N_5017);
and U5233 (N_5233,N_5146,N_5101);
xor U5234 (N_5234,N_5084,N_5187);
nand U5235 (N_5235,N_5114,N_5177);
and U5236 (N_5236,N_5000,N_5173);
or U5237 (N_5237,N_5043,N_5129);
and U5238 (N_5238,N_5081,N_5142);
and U5239 (N_5239,N_5170,N_5032);
xor U5240 (N_5240,N_5152,N_5150);
xnor U5241 (N_5241,N_5053,N_5158);
or U5242 (N_5242,N_5048,N_5097);
nor U5243 (N_5243,N_5025,N_5076);
or U5244 (N_5244,N_5023,N_5153);
and U5245 (N_5245,N_5073,N_5181);
nand U5246 (N_5246,N_5156,N_5154);
nor U5247 (N_5247,N_5030,N_5060);
or U5248 (N_5248,N_5016,N_5115);
and U5249 (N_5249,N_5194,N_5121);
nand U5250 (N_5250,N_5031,N_5044);
or U5251 (N_5251,N_5042,N_5035);
xnor U5252 (N_5252,N_5040,N_5119);
nor U5253 (N_5253,N_5174,N_5133);
nor U5254 (N_5254,N_5092,N_5116);
or U5255 (N_5255,N_5059,N_5019);
or U5256 (N_5256,N_5172,N_5034);
nand U5257 (N_5257,N_5157,N_5109);
and U5258 (N_5258,N_5134,N_5118);
xnor U5259 (N_5259,N_5055,N_5013);
xor U5260 (N_5260,N_5012,N_5083);
xnor U5261 (N_5261,N_5199,N_5052);
nand U5262 (N_5262,N_5096,N_5064);
or U5263 (N_5263,N_5197,N_5068);
and U5264 (N_5264,N_5102,N_5005);
xnor U5265 (N_5265,N_5175,N_5075);
nor U5266 (N_5266,N_5028,N_5038);
nand U5267 (N_5267,N_5002,N_5122);
or U5268 (N_5268,N_5026,N_5147);
or U5269 (N_5269,N_5051,N_5130);
nand U5270 (N_5270,N_5143,N_5089);
and U5271 (N_5271,N_5155,N_5004);
nor U5272 (N_5272,N_5001,N_5029);
nor U5273 (N_5273,N_5071,N_5100);
or U5274 (N_5274,N_5080,N_5041);
xor U5275 (N_5275,N_5189,N_5128);
nor U5276 (N_5276,N_5037,N_5091);
and U5277 (N_5277,N_5014,N_5191);
nand U5278 (N_5278,N_5067,N_5007);
xnor U5279 (N_5279,N_5078,N_5069);
xnor U5280 (N_5280,N_5171,N_5162);
xnor U5281 (N_5281,N_5178,N_5104);
nand U5282 (N_5282,N_5086,N_5006);
and U5283 (N_5283,N_5077,N_5149);
and U5284 (N_5284,N_5167,N_5151);
nand U5285 (N_5285,N_5184,N_5015);
nand U5286 (N_5286,N_5168,N_5179);
or U5287 (N_5287,N_5164,N_5074);
or U5288 (N_5288,N_5046,N_5166);
xor U5289 (N_5289,N_5140,N_5061);
nand U5290 (N_5290,N_5124,N_5160);
nand U5291 (N_5291,N_5021,N_5198);
or U5292 (N_5292,N_5049,N_5036);
or U5293 (N_5293,N_5190,N_5079);
nand U5294 (N_5294,N_5050,N_5193);
nand U5295 (N_5295,N_5123,N_5126);
and U5296 (N_5296,N_5117,N_5182);
xnor U5297 (N_5297,N_5125,N_5003);
and U5298 (N_5298,N_5010,N_5054);
or U5299 (N_5299,N_5062,N_5169);
xor U5300 (N_5300,N_5073,N_5123);
nor U5301 (N_5301,N_5013,N_5102);
and U5302 (N_5302,N_5062,N_5161);
and U5303 (N_5303,N_5094,N_5183);
nor U5304 (N_5304,N_5164,N_5049);
nor U5305 (N_5305,N_5083,N_5132);
nor U5306 (N_5306,N_5120,N_5114);
nor U5307 (N_5307,N_5063,N_5131);
and U5308 (N_5308,N_5174,N_5182);
and U5309 (N_5309,N_5078,N_5089);
nor U5310 (N_5310,N_5086,N_5032);
nor U5311 (N_5311,N_5002,N_5088);
nor U5312 (N_5312,N_5032,N_5166);
xnor U5313 (N_5313,N_5035,N_5076);
or U5314 (N_5314,N_5102,N_5144);
and U5315 (N_5315,N_5047,N_5185);
xor U5316 (N_5316,N_5065,N_5036);
or U5317 (N_5317,N_5090,N_5071);
nor U5318 (N_5318,N_5075,N_5024);
and U5319 (N_5319,N_5163,N_5025);
and U5320 (N_5320,N_5032,N_5135);
or U5321 (N_5321,N_5133,N_5187);
xnor U5322 (N_5322,N_5027,N_5044);
xor U5323 (N_5323,N_5115,N_5181);
nand U5324 (N_5324,N_5110,N_5107);
nor U5325 (N_5325,N_5016,N_5105);
or U5326 (N_5326,N_5151,N_5107);
nand U5327 (N_5327,N_5007,N_5083);
nand U5328 (N_5328,N_5019,N_5098);
nand U5329 (N_5329,N_5172,N_5117);
or U5330 (N_5330,N_5046,N_5155);
and U5331 (N_5331,N_5089,N_5186);
nor U5332 (N_5332,N_5180,N_5198);
or U5333 (N_5333,N_5115,N_5002);
or U5334 (N_5334,N_5022,N_5005);
and U5335 (N_5335,N_5064,N_5118);
and U5336 (N_5336,N_5162,N_5064);
xnor U5337 (N_5337,N_5031,N_5158);
xnor U5338 (N_5338,N_5031,N_5077);
xor U5339 (N_5339,N_5164,N_5121);
xor U5340 (N_5340,N_5138,N_5133);
nor U5341 (N_5341,N_5038,N_5085);
or U5342 (N_5342,N_5171,N_5132);
nand U5343 (N_5343,N_5032,N_5088);
xor U5344 (N_5344,N_5151,N_5044);
xor U5345 (N_5345,N_5196,N_5167);
xor U5346 (N_5346,N_5117,N_5053);
and U5347 (N_5347,N_5140,N_5037);
xor U5348 (N_5348,N_5199,N_5161);
and U5349 (N_5349,N_5150,N_5025);
xnor U5350 (N_5350,N_5073,N_5148);
nand U5351 (N_5351,N_5075,N_5138);
nor U5352 (N_5352,N_5077,N_5025);
nand U5353 (N_5353,N_5180,N_5151);
xnor U5354 (N_5354,N_5179,N_5189);
or U5355 (N_5355,N_5041,N_5024);
nor U5356 (N_5356,N_5101,N_5173);
nand U5357 (N_5357,N_5152,N_5084);
xor U5358 (N_5358,N_5001,N_5114);
nand U5359 (N_5359,N_5162,N_5052);
or U5360 (N_5360,N_5119,N_5194);
xor U5361 (N_5361,N_5012,N_5015);
and U5362 (N_5362,N_5064,N_5180);
or U5363 (N_5363,N_5118,N_5082);
and U5364 (N_5364,N_5167,N_5047);
xor U5365 (N_5365,N_5196,N_5009);
or U5366 (N_5366,N_5015,N_5175);
nor U5367 (N_5367,N_5000,N_5096);
and U5368 (N_5368,N_5131,N_5104);
or U5369 (N_5369,N_5148,N_5071);
or U5370 (N_5370,N_5112,N_5068);
xor U5371 (N_5371,N_5036,N_5034);
xor U5372 (N_5372,N_5115,N_5006);
nor U5373 (N_5373,N_5102,N_5163);
xnor U5374 (N_5374,N_5108,N_5115);
and U5375 (N_5375,N_5047,N_5190);
or U5376 (N_5376,N_5127,N_5064);
xor U5377 (N_5377,N_5117,N_5023);
xnor U5378 (N_5378,N_5121,N_5124);
or U5379 (N_5379,N_5080,N_5014);
nor U5380 (N_5380,N_5088,N_5145);
and U5381 (N_5381,N_5008,N_5025);
or U5382 (N_5382,N_5117,N_5065);
nand U5383 (N_5383,N_5034,N_5125);
and U5384 (N_5384,N_5097,N_5040);
or U5385 (N_5385,N_5011,N_5047);
nand U5386 (N_5386,N_5052,N_5093);
or U5387 (N_5387,N_5072,N_5140);
or U5388 (N_5388,N_5041,N_5179);
nand U5389 (N_5389,N_5016,N_5011);
or U5390 (N_5390,N_5152,N_5179);
and U5391 (N_5391,N_5084,N_5151);
or U5392 (N_5392,N_5054,N_5125);
nand U5393 (N_5393,N_5121,N_5027);
xnor U5394 (N_5394,N_5171,N_5199);
nor U5395 (N_5395,N_5152,N_5043);
and U5396 (N_5396,N_5048,N_5124);
nand U5397 (N_5397,N_5070,N_5117);
or U5398 (N_5398,N_5019,N_5054);
and U5399 (N_5399,N_5192,N_5011);
or U5400 (N_5400,N_5322,N_5205);
or U5401 (N_5401,N_5357,N_5272);
or U5402 (N_5402,N_5333,N_5312);
xnor U5403 (N_5403,N_5391,N_5337);
or U5404 (N_5404,N_5202,N_5327);
nand U5405 (N_5405,N_5323,N_5378);
or U5406 (N_5406,N_5267,N_5225);
and U5407 (N_5407,N_5289,N_5223);
and U5408 (N_5408,N_5372,N_5282);
nor U5409 (N_5409,N_5286,N_5249);
or U5410 (N_5410,N_5243,N_5371);
or U5411 (N_5411,N_5277,N_5342);
xor U5412 (N_5412,N_5293,N_5311);
and U5413 (N_5413,N_5360,N_5216);
nand U5414 (N_5414,N_5398,N_5339);
nand U5415 (N_5415,N_5305,N_5259);
xor U5416 (N_5416,N_5228,N_5231);
nand U5417 (N_5417,N_5392,N_5278);
or U5418 (N_5418,N_5353,N_5344);
xnor U5419 (N_5419,N_5363,N_5247);
nor U5420 (N_5420,N_5257,N_5276);
nor U5421 (N_5421,N_5300,N_5307);
or U5422 (N_5422,N_5358,N_5214);
or U5423 (N_5423,N_5332,N_5330);
nand U5424 (N_5424,N_5366,N_5241);
and U5425 (N_5425,N_5274,N_5294);
nand U5426 (N_5426,N_5343,N_5291);
and U5427 (N_5427,N_5244,N_5220);
or U5428 (N_5428,N_5380,N_5369);
nor U5429 (N_5429,N_5310,N_5329);
nor U5430 (N_5430,N_5376,N_5203);
nand U5431 (N_5431,N_5387,N_5298);
nand U5432 (N_5432,N_5348,N_5385);
nor U5433 (N_5433,N_5386,N_5265);
or U5434 (N_5434,N_5389,N_5271);
nand U5435 (N_5435,N_5219,N_5364);
and U5436 (N_5436,N_5347,N_5253);
nand U5437 (N_5437,N_5368,N_5308);
or U5438 (N_5438,N_5258,N_5230);
nand U5439 (N_5439,N_5250,N_5356);
and U5440 (N_5440,N_5263,N_5284);
nor U5441 (N_5441,N_5299,N_5240);
or U5442 (N_5442,N_5224,N_5221);
nor U5443 (N_5443,N_5381,N_5396);
xor U5444 (N_5444,N_5229,N_5367);
or U5445 (N_5445,N_5237,N_5248);
nand U5446 (N_5446,N_5251,N_5236);
or U5447 (N_5447,N_5331,N_5317);
or U5448 (N_5448,N_5313,N_5399);
and U5449 (N_5449,N_5288,N_5269);
or U5450 (N_5450,N_5315,N_5346);
or U5451 (N_5451,N_5296,N_5255);
nor U5452 (N_5452,N_5379,N_5297);
and U5453 (N_5453,N_5314,N_5309);
and U5454 (N_5454,N_5361,N_5377);
nor U5455 (N_5455,N_5384,N_5316);
xnor U5456 (N_5456,N_5355,N_5335);
nand U5457 (N_5457,N_5318,N_5390);
nand U5458 (N_5458,N_5204,N_5340);
nand U5459 (N_5459,N_5280,N_5319);
nor U5460 (N_5460,N_5351,N_5232);
or U5461 (N_5461,N_5382,N_5210);
and U5462 (N_5462,N_5375,N_5227);
or U5463 (N_5463,N_5273,N_5207);
xor U5464 (N_5464,N_5295,N_5206);
and U5465 (N_5465,N_5270,N_5336);
nand U5466 (N_5466,N_5254,N_5359);
or U5467 (N_5467,N_5261,N_5242);
and U5468 (N_5468,N_5283,N_5362);
xnor U5469 (N_5469,N_5338,N_5373);
and U5470 (N_5470,N_5302,N_5306);
nand U5471 (N_5471,N_5208,N_5354);
and U5472 (N_5472,N_5321,N_5324);
nor U5473 (N_5473,N_5303,N_5235);
or U5474 (N_5474,N_5320,N_5349);
nor U5475 (N_5475,N_5365,N_5304);
or U5476 (N_5476,N_5226,N_5301);
nor U5477 (N_5477,N_5334,N_5370);
nor U5478 (N_5478,N_5234,N_5352);
and U5479 (N_5479,N_5211,N_5292);
nor U5480 (N_5480,N_5279,N_5256);
nor U5481 (N_5481,N_5260,N_5201);
xor U5482 (N_5482,N_5328,N_5287);
and U5483 (N_5483,N_5200,N_5212);
xor U5484 (N_5484,N_5233,N_5222);
and U5485 (N_5485,N_5218,N_5374);
xnor U5486 (N_5486,N_5239,N_5238);
nor U5487 (N_5487,N_5281,N_5262);
xnor U5488 (N_5488,N_5341,N_5326);
nand U5489 (N_5489,N_5394,N_5290);
and U5490 (N_5490,N_5397,N_5209);
or U5491 (N_5491,N_5268,N_5264);
or U5492 (N_5492,N_5345,N_5383);
xor U5493 (N_5493,N_5285,N_5350);
or U5494 (N_5494,N_5213,N_5252);
or U5495 (N_5495,N_5266,N_5245);
and U5496 (N_5496,N_5395,N_5217);
or U5497 (N_5497,N_5325,N_5275);
xor U5498 (N_5498,N_5393,N_5388);
nor U5499 (N_5499,N_5246,N_5215);
and U5500 (N_5500,N_5371,N_5271);
and U5501 (N_5501,N_5362,N_5304);
nand U5502 (N_5502,N_5320,N_5350);
and U5503 (N_5503,N_5264,N_5257);
nand U5504 (N_5504,N_5266,N_5202);
and U5505 (N_5505,N_5264,N_5218);
xnor U5506 (N_5506,N_5261,N_5237);
nand U5507 (N_5507,N_5202,N_5386);
and U5508 (N_5508,N_5204,N_5341);
nor U5509 (N_5509,N_5328,N_5201);
nor U5510 (N_5510,N_5240,N_5201);
xnor U5511 (N_5511,N_5207,N_5314);
xnor U5512 (N_5512,N_5272,N_5260);
nand U5513 (N_5513,N_5356,N_5263);
xor U5514 (N_5514,N_5280,N_5314);
nand U5515 (N_5515,N_5309,N_5358);
and U5516 (N_5516,N_5342,N_5202);
nor U5517 (N_5517,N_5368,N_5318);
xnor U5518 (N_5518,N_5309,N_5384);
nor U5519 (N_5519,N_5283,N_5203);
and U5520 (N_5520,N_5236,N_5364);
xor U5521 (N_5521,N_5394,N_5379);
nor U5522 (N_5522,N_5322,N_5244);
or U5523 (N_5523,N_5211,N_5348);
or U5524 (N_5524,N_5328,N_5308);
or U5525 (N_5525,N_5313,N_5352);
or U5526 (N_5526,N_5288,N_5346);
nand U5527 (N_5527,N_5263,N_5210);
nand U5528 (N_5528,N_5294,N_5376);
nor U5529 (N_5529,N_5286,N_5383);
nand U5530 (N_5530,N_5208,N_5255);
xnor U5531 (N_5531,N_5238,N_5272);
or U5532 (N_5532,N_5279,N_5327);
and U5533 (N_5533,N_5300,N_5368);
or U5534 (N_5534,N_5344,N_5312);
or U5535 (N_5535,N_5394,N_5324);
nor U5536 (N_5536,N_5284,N_5391);
or U5537 (N_5537,N_5339,N_5262);
nor U5538 (N_5538,N_5371,N_5381);
nor U5539 (N_5539,N_5311,N_5223);
xor U5540 (N_5540,N_5350,N_5340);
xnor U5541 (N_5541,N_5309,N_5250);
or U5542 (N_5542,N_5207,N_5381);
or U5543 (N_5543,N_5271,N_5295);
nand U5544 (N_5544,N_5367,N_5363);
nor U5545 (N_5545,N_5241,N_5354);
nand U5546 (N_5546,N_5273,N_5301);
nand U5547 (N_5547,N_5229,N_5329);
xnor U5548 (N_5548,N_5252,N_5339);
and U5549 (N_5549,N_5302,N_5328);
xnor U5550 (N_5550,N_5281,N_5239);
nand U5551 (N_5551,N_5224,N_5222);
or U5552 (N_5552,N_5371,N_5259);
and U5553 (N_5553,N_5226,N_5317);
nand U5554 (N_5554,N_5244,N_5330);
or U5555 (N_5555,N_5300,N_5215);
nand U5556 (N_5556,N_5334,N_5353);
or U5557 (N_5557,N_5391,N_5316);
and U5558 (N_5558,N_5352,N_5206);
xor U5559 (N_5559,N_5252,N_5260);
nor U5560 (N_5560,N_5236,N_5273);
nand U5561 (N_5561,N_5335,N_5238);
xnor U5562 (N_5562,N_5359,N_5268);
nand U5563 (N_5563,N_5200,N_5354);
or U5564 (N_5564,N_5217,N_5382);
and U5565 (N_5565,N_5380,N_5219);
nor U5566 (N_5566,N_5264,N_5213);
nand U5567 (N_5567,N_5365,N_5398);
xnor U5568 (N_5568,N_5206,N_5223);
xnor U5569 (N_5569,N_5292,N_5273);
or U5570 (N_5570,N_5381,N_5318);
nand U5571 (N_5571,N_5203,N_5399);
nand U5572 (N_5572,N_5241,N_5271);
nor U5573 (N_5573,N_5277,N_5313);
nor U5574 (N_5574,N_5244,N_5378);
or U5575 (N_5575,N_5355,N_5348);
nand U5576 (N_5576,N_5340,N_5330);
nor U5577 (N_5577,N_5221,N_5381);
and U5578 (N_5578,N_5286,N_5202);
and U5579 (N_5579,N_5230,N_5221);
nor U5580 (N_5580,N_5294,N_5379);
or U5581 (N_5581,N_5312,N_5218);
and U5582 (N_5582,N_5255,N_5251);
nand U5583 (N_5583,N_5247,N_5310);
nor U5584 (N_5584,N_5297,N_5395);
or U5585 (N_5585,N_5243,N_5228);
nand U5586 (N_5586,N_5229,N_5341);
xnor U5587 (N_5587,N_5284,N_5361);
xnor U5588 (N_5588,N_5308,N_5211);
xnor U5589 (N_5589,N_5216,N_5262);
nand U5590 (N_5590,N_5389,N_5250);
nand U5591 (N_5591,N_5300,N_5211);
nor U5592 (N_5592,N_5232,N_5256);
or U5593 (N_5593,N_5293,N_5234);
xor U5594 (N_5594,N_5277,N_5251);
nand U5595 (N_5595,N_5306,N_5275);
xor U5596 (N_5596,N_5316,N_5282);
nor U5597 (N_5597,N_5393,N_5216);
xnor U5598 (N_5598,N_5390,N_5203);
or U5599 (N_5599,N_5393,N_5378);
nor U5600 (N_5600,N_5564,N_5543);
nor U5601 (N_5601,N_5512,N_5447);
nand U5602 (N_5602,N_5595,N_5466);
nand U5603 (N_5603,N_5575,N_5486);
xor U5604 (N_5604,N_5433,N_5468);
nor U5605 (N_5605,N_5412,N_5403);
nand U5606 (N_5606,N_5505,N_5509);
xor U5607 (N_5607,N_5407,N_5405);
nor U5608 (N_5608,N_5553,N_5589);
nor U5609 (N_5609,N_5503,N_5582);
and U5610 (N_5610,N_5415,N_5540);
and U5611 (N_5611,N_5484,N_5411);
or U5612 (N_5612,N_5496,N_5429);
nor U5613 (N_5613,N_5404,N_5443);
xnor U5614 (N_5614,N_5401,N_5545);
nand U5615 (N_5615,N_5520,N_5470);
or U5616 (N_5616,N_5559,N_5514);
xor U5617 (N_5617,N_5421,N_5416);
or U5618 (N_5618,N_5464,N_5473);
xor U5619 (N_5619,N_5471,N_5532);
or U5620 (N_5620,N_5577,N_5555);
or U5621 (N_5621,N_5534,N_5598);
nand U5622 (N_5622,N_5574,N_5506);
and U5623 (N_5623,N_5568,N_5501);
xor U5624 (N_5624,N_5583,N_5406);
nor U5625 (N_5625,N_5573,N_5511);
nor U5626 (N_5626,N_5402,N_5525);
xor U5627 (N_5627,N_5565,N_5502);
nand U5628 (N_5628,N_5436,N_5454);
xnor U5629 (N_5629,N_5596,N_5523);
nand U5630 (N_5630,N_5556,N_5586);
nor U5631 (N_5631,N_5594,N_5458);
or U5632 (N_5632,N_5439,N_5580);
nand U5633 (N_5633,N_5477,N_5495);
nor U5634 (N_5634,N_5578,N_5519);
and U5635 (N_5635,N_5446,N_5461);
nor U5636 (N_5636,N_5499,N_5418);
xor U5637 (N_5637,N_5526,N_5452);
and U5638 (N_5638,N_5490,N_5417);
and U5639 (N_5639,N_5541,N_5562);
and U5640 (N_5640,N_5524,N_5537);
nand U5641 (N_5641,N_5434,N_5529);
nor U5642 (N_5642,N_5467,N_5409);
nor U5643 (N_5643,N_5561,N_5542);
xor U5644 (N_5644,N_5535,N_5530);
and U5645 (N_5645,N_5493,N_5420);
or U5646 (N_5646,N_5475,N_5581);
nand U5647 (N_5647,N_5451,N_5552);
or U5648 (N_5648,N_5482,N_5547);
xnor U5649 (N_5649,N_5538,N_5522);
nand U5650 (N_5650,N_5597,N_5527);
and U5651 (N_5651,N_5587,N_5460);
nor U5652 (N_5652,N_5437,N_5428);
or U5653 (N_5653,N_5485,N_5593);
and U5654 (N_5654,N_5450,N_5444);
xor U5655 (N_5655,N_5408,N_5585);
xor U5656 (N_5656,N_5518,N_5576);
or U5657 (N_5657,N_5424,N_5492);
xnor U5658 (N_5658,N_5413,N_5513);
nor U5659 (N_5659,N_5504,N_5441);
or U5660 (N_5660,N_5572,N_5557);
xor U5661 (N_5661,N_5423,N_5558);
or U5662 (N_5662,N_5456,N_5435);
nor U5663 (N_5663,N_5491,N_5531);
nor U5664 (N_5664,N_5469,N_5570);
or U5665 (N_5665,N_5549,N_5480);
xnor U5666 (N_5666,N_5481,N_5442);
nor U5667 (N_5667,N_5425,N_5571);
and U5668 (N_5668,N_5533,N_5489);
xnor U5669 (N_5669,N_5426,N_5498);
and U5670 (N_5670,N_5474,N_5515);
nor U5671 (N_5671,N_5591,N_5528);
xor U5672 (N_5672,N_5599,N_5445);
or U5673 (N_5673,N_5462,N_5507);
xnor U5674 (N_5674,N_5516,N_5419);
and U5675 (N_5675,N_5592,N_5448);
xnor U5676 (N_5676,N_5432,N_5497);
nor U5677 (N_5677,N_5430,N_5422);
xor U5678 (N_5678,N_5400,N_5551);
and U5679 (N_5679,N_5494,N_5463);
or U5680 (N_5680,N_5539,N_5546);
or U5681 (N_5681,N_5476,N_5550);
or U5682 (N_5682,N_5479,N_5453);
xnor U5683 (N_5683,N_5579,N_5472);
and U5684 (N_5684,N_5500,N_5569);
or U5685 (N_5685,N_5410,N_5455);
nor U5686 (N_5686,N_5487,N_5560);
nand U5687 (N_5687,N_5517,N_5440);
nand U5688 (N_5688,N_5563,N_5567);
or U5689 (N_5689,N_5588,N_5427);
or U5690 (N_5690,N_5431,N_5438);
nand U5691 (N_5691,N_5566,N_5544);
nor U5692 (N_5692,N_5483,N_5508);
nand U5693 (N_5693,N_5459,N_5554);
nand U5694 (N_5694,N_5457,N_5548);
or U5695 (N_5695,N_5414,N_5521);
or U5696 (N_5696,N_5584,N_5465);
or U5697 (N_5697,N_5590,N_5478);
nor U5698 (N_5698,N_5536,N_5488);
or U5699 (N_5699,N_5449,N_5510);
or U5700 (N_5700,N_5448,N_5493);
and U5701 (N_5701,N_5461,N_5572);
or U5702 (N_5702,N_5493,N_5562);
nor U5703 (N_5703,N_5421,N_5406);
nor U5704 (N_5704,N_5445,N_5593);
nand U5705 (N_5705,N_5467,N_5417);
xnor U5706 (N_5706,N_5489,N_5577);
nand U5707 (N_5707,N_5491,N_5408);
nor U5708 (N_5708,N_5544,N_5447);
nand U5709 (N_5709,N_5471,N_5567);
and U5710 (N_5710,N_5493,N_5519);
nor U5711 (N_5711,N_5567,N_5560);
nor U5712 (N_5712,N_5533,N_5420);
nor U5713 (N_5713,N_5465,N_5474);
and U5714 (N_5714,N_5471,N_5531);
or U5715 (N_5715,N_5518,N_5598);
or U5716 (N_5716,N_5502,N_5402);
xnor U5717 (N_5717,N_5583,N_5542);
or U5718 (N_5718,N_5424,N_5425);
or U5719 (N_5719,N_5513,N_5485);
xnor U5720 (N_5720,N_5454,N_5529);
and U5721 (N_5721,N_5419,N_5445);
xnor U5722 (N_5722,N_5450,N_5590);
nand U5723 (N_5723,N_5462,N_5459);
nand U5724 (N_5724,N_5545,N_5433);
or U5725 (N_5725,N_5593,N_5424);
xor U5726 (N_5726,N_5547,N_5555);
and U5727 (N_5727,N_5572,N_5410);
xor U5728 (N_5728,N_5509,N_5558);
nand U5729 (N_5729,N_5469,N_5586);
and U5730 (N_5730,N_5444,N_5497);
nor U5731 (N_5731,N_5457,N_5516);
xor U5732 (N_5732,N_5430,N_5532);
xor U5733 (N_5733,N_5554,N_5521);
xnor U5734 (N_5734,N_5463,N_5531);
xor U5735 (N_5735,N_5484,N_5518);
or U5736 (N_5736,N_5464,N_5579);
nor U5737 (N_5737,N_5511,N_5566);
xnor U5738 (N_5738,N_5594,N_5502);
or U5739 (N_5739,N_5515,N_5412);
nand U5740 (N_5740,N_5450,N_5522);
xnor U5741 (N_5741,N_5498,N_5577);
and U5742 (N_5742,N_5405,N_5402);
or U5743 (N_5743,N_5479,N_5480);
and U5744 (N_5744,N_5466,N_5422);
and U5745 (N_5745,N_5404,N_5492);
and U5746 (N_5746,N_5559,N_5413);
nor U5747 (N_5747,N_5451,N_5423);
xor U5748 (N_5748,N_5417,N_5513);
xor U5749 (N_5749,N_5405,N_5581);
and U5750 (N_5750,N_5472,N_5408);
nand U5751 (N_5751,N_5581,N_5442);
or U5752 (N_5752,N_5458,N_5466);
nor U5753 (N_5753,N_5556,N_5497);
and U5754 (N_5754,N_5491,N_5548);
xor U5755 (N_5755,N_5434,N_5411);
nor U5756 (N_5756,N_5427,N_5527);
xor U5757 (N_5757,N_5493,N_5585);
and U5758 (N_5758,N_5543,N_5572);
and U5759 (N_5759,N_5421,N_5485);
or U5760 (N_5760,N_5455,N_5504);
or U5761 (N_5761,N_5450,N_5516);
xor U5762 (N_5762,N_5449,N_5590);
nor U5763 (N_5763,N_5563,N_5484);
nand U5764 (N_5764,N_5517,N_5558);
xnor U5765 (N_5765,N_5494,N_5450);
and U5766 (N_5766,N_5517,N_5433);
or U5767 (N_5767,N_5549,N_5537);
and U5768 (N_5768,N_5557,N_5410);
and U5769 (N_5769,N_5554,N_5525);
nor U5770 (N_5770,N_5440,N_5456);
or U5771 (N_5771,N_5581,N_5510);
xor U5772 (N_5772,N_5474,N_5527);
or U5773 (N_5773,N_5400,N_5535);
or U5774 (N_5774,N_5532,N_5469);
xor U5775 (N_5775,N_5451,N_5516);
and U5776 (N_5776,N_5588,N_5564);
xnor U5777 (N_5777,N_5525,N_5408);
xnor U5778 (N_5778,N_5454,N_5572);
nand U5779 (N_5779,N_5490,N_5474);
xor U5780 (N_5780,N_5423,N_5411);
and U5781 (N_5781,N_5526,N_5511);
xor U5782 (N_5782,N_5508,N_5513);
or U5783 (N_5783,N_5487,N_5425);
and U5784 (N_5784,N_5469,N_5582);
or U5785 (N_5785,N_5529,N_5405);
nand U5786 (N_5786,N_5491,N_5485);
and U5787 (N_5787,N_5438,N_5464);
nor U5788 (N_5788,N_5508,N_5553);
xnor U5789 (N_5789,N_5570,N_5534);
or U5790 (N_5790,N_5531,N_5470);
and U5791 (N_5791,N_5456,N_5549);
nand U5792 (N_5792,N_5404,N_5537);
nor U5793 (N_5793,N_5455,N_5493);
nand U5794 (N_5794,N_5509,N_5522);
nand U5795 (N_5795,N_5596,N_5545);
nor U5796 (N_5796,N_5512,N_5480);
nor U5797 (N_5797,N_5520,N_5480);
xor U5798 (N_5798,N_5582,N_5474);
xnor U5799 (N_5799,N_5520,N_5406);
nor U5800 (N_5800,N_5609,N_5765);
xnor U5801 (N_5801,N_5711,N_5764);
xnor U5802 (N_5802,N_5712,N_5730);
nand U5803 (N_5803,N_5724,N_5625);
xnor U5804 (N_5804,N_5792,N_5601);
and U5805 (N_5805,N_5789,N_5731);
nand U5806 (N_5806,N_5714,N_5617);
nand U5807 (N_5807,N_5605,N_5706);
or U5808 (N_5808,N_5787,N_5780);
and U5809 (N_5809,N_5746,N_5702);
nor U5810 (N_5810,N_5635,N_5784);
xor U5811 (N_5811,N_5690,N_5620);
nand U5812 (N_5812,N_5685,N_5632);
and U5813 (N_5813,N_5783,N_5713);
nand U5814 (N_5814,N_5687,N_5782);
or U5815 (N_5815,N_5602,N_5623);
and U5816 (N_5816,N_5618,N_5663);
and U5817 (N_5817,N_5697,N_5600);
nor U5818 (N_5818,N_5752,N_5686);
nor U5819 (N_5819,N_5722,N_5734);
nor U5820 (N_5820,N_5732,N_5680);
nor U5821 (N_5821,N_5776,N_5791);
nor U5822 (N_5822,N_5646,N_5626);
or U5823 (N_5823,N_5645,N_5629);
nor U5824 (N_5824,N_5628,N_5676);
nand U5825 (N_5825,N_5723,N_5772);
nand U5826 (N_5826,N_5736,N_5665);
nand U5827 (N_5827,N_5766,N_5774);
nor U5828 (N_5828,N_5673,N_5643);
nand U5829 (N_5829,N_5651,N_5788);
xor U5830 (N_5830,N_5640,N_5684);
and U5831 (N_5831,N_5682,N_5619);
nor U5832 (N_5832,N_5708,N_5747);
and U5833 (N_5833,N_5677,N_5700);
nand U5834 (N_5834,N_5654,N_5761);
nor U5835 (N_5835,N_5727,N_5611);
or U5836 (N_5836,N_5785,N_5715);
nand U5837 (N_5837,N_5672,N_5777);
nand U5838 (N_5838,N_5769,N_5668);
and U5839 (N_5839,N_5705,N_5657);
or U5840 (N_5840,N_5666,N_5737);
and U5841 (N_5841,N_5610,N_5678);
or U5842 (N_5842,N_5768,N_5603);
and U5843 (N_5843,N_5671,N_5775);
nor U5844 (N_5844,N_5795,N_5650);
xnor U5845 (N_5845,N_5659,N_5797);
xor U5846 (N_5846,N_5660,N_5689);
nor U5847 (N_5847,N_5630,N_5720);
xor U5848 (N_5848,N_5698,N_5637);
and U5849 (N_5849,N_5779,N_5631);
nor U5850 (N_5850,N_5633,N_5622);
nor U5851 (N_5851,N_5621,N_5616);
and U5852 (N_5852,N_5790,N_5652);
and U5853 (N_5853,N_5710,N_5741);
xnor U5854 (N_5854,N_5675,N_5771);
nor U5855 (N_5855,N_5721,N_5679);
nand U5856 (N_5856,N_5745,N_5613);
and U5857 (N_5857,N_5716,N_5607);
nand U5858 (N_5858,N_5642,N_5692);
nand U5859 (N_5859,N_5608,N_5674);
or U5860 (N_5860,N_5756,N_5624);
and U5861 (N_5861,N_5755,N_5604);
and U5862 (N_5862,N_5770,N_5653);
nand U5863 (N_5863,N_5606,N_5728);
nor U5864 (N_5864,N_5641,N_5742);
nand U5865 (N_5865,N_5719,N_5762);
nor U5866 (N_5866,N_5786,N_5738);
and U5867 (N_5867,N_5636,N_5753);
or U5868 (N_5868,N_5662,N_5758);
or U5869 (N_5869,N_5773,N_5656);
xnor U5870 (N_5870,N_5717,N_5749);
and U5871 (N_5871,N_5699,N_5655);
and U5872 (N_5872,N_5794,N_5759);
and U5873 (N_5873,N_5735,N_5683);
nor U5874 (N_5874,N_5661,N_5647);
nand U5875 (N_5875,N_5740,N_5694);
xnor U5876 (N_5876,N_5688,N_5778);
xnor U5877 (N_5877,N_5703,N_5658);
nor U5878 (N_5878,N_5681,N_5781);
or U5879 (N_5879,N_5648,N_5615);
or U5880 (N_5880,N_5751,N_5739);
and U5881 (N_5881,N_5644,N_5744);
xor U5882 (N_5882,N_5767,N_5670);
xnor U5883 (N_5883,N_5743,N_5733);
nor U5884 (N_5884,N_5707,N_5709);
xnor U5885 (N_5885,N_5614,N_5669);
or U5886 (N_5886,N_5649,N_5750);
and U5887 (N_5887,N_5760,N_5664);
nand U5888 (N_5888,N_5627,N_5729);
nor U5889 (N_5889,N_5726,N_5701);
and U5890 (N_5890,N_5638,N_5757);
nor U5891 (N_5891,N_5725,N_5718);
nand U5892 (N_5892,N_5796,N_5639);
nor U5893 (N_5893,N_5763,N_5612);
and U5894 (N_5894,N_5691,N_5695);
nand U5895 (N_5895,N_5793,N_5799);
or U5896 (N_5896,N_5693,N_5704);
and U5897 (N_5897,N_5798,N_5754);
nor U5898 (N_5898,N_5748,N_5696);
nand U5899 (N_5899,N_5667,N_5634);
xor U5900 (N_5900,N_5620,N_5631);
or U5901 (N_5901,N_5784,N_5792);
xor U5902 (N_5902,N_5769,N_5775);
nand U5903 (N_5903,N_5778,N_5771);
nor U5904 (N_5904,N_5770,N_5606);
xor U5905 (N_5905,N_5674,N_5717);
xor U5906 (N_5906,N_5673,N_5602);
nor U5907 (N_5907,N_5725,N_5684);
xnor U5908 (N_5908,N_5777,N_5641);
or U5909 (N_5909,N_5698,N_5709);
and U5910 (N_5910,N_5656,N_5642);
and U5911 (N_5911,N_5703,N_5711);
or U5912 (N_5912,N_5683,N_5607);
nor U5913 (N_5913,N_5685,N_5710);
nor U5914 (N_5914,N_5719,N_5685);
nand U5915 (N_5915,N_5790,N_5776);
nand U5916 (N_5916,N_5608,N_5613);
nand U5917 (N_5917,N_5693,N_5782);
and U5918 (N_5918,N_5795,N_5710);
nor U5919 (N_5919,N_5678,N_5719);
or U5920 (N_5920,N_5645,N_5616);
nor U5921 (N_5921,N_5726,N_5621);
nor U5922 (N_5922,N_5607,N_5750);
nand U5923 (N_5923,N_5617,N_5767);
nand U5924 (N_5924,N_5718,N_5710);
xor U5925 (N_5925,N_5797,N_5605);
xor U5926 (N_5926,N_5632,N_5718);
xor U5927 (N_5927,N_5665,N_5690);
or U5928 (N_5928,N_5738,N_5773);
and U5929 (N_5929,N_5768,N_5749);
nor U5930 (N_5930,N_5780,N_5613);
xor U5931 (N_5931,N_5611,N_5631);
or U5932 (N_5932,N_5779,N_5609);
nand U5933 (N_5933,N_5749,N_5606);
nand U5934 (N_5934,N_5738,N_5747);
or U5935 (N_5935,N_5736,N_5698);
nand U5936 (N_5936,N_5761,N_5662);
xnor U5937 (N_5937,N_5668,N_5739);
nor U5938 (N_5938,N_5745,N_5794);
nor U5939 (N_5939,N_5708,N_5690);
nand U5940 (N_5940,N_5725,N_5795);
xor U5941 (N_5941,N_5624,N_5694);
xor U5942 (N_5942,N_5648,N_5607);
and U5943 (N_5943,N_5722,N_5659);
or U5944 (N_5944,N_5733,N_5677);
nor U5945 (N_5945,N_5778,N_5611);
nand U5946 (N_5946,N_5691,N_5665);
xnor U5947 (N_5947,N_5687,N_5625);
or U5948 (N_5948,N_5749,N_5688);
and U5949 (N_5949,N_5715,N_5756);
or U5950 (N_5950,N_5758,N_5667);
nand U5951 (N_5951,N_5665,N_5744);
nand U5952 (N_5952,N_5730,N_5745);
or U5953 (N_5953,N_5640,N_5696);
or U5954 (N_5954,N_5607,N_5747);
nand U5955 (N_5955,N_5678,N_5687);
and U5956 (N_5956,N_5751,N_5669);
nor U5957 (N_5957,N_5604,N_5715);
nor U5958 (N_5958,N_5778,N_5681);
nor U5959 (N_5959,N_5634,N_5651);
or U5960 (N_5960,N_5679,N_5758);
nand U5961 (N_5961,N_5712,N_5629);
and U5962 (N_5962,N_5686,N_5750);
and U5963 (N_5963,N_5613,N_5666);
and U5964 (N_5964,N_5651,N_5764);
and U5965 (N_5965,N_5724,N_5627);
or U5966 (N_5966,N_5613,N_5717);
nand U5967 (N_5967,N_5700,N_5686);
and U5968 (N_5968,N_5603,N_5683);
nor U5969 (N_5969,N_5655,N_5691);
nor U5970 (N_5970,N_5608,N_5662);
and U5971 (N_5971,N_5786,N_5777);
xor U5972 (N_5972,N_5681,N_5766);
nand U5973 (N_5973,N_5691,N_5727);
and U5974 (N_5974,N_5702,N_5773);
xor U5975 (N_5975,N_5704,N_5672);
and U5976 (N_5976,N_5735,N_5679);
and U5977 (N_5977,N_5671,N_5633);
nand U5978 (N_5978,N_5627,N_5687);
xor U5979 (N_5979,N_5661,N_5737);
or U5980 (N_5980,N_5659,N_5698);
xor U5981 (N_5981,N_5780,N_5693);
and U5982 (N_5982,N_5785,N_5773);
xor U5983 (N_5983,N_5655,N_5711);
xnor U5984 (N_5984,N_5674,N_5699);
or U5985 (N_5985,N_5798,N_5661);
nand U5986 (N_5986,N_5774,N_5713);
xnor U5987 (N_5987,N_5617,N_5741);
xor U5988 (N_5988,N_5752,N_5798);
and U5989 (N_5989,N_5764,N_5605);
xnor U5990 (N_5990,N_5786,N_5707);
xnor U5991 (N_5991,N_5725,N_5769);
nor U5992 (N_5992,N_5612,N_5783);
and U5993 (N_5993,N_5660,N_5659);
nor U5994 (N_5994,N_5678,N_5629);
nand U5995 (N_5995,N_5697,N_5716);
or U5996 (N_5996,N_5747,N_5663);
or U5997 (N_5997,N_5603,N_5681);
xnor U5998 (N_5998,N_5676,N_5707);
xor U5999 (N_5999,N_5633,N_5685);
or U6000 (N_6000,N_5977,N_5934);
xnor U6001 (N_6001,N_5987,N_5899);
nand U6002 (N_6002,N_5989,N_5928);
or U6003 (N_6003,N_5932,N_5848);
or U6004 (N_6004,N_5971,N_5801);
nor U6005 (N_6005,N_5978,N_5804);
nor U6006 (N_6006,N_5853,N_5823);
nand U6007 (N_6007,N_5884,N_5918);
xor U6008 (N_6008,N_5850,N_5845);
and U6009 (N_6009,N_5811,N_5908);
nand U6010 (N_6010,N_5923,N_5861);
xor U6011 (N_6011,N_5844,N_5967);
and U6012 (N_6012,N_5951,N_5873);
xor U6013 (N_6013,N_5947,N_5935);
xnor U6014 (N_6014,N_5907,N_5886);
and U6015 (N_6015,N_5930,N_5986);
xnor U6016 (N_6016,N_5803,N_5877);
nor U6017 (N_6017,N_5810,N_5821);
or U6018 (N_6018,N_5917,N_5966);
xnor U6019 (N_6019,N_5852,N_5879);
xnor U6020 (N_6020,N_5817,N_5965);
nand U6021 (N_6021,N_5862,N_5842);
nor U6022 (N_6022,N_5936,N_5996);
nand U6023 (N_6023,N_5805,N_5968);
and U6024 (N_6024,N_5833,N_5822);
and U6025 (N_6025,N_5808,N_5984);
nor U6026 (N_6026,N_5855,N_5888);
nor U6027 (N_6027,N_5829,N_5800);
and U6028 (N_6028,N_5969,N_5938);
nand U6029 (N_6029,N_5948,N_5871);
or U6030 (N_6030,N_5913,N_5815);
xnor U6031 (N_6031,N_5953,N_5856);
nand U6032 (N_6032,N_5880,N_5919);
nand U6033 (N_6033,N_5992,N_5806);
or U6034 (N_6034,N_5922,N_5870);
nor U6035 (N_6035,N_5903,N_5997);
and U6036 (N_6036,N_5863,N_5854);
nand U6037 (N_6037,N_5824,N_5878);
or U6038 (N_6038,N_5820,N_5921);
nand U6039 (N_6039,N_5875,N_5836);
and U6040 (N_6040,N_5894,N_5991);
xor U6041 (N_6041,N_5892,N_5939);
or U6042 (N_6042,N_5976,N_5958);
nand U6043 (N_6043,N_5995,N_5979);
or U6044 (N_6044,N_5846,N_5883);
nand U6045 (N_6045,N_5956,N_5898);
nand U6046 (N_6046,N_5895,N_5905);
or U6047 (N_6047,N_5982,N_5999);
and U6048 (N_6048,N_5945,N_5837);
or U6049 (N_6049,N_5868,N_5915);
xnor U6050 (N_6050,N_5927,N_5835);
or U6051 (N_6051,N_5818,N_5857);
and U6052 (N_6052,N_5920,N_5813);
and U6053 (N_6053,N_5890,N_5866);
and U6054 (N_6054,N_5831,N_5975);
nor U6055 (N_6055,N_5906,N_5826);
nor U6056 (N_6056,N_5937,N_5802);
xnor U6057 (N_6057,N_5961,N_5942);
nand U6058 (N_6058,N_5914,N_5851);
nand U6059 (N_6059,N_5985,N_5974);
nor U6060 (N_6060,N_5893,N_5825);
and U6061 (N_6061,N_5944,N_5946);
xnor U6062 (N_6062,N_5807,N_5912);
nor U6063 (N_6063,N_5950,N_5859);
or U6064 (N_6064,N_5916,N_5839);
or U6065 (N_6065,N_5925,N_5955);
nor U6066 (N_6066,N_5902,N_5840);
or U6067 (N_6067,N_5819,N_5929);
or U6068 (N_6068,N_5973,N_5901);
nor U6069 (N_6069,N_5994,N_5891);
and U6070 (N_6070,N_5834,N_5876);
xor U6071 (N_6071,N_5943,N_5830);
nand U6072 (N_6072,N_5952,N_5954);
nor U6073 (N_6073,N_5972,N_5812);
and U6074 (N_6074,N_5814,N_5896);
xor U6075 (N_6075,N_5867,N_5990);
nand U6076 (N_6076,N_5869,N_5897);
nand U6077 (N_6077,N_5838,N_5887);
nand U6078 (N_6078,N_5963,N_5911);
and U6079 (N_6079,N_5988,N_5881);
xor U6080 (N_6080,N_5865,N_5832);
nor U6081 (N_6081,N_5885,N_5931);
nor U6082 (N_6082,N_5998,N_5981);
nor U6083 (N_6083,N_5809,N_5910);
nor U6084 (N_6084,N_5941,N_5860);
and U6085 (N_6085,N_5909,N_5957);
or U6086 (N_6086,N_5900,N_5864);
nand U6087 (N_6087,N_5827,N_5933);
nand U6088 (N_6088,N_5889,N_5959);
or U6089 (N_6089,N_5904,N_5847);
nand U6090 (N_6090,N_5962,N_5924);
nor U6091 (N_6091,N_5816,N_5858);
xnor U6092 (N_6092,N_5841,N_5882);
nor U6093 (N_6093,N_5960,N_5980);
or U6094 (N_6094,N_5828,N_5983);
nor U6095 (N_6095,N_5874,N_5970);
xnor U6096 (N_6096,N_5872,N_5843);
nand U6097 (N_6097,N_5993,N_5964);
and U6098 (N_6098,N_5940,N_5926);
nand U6099 (N_6099,N_5849,N_5949);
nor U6100 (N_6100,N_5932,N_5927);
nand U6101 (N_6101,N_5867,N_5974);
nor U6102 (N_6102,N_5940,N_5946);
xnor U6103 (N_6103,N_5977,N_5833);
nand U6104 (N_6104,N_5904,N_5956);
or U6105 (N_6105,N_5985,N_5971);
nand U6106 (N_6106,N_5982,N_5889);
and U6107 (N_6107,N_5928,N_5990);
and U6108 (N_6108,N_5939,N_5802);
or U6109 (N_6109,N_5832,N_5930);
or U6110 (N_6110,N_5855,N_5983);
and U6111 (N_6111,N_5821,N_5960);
xnor U6112 (N_6112,N_5970,N_5883);
nor U6113 (N_6113,N_5947,N_5905);
xnor U6114 (N_6114,N_5878,N_5816);
nor U6115 (N_6115,N_5947,N_5948);
or U6116 (N_6116,N_5918,N_5925);
or U6117 (N_6117,N_5929,N_5877);
or U6118 (N_6118,N_5881,N_5989);
and U6119 (N_6119,N_5883,N_5811);
xnor U6120 (N_6120,N_5927,N_5861);
or U6121 (N_6121,N_5878,N_5989);
and U6122 (N_6122,N_5967,N_5822);
or U6123 (N_6123,N_5975,N_5865);
xor U6124 (N_6124,N_5973,N_5869);
nor U6125 (N_6125,N_5840,N_5935);
nor U6126 (N_6126,N_5943,N_5850);
xnor U6127 (N_6127,N_5941,N_5844);
xor U6128 (N_6128,N_5935,N_5960);
and U6129 (N_6129,N_5998,N_5956);
and U6130 (N_6130,N_5923,N_5855);
or U6131 (N_6131,N_5829,N_5833);
nor U6132 (N_6132,N_5843,N_5988);
xnor U6133 (N_6133,N_5911,N_5993);
nand U6134 (N_6134,N_5937,N_5854);
and U6135 (N_6135,N_5866,N_5961);
and U6136 (N_6136,N_5955,N_5891);
xor U6137 (N_6137,N_5903,N_5917);
and U6138 (N_6138,N_5980,N_5986);
xnor U6139 (N_6139,N_5918,N_5934);
or U6140 (N_6140,N_5842,N_5899);
nand U6141 (N_6141,N_5822,N_5968);
and U6142 (N_6142,N_5805,N_5918);
and U6143 (N_6143,N_5977,N_5921);
nor U6144 (N_6144,N_5918,N_5814);
xor U6145 (N_6145,N_5825,N_5826);
xnor U6146 (N_6146,N_5813,N_5967);
nor U6147 (N_6147,N_5964,N_5844);
or U6148 (N_6148,N_5870,N_5891);
or U6149 (N_6149,N_5908,N_5857);
or U6150 (N_6150,N_5851,N_5936);
nor U6151 (N_6151,N_5807,N_5842);
nand U6152 (N_6152,N_5943,N_5867);
or U6153 (N_6153,N_5836,N_5876);
nand U6154 (N_6154,N_5860,N_5967);
and U6155 (N_6155,N_5943,N_5861);
and U6156 (N_6156,N_5956,N_5873);
nor U6157 (N_6157,N_5948,N_5998);
or U6158 (N_6158,N_5963,N_5939);
xor U6159 (N_6159,N_5820,N_5968);
or U6160 (N_6160,N_5801,N_5897);
or U6161 (N_6161,N_5923,N_5842);
nand U6162 (N_6162,N_5836,N_5890);
nand U6163 (N_6163,N_5853,N_5943);
and U6164 (N_6164,N_5853,N_5978);
and U6165 (N_6165,N_5853,N_5882);
and U6166 (N_6166,N_5860,N_5985);
xor U6167 (N_6167,N_5924,N_5857);
nand U6168 (N_6168,N_5886,N_5815);
and U6169 (N_6169,N_5822,N_5940);
and U6170 (N_6170,N_5900,N_5948);
nand U6171 (N_6171,N_5907,N_5998);
xor U6172 (N_6172,N_5903,N_5867);
or U6173 (N_6173,N_5867,N_5936);
nor U6174 (N_6174,N_5956,N_5841);
or U6175 (N_6175,N_5895,N_5808);
and U6176 (N_6176,N_5812,N_5956);
and U6177 (N_6177,N_5887,N_5807);
or U6178 (N_6178,N_5959,N_5848);
xnor U6179 (N_6179,N_5889,N_5868);
xnor U6180 (N_6180,N_5974,N_5865);
or U6181 (N_6181,N_5815,N_5963);
or U6182 (N_6182,N_5828,N_5848);
and U6183 (N_6183,N_5951,N_5801);
xor U6184 (N_6184,N_5893,N_5818);
nor U6185 (N_6185,N_5883,N_5937);
xnor U6186 (N_6186,N_5960,N_5996);
and U6187 (N_6187,N_5928,N_5821);
or U6188 (N_6188,N_5839,N_5800);
or U6189 (N_6189,N_5921,N_5817);
and U6190 (N_6190,N_5985,N_5818);
and U6191 (N_6191,N_5829,N_5968);
and U6192 (N_6192,N_5916,N_5803);
nor U6193 (N_6193,N_5808,N_5829);
and U6194 (N_6194,N_5845,N_5852);
or U6195 (N_6195,N_5872,N_5937);
nand U6196 (N_6196,N_5803,N_5940);
or U6197 (N_6197,N_5865,N_5914);
and U6198 (N_6198,N_5998,N_5852);
or U6199 (N_6199,N_5987,N_5901);
and U6200 (N_6200,N_6199,N_6073);
xnor U6201 (N_6201,N_6192,N_6191);
and U6202 (N_6202,N_6197,N_6116);
nand U6203 (N_6203,N_6034,N_6055);
nor U6204 (N_6204,N_6047,N_6112);
and U6205 (N_6205,N_6157,N_6097);
nand U6206 (N_6206,N_6148,N_6011);
or U6207 (N_6207,N_6059,N_6051);
or U6208 (N_6208,N_6198,N_6018);
or U6209 (N_6209,N_6124,N_6026);
and U6210 (N_6210,N_6162,N_6042);
and U6211 (N_6211,N_6096,N_6058);
and U6212 (N_6212,N_6091,N_6120);
nor U6213 (N_6213,N_6175,N_6138);
or U6214 (N_6214,N_6039,N_6159);
nand U6215 (N_6215,N_6040,N_6095);
xnor U6216 (N_6216,N_6065,N_6074);
or U6217 (N_6217,N_6114,N_6196);
nor U6218 (N_6218,N_6090,N_6113);
nor U6219 (N_6219,N_6105,N_6088);
nand U6220 (N_6220,N_6182,N_6109);
or U6221 (N_6221,N_6024,N_6083);
or U6222 (N_6222,N_6012,N_6045);
and U6223 (N_6223,N_6069,N_6160);
or U6224 (N_6224,N_6156,N_6053);
or U6225 (N_6225,N_6131,N_6004);
nand U6226 (N_6226,N_6079,N_6111);
nor U6227 (N_6227,N_6110,N_6136);
nor U6228 (N_6228,N_6032,N_6103);
nand U6229 (N_6229,N_6108,N_6021);
xor U6230 (N_6230,N_6005,N_6187);
nand U6231 (N_6231,N_6002,N_6128);
or U6232 (N_6232,N_6098,N_6019);
nand U6233 (N_6233,N_6142,N_6193);
and U6234 (N_6234,N_6106,N_6144);
xor U6235 (N_6235,N_6190,N_6031);
nor U6236 (N_6236,N_6117,N_6023);
or U6237 (N_6237,N_6094,N_6081);
xnor U6238 (N_6238,N_6022,N_6014);
or U6239 (N_6239,N_6037,N_6164);
nand U6240 (N_6240,N_6194,N_6089);
nor U6241 (N_6241,N_6028,N_6188);
or U6242 (N_6242,N_6167,N_6139);
nand U6243 (N_6243,N_6007,N_6183);
and U6244 (N_6244,N_6184,N_6086);
nand U6245 (N_6245,N_6102,N_6046);
and U6246 (N_6246,N_6115,N_6078);
xnor U6247 (N_6247,N_6072,N_6009);
and U6248 (N_6248,N_6177,N_6033);
and U6249 (N_6249,N_6143,N_6008);
xor U6250 (N_6250,N_6087,N_6010);
or U6251 (N_6251,N_6071,N_6025);
nand U6252 (N_6252,N_6101,N_6075);
or U6253 (N_6253,N_6125,N_6150);
or U6254 (N_6254,N_6063,N_6027);
xnor U6255 (N_6255,N_6048,N_6161);
nor U6256 (N_6256,N_6050,N_6153);
xnor U6257 (N_6257,N_6056,N_6186);
and U6258 (N_6258,N_6107,N_6060);
or U6259 (N_6259,N_6104,N_6080);
xnor U6260 (N_6260,N_6172,N_6146);
nor U6261 (N_6261,N_6171,N_6043);
xor U6262 (N_6262,N_6155,N_6070);
and U6263 (N_6263,N_6029,N_6154);
nor U6264 (N_6264,N_6038,N_6122);
or U6265 (N_6265,N_6147,N_6044);
nand U6266 (N_6266,N_6067,N_6126);
xor U6267 (N_6267,N_6016,N_6145);
nand U6268 (N_6268,N_6015,N_6163);
nand U6269 (N_6269,N_6176,N_6185);
xnor U6270 (N_6270,N_6030,N_6173);
and U6271 (N_6271,N_6179,N_6178);
nor U6272 (N_6272,N_6130,N_6062);
or U6273 (N_6273,N_6052,N_6166);
nor U6274 (N_6274,N_6001,N_6168);
nand U6275 (N_6275,N_6169,N_6100);
xor U6276 (N_6276,N_6049,N_6066);
nor U6277 (N_6277,N_6017,N_6134);
nor U6278 (N_6278,N_6123,N_6129);
xor U6279 (N_6279,N_6061,N_6180);
nand U6280 (N_6280,N_6174,N_6013);
nor U6281 (N_6281,N_6020,N_6152);
nor U6282 (N_6282,N_6127,N_6121);
or U6283 (N_6283,N_6170,N_6165);
or U6284 (N_6284,N_6141,N_6000);
or U6285 (N_6285,N_6064,N_6133);
or U6286 (N_6286,N_6099,N_6132);
and U6287 (N_6287,N_6093,N_6006);
nand U6288 (N_6288,N_6035,N_6092);
xor U6289 (N_6289,N_6054,N_6149);
nor U6290 (N_6290,N_6181,N_6189);
xnor U6291 (N_6291,N_6077,N_6151);
nor U6292 (N_6292,N_6003,N_6084);
xnor U6293 (N_6293,N_6036,N_6068);
nand U6294 (N_6294,N_6076,N_6085);
nor U6295 (N_6295,N_6119,N_6135);
xor U6296 (N_6296,N_6158,N_6118);
xnor U6297 (N_6297,N_6140,N_6137);
xnor U6298 (N_6298,N_6195,N_6082);
and U6299 (N_6299,N_6057,N_6041);
and U6300 (N_6300,N_6022,N_6092);
or U6301 (N_6301,N_6170,N_6041);
xor U6302 (N_6302,N_6175,N_6089);
xor U6303 (N_6303,N_6106,N_6146);
or U6304 (N_6304,N_6041,N_6075);
nand U6305 (N_6305,N_6069,N_6140);
nand U6306 (N_6306,N_6175,N_6158);
nor U6307 (N_6307,N_6071,N_6069);
or U6308 (N_6308,N_6050,N_6076);
nand U6309 (N_6309,N_6036,N_6075);
or U6310 (N_6310,N_6072,N_6136);
xnor U6311 (N_6311,N_6138,N_6107);
nor U6312 (N_6312,N_6078,N_6094);
nor U6313 (N_6313,N_6085,N_6082);
xor U6314 (N_6314,N_6106,N_6031);
and U6315 (N_6315,N_6128,N_6176);
and U6316 (N_6316,N_6146,N_6081);
and U6317 (N_6317,N_6015,N_6006);
nand U6318 (N_6318,N_6097,N_6047);
nor U6319 (N_6319,N_6089,N_6061);
nor U6320 (N_6320,N_6047,N_6039);
nor U6321 (N_6321,N_6102,N_6157);
nand U6322 (N_6322,N_6162,N_6012);
or U6323 (N_6323,N_6134,N_6075);
nand U6324 (N_6324,N_6038,N_6138);
and U6325 (N_6325,N_6196,N_6075);
and U6326 (N_6326,N_6046,N_6139);
xnor U6327 (N_6327,N_6078,N_6026);
and U6328 (N_6328,N_6060,N_6017);
and U6329 (N_6329,N_6152,N_6051);
xnor U6330 (N_6330,N_6125,N_6017);
nand U6331 (N_6331,N_6147,N_6011);
nand U6332 (N_6332,N_6018,N_6185);
nand U6333 (N_6333,N_6164,N_6170);
nor U6334 (N_6334,N_6054,N_6040);
nor U6335 (N_6335,N_6156,N_6040);
or U6336 (N_6336,N_6185,N_6074);
nor U6337 (N_6337,N_6090,N_6104);
xor U6338 (N_6338,N_6150,N_6073);
and U6339 (N_6339,N_6045,N_6189);
and U6340 (N_6340,N_6024,N_6181);
or U6341 (N_6341,N_6127,N_6186);
and U6342 (N_6342,N_6112,N_6067);
nor U6343 (N_6343,N_6071,N_6099);
xnor U6344 (N_6344,N_6131,N_6108);
and U6345 (N_6345,N_6153,N_6193);
xor U6346 (N_6346,N_6018,N_6088);
and U6347 (N_6347,N_6108,N_6050);
xnor U6348 (N_6348,N_6160,N_6166);
xnor U6349 (N_6349,N_6043,N_6090);
nor U6350 (N_6350,N_6063,N_6121);
or U6351 (N_6351,N_6192,N_6120);
or U6352 (N_6352,N_6047,N_6079);
nor U6353 (N_6353,N_6042,N_6093);
or U6354 (N_6354,N_6187,N_6032);
nand U6355 (N_6355,N_6167,N_6105);
or U6356 (N_6356,N_6163,N_6060);
nand U6357 (N_6357,N_6095,N_6193);
xnor U6358 (N_6358,N_6187,N_6139);
or U6359 (N_6359,N_6118,N_6192);
nand U6360 (N_6360,N_6132,N_6017);
nor U6361 (N_6361,N_6097,N_6144);
xnor U6362 (N_6362,N_6177,N_6083);
nor U6363 (N_6363,N_6073,N_6078);
xor U6364 (N_6364,N_6033,N_6094);
nor U6365 (N_6365,N_6147,N_6136);
xnor U6366 (N_6366,N_6129,N_6131);
nor U6367 (N_6367,N_6091,N_6002);
nand U6368 (N_6368,N_6130,N_6097);
nand U6369 (N_6369,N_6035,N_6093);
nor U6370 (N_6370,N_6048,N_6143);
nand U6371 (N_6371,N_6067,N_6014);
nand U6372 (N_6372,N_6021,N_6036);
or U6373 (N_6373,N_6160,N_6097);
nor U6374 (N_6374,N_6107,N_6156);
xnor U6375 (N_6375,N_6153,N_6163);
xnor U6376 (N_6376,N_6101,N_6019);
or U6377 (N_6377,N_6073,N_6138);
or U6378 (N_6378,N_6091,N_6197);
or U6379 (N_6379,N_6124,N_6054);
xnor U6380 (N_6380,N_6110,N_6117);
nor U6381 (N_6381,N_6123,N_6131);
nor U6382 (N_6382,N_6079,N_6013);
or U6383 (N_6383,N_6058,N_6130);
or U6384 (N_6384,N_6105,N_6193);
nor U6385 (N_6385,N_6047,N_6003);
nand U6386 (N_6386,N_6044,N_6111);
nand U6387 (N_6387,N_6130,N_6169);
or U6388 (N_6388,N_6099,N_6138);
or U6389 (N_6389,N_6119,N_6130);
or U6390 (N_6390,N_6148,N_6125);
nor U6391 (N_6391,N_6058,N_6044);
nor U6392 (N_6392,N_6121,N_6034);
or U6393 (N_6393,N_6101,N_6011);
xnor U6394 (N_6394,N_6107,N_6093);
nor U6395 (N_6395,N_6009,N_6063);
or U6396 (N_6396,N_6067,N_6108);
nand U6397 (N_6397,N_6045,N_6164);
xnor U6398 (N_6398,N_6119,N_6180);
nor U6399 (N_6399,N_6001,N_6151);
nand U6400 (N_6400,N_6351,N_6328);
nand U6401 (N_6401,N_6319,N_6338);
nor U6402 (N_6402,N_6244,N_6288);
or U6403 (N_6403,N_6321,N_6301);
nor U6404 (N_6404,N_6341,N_6245);
xor U6405 (N_6405,N_6370,N_6339);
and U6406 (N_6406,N_6377,N_6355);
nor U6407 (N_6407,N_6369,N_6205);
xor U6408 (N_6408,N_6248,N_6382);
and U6409 (N_6409,N_6327,N_6211);
nand U6410 (N_6410,N_6318,N_6208);
nor U6411 (N_6411,N_6395,N_6389);
nand U6412 (N_6412,N_6334,N_6232);
xnor U6413 (N_6413,N_6219,N_6368);
and U6414 (N_6414,N_6397,N_6345);
nor U6415 (N_6415,N_6293,N_6272);
nand U6416 (N_6416,N_6295,N_6216);
or U6417 (N_6417,N_6342,N_6343);
xor U6418 (N_6418,N_6383,N_6296);
nand U6419 (N_6419,N_6262,N_6267);
xnor U6420 (N_6420,N_6300,N_6200);
nor U6421 (N_6421,N_6276,N_6206);
or U6422 (N_6422,N_6354,N_6265);
xor U6423 (N_6423,N_6253,N_6239);
and U6424 (N_6424,N_6224,N_6212);
and U6425 (N_6425,N_6213,N_6278);
or U6426 (N_6426,N_6387,N_6376);
and U6427 (N_6427,N_6350,N_6258);
xnor U6428 (N_6428,N_6305,N_6357);
and U6429 (N_6429,N_6263,N_6203);
and U6430 (N_6430,N_6230,N_6303);
nand U6431 (N_6431,N_6307,N_6352);
nand U6432 (N_6432,N_6393,N_6252);
xnor U6433 (N_6433,N_6241,N_6392);
or U6434 (N_6434,N_6346,N_6375);
nand U6435 (N_6435,N_6283,N_6225);
xnor U6436 (N_6436,N_6396,N_6234);
nand U6437 (N_6437,N_6372,N_6240);
nand U6438 (N_6438,N_6201,N_6237);
and U6439 (N_6439,N_6246,N_6322);
and U6440 (N_6440,N_6209,N_6329);
or U6441 (N_6441,N_6381,N_6228);
and U6442 (N_6442,N_6227,N_6279);
or U6443 (N_6443,N_6259,N_6347);
or U6444 (N_6444,N_6348,N_6233);
and U6445 (N_6445,N_6226,N_6254);
nor U6446 (N_6446,N_6284,N_6344);
xor U6447 (N_6447,N_6380,N_6317);
nand U6448 (N_6448,N_6379,N_6310);
nand U6449 (N_6449,N_6314,N_6257);
nand U6450 (N_6450,N_6289,N_6332);
and U6451 (N_6451,N_6299,N_6269);
nand U6452 (N_6452,N_6362,N_6378);
or U6453 (N_6453,N_6371,N_6222);
xor U6454 (N_6454,N_6231,N_6330);
xnor U6455 (N_6455,N_6250,N_6353);
xor U6456 (N_6456,N_6275,N_6336);
nand U6457 (N_6457,N_6202,N_6360);
nand U6458 (N_6458,N_6210,N_6312);
or U6459 (N_6459,N_6358,N_6385);
xnor U6460 (N_6460,N_6294,N_6316);
nand U6461 (N_6461,N_6256,N_6242);
nor U6462 (N_6462,N_6388,N_6290);
nand U6463 (N_6463,N_6235,N_6308);
or U6464 (N_6464,N_6356,N_6217);
nor U6465 (N_6465,N_6340,N_6398);
xor U6466 (N_6466,N_6297,N_6333);
xor U6467 (N_6467,N_6298,N_6287);
or U6468 (N_6468,N_6249,N_6271);
or U6469 (N_6469,N_6320,N_6313);
or U6470 (N_6470,N_6363,N_6277);
or U6471 (N_6471,N_6238,N_6306);
xor U6472 (N_6472,N_6311,N_6280);
xor U6473 (N_6473,N_6251,N_6302);
and U6474 (N_6474,N_6266,N_6247);
or U6475 (N_6475,N_6325,N_6386);
nor U6476 (N_6476,N_6394,N_6229);
and U6477 (N_6477,N_6323,N_6391);
xnor U6478 (N_6478,N_6365,N_6291);
xnor U6479 (N_6479,N_6218,N_6292);
or U6480 (N_6480,N_6337,N_6282);
nand U6481 (N_6481,N_6373,N_6304);
and U6482 (N_6482,N_6207,N_6214);
nor U6483 (N_6483,N_6268,N_6384);
nor U6484 (N_6484,N_6309,N_6285);
and U6485 (N_6485,N_6215,N_6286);
or U6486 (N_6486,N_6335,N_6260);
or U6487 (N_6487,N_6255,N_6326);
nor U6488 (N_6488,N_6364,N_6243);
nand U6489 (N_6489,N_6361,N_6220);
nor U6490 (N_6490,N_6273,N_6270);
and U6491 (N_6491,N_6264,N_6324);
and U6492 (N_6492,N_6331,N_6390);
xor U6493 (N_6493,N_6349,N_6223);
xnor U6494 (N_6494,N_6261,N_6399);
xnor U6495 (N_6495,N_6374,N_6274);
and U6496 (N_6496,N_6315,N_6367);
nand U6497 (N_6497,N_6366,N_6281);
or U6498 (N_6498,N_6359,N_6236);
xor U6499 (N_6499,N_6221,N_6204);
xnor U6500 (N_6500,N_6301,N_6392);
nor U6501 (N_6501,N_6348,N_6388);
nand U6502 (N_6502,N_6307,N_6302);
xor U6503 (N_6503,N_6300,N_6236);
or U6504 (N_6504,N_6394,N_6248);
or U6505 (N_6505,N_6234,N_6229);
nor U6506 (N_6506,N_6334,N_6390);
nand U6507 (N_6507,N_6328,N_6378);
or U6508 (N_6508,N_6232,N_6363);
nor U6509 (N_6509,N_6259,N_6210);
nand U6510 (N_6510,N_6376,N_6213);
nor U6511 (N_6511,N_6207,N_6387);
and U6512 (N_6512,N_6270,N_6220);
or U6513 (N_6513,N_6313,N_6312);
nand U6514 (N_6514,N_6288,N_6366);
nor U6515 (N_6515,N_6264,N_6260);
nor U6516 (N_6516,N_6246,N_6332);
nor U6517 (N_6517,N_6333,N_6291);
nand U6518 (N_6518,N_6289,N_6229);
nand U6519 (N_6519,N_6291,N_6367);
xnor U6520 (N_6520,N_6375,N_6202);
and U6521 (N_6521,N_6258,N_6319);
nand U6522 (N_6522,N_6245,N_6292);
nor U6523 (N_6523,N_6303,N_6247);
xnor U6524 (N_6524,N_6273,N_6309);
and U6525 (N_6525,N_6305,N_6211);
xnor U6526 (N_6526,N_6211,N_6291);
nand U6527 (N_6527,N_6283,N_6246);
and U6528 (N_6528,N_6285,N_6303);
and U6529 (N_6529,N_6383,N_6328);
nand U6530 (N_6530,N_6290,N_6377);
and U6531 (N_6531,N_6248,N_6299);
xor U6532 (N_6532,N_6213,N_6342);
and U6533 (N_6533,N_6333,N_6316);
or U6534 (N_6534,N_6248,N_6334);
xnor U6535 (N_6535,N_6305,N_6208);
or U6536 (N_6536,N_6363,N_6348);
and U6537 (N_6537,N_6336,N_6295);
or U6538 (N_6538,N_6257,N_6234);
and U6539 (N_6539,N_6322,N_6326);
and U6540 (N_6540,N_6271,N_6216);
nor U6541 (N_6541,N_6286,N_6219);
and U6542 (N_6542,N_6221,N_6313);
nor U6543 (N_6543,N_6254,N_6386);
nand U6544 (N_6544,N_6363,N_6203);
nand U6545 (N_6545,N_6381,N_6274);
nand U6546 (N_6546,N_6355,N_6252);
nor U6547 (N_6547,N_6372,N_6296);
or U6548 (N_6548,N_6292,N_6210);
xnor U6549 (N_6549,N_6280,N_6220);
nor U6550 (N_6550,N_6369,N_6331);
xnor U6551 (N_6551,N_6336,N_6351);
and U6552 (N_6552,N_6336,N_6342);
or U6553 (N_6553,N_6303,N_6301);
and U6554 (N_6554,N_6218,N_6397);
nand U6555 (N_6555,N_6376,N_6243);
nor U6556 (N_6556,N_6306,N_6200);
and U6557 (N_6557,N_6297,N_6235);
and U6558 (N_6558,N_6375,N_6252);
nor U6559 (N_6559,N_6278,N_6382);
xor U6560 (N_6560,N_6377,N_6261);
nor U6561 (N_6561,N_6350,N_6375);
nor U6562 (N_6562,N_6362,N_6268);
nand U6563 (N_6563,N_6344,N_6210);
or U6564 (N_6564,N_6252,N_6295);
or U6565 (N_6565,N_6296,N_6371);
nand U6566 (N_6566,N_6259,N_6215);
nor U6567 (N_6567,N_6381,N_6233);
nand U6568 (N_6568,N_6224,N_6259);
nor U6569 (N_6569,N_6392,N_6319);
and U6570 (N_6570,N_6360,N_6358);
xor U6571 (N_6571,N_6268,N_6228);
nand U6572 (N_6572,N_6201,N_6271);
and U6573 (N_6573,N_6260,N_6390);
nor U6574 (N_6574,N_6290,N_6246);
or U6575 (N_6575,N_6374,N_6264);
xor U6576 (N_6576,N_6338,N_6259);
or U6577 (N_6577,N_6235,N_6204);
and U6578 (N_6578,N_6281,N_6207);
or U6579 (N_6579,N_6399,N_6300);
and U6580 (N_6580,N_6397,N_6371);
and U6581 (N_6581,N_6215,N_6228);
or U6582 (N_6582,N_6236,N_6336);
nand U6583 (N_6583,N_6212,N_6213);
nand U6584 (N_6584,N_6217,N_6204);
and U6585 (N_6585,N_6383,N_6330);
nor U6586 (N_6586,N_6265,N_6209);
nor U6587 (N_6587,N_6261,N_6255);
xnor U6588 (N_6588,N_6365,N_6230);
nand U6589 (N_6589,N_6354,N_6344);
nor U6590 (N_6590,N_6214,N_6363);
nand U6591 (N_6591,N_6224,N_6314);
nor U6592 (N_6592,N_6368,N_6338);
nor U6593 (N_6593,N_6395,N_6398);
nand U6594 (N_6594,N_6339,N_6262);
and U6595 (N_6595,N_6285,N_6282);
and U6596 (N_6596,N_6258,N_6378);
xnor U6597 (N_6597,N_6273,N_6259);
nand U6598 (N_6598,N_6230,N_6367);
and U6599 (N_6599,N_6316,N_6370);
xor U6600 (N_6600,N_6494,N_6537);
or U6601 (N_6601,N_6485,N_6502);
and U6602 (N_6602,N_6512,N_6416);
nand U6603 (N_6603,N_6409,N_6520);
or U6604 (N_6604,N_6463,N_6572);
nor U6605 (N_6605,N_6513,N_6426);
nand U6606 (N_6606,N_6548,N_6473);
or U6607 (N_6607,N_6497,N_6425);
xnor U6608 (N_6608,N_6431,N_6533);
nor U6609 (N_6609,N_6436,N_6449);
nor U6610 (N_6610,N_6508,N_6484);
and U6611 (N_6611,N_6458,N_6408);
or U6612 (N_6612,N_6529,N_6570);
xnor U6613 (N_6613,N_6596,N_6546);
nand U6614 (N_6614,N_6454,N_6551);
xor U6615 (N_6615,N_6578,N_6510);
or U6616 (N_6616,N_6523,N_6585);
or U6617 (N_6617,N_6465,N_6536);
and U6618 (N_6618,N_6500,N_6450);
and U6619 (N_6619,N_6507,N_6549);
nand U6620 (N_6620,N_6437,N_6555);
xor U6621 (N_6621,N_6595,N_6525);
nor U6622 (N_6622,N_6453,N_6574);
xnor U6623 (N_6623,N_6582,N_6417);
nor U6624 (N_6624,N_6557,N_6519);
or U6625 (N_6625,N_6486,N_6491);
xnor U6626 (N_6626,N_6418,N_6407);
xor U6627 (N_6627,N_6489,N_6438);
nand U6628 (N_6628,N_6590,N_6569);
xor U6629 (N_6629,N_6597,N_6580);
xor U6630 (N_6630,N_6543,N_6444);
nor U6631 (N_6631,N_6492,N_6400);
xnor U6632 (N_6632,N_6581,N_6579);
and U6633 (N_6633,N_6565,N_6493);
nor U6634 (N_6634,N_6411,N_6477);
xnor U6635 (N_6635,N_6479,N_6427);
nor U6636 (N_6636,N_6464,N_6552);
and U6637 (N_6637,N_6499,N_6422);
nand U6638 (N_6638,N_6506,N_6560);
nor U6639 (N_6639,N_6440,N_6429);
or U6640 (N_6640,N_6448,N_6592);
xor U6641 (N_6641,N_6490,N_6526);
or U6642 (N_6642,N_6412,N_6594);
and U6643 (N_6643,N_6583,N_6511);
and U6644 (N_6644,N_6474,N_6577);
nor U6645 (N_6645,N_6567,N_6547);
nor U6646 (N_6646,N_6562,N_6466);
or U6647 (N_6647,N_6591,N_6470);
xnor U6648 (N_6648,N_6521,N_6472);
and U6649 (N_6649,N_6541,N_6455);
or U6650 (N_6650,N_6535,N_6446);
or U6651 (N_6651,N_6419,N_6542);
or U6652 (N_6652,N_6584,N_6403);
or U6653 (N_6653,N_6530,N_6401);
nor U6654 (N_6654,N_6563,N_6517);
nand U6655 (N_6655,N_6571,N_6532);
or U6656 (N_6656,N_6435,N_6404);
nor U6657 (N_6657,N_6524,N_6568);
or U6658 (N_6658,N_6576,N_6516);
xnor U6659 (N_6659,N_6468,N_6588);
and U6660 (N_6660,N_6566,N_6545);
and U6661 (N_6661,N_6573,N_6503);
xor U6662 (N_6662,N_6564,N_6456);
nand U6663 (N_6663,N_6501,N_6505);
nor U6664 (N_6664,N_6405,N_6406);
and U6665 (N_6665,N_6462,N_6522);
nor U6666 (N_6666,N_6561,N_6527);
nor U6667 (N_6667,N_6488,N_6553);
or U6668 (N_6668,N_6586,N_6478);
nor U6669 (N_6669,N_6447,N_6498);
xnor U6670 (N_6670,N_6460,N_6558);
nor U6671 (N_6671,N_6415,N_6487);
xor U6672 (N_6672,N_6504,N_6480);
or U6673 (N_6673,N_6424,N_6538);
or U6674 (N_6674,N_6593,N_6413);
nor U6675 (N_6675,N_6589,N_6481);
nor U6676 (N_6676,N_6534,N_6539);
nor U6677 (N_6677,N_6528,N_6559);
xnor U6678 (N_6678,N_6442,N_6515);
and U6679 (N_6679,N_6414,N_6475);
or U6680 (N_6680,N_6482,N_6509);
nand U6681 (N_6681,N_6430,N_6439);
nand U6682 (N_6682,N_6434,N_6518);
nor U6683 (N_6683,N_6445,N_6540);
nand U6684 (N_6684,N_6495,N_6459);
nand U6685 (N_6685,N_6469,N_6467);
xnor U6686 (N_6686,N_6441,N_6575);
xnor U6687 (N_6687,N_6420,N_6514);
nor U6688 (N_6688,N_6457,N_6421);
nand U6689 (N_6689,N_6554,N_6550);
or U6690 (N_6690,N_6443,N_6428);
nand U6691 (N_6691,N_6476,N_6483);
xnor U6692 (N_6692,N_6471,N_6461);
or U6693 (N_6693,N_6587,N_6531);
nand U6694 (N_6694,N_6599,N_6598);
or U6695 (N_6695,N_6496,N_6433);
nand U6696 (N_6696,N_6432,N_6451);
nand U6697 (N_6697,N_6402,N_6544);
xor U6698 (N_6698,N_6423,N_6410);
or U6699 (N_6699,N_6452,N_6556);
xnor U6700 (N_6700,N_6513,N_6526);
or U6701 (N_6701,N_6576,N_6424);
nor U6702 (N_6702,N_6417,N_6465);
or U6703 (N_6703,N_6478,N_6444);
nor U6704 (N_6704,N_6575,N_6570);
and U6705 (N_6705,N_6569,N_6424);
or U6706 (N_6706,N_6557,N_6461);
nor U6707 (N_6707,N_6507,N_6438);
nor U6708 (N_6708,N_6490,N_6458);
or U6709 (N_6709,N_6420,N_6435);
xor U6710 (N_6710,N_6506,N_6492);
and U6711 (N_6711,N_6549,N_6476);
and U6712 (N_6712,N_6557,N_6507);
xor U6713 (N_6713,N_6578,N_6522);
and U6714 (N_6714,N_6542,N_6566);
xor U6715 (N_6715,N_6532,N_6410);
or U6716 (N_6716,N_6488,N_6538);
or U6717 (N_6717,N_6566,N_6498);
nand U6718 (N_6718,N_6419,N_6493);
nand U6719 (N_6719,N_6496,N_6516);
nand U6720 (N_6720,N_6461,N_6457);
nor U6721 (N_6721,N_6460,N_6458);
nand U6722 (N_6722,N_6497,N_6586);
xnor U6723 (N_6723,N_6457,N_6433);
or U6724 (N_6724,N_6484,N_6549);
and U6725 (N_6725,N_6555,N_6451);
nand U6726 (N_6726,N_6579,N_6573);
or U6727 (N_6727,N_6504,N_6521);
and U6728 (N_6728,N_6571,N_6512);
xor U6729 (N_6729,N_6467,N_6516);
or U6730 (N_6730,N_6526,N_6546);
nand U6731 (N_6731,N_6483,N_6529);
or U6732 (N_6732,N_6534,N_6552);
xor U6733 (N_6733,N_6515,N_6478);
nand U6734 (N_6734,N_6439,N_6464);
nand U6735 (N_6735,N_6566,N_6534);
nor U6736 (N_6736,N_6584,N_6423);
or U6737 (N_6737,N_6403,N_6506);
nand U6738 (N_6738,N_6521,N_6482);
xor U6739 (N_6739,N_6467,N_6542);
nor U6740 (N_6740,N_6518,N_6425);
nor U6741 (N_6741,N_6582,N_6599);
or U6742 (N_6742,N_6447,N_6516);
nor U6743 (N_6743,N_6471,N_6513);
xnor U6744 (N_6744,N_6492,N_6508);
nand U6745 (N_6745,N_6453,N_6580);
nor U6746 (N_6746,N_6579,N_6421);
nand U6747 (N_6747,N_6539,N_6443);
nor U6748 (N_6748,N_6415,N_6458);
and U6749 (N_6749,N_6451,N_6429);
and U6750 (N_6750,N_6472,N_6542);
and U6751 (N_6751,N_6538,N_6465);
nor U6752 (N_6752,N_6430,N_6402);
nand U6753 (N_6753,N_6523,N_6427);
nand U6754 (N_6754,N_6449,N_6493);
nor U6755 (N_6755,N_6566,N_6403);
xnor U6756 (N_6756,N_6469,N_6422);
and U6757 (N_6757,N_6515,N_6422);
nand U6758 (N_6758,N_6566,N_6453);
nor U6759 (N_6759,N_6591,N_6435);
or U6760 (N_6760,N_6402,N_6462);
and U6761 (N_6761,N_6599,N_6436);
nor U6762 (N_6762,N_6545,N_6528);
or U6763 (N_6763,N_6440,N_6435);
nand U6764 (N_6764,N_6476,N_6502);
or U6765 (N_6765,N_6494,N_6473);
and U6766 (N_6766,N_6504,N_6454);
or U6767 (N_6767,N_6595,N_6506);
nand U6768 (N_6768,N_6430,N_6499);
nor U6769 (N_6769,N_6592,N_6462);
or U6770 (N_6770,N_6537,N_6459);
xnor U6771 (N_6771,N_6535,N_6519);
nand U6772 (N_6772,N_6462,N_6575);
and U6773 (N_6773,N_6470,N_6482);
and U6774 (N_6774,N_6553,N_6521);
and U6775 (N_6775,N_6543,N_6552);
nand U6776 (N_6776,N_6434,N_6503);
nand U6777 (N_6777,N_6525,N_6484);
and U6778 (N_6778,N_6492,N_6523);
and U6779 (N_6779,N_6477,N_6573);
or U6780 (N_6780,N_6404,N_6414);
nor U6781 (N_6781,N_6550,N_6473);
nand U6782 (N_6782,N_6437,N_6567);
nand U6783 (N_6783,N_6557,N_6411);
nand U6784 (N_6784,N_6521,N_6544);
and U6785 (N_6785,N_6481,N_6568);
and U6786 (N_6786,N_6439,N_6451);
and U6787 (N_6787,N_6491,N_6448);
nor U6788 (N_6788,N_6460,N_6438);
nand U6789 (N_6789,N_6462,N_6596);
nand U6790 (N_6790,N_6595,N_6519);
nand U6791 (N_6791,N_6466,N_6504);
nor U6792 (N_6792,N_6496,N_6464);
xor U6793 (N_6793,N_6435,N_6521);
nand U6794 (N_6794,N_6576,N_6401);
or U6795 (N_6795,N_6540,N_6511);
nor U6796 (N_6796,N_6499,N_6445);
xor U6797 (N_6797,N_6439,N_6542);
nand U6798 (N_6798,N_6550,N_6423);
or U6799 (N_6799,N_6488,N_6591);
nor U6800 (N_6800,N_6774,N_6655);
xor U6801 (N_6801,N_6668,N_6612);
nor U6802 (N_6802,N_6769,N_6605);
xnor U6803 (N_6803,N_6737,N_6681);
nand U6804 (N_6804,N_6758,N_6771);
nand U6805 (N_6805,N_6635,N_6709);
or U6806 (N_6806,N_6613,N_6706);
nand U6807 (N_6807,N_6784,N_6670);
xor U6808 (N_6808,N_6671,N_6763);
nor U6809 (N_6809,N_6750,N_6632);
or U6810 (N_6810,N_6779,N_6694);
and U6811 (N_6811,N_6646,N_6625);
and U6812 (N_6812,N_6678,N_6796);
xnor U6813 (N_6813,N_6778,N_6773);
and U6814 (N_6814,N_6744,N_6777);
nor U6815 (N_6815,N_6700,N_6759);
and U6816 (N_6816,N_6720,N_6661);
nand U6817 (N_6817,N_6703,N_6718);
and U6818 (N_6818,N_6667,N_6641);
nand U6819 (N_6819,N_6740,N_6716);
xnor U6820 (N_6820,N_6672,N_6757);
nor U6821 (N_6821,N_6658,N_6696);
xnor U6822 (N_6822,N_6618,N_6787);
nor U6823 (N_6823,N_6653,N_6620);
and U6824 (N_6824,N_6719,N_6747);
nor U6825 (N_6825,N_6637,N_6665);
nand U6826 (N_6826,N_6776,N_6765);
nand U6827 (N_6827,N_6639,N_6663);
and U6828 (N_6828,N_6725,N_6628);
nand U6829 (N_6829,N_6659,N_6664);
nand U6830 (N_6830,N_6697,N_6735);
nor U6831 (N_6831,N_6723,N_6752);
or U6832 (N_6832,N_6600,N_6794);
nor U6833 (N_6833,N_6617,N_6609);
xnor U6834 (N_6834,N_6698,N_6679);
and U6835 (N_6835,N_6680,N_6645);
or U6836 (N_6836,N_6644,N_6691);
nand U6837 (N_6837,N_6627,N_6614);
nand U6838 (N_6838,N_6756,N_6767);
xnor U6839 (N_6839,N_6751,N_6669);
xnor U6840 (N_6840,N_6781,N_6733);
nand U6841 (N_6841,N_6676,N_6687);
or U6842 (N_6842,N_6761,N_6651);
nand U6843 (N_6843,N_6768,N_6708);
or U6844 (N_6844,N_6713,N_6690);
nor U6845 (N_6845,N_6638,N_6604);
nor U6846 (N_6846,N_6660,N_6746);
and U6847 (N_6847,N_6795,N_6792);
or U6848 (N_6848,N_6607,N_6724);
or U6849 (N_6849,N_6775,N_6707);
and U6850 (N_6850,N_6657,N_6745);
or U6851 (N_6851,N_6754,N_6630);
or U6852 (N_6852,N_6726,N_6710);
nor U6853 (N_6853,N_6755,N_6610);
xor U6854 (N_6854,N_6608,N_6730);
and U6855 (N_6855,N_6798,N_6729);
xnor U6856 (N_6856,N_6674,N_6673);
or U6857 (N_6857,N_6712,N_6626);
xor U6858 (N_6858,N_6647,N_6788);
and U6859 (N_6859,N_6766,N_6743);
xnor U6860 (N_6860,N_6685,N_6602);
nand U6861 (N_6861,N_6714,N_6790);
and U6862 (N_6862,N_6783,N_6749);
or U6863 (N_6863,N_6722,N_6793);
xor U6864 (N_6864,N_6616,N_6705);
or U6865 (N_6865,N_6699,N_6686);
nand U6866 (N_6866,N_6736,N_6636);
or U6867 (N_6867,N_6677,N_6715);
or U6868 (N_6868,N_6601,N_6643);
nand U6869 (N_6869,N_6764,N_6684);
or U6870 (N_6870,N_6695,N_6654);
or U6871 (N_6871,N_6634,N_6799);
xor U6872 (N_6872,N_6770,N_6782);
nor U6873 (N_6873,N_6739,N_6619);
nor U6874 (N_6874,N_6785,N_6762);
xor U6875 (N_6875,N_6732,N_6615);
and U6876 (N_6876,N_6780,N_6622);
or U6877 (N_6877,N_6675,N_6689);
nand U6878 (N_6878,N_6742,N_6666);
xnor U6879 (N_6879,N_6789,N_6649);
and U6880 (N_6880,N_6760,N_6688);
xnor U6881 (N_6881,N_6711,N_6631);
or U6882 (N_6882,N_6721,N_6734);
nor U6883 (N_6883,N_6731,N_6648);
and U6884 (N_6884,N_6603,N_6797);
xor U6885 (N_6885,N_6623,N_6633);
or U6886 (N_6886,N_6692,N_6704);
and U6887 (N_6887,N_6683,N_6786);
nand U6888 (N_6888,N_6753,N_6642);
and U6889 (N_6889,N_6741,N_6640);
nor U6890 (N_6890,N_6702,N_6791);
nor U6891 (N_6891,N_6728,N_6727);
nand U6892 (N_6892,N_6772,N_6717);
and U6893 (N_6893,N_6606,N_6611);
or U6894 (N_6894,N_6738,N_6652);
nand U6895 (N_6895,N_6650,N_6748);
xnor U6896 (N_6896,N_6656,N_6629);
nor U6897 (N_6897,N_6624,N_6682);
and U6898 (N_6898,N_6621,N_6701);
or U6899 (N_6899,N_6693,N_6662);
or U6900 (N_6900,N_6673,N_6775);
and U6901 (N_6901,N_6741,N_6687);
xnor U6902 (N_6902,N_6630,N_6658);
nor U6903 (N_6903,N_6677,N_6763);
and U6904 (N_6904,N_6766,N_6741);
nor U6905 (N_6905,N_6766,N_6670);
or U6906 (N_6906,N_6706,N_6737);
or U6907 (N_6907,N_6610,N_6762);
and U6908 (N_6908,N_6783,N_6710);
or U6909 (N_6909,N_6625,N_6618);
or U6910 (N_6910,N_6694,N_6728);
and U6911 (N_6911,N_6798,N_6762);
or U6912 (N_6912,N_6662,N_6730);
nor U6913 (N_6913,N_6763,N_6675);
nor U6914 (N_6914,N_6744,N_6654);
or U6915 (N_6915,N_6758,N_6687);
or U6916 (N_6916,N_6642,N_6776);
and U6917 (N_6917,N_6637,N_6730);
nor U6918 (N_6918,N_6679,N_6660);
nor U6919 (N_6919,N_6626,N_6708);
xor U6920 (N_6920,N_6749,N_6686);
xor U6921 (N_6921,N_6755,N_6699);
nor U6922 (N_6922,N_6681,N_6643);
or U6923 (N_6923,N_6629,N_6610);
and U6924 (N_6924,N_6762,N_6615);
nor U6925 (N_6925,N_6618,N_6679);
nand U6926 (N_6926,N_6755,N_6739);
nor U6927 (N_6927,N_6784,N_6794);
or U6928 (N_6928,N_6720,N_6642);
nor U6929 (N_6929,N_6678,N_6784);
and U6930 (N_6930,N_6768,N_6747);
nand U6931 (N_6931,N_6742,N_6637);
nor U6932 (N_6932,N_6737,N_6779);
and U6933 (N_6933,N_6799,N_6731);
or U6934 (N_6934,N_6764,N_6624);
or U6935 (N_6935,N_6707,N_6756);
or U6936 (N_6936,N_6637,N_6649);
and U6937 (N_6937,N_6632,N_6615);
and U6938 (N_6938,N_6629,N_6766);
or U6939 (N_6939,N_6786,N_6678);
nor U6940 (N_6940,N_6782,N_6748);
or U6941 (N_6941,N_6713,N_6781);
and U6942 (N_6942,N_6728,N_6609);
xor U6943 (N_6943,N_6719,N_6623);
and U6944 (N_6944,N_6617,N_6661);
nor U6945 (N_6945,N_6783,N_6773);
or U6946 (N_6946,N_6687,N_6772);
nor U6947 (N_6947,N_6795,N_6713);
nor U6948 (N_6948,N_6688,N_6602);
xnor U6949 (N_6949,N_6733,N_6729);
nor U6950 (N_6950,N_6620,N_6693);
nand U6951 (N_6951,N_6642,N_6728);
or U6952 (N_6952,N_6670,N_6688);
nor U6953 (N_6953,N_6778,N_6704);
xor U6954 (N_6954,N_6796,N_6753);
or U6955 (N_6955,N_6757,N_6713);
xnor U6956 (N_6956,N_6761,N_6779);
nand U6957 (N_6957,N_6709,N_6741);
xnor U6958 (N_6958,N_6778,N_6692);
nand U6959 (N_6959,N_6600,N_6646);
or U6960 (N_6960,N_6775,N_6727);
nand U6961 (N_6961,N_6671,N_6701);
and U6962 (N_6962,N_6743,N_6685);
or U6963 (N_6963,N_6655,N_6730);
or U6964 (N_6964,N_6644,N_6635);
xor U6965 (N_6965,N_6610,N_6627);
xor U6966 (N_6966,N_6620,N_6692);
nand U6967 (N_6967,N_6735,N_6765);
nand U6968 (N_6968,N_6683,N_6600);
nor U6969 (N_6969,N_6723,N_6748);
or U6970 (N_6970,N_6697,N_6798);
nor U6971 (N_6971,N_6620,N_6783);
nand U6972 (N_6972,N_6696,N_6793);
and U6973 (N_6973,N_6729,N_6751);
and U6974 (N_6974,N_6709,N_6752);
xnor U6975 (N_6975,N_6752,N_6757);
nor U6976 (N_6976,N_6613,N_6754);
nor U6977 (N_6977,N_6750,N_6759);
and U6978 (N_6978,N_6655,N_6639);
and U6979 (N_6979,N_6603,N_6657);
nand U6980 (N_6980,N_6644,N_6679);
xor U6981 (N_6981,N_6660,N_6771);
nor U6982 (N_6982,N_6762,N_6651);
nor U6983 (N_6983,N_6744,N_6670);
xor U6984 (N_6984,N_6612,N_6721);
nor U6985 (N_6985,N_6726,N_6773);
xor U6986 (N_6986,N_6738,N_6719);
or U6987 (N_6987,N_6662,N_6631);
and U6988 (N_6988,N_6674,N_6749);
xnor U6989 (N_6989,N_6791,N_6795);
and U6990 (N_6990,N_6663,N_6733);
nand U6991 (N_6991,N_6657,N_6795);
or U6992 (N_6992,N_6626,N_6655);
and U6993 (N_6993,N_6708,N_6667);
nor U6994 (N_6994,N_6630,N_6611);
xor U6995 (N_6995,N_6683,N_6729);
nand U6996 (N_6996,N_6784,N_6756);
nor U6997 (N_6997,N_6631,N_6796);
or U6998 (N_6998,N_6632,N_6635);
nor U6999 (N_6999,N_6602,N_6708);
xnor U7000 (N_7000,N_6955,N_6985);
nand U7001 (N_7001,N_6853,N_6967);
xnor U7002 (N_7002,N_6929,N_6839);
or U7003 (N_7003,N_6976,N_6942);
and U7004 (N_7004,N_6886,N_6810);
nand U7005 (N_7005,N_6861,N_6895);
or U7006 (N_7006,N_6969,N_6872);
and U7007 (N_7007,N_6952,N_6892);
or U7008 (N_7008,N_6846,N_6877);
nor U7009 (N_7009,N_6897,N_6937);
nand U7010 (N_7010,N_6960,N_6978);
or U7011 (N_7011,N_6984,N_6820);
xor U7012 (N_7012,N_6857,N_6855);
and U7013 (N_7013,N_6873,N_6858);
or U7014 (N_7014,N_6815,N_6860);
and U7015 (N_7015,N_6808,N_6830);
xnor U7016 (N_7016,N_6849,N_6851);
or U7017 (N_7017,N_6874,N_6871);
and U7018 (N_7018,N_6946,N_6910);
nand U7019 (N_7019,N_6829,N_6993);
and U7020 (N_7020,N_6866,N_6932);
and U7021 (N_7021,N_6826,N_6896);
or U7022 (N_7022,N_6919,N_6838);
xnor U7023 (N_7023,N_6828,N_6922);
or U7024 (N_7024,N_6903,N_6887);
nor U7025 (N_7025,N_6805,N_6876);
xor U7026 (N_7026,N_6834,N_6819);
nor U7027 (N_7027,N_6804,N_6814);
and U7028 (N_7028,N_6812,N_6987);
and U7029 (N_7029,N_6974,N_6850);
xor U7030 (N_7030,N_6862,N_6962);
or U7031 (N_7031,N_6904,N_6990);
xnor U7032 (N_7032,N_6822,N_6816);
xor U7033 (N_7033,N_6881,N_6868);
or U7034 (N_7034,N_6807,N_6856);
nand U7035 (N_7035,N_6923,N_6931);
and U7036 (N_7036,N_6833,N_6803);
and U7037 (N_7037,N_6912,N_6977);
xor U7038 (N_7038,N_6933,N_6940);
nor U7039 (N_7039,N_6869,N_6949);
nand U7040 (N_7040,N_6813,N_6864);
nor U7041 (N_7041,N_6821,N_6840);
nor U7042 (N_7042,N_6885,N_6883);
nor U7043 (N_7043,N_6947,N_6843);
nor U7044 (N_7044,N_6842,N_6863);
or U7045 (N_7045,N_6859,N_6806);
nor U7046 (N_7046,N_6844,N_6920);
xor U7047 (N_7047,N_6953,N_6988);
or U7048 (N_7048,N_6907,N_6818);
xnor U7049 (N_7049,N_6802,N_6957);
nor U7050 (N_7050,N_6964,N_6831);
nor U7051 (N_7051,N_6894,N_6956);
and U7052 (N_7052,N_6837,N_6906);
or U7053 (N_7053,N_6884,N_6888);
xnor U7054 (N_7054,N_6971,N_6836);
nor U7055 (N_7055,N_6994,N_6898);
or U7056 (N_7056,N_6880,N_6824);
xnor U7057 (N_7057,N_6823,N_6916);
and U7058 (N_7058,N_6944,N_6909);
xnor U7059 (N_7059,N_6961,N_6914);
or U7060 (N_7060,N_6878,N_6954);
xnor U7061 (N_7061,N_6986,N_6998);
nand U7062 (N_7062,N_6867,N_6926);
and U7063 (N_7063,N_6958,N_6845);
and U7064 (N_7064,N_6983,N_6973);
and U7065 (N_7065,N_6852,N_6827);
and U7066 (N_7066,N_6901,N_6848);
and U7067 (N_7067,N_6975,N_6902);
nand U7068 (N_7068,N_6948,N_6825);
and U7069 (N_7069,N_6832,N_6917);
or U7070 (N_7070,N_6911,N_6970);
nand U7071 (N_7071,N_6999,N_6890);
and U7072 (N_7072,N_6870,N_6968);
and U7073 (N_7073,N_6879,N_6981);
nor U7074 (N_7074,N_6889,N_6924);
or U7075 (N_7075,N_6921,N_6801);
nand U7076 (N_7076,N_6927,N_6979);
and U7077 (N_7077,N_6972,N_6966);
nor U7078 (N_7078,N_6905,N_6908);
and U7079 (N_7079,N_6800,N_6930);
nand U7080 (N_7080,N_6959,N_6939);
xnor U7081 (N_7081,N_6950,N_6951);
or U7082 (N_7082,N_6915,N_6963);
nand U7083 (N_7083,N_6945,N_6989);
xor U7084 (N_7084,N_6900,N_6817);
nand U7085 (N_7085,N_6882,N_6925);
nor U7086 (N_7086,N_6982,N_6891);
nor U7087 (N_7087,N_6928,N_6943);
or U7088 (N_7088,N_6899,N_6835);
nand U7089 (N_7089,N_6865,N_6938);
nand U7090 (N_7090,N_6991,N_6847);
nand U7091 (N_7091,N_6997,N_6809);
and U7092 (N_7092,N_6995,N_6996);
xor U7093 (N_7093,N_6980,N_6841);
and U7094 (N_7094,N_6854,N_6935);
xor U7095 (N_7095,N_6811,N_6936);
xnor U7096 (N_7096,N_6893,N_6875);
and U7097 (N_7097,N_6918,N_6941);
nand U7098 (N_7098,N_6992,N_6965);
nand U7099 (N_7099,N_6913,N_6934);
xnor U7100 (N_7100,N_6875,N_6902);
nand U7101 (N_7101,N_6973,N_6961);
nand U7102 (N_7102,N_6947,N_6933);
nand U7103 (N_7103,N_6921,N_6915);
nor U7104 (N_7104,N_6802,N_6923);
nor U7105 (N_7105,N_6844,N_6956);
nor U7106 (N_7106,N_6972,N_6881);
nand U7107 (N_7107,N_6898,N_6852);
nand U7108 (N_7108,N_6806,N_6878);
or U7109 (N_7109,N_6965,N_6976);
nor U7110 (N_7110,N_6911,N_6856);
nand U7111 (N_7111,N_6894,N_6846);
xnor U7112 (N_7112,N_6841,N_6985);
nor U7113 (N_7113,N_6837,N_6926);
nand U7114 (N_7114,N_6889,N_6963);
or U7115 (N_7115,N_6957,N_6874);
or U7116 (N_7116,N_6992,N_6804);
nand U7117 (N_7117,N_6898,N_6930);
nor U7118 (N_7118,N_6878,N_6873);
and U7119 (N_7119,N_6966,N_6825);
and U7120 (N_7120,N_6885,N_6931);
nor U7121 (N_7121,N_6952,N_6956);
nor U7122 (N_7122,N_6976,N_6883);
xnor U7123 (N_7123,N_6805,N_6964);
or U7124 (N_7124,N_6895,N_6823);
or U7125 (N_7125,N_6991,N_6958);
xnor U7126 (N_7126,N_6942,N_6840);
or U7127 (N_7127,N_6937,N_6979);
nor U7128 (N_7128,N_6902,N_6834);
xor U7129 (N_7129,N_6956,N_6805);
nor U7130 (N_7130,N_6862,N_6924);
and U7131 (N_7131,N_6831,N_6941);
or U7132 (N_7132,N_6979,N_6862);
or U7133 (N_7133,N_6823,N_6901);
nor U7134 (N_7134,N_6992,N_6978);
nor U7135 (N_7135,N_6905,N_6987);
or U7136 (N_7136,N_6931,N_6984);
and U7137 (N_7137,N_6812,N_6879);
nor U7138 (N_7138,N_6960,N_6830);
nor U7139 (N_7139,N_6874,N_6816);
and U7140 (N_7140,N_6830,N_6880);
xnor U7141 (N_7141,N_6871,N_6971);
and U7142 (N_7142,N_6912,N_6836);
and U7143 (N_7143,N_6874,N_6869);
and U7144 (N_7144,N_6925,N_6872);
or U7145 (N_7145,N_6887,N_6949);
or U7146 (N_7146,N_6871,N_6826);
and U7147 (N_7147,N_6908,N_6854);
xor U7148 (N_7148,N_6967,N_6806);
or U7149 (N_7149,N_6931,N_6985);
or U7150 (N_7150,N_6959,N_6981);
nand U7151 (N_7151,N_6984,N_6807);
nor U7152 (N_7152,N_6901,N_6999);
or U7153 (N_7153,N_6866,N_6906);
xor U7154 (N_7154,N_6829,N_6823);
xnor U7155 (N_7155,N_6945,N_6809);
nor U7156 (N_7156,N_6805,N_6940);
xnor U7157 (N_7157,N_6906,N_6805);
xor U7158 (N_7158,N_6911,N_6893);
nand U7159 (N_7159,N_6964,N_6838);
or U7160 (N_7160,N_6836,N_6842);
xnor U7161 (N_7161,N_6906,N_6910);
nor U7162 (N_7162,N_6984,N_6883);
xor U7163 (N_7163,N_6809,N_6916);
and U7164 (N_7164,N_6825,N_6855);
nor U7165 (N_7165,N_6953,N_6997);
and U7166 (N_7166,N_6919,N_6961);
xor U7167 (N_7167,N_6954,N_6879);
or U7168 (N_7168,N_6880,N_6848);
or U7169 (N_7169,N_6877,N_6821);
or U7170 (N_7170,N_6997,N_6982);
xor U7171 (N_7171,N_6856,N_6855);
nor U7172 (N_7172,N_6949,N_6802);
nand U7173 (N_7173,N_6882,N_6922);
nor U7174 (N_7174,N_6844,N_6899);
xor U7175 (N_7175,N_6913,N_6976);
xor U7176 (N_7176,N_6864,N_6963);
nor U7177 (N_7177,N_6843,N_6822);
nand U7178 (N_7178,N_6979,N_6879);
and U7179 (N_7179,N_6901,N_6910);
or U7180 (N_7180,N_6894,N_6822);
xnor U7181 (N_7181,N_6860,N_6865);
or U7182 (N_7182,N_6975,N_6992);
nand U7183 (N_7183,N_6884,N_6840);
nor U7184 (N_7184,N_6976,N_6848);
and U7185 (N_7185,N_6802,N_6997);
nor U7186 (N_7186,N_6842,N_6965);
or U7187 (N_7187,N_6811,N_6804);
and U7188 (N_7188,N_6819,N_6860);
and U7189 (N_7189,N_6931,N_6827);
xor U7190 (N_7190,N_6882,N_6860);
xnor U7191 (N_7191,N_6986,N_6857);
xnor U7192 (N_7192,N_6861,N_6857);
xor U7193 (N_7193,N_6940,N_6963);
or U7194 (N_7194,N_6920,N_6840);
xnor U7195 (N_7195,N_6830,N_6946);
nand U7196 (N_7196,N_6918,N_6930);
nand U7197 (N_7197,N_6957,N_6972);
nand U7198 (N_7198,N_6969,N_6886);
xor U7199 (N_7199,N_6898,N_6965);
or U7200 (N_7200,N_7030,N_7158);
xor U7201 (N_7201,N_7004,N_7054);
xnor U7202 (N_7202,N_7083,N_7039);
and U7203 (N_7203,N_7124,N_7063);
xnor U7204 (N_7204,N_7103,N_7150);
or U7205 (N_7205,N_7025,N_7107);
nor U7206 (N_7206,N_7147,N_7168);
nor U7207 (N_7207,N_7024,N_7172);
or U7208 (N_7208,N_7197,N_7196);
xor U7209 (N_7209,N_7178,N_7156);
or U7210 (N_7210,N_7183,N_7174);
and U7211 (N_7211,N_7097,N_7072);
xor U7212 (N_7212,N_7073,N_7036);
or U7213 (N_7213,N_7042,N_7060);
nand U7214 (N_7214,N_7023,N_7017);
and U7215 (N_7215,N_7151,N_7116);
nor U7216 (N_7216,N_7110,N_7049);
or U7217 (N_7217,N_7018,N_7099);
and U7218 (N_7218,N_7000,N_7062);
nor U7219 (N_7219,N_7096,N_7015);
nor U7220 (N_7220,N_7132,N_7081);
xnor U7221 (N_7221,N_7167,N_7155);
and U7222 (N_7222,N_7198,N_7053);
nor U7223 (N_7223,N_7087,N_7058);
xor U7224 (N_7224,N_7006,N_7077);
nand U7225 (N_7225,N_7045,N_7061);
nand U7226 (N_7226,N_7080,N_7127);
nand U7227 (N_7227,N_7123,N_7090);
xor U7228 (N_7228,N_7192,N_7120);
or U7229 (N_7229,N_7057,N_7101);
nor U7230 (N_7230,N_7069,N_7138);
and U7231 (N_7231,N_7068,N_7171);
xor U7232 (N_7232,N_7041,N_7095);
or U7233 (N_7233,N_7162,N_7008);
xor U7234 (N_7234,N_7010,N_7142);
and U7235 (N_7235,N_7133,N_7022);
nand U7236 (N_7236,N_7126,N_7164);
or U7237 (N_7237,N_7082,N_7009);
and U7238 (N_7238,N_7046,N_7102);
nand U7239 (N_7239,N_7003,N_7074);
nand U7240 (N_7240,N_7013,N_7169);
nor U7241 (N_7241,N_7109,N_7056);
nor U7242 (N_7242,N_7076,N_7014);
or U7243 (N_7243,N_7148,N_7149);
and U7244 (N_7244,N_7152,N_7121);
or U7245 (N_7245,N_7134,N_7002);
xnor U7246 (N_7246,N_7199,N_7078);
and U7247 (N_7247,N_7188,N_7108);
nand U7248 (N_7248,N_7001,N_7092);
xnor U7249 (N_7249,N_7091,N_7035);
nand U7250 (N_7250,N_7166,N_7055);
and U7251 (N_7251,N_7160,N_7159);
nor U7252 (N_7252,N_7043,N_7193);
nand U7253 (N_7253,N_7106,N_7098);
or U7254 (N_7254,N_7071,N_7011);
and U7255 (N_7255,N_7031,N_7154);
xor U7256 (N_7256,N_7115,N_7066);
xor U7257 (N_7257,N_7165,N_7117);
nor U7258 (N_7258,N_7007,N_7027);
nand U7259 (N_7259,N_7146,N_7187);
xor U7260 (N_7260,N_7163,N_7033);
or U7261 (N_7261,N_7005,N_7191);
nor U7262 (N_7262,N_7021,N_7026);
nor U7263 (N_7263,N_7125,N_7179);
nor U7264 (N_7264,N_7089,N_7016);
nand U7265 (N_7265,N_7190,N_7051);
xnor U7266 (N_7266,N_7044,N_7064);
xnor U7267 (N_7267,N_7028,N_7177);
xnor U7268 (N_7268,N_7100,N_7047);
nor U7269 (N_7269,N_7111,N_7094);
or U7270 (N_7270,N_7185,N_7075);
and U7271 (N_7271,N_7070,N_7038);
nor U7272 (N_7272,N_7048,N_7194);
and U7273 (N_7273,N_7135,N_7122);
or U7274 (N_7274,N_7182,N_7144);
or U7275 (N_7275,N_7052,N_7065);
xnor U7276 (N_7276,N_7093,N_7173);
nor U7277 (N_7277,N_7140,N_7175);
nor U7278 (N_7278,N_7088,N_7119);
or U7279 (N_7279,N_7032,N_7050);
nand U7280 (N_7280,N_7130,N_7129);
nand U7281 (N_7281,N_7029,N_7180);
and U7282 (N_7282,N_7034,N_7114);
xor U7283 (N_7283,N_7086,N_7067);
nor U7284 (N_7284,N_7141,N_7143);
or U7285 (N_7285,N_7139,N_7105);
nor U7286 (N_7286,N_7170,N_7189);
nor U7287 (N_7287,N_7112,N_7131);
or U7288 (N_7288,N_7020,N_7113);
nor U7289 (N_7289,N_7195,N_7176);
and U7290 (N_7290,N_7085,N_7084);
nand U7291 (N_7291,N_7186,N_7012);
nor U7292 (N_7292,N_7040,N_7128);
nand U7293 (N_7293,N_7037,N_7118);
and U7294 (N_7294,N_7137,N_7184);
xnor U7295 (N_7295,N_7059,N_7181);
or U7296 (N_7296,N_7157,N_7136);
nor U7297 (N_7297,N_7161,N_7019);
nor U7298 (N_7298,N_7145,N_7104);
xor U7299 (N_7299,N_7079,N_7153);
xnor U7300 (N_7300,N_7170,N_7146);
and U7301 (N_7301,N_7116,N_7038);
or U7302 (N_7302,N_7196,N_7005);
xnor U7303 (N_7303,N_7167,N_7074);
nor U7304 (N_7304,N_7088,N_7055);
or U7305 (N_7305,N_7086,N_7125);
nor U7306 (N_7306,N_7101,N_7080);
and U7307 (N_7307,N_7007,N_7094);
and U7308 (N_7308,N_7168,N_7198);
nor U7309 (N_7309,N_7146,N_7054);
nor U7310 (N_7310,N_7008,N_7127);
or U7311 (N_7311,N_7104,N_7029);
nand U7312 (N_7312,N_7165,N_7010);
nor U7313 (N_7313,N_7129,N_7087);
nand U7314 (N_7314,N_7100,N_7165);
nor U7315 (N_7315,N_7053,N_7127);
nor U7316 (N_7316,N_7047,N_7134);
nand U7317 (N_7317,N_7025,N_7056);
nor U7318 (N_7318,N_7133,N_7000);
and U7319 (N_7319,N_7178,N_7089);
and U7320 (N_7320,N_7110,N_7028);
nand U7321 (N_7321,N_7048,N_7108);
or U7322 (N_7322,N_7134,N_7172);
nor U7323 (N_7323,N_7135,N_7155);
and U7324 (N_7324,N_7108,N_7157);
and U7325 (N_7325,N_7142,N_7166);
xor U7326 (N_7326,N_7139,N_7026);
nor U7327 (N_7327,N_7065,N_7060);
and U7328 (N_7328,N_7026,N_7096);
nand U7329 (N_7329,N_7153,N_7148);
and U7330 (N_7330,N_7007,N_7024);
nor U7331 (N_7331,N_7131,N_7070);
and U7332 (N_7332,N_7024,N_7169);
or U7333 (N_7333,N_7025,N_7086);
nand U7334 (N_7334,N_7146,N_7195);
or U7335 (N_7335,N_7097,N_7077);
and U7336 (N_7336,N_7127,N_7103);
nand U7337 (N_7337,N_7003,N_7055);
nor U7338 (N_7338,N_7102,N_7070);
nand U7339 (N_7339,N_7138,N_7040);
nor U7340 (N_7340,N_7115,N_7141);
and U7341 (N_7341,N_7132,N_7186);
or U7342 (N_7342,N_7099,N_7183);
nand U7343 (N_7343,N_7118,N_7091);
or U7344 (N_7344,N_7066,N_7131);
or U7345 (N_7345,N_7186,N_7141);
or U7346 (N_7346,N_7195,N_7016);
nor U7347 (N_7347,N_7188,N_7038);
or U7348 (N_7348,N_7102,N_7190);
xnor U7349 (N_7349,N_7005,N_7177);
nand U7350 (N_7350,N_7182,N_7140);
nand U7351 (N_7351,N_7177,N_7098);
xor U7352 (N_7352,N_7036,N_7087);
nor U7353 (N_7353,N_7080,N_7103);
and U7354 (N_7354,N_7163,N_7006);
nand U7355 (N_7355,N_7107,N_7037);
xnor U7356 (N_7356,N_7178,N_7073);
or U7357 (N_7357,N_7075,N_7032);
xnor U7358 (N_7358,N_7185,N_7192);
nand U7359 (N_7359,N_7153,N_7130);
xor U7360 (N_7360,N_7159,N_7014);
nand U7361 (N_7361,N_7059,N_7021);
nand U7362 (N_7362,N_7188,N_7120);
nor U7363 (N_7363,N_7088,N_7184);
and U7364 (N_7364,N_7027,N_7101);
or U7365 (N_7365,N_7087,N_7004);
xnor U7366 (N_7366,N_7148,N_7152);
and U7367 (N_7367,N_7151,N_7103);
nand U7368 (N_7368,N_7088,N_7133);
xnor U7369 (N_7369,N_7043,N_7169);
and U7370 (N_7370,N_7060,N_7045);
or U7371 (N_7371,N_7072,N_7012);
and U7372 (N_7372,N_7089,N_7158);
and U7373 (N_7373,N_7057,N_7138);
or U7374 (N_7374,N_7044,N_7194);
or U7375 (N_7375,N_7095,N_7065);
and U7376 (N_7376,N_7196,N_7079);
or U7377 (N_7377,N_7173,N_7067);
xnor U7378 (N_7378,N_7154,N_7016);
nor U7379 (N_7379,N_7102,N_7143);
nor U7380 (N_7380,N_7053,N_7166);
nor U7381 (N_7381,N_7128,N_7192);
and U7382 (N_7382,N_7124,N_7034);
or U7383 (N_7383,N_7004,N_7057);
nor U7384 (N_7384,N_7046,N_7167);
nand U7385 (N_7385,N_7016,N_7052);
xor U7386 (N_7386,N_7195,N_7031);
nor U7387 (N_7387,N_7199,N_7044);
xnor U7388 (N_7388,N_7106,N_7073);
nor U7389 (N_7389,N_7047,N_7142);
nor U7390 (N_7390,N_7053,N_7173);
xnor U7391 (N_7391,N_7114,N_7082);
nand U7392 (N_7392,N_7067,N_7128);
nor U7393 (N_7393,N_7185,N_7048);
and U7394 (N_7394,N_7102,N_7021);
xor U7395 (N_7395,N_7047,N_7028);
nand U7396 (N_7396,N_7023,N_7186);
and U7397 (N_7397,N_7193,N_7091);
nor U7398 (N_7398,N_7151,N_7168);
or U7399 (N_7399,N_7076,N_7031);
and U7400 (N_7400,N_7246,N_7225);
nand U7401 (N_7401,N_7250,N_7304);
and U7402 (N_7402,N_7348,N_7268);
and U7403 (N_7403,N_7292,N_7286);
nor U7404 (N_7404,N_7315,N_7293);
nand U7405 (N_7405,N_7309,N_7308);
and U7406 (N_7406,N_7326,N_7206);
nor U7407 (N_7407,N_7272,N_7366);
and U7408 (N_7408,N_7334,N_7237);
and U7409 (N_7409,N_7345,N_7257);
xnor U7410 (N_7410,N_7393,N_7310);
nand U7411 (N_7411,N_7261,N_7306);
or U7412 (N_7412,N_7288,N_7359);
nor U7413 (N_7413,N_7244,N_7385);
or U7414 (N_7414,N_7220,N_7396);
and U7415 (N_7415,N_7295,N_7373);
or U7416 (N_7416,N_7266,N_7296);
nand U7417 (N_7417,N_7389,N_7277);
nand U7418 (N_7418,N_7355,N_7242);
or U7419 (N_7419,N_7352,N_7379);
xor U7420 (N_7420,N_7204,N_7320);
and U7421 (N_7421,N_7201,N_7298);
and U7422 (N_7422,N_7251,N_7336);
and U7423 (N_7423,N_7314,N_7229);
and U7424 (N_7424,N_7354,N_7331);
xnor U7425 (N_7425,N_7262,N_7369);
or U7426 (N_7426,N_7273,N_7233);
or U7427 (N_7427,N_7205,N_7221);
nor U7428 (N_7428,N_7323,N_7260);
xnor U7429 (N_7429,N_7285,N_7353);
or U7430 (N_7430,N_7207,N_7371);
or U7431 (N_7431,N_7226,N_7243);
and U7432 (N_7432,N_7215,N_7387);
xnor U7433 (N_7433,N_7344,N_7335);
nor U7434 (N_7434,N_7208,N_7301);
and U7435 (N_7435,N_7356,N_7375);
nor U7436 (N_7436,N_7275,N_7287);
xnor U7437 (N_7437,N_7380,N_7318);
nor U7438 (N_7438,N_7202,N_7383);
nor U7439 (N_7439,N_7329,N_7311);
nor U7440 (N_7440,N_7305,N_7327);
or U7441 (N_7441,N_7222,N_7280);
or U7442 (N_7442,N_7322,N_7264);
nand U7443 (N_7443,N_7328,N_7211);
and U7444 (N_7444,N_7399,N_7367);
xnor U7445 (N_7445,N_7363,N_7346);
nand U7446 (N_7446,N_7394,N_7370);
nor U7447 (N_7447,N_7300,N_7281);
nor U7448 (N_7448,N_7256,N_7240);
xnor U7449 (N_7449,N_7342,N_7319);
nand U7450 (N_7450,N_7384,N_7269);
or U7451 (N_7451,N_7239,N_7231);
nand U7452 (N_7452,N_7361,N_7247);
nor U7453 (N_7453,N_7234,N_7294);
or U7454 (N_7454,N_7282,N_7357);
nor U7455 (N_7455,N_7249,N_7238);
nand U7456 (N_7456,N_7253,N_7332);
nor U7457 (N_7457,N_7321,N_7218);
nand U7458 (N_7458,N_7325,N_7398);
or U7459 (N_7459,N_7391,N_7377);
or U7460 (N_7460,N_7224,N_7284);
nor U7461 (N_7461,N_7252,N_7397);
or U7462 (N_7462,N_7364,N_7337);
and U7463 (N_7463,N_7245,N_7232);
nand U7464 (N_7464,N_7223,N_7248);
xor U7465 (N_7465,N_7302,N_7265);
xnor U7466 (N_7466,N_7330,N_7279);
nand U7467 (N_7467,N_7227,N_7230);
and U7468 (N_7468,N_7289,N_7358);
and U7469 (N_7469,N_7219,N_7235);
and U7470 (N_7470,N_7203,N_7381);
nand U7471 (N_7471,N_7267,N_7341);
or U7472 (N_7472,N_7349,N_7339);
xnor U7473 (N_7473,N_7217,N_7362);
nor U7474 (N_7474,N_7210,N_7386);
and U7475 (N_7475,N_7270,N_7297);
and U7476 (N_7476,N_7213,N_7340);
or U7477 (N_7477,N_7241,N_7271);
xnor U7478 (N_7478,N_7274,N_7372);
nor U7479 (N_7479,N_7333,N_7365);
nor U7480 (N_7480,N_7378,N_7212);
nand U7481 (N_7481,N_7258,N_7350);
nor U7482 (N_7482,N_7324,N_7360);
and U7483 (N_7483,N_7343,N_7228);
or U7484 (N_7484,N_7200,N_7291);
or U7485 (N_7485,N_7338,N_7390);
and U7486 (N_7486,N_7259,N_7278);
or U7487 (N_7487,N_7351,N_7382);
nor U7488 (N_7488,N_7216,N_7255);
nor U7489 (N_7489,N_7376,N_7395);
nor U7490 (N_7490,N_7303,N_7316);
or U7491 (N_7491,N_7290,N_7283);
nor U7492 (N_7492,N_7254,N_7374);
and U7493 (N_7493,N_7312,N_7313);
nand U7494 (N_7494,N_7392,N_7299);
nor U7495 (N_7495,N_7214,N_7307);
or U7496 (N_7496,N_7263,N_7317);
and U7497 (N_7497,N_7368,N_7276);
xor U7498 (N_7498,N_7236,N_7347);
nor U7499 (N_7499,N_7388,N_7209);
nand U7500 (N_7500,N_7317,N_7314);
nand U7501 (N_7501,N_7240,N_7354);
nand U7502 (N_7502,N_7374,N_7226);
xnor U7503 (N_7503,N_7266,N_7314);
and U7504 (N_7504,N_7331,N_7248);
or U7505 (N_7505,N_7399,N_7398);
or U7506 (N_7506,N_7354,N_7373);
or U7507 (N_7507,N_7338,N_7373);
xnor U7508 (N_7508,N_7275,N_7241);
and U7509 (N_7509,N_7361,N_7268);
and U7510 (N_7510,N_7274,N_7270);
or U7511 (N_7511,N_7234,N_7273);
nand U7512 (N_7512,N_7333,N_7336);
or U7513 (N_7513,N_7355,N_7368);
or U7514 (N_7514,N_7389,N_7282);
nor U7515 (N_7515,N_7312,N_7252);
xor U7516 (N_7516,N_7319,N_7305);
nor U7517 (N_7517,N_7366,N_7376);
nor U7518 (N_7518,N_7377,N_7349);
nand U7519 (N_7519,N_7238,N_7365);
nor U7520 (N_7520,N_7257,N_7285);
nand U7521 (N_7521,N_7337,N_7296);
and U7522 (N_7522,N_7352,N_7296);
or U7523 (N_7523,N_7386,N_7393);
nor U7524 (N_7524,N_7282,N_7313);
and U7525 (N_7525,N_7382,N_7347);
xnor U7526 (N_7526,N_7305,N_7256);
or U7527 (N_7527,N_7328,N_7366);
and U7528 (N_7528,N_7394,N_7338);
and U7529 (N_7529,N_7298,N_7370);
nand U7530 (N_7530,N_7355,N_7399);
xor U7531 (N_7531,N_7280,N_7391);
and U7532 (N_7532,N_7323,N_7360);
or U7533 (N_7533,N_7315,N_7290);
and U7534 (N_7534,N_7285,N_7312);
and U7535 (N_7535,N_7347,N_7200);
nor U7536 (N_7536,N_7361,N_7358);
or U7537 (N_7537,N_7202,N_7221);
nand U7538 (N_7538,N_7261,N_7376);
and U7539 (N_7539,N_7375,N_7317);
nor U7540 (N_7540,N_7390,N_7372);
xor U7541 (N_7541,N_7281,N_7390);
nor U7542 (N_7542,N_7263,N_7235);
xor U7543 (N_7543,N_7349,N_7328);
nand U7544 (N_7544,N_7222,N_7366);
xor U7545 (N_7545,N_7322,N_7357);
xor U7546 (N_7546,N_7292,N_7217);
nor U7547 (N_7547,N_7299,N_7355);
xnor U7548 (N_7548,N_7208,N_7337);
nand U7549 (N_7549,N_7339,N_7305);
and U7550 (N_7550,N_7226,N_7346);
nand U7551 (N_7551,N_7387,N_7262);
or U7552 (N_7552,N_7273,N_7382);
xnor U7553 (N_7553,N_7301,N_7219);
xnor U7554 (N_7554,N_7221,N_7245);
and U7555 (N_7555,N_7200,N_7380);
or U7556 (N_7556,N_7325,N_7366);
nor U7557 (N_7557,N_7332,N_7377);
nand U7558 (N_7558,N_7204,N_7220);
or U7559 (N_7559,N_7340,N_7283);
and U7560 (N_7560,N_7343,N_7349);
nor U7561 (N_7561,N_7362,N_7372);
xor U7562 (N_7562,N_7237,N_7207);
xor U7563 (N_7563,N_7204,N_7343);
and U7564 (N_7564,N_7262,N_7394);
and U7565 (N_7565,N_7385,N_7302);
xor U7566 (N_7566,N_7287,N_7299);
xnor U7567 (N_7567,N_7270,N_7352);
and U7568 (N_7568,N_7204,N_7266);
nor U7569 (N_7569,N_7355,N_7233);
nand U7570 (N_7570,N_7323,N_7363);
or U7571 (N_7571,N_7331,N_7215);
nand U7572 (N_7572,N_7320,N_7321);
nor U7573 (N_7573,N_7337,N_7306);
nand U7574 (N_7574,N_7307,N_7355);
nand U7575 (N_7575,N_7277,N_7201);
or U7576 (N_7576,N_7276,N_7302);
and U7577 (N_7577,N_7243,N_7266);
nand U7578 (N_7578,N_7253,N_7264);
and U7579 (N_7579,N_7354,N_7258);
or U7580 (N_7580,N_7248,N_7301);
nand U7581 (N_7581,N_7200,N_7313);
or U7582 (N_7582,N_7291,N_7299);
or U7583 (N_7583,N_7334,N_7274);
xnor U7584 (N_7584,N_7251,N_7333);
xor U7585 (N_7585,N_7399,N_7284);
nor U7586 (N_7586,N_7393,N_7379);
xnor U7587 (N_7587,N_7295,N_7267);
nand U7588 (N_7588,N_7265,N_7393);
and U7589 (N_7589,N_7360,N_7291);
xnor U7590 (N_7590,N_7235,N_7295);
and U7591 (N_7591,N_7240,N_7243);
xor U7592 (N_7592,N_7321,N_7244);
nand U7593 (N_7593,N_7370,N_7299);
nor U7594 (N_7594,N_7272,N_7288);
xnor U7595 (N_7595,N_7351,N_7214);
and U7596 (N_7596,N_7232,N_7282);
nand U7597 (N_7597,N_7221,N_7360);
xor U7598 (N_7598,N_7353,N_7307);
or U7599 (N_7599,N_7332,N_7391);
or U7600 (N_7600,N_7441,N_7589);
xnor U7601 (N_7601,N_7474,N_7442);
or U7602 (N_7602,N_7590,N_7453);
or U7603 (N_7603,N_7537,N_7489);
nand U7604 (N_7604,N_7558,N_7405);
nand U7605 (N_7605,N_7559,N_7436);
nand U7606 (N_7606,N_7426,N_7499);
xor U7607 (N_7607,N_7432,N_7502);
and U7608 (N_7608,N_7587,N_7579);
or U7609 (N_7609,N_7512,N_7532);
xnor U7610 (N_7610,N_7524,N_7594);
nand U7611 (N_7611,N_7509,N_7554);
nor U7612 (N_7612,N_7572,N_7550);
xnor U7613 (N_7613,N_7497,N_7531);
nand U7614 (N_7614,N_7469,N_7565);
nor U7615 (N_7615,N_7404,N_7494);
or U7616 (N_7616,N_7526,N_7408);
xor U7617 (N_7617,N_7501,N_7460);
xnor U7618 (N_7618,N_7403,N_7451);
xnor U7619 (N_7619,N_7575,N_7539);
and U7620 (N_7620,N_7447,N_7529);
xnor U7621 (N_7621,N_7419,N_7566);
nor U7622 (N_7622,N_7576,N_7569);
or U7623 (N_7623,N_7452,N_7522);
xnor U7624 (N_7624,N_7544,N_7515);
xor U7625 (N_7625,N_7472,N_7567);
nor U7626 (N_7626,N_7454,N_7400);
nor U7627 (N_7627,N_7496,N_7508);
xor U7628 (N_7628,N_7483,N_7493);
nor U7629 (N_7629,N_7479,N_7412);
xnor U7630 (N_7630,N_7578,N_7401);
nor U7631 (N_7631,N_7520,N_7563);
xor U7632 (N_7632,N_7431,N_7504);
and U7633 (N_7633,N_7481,N_7530);
and U7634 (N_7634,N_7477,N_7488);
nor U7635 (N_7635,N_7402,N_7407);
xnor U7636 (N_7636,N_7592,N_7444);
nor U7637 (N_7637,N_7434,N_7410);
xnor U7638 (N_7638,N_7588,N_7503);
and U7639 (N_7639,N_7551,N_7549);
or U7640 (N_7640,N_7471,N_7450);
nand U7641 (N_7641,N_7409,N_7429);
xnor U7642 (N_7642,N_7495,N_7593);
or U7643 (N_7643,N_7425,N_7500);
xnor U7644 (N_7644,N_7555,N_7475);
and U7645 (N_7645,N_7448,N_7421);
or U7646 (N_7646,N_7518,N_7548);
nand U7647 (N_7647,N_7585,N_7513);
and U7648 (N_7648,N_7540,N_7577);
nand U7649 (N_7649,N_7461,N_7418);
nand U7650 (N_7650,N_7464,N_7511);
nor U7651 (N_7651,N_7416,N_7424);
xor U7652 (N_7652,N_7553,N_7599);
and U7653 (N_7653,N_7462,N_7580);
and U7654 (N_7654,N_7591,N_7568);
or U7655 (N_7655,N_7492,N_7428);
xnor U7656 (N_7656,N_7560,N_7423);
xor U7657 (N_7657,N_7420,N_7427);
or U7658 (N_7658,N_7552,N_7417);
or U7659 (N_7659,N_7571,N_7422);
nand U7660 (N_7660,N_7485,N_7598);
nor U7661 (N_7661,N_7573,N_7525);
and U7662 (N_7662,N_7542,N_7467);
nand U7663 (N_7663,N_7468,N_7574);
nand U7664 (N_7664,N_7445,N_7581);
or U7665 (N_7665,N_7536,N_7545);
xor U7666 (N_7666,N_7480,N_7438);
or U7667 (N_7667,N_7487,N_7463);
or U7668 (N_7668,N_7586,N_7411);
nor U7669 (N_7669,N_7557,N_7456);
xnor U7670 (N_7670,N_7533,N_7583);
or U7671 (N_7671,N_7523,N_7439);
nor U7672 (N_7672,N_7478,N_7455);
xnor U7673 (N_7673,N_7459,N_7470);
nand U7674 (N_7674,N_7570,N_7516);
xnor U7675 (N_7675,N_7561,N_7519);
nand U7676 (N_7676,N_7498,N_7534);
nor U7677 (N_7677,N_7484,N_7482);
and U7678 (N_7678,N_7597,N_7505);
and U7679 (N_7679,N_7507,N_7490);
and U7680 (N_7680,N_7465,N_7541);
and U7681 (N_7681,N_7457,N_7486);
nor U7682 (N_7682,N_7415,N_7491);
nand U7683 (N_7683,N_7458,N_7406);
nand U7684 (N_7684,N_7517,N_7476);
nand U7685 (N_7685,N_7413,N_7437);
xnor U7686 (N_7686,N_7595,N_7433);
nand U7687 (N_7687,N_7446,N_7538);
nand U7688 (N_7688,N_7556,N_7527);
and U7689 (N_7689,N_7543,N_7546);
nor U7690 (N_7690,N_7440,N_7414);
or U7691 (N_7691,N_7582,N_7562);
and U7692 (N_7692,N_7528,N_7547);
nand U7693 (N_7693,N_7449,N_7514);
xnor U7694 (N_7694,N_7443,N_7596);
nand U7695 (N_7695,N_7564,N_7535);
xnor U7696 (N_7696,N_7430,N_7584);
xnor U7697 (N_7697,N_7466,N_7521);
xor U7698 (N_7698,N_7435,N_7506);
or U7699 (N_7699,N_7510,N_7473);
nor U7700 (N_7700,N_7560,N_7516);
nand U7701 (N_7701,N_7475,N_7554);
or U7702 (N_7702,N_7454,N_7408);
and U7703 (N_7703,N_7512,N_7432);
nand U7704 (N_7704,N_7472,N_7442);
nand U7705 (N_7705,N_7478,N_7474);
nor U7706 (N_7706,N_7472,N_7451);
xor U7707 (N_7707,N_7537,N_7444);
xor U7708 (N_7708,N_7567,N_7526);
nand U7709 (N_7709,N_7544,N_7546);
nor U7710 (N_7710,N_7530,N_7424);
or U7711 (N_7711,N_7488,N_7504);
or U7712 (N_7712,N_7441,N_7400);
and U7713 (N_7713,N_7533,N_7414);
xor U7714 (N_7714,N_7598,N_7532);
or U7715 (N_7715,N_7547,N_7524);
xor U7716 (N_7716,N_7575,N_7438);
or U7717 (N_7717,N_7561,N_7412);
nor U7718 (N_7718,N_7487,N_7584);
and U7719 (N_7719,N_7458,N_7598);
or U7720 (N_7720,N_7573,N_7520);
and U7721 (N_7721,N_7524,N_7488);
or U7722 (N_7722,N_7550,N_7579);
nand U7723 (N_7723,N_7458,N_7563);
or U7724 (N_7724,N_7434,N_7472);
nand U7725 (N_7725,N_7556,N_7524);
nor U7726 (N_7726,N_7582,N_7586);
nand U7727 (N_7727,N_7500,N_7555);
or U7728 (N_7728,N_7559,N_7513);
nand U7729 (N_7729,N_7521,N_7414);
nand U7730 (N_7730,N_7499,N_7575);
or U7731 (N_7731,N_7485,N_7564);
and U7732 (N_7732,N_7580,N_7598);
and U7733 (N_7733,N_7525,N_7429);
and U7734 (N_7734,N_7543,N_7414);
nor U7735 (N_7735,N_7529,N_7512);
and U7736 (N_7736,N_7411,N_7447);
nand U7737 (N_7737,N_7446,N_7486);
and U7738 (N_7738,N_7457,N_7430);
or U7739 (N_7739,N_7558,N_7455);
nor U7740 (N_7740,N_7555,N_7466);
or U7741 (N_7741,N_7559,N_7596);
or U7742 (N_7742,N_7441,N_7518);
and U7743 (N_7743,N_7512,N_7558);
xor U7744 (N_7744,N_7550,N_7566);
and U7745 (N_7745,N_7595,N_7409);
and U7746 (N_7746,N_7491,N_7444);
nand U7747 (N_7747,N_7405,N_7487);
xnor U7748 (N_7748,N_7424,N_7523);
xnor U7749 (N_7749,N_7430,N_7495);
nand U7750 (N_7750,N_7529,N_7405);
nand U7751 (N_7751,N_7530,N_7462);
or U7752 (N_7752,N_7403,N_7506);
nor U7753 (N_7753,N_7569,N_7562);
and U7754 (N_7754,N_7428,N_7470);
nor U7755 (N_7755,N_7566,N_7571);
nand U7756 (N_7756,N_7597,N_7410);
or U7757 (N_7757,N_7577,N_7486);
and U7758 (N_7758,N_7596,N_7515);
nand U7759 (N_7759,N_7441,N_7410);
nor U7760 (N_7760,N_7475,N_7560);
nand U7761 (N_7761,N_7444,N_7568);
xnor U7762 (N_7762,N_7429,N_7563);
nor U7763 (N_7763,N_7579,N_7569);
or U7764 (N_7764,N_7497,N_7552);
and U7765 (N_7765,N_7575,N_7478);
nor U7766 (N_7766,N_7516,N_7538);
and U7767 (N_7767,N_7485,N_7444);
xnor U7768 (N_7768,N_7566,N_7528);
or U7769 (N_7769,N_7458,N_7460);
xnor U7770 (N_7770,N_7564,N_7558);
nand U7771 (N_7771,N_7538,N_7591);
nor U7772 (N_7772,N_7411,N_7518);
xnor U7773 (N_7773,N_7531,N_7443);
xnor U7774 (N_7774,N_7505,N_7583);
and U7775 (N_7775,N_7568,N_7537);
nand U7776 (N_7776,N_7553,N_7420);
nand U7777 (N_7777,N_7589,N_7498);
nand U7778 (N_7778,N_7517,N_7590);
xnor U7779 (N_7779,N_7553,N_7476);
xnor U7780 (N_7780,N_7570,N_7495);
nor U7781 (N_7781,N_7587,N_7534);
nor U7782 (N_7782,N_7475,N_7563);
nand U7783 (N_7783,N_7404,N_7538);
nand U7784 (N_7784,N_7481,N_7506);
nor U7785 (N_7785,N_7438,N_7598);
or U7786 (N_7786,N_7504,N_7589);
nor U7787 (N_7787,N_7498,N_7557);
and U7788 (N_7788,N_7491,N_7452);
or U7789 (N_7789,N_7470,N_7469);
and U7790 (N_7790,N_7411,N_7449);
or U7791 (N_7791,N_7573,N_7406);
xor U7792 (N_7792,N_7470,N_7430);
or U7793 (N_7793,N_7562,N_7485);
or U7794 (N_7794,N_7495,N_7554);
nand U7795 (N_7795,N_7590,N_7537);
and U7796 (N_7796,N_7438,N_7514);
or U7797 (N_7797,N_7458,N_7508);
and U7798 (N_7798,N_7517,N_7441);
nor U7799 (N_7799,N_7559,N_7491);
or U7800 (N_7800,N_7647,N_7625);
xor U7801 (N_7801,N_7796,N_7786);
and U7802 (N_7802,N_7742,N_7606);
and U7803 (N_7803,N_7782,N_7652);
xor U7804 (N_7804,N_7667,N_7669);
nand U7805 (N_7805,N_7602,N_7720);
and U7806 (N_7806,N_7722,N_7632);
or U7807 (N_7807,N_7662,N_7791);
and U7808 (N_7808,N_7658,N_7609);
and U7809 (N_7809,N_7765,N_7628);
nand U7810 (N_7810,N_7728,N_7682);
or U7811 (N_7811,N_7741,N_7610);
nand U7812 (N_7812,N_7706,N_7649);
nor U7813 (N_7813,N_7622,N_7672);
nor U7814 (N_7814,N_7729,N_7758);
nand U7815 (N_7815,N_7618,N_7670);
nor U7816 (N_7816,N_7707,N_7760);
nand U7817 (N_7817,N_7642,N_7736);
nor U7818 (N_7818,N_7636,N_7779);
xnor U7819 (N_7819,N_7650,N_7626);
or U7820 (N_7820,N_7689,N_7619);
nand U7821 (N_7821,N_7620,N_7603);
nor U7822 (N_7822,N_7709,N_7790);
and U7823 (N_7823,N_7695,N_7711);
or U7824 (N_7824,N_7778,N_7771);
or U7825 (N_7825,N_7681,N_7677);
and U7826 (N_7826,N_7735,N_7661);
and U7827 (N_7827,N_7692,N_7785);
nor U7828 (N_7828,N_7768,N_7750);
and U7829 (N_7829,N_7713,N_7724);
nor U7830 (N_7830,N_7687,N_7717);
or U7831 (N_7831,N_7726,N_7653);
xor U7832 (N_7832,N_7607,N_7769);
or U7833 (N_7833,N_7799,N_7748);
and U7834 (N_7834,N_7775,N_7648);
nor U7835 (N_7835,N_7698,N_7755);
nor U7836 (N_7836,N_7732,N_7757);
nor U7837 (N_7837,N_7754,N_7639);
nand U7838 (N_7838,N_7731,N_7671);
nand U7839 (N_7839,N_7756,N_7614);
nand U7840 (N_7840,N_7705,N_7676);
xor U7841 (N_7841,N_7691,N_7657);
nor U7842 (N_7842,N_7714,N_7787);
nand U7843 (N_7843,N_7710,N_7673);
xor U7844 (N_7844,N_7767,N_7699);
or U7845 (N_7845,N_7702,N_7633);
and U7846 (N_7846,N_7747,N_7645);
nor U7847 (N_7847,N_7612,N_7646);
or U7848 (N_7848,N_7762,N_7737);
nand U7849 (N_7849,N_7763,N_7621);
and U7850 (N_7850,N_7680,N_7694);
nor U7851 (N_7851,N_7793,N_7688);
and U7852 (N_7852,N_7746,N_7745);
and U7853 (N_7853,N_7627,N_7733);
nand U7854 (N_7854,N_7774,N_7708);
or U7855 (N_7855,N_7770,N_7751);
and U7856 (N_7856,N_7684,N_7660);
nor U7857 (N_7857,N_7761,N_7604);
nor U7858 (N_7858,N_7685,N_7654);
nor U7859 (N_7859,N_7629,N_7739);
and U7860 (N_7860,N_7656,N_7712);
nor U7861 (N_7861,N_7601,N_7697);
xnor U7862 (N_7862,N_7792,N_7723);
xor U7863 (N_7863,N_7752,N_7701);
or U7864 (N_7864,N_7730,N_7740);
and U7865 (N_7865,N_7663,N_7666);
nand U7866 (N_7866,N_7679,N_7623);
xnor U7867 (N_7867,N_7624,N_7783);
and U7868 (N_7868,N_7703,N_7615);
or U7869 (N_7869,N_7696,N_7664);
nor U7870 (N_7870,N_7716,N_7797);
nand U7871 (N_7871,N_7608,N_7749);
nand U7872 (N_7872,N_7659,N_7776);
nand U7873 (N_7873,N_7788,N_7743);
and U7874 (N_7874,N_7780,N_7616);
xnor U7875 (N_7875,N_7700,N_7718);
xnor U7876 (N_7876,N_7798,N_7631);
nand U7877 (N_7877,N_7675,N_7605);
or U7878 (N_7878,N_7635,N_7738);
and U7879 (N_7879,N_7773,N_7678);
nand U7880 (N_7880,N_7704,N_7744);
nand U7881 (N_7881,N_7719,N_7725);
or U7882 (N_7882,N_7683,N_7674);
nor U7883 (N_7883,N_7795,N_7644);
and U7884 (N_7884,N_7611,N_7686);
xor U7885 (N_7885,N_7630,N_7668);
nand U7886 (N_7886,N_7600,N_7637);
xnor U7887 (N_7887,N_7651,N_7665);
and U7888 (N_7888,N_7766,N_7784);
xor U7889 (N_7889,N_7734,N_7634);
xor U7890 (N_7890,N_7641,N_7721);
xor U7891 (N_7891,N_7781,N_7715);
xor U7892 (N_7892,N_7693,N_7764);
and U7893 (N_7893,N_7772,N_7655);
xnor U7894 (N_7894,N_7727,N_7794);
nor U7895 (N_7895,N_7638,N_7789);
nand U7896 (N_7896,N_7777,N_7753);
and U7897 (N_7897,N_7617,N_7759);
and U7898 (N_7898,N_7613,N_7640);
xnor U7899 (N_7899,N_7690,N_7643);
and U7900 (N_7900,N_7659,N_7685);
and U7901 (N_7901,N_7678,N_7685);
xnor U7902 (N_7902,N_7649,N_7795);
nand U7903 (N_7903,N_7733,N_7668);
and U7904 (N_7904,N_7611,N_7672);
or U7905 (N_7905,N_7691,N_7717);
and U7906 (N_7906,N_7705,N_7700);
xnor U7907 (N_7907,N_7668,N_7764);
nand U7908 (N_7908,N_7789,N_7615);
or U7909 (N_7909,N_7635,N_7643);
xor U7910 (N_7910,N_7783,N_7604);
nor U7911 (N_7911,N_7620,N_7768);
and U7912 (N_7912,N_7627,N_7791);
nor U7913 (N_7913,N_7773,N_7745);
and U7914 (N_7914,N_7700,N_7760);
and U7915 (N_7915,N_7671,N_7610);
nor U7916 (N_7916,N_7603,N_7731);
nor U7917 (N_7917,N_7672,N_7719);
xor U7918 (N_7918,N_7691,N_7682);
nand U7919 (N_7919,N_7616,N_7798);
nand U7920 (N_7920,N_7622,N_7745);
nor U7921 (N_7921,N_7646,N_7706);
or U7922 (N_7922,N_7792,N_7623);
or U7923 (N_7923,N_7671,N_7600);
or U7924 (N_7924,N_7737,N_7623);
nor U7925 (N_7925,N_7628,N_7698);
xnor U7926 (N_7926,N_7785,N_7748);
nand U7927 (N_7927,N_7696,N_7609);
nand U7928 (N_7928,N_7696,N_7786);
nor U7929 (N_7929,N_7739,N_7600);
or U7930 (N_7930,N_7700,N_7666);
xor U7931 (N_7931,N_7648,N_7672);
or U7932 (N_7932,N_7606,N_7680);
or U7933 (N_7933,N_7753,N_7711);
nor U7934 (N_7934,N_7749,N_7796);
or U7935 (N_7935,N_7636,N_7616);
nor U7936 (N_7936,N_7715,N_7711);
nand U7937 (N_7937,N_7705,N_7779);
and U7938 (N_7938,N_7684,N_7657);
or U7939 (N_7939,N_7788,N_7766);
nand U7940 (N_7940,N_7640,N_7607);
nor U7941 (N_7941,N_7689,N_7719);
xnor U7942 (N_7942,N_7689,N_7776);
nor U7943 (N_7943,N_7766,N_7684);
nand U7944 (N_7944,N_7703,N_7712);
nand U7945 (N_7945,N_7740,N_7768);
xnor U7946 (N_7946,N_7796,N_7769);
or U7947 (N_7947,N_7610,N_7664);
xor U7948 (N_7948,N_7787,N_7639);
or U7949 (N_7949,N_7704,N_7785);
nand U7950 (N_7950,N_7776,N_7674);
or U7951 (N_7951,N_7600,N_7742);
or U7952 (N_7952,N_7638,N_7773);
or U7953 (N_7953,N_7607,N_7782);
xor U7954 (N_7954,N_7798,N_7766);
nor U7955 (N_7955,N_7711,N_7728);
and U7956 (N_7956,N_7665,N_7634);
nor U7957 (N_7957,N_7747,N_7671);
or U7958 (N_7958,N_7607,N_7717);
and U7959 (N_7959,N_7604,N_7796);
xor U7960 (N_7960,N_7652,N_7638);
nand U7961 (N_7961,N_7639,N_7740);
nor U7962 (N_7962,N_7697,N_7773);
or U7963 (N_7963,N_7788,N_7716);
xor U7964 (N_7964,N_7756,N_7782);
nand U7965 (N_7965,N_7678,N_7614);
or U7966 (N_7966,N_7795,N_7642);
or U7967 (N_7967,N_7727,N_7654);
nand U7968 (N_7968,N_7751,N_7726);
xor U7969 (N_7969,N_7770,N_7714);
nor U7970 (N_7970,N_7736,N_7721);
xor U7971 (N_7971,N_7750,N_7747);
nand U7972 (N_7972,N_7764,N_7704);
nor U7973 (N_7973,N_7750,N_7686);
xnor U7974 (N_7974,N_7620,N_7750);
and U7975 (N_7975,N_7669,N_7624);
and U7976 (N_7976,N_7622,N_7661);
or U7977 (N_7977,N_7713,N_7778);
nand U7978 (N_7978,N_7619,N_7603);
and U7979 (N_7979,N_7717,N_7634);
nor U7980 (N_7980,N_7712,N_7623);
and U7981 (N_7981,N_7675,N_7768);
nor U7982 (N_7982,N_7604,N_7756);
nand U7983 (N_7983,N_7745,N_7623);
or U7984 (N_7984,N_7685,N_7791);
nand U7985 (N_7985,N_7731,N_7696);
or U7986 (N_7986,N_7679,N_7782);
nand U7987 (N_7987,N_7695,N_7666);
nor U7988 (N_7988,N_7626,N_7623);
or U7989 (N_7989,N_7703,N_7625);
and U7990 (N_7990,N_7757,N_7740);
or U7991 (N_7991,N_7602,N_7736);
xor U7992 (N_7992,N_7741,N_7782);
and U7993 (N_7993,N_7646,N_7666);
xnor U7994 (N_7994,N_7659,N_7663);
nand U7995 (N_7995,N_7602,N_7662);
and U7996 (N_7996,N_7694,N_7768);
and U7997 (N_7997,N_7672,N_7772);
xnor U7998 (N_7998,N_7629,N_7729);
or U7999 (N_7999,N_7606,N_7746);
nand U8000 (N_8000,N_7924,N_7895);
xnor U8001 (N_8001,N_7880,N_7909);
xnor U8002 (N_8002,N_7965,N_7801);
xor U8003 (N_8003,N_7874,N_7985);
nand U8004 (N_8004,N_7848,N_7803);
and U8005 (N_8005,N_7980,N_7818);
or U8006 (N_8006,N_7926,N_7897);
or U8007 (N_8007,N_7960,N_7853);
and U8008 (N_8008,N_7968,N_7964);
and U8009 (N_8009,N_7949,N_7870);
nor U8010 (N_8010,N_7809,N_7877);
nand U8011 (N_8011,N_7971,N_7952);
or U8012 (N_8012,N_7810,N_7961);
xor U8013 (N_8013,N_7813,N_7804);
and U8014 (N_8014,N_7939,N_7811);
or U8015 (N_8015,N_7879,N_7955);
nand U8016 (N_8016,N_7963,N_7925);
nor U8017 (N_8017,N_7823,N_7982);
or U8018 (N_8018,N_7852,N_7993);
or U8019 (N_8019,N_7862,N_7966);
and U8020 (N_8020,N_7987,N_7934);
nand U8021 (N_8021,N_7986,N_7900);
or U8022 (N_8022,N_7995,N_7962);
or U8023 (N_8023,N_7802,N_7994);
and U8024 (N_8024,N_7891,N_7857);
xor U8025 (N_8025,N_7854,N_7855);
nor U8026 (N_8026,N_7953,N_7808);
xor U8027 (N_8027,N_7945,N_7951);
and U8028 (N_8028,N_7830,N_7930);
xor U8029 (N_8029,N_7988,N_7819);
nor U8030 (N_8030,N_7827,N_7841);
and U8031 (N_8031,N_7832,N_7817);
or U8032 (N_8032,N_7884,N_7881);
or U8033 (N_8033,N_7866,N_7999);
nand U8034 (N_8034,N_7834,N_7836);
xor U8035 (N_8035,N_7858,N_7878);
xor U8036 (N_8036,N_7947,N_7919);
or U8037 (N_8037,N_7846,N_7969);
xnor U8038 (N_8038,N_7814,N_7928);
xnor U8039 (N_8039,N_7888,N_7840);
nand U8040 (N_8040,N_7931,N_7869);
and U8041 (N_8041,N_7973,N_7896);
nand U8042 (N_8042,N_7917,N_7937);
nand U8043 (N_8043,N_7893,N_7938);
xor U8044 (N_8044,N_7867,N_7800);
or U8045 (N_8045,N_7815,N_7860);
or U8046 (N_8046,N_7898,N_7875);
nor U8047 (N_8047,N_7863,N_7807);
nand U8048 (N_8048,N_7967,N_7890);
xor U8049 (N_8049,N_7886,N_7916);
xnor U8050 (N_8050,N_7899,N_7956);
or U8051 (N_8051,N_7833,N_7972);
nor U8052 (N_8052,N_7842,N_7865);
xnor U8053 (N_8053,N_7977,N_7816);
nand U8054 (N_8054,N_7911,N_7844);
and U8055 (N_8055,N_7943,N_7824);
nand U8056 (N_8056,N_7856,N_7929);
or U8057 (N_8057,N_7997,N_7970);
or U8058 (N_8058,N_7826,N_7923);
xnor U8059 (N_8059,N_7825,N_7903);
nand U8060 (N_8060,N_7901,N_7910);
nand U8061 (N_8061,N_7912,N_7847);
or U8062 (N_8062,N_7941,N_7837);
and U8063 (N_8063,N_7992,N_7828);
xor U8064 (N_8064,N_7873,N_7889);
nor U8065 (N_8065,N_7864,N_7996);
xor U8066 (N_8066,N_7976,N_7871);
nor U8067 (N_8067,N_7843,N_7820);
nand U8068 (N_8068,N_7876,N_7835);
nand U8069 (N_8069,N_7915,N_7906);
or U8070 (N_8070,N_7905,N_7908);
or U8071 (N_8071,N_7932,N_7892);
and U8072 (N_8072,N_7839,N_7922);
and U8073 (N_8073,N_7882,N_7904);
nor U8074 (N_8074,N_7885,N_7984);
nand U8075 (N_8075,N_7990,N_7991);
and U8076 (N_8076,N_7975,N_7806);
and U8077 (N_8077,N_7859,N_7920);
xor U8078 (N_8078,N_7902,N_7812);
and U8079 (N_8079,N_7942,N_7954);
nor U8080 (N_8080,N_7821,N_7894);
nand U8081 (N_8081,N_7872,N_7849);
nand U8082 (N_8082,N_7822,N_7851);
and U8083 (N_8083,N_7887,N_7940);
nor U8084 (N_8084,N_7989,N_7933);
or U8085 (N_8085,N_7913,N_7981);
nand U8086 (N_8086,N_7983,N_7845);
nor U8087 (N_8087,N_7829,N_7946);
nand U8088 (N_8088,N_7978,N_7936);
and U8089 (N_8089,N_7935,N_7805);
or U8090 (N_8090,N_7974,N_7918);
and U8091 (N_8091,N_7950,N_7948);
xnor U8092 (N_8092,N_7979,N_7838);
and U8093 (N_8093,N_7921,N_7998);
and U8094 (N_8094,N_7861,N_7927);
or U8095 (N_8095,N_7883,N_7957);
nand U8096 (N_8096,N_7944,N_7907);
and U8097 (N_8097,N_7958,N_7831);
or U8098 (N_8098,N_7914,N_7868);
xnor U8099 (N_8099,N_7850,N_7959);
nand U8100 (N_8100,N_7869,N_7929);
nor U8101 (N_8101,N_7926,N_7864);
or U8102 (N_8102,N_7806,N_7943);
nand U8103 (N_8103,N_7977,N_7875);
nor U8104 (N_8104,N_7853,N_7979);
xnor U8105 (N_8105,N_7954,N_7847);
xor U8106 (N_8106,N_7806,N_7945);
nor U8107 (N_8107,N_7995,N_7895);
nand U8108 (N_8108,N_7972,N_7958);
xor U8109 (N_8109,N_7871,N_7930);
nor U8110 (N_8110,N_7994,N_7830);
nand U8111 (N_8111,N_7939,N_7959);
nor U8112 (N_8112,N_7908,N_7901);
and U8113 (N_8113,N_7890,N_7995);
xnor U8114 (N_8114,N_7850,N_7820);
and U8115 (N_8115,N_7801,N_7902);
xnor U8116 (N_8116,N_7813,N_7935);
nand U8117 (N_8117,N_7955,N_7908);
nand U8118 (N_8118,N_7956,N_7832);
nand U8119 (N_8119,N_7855,N_7944);
or U8120 (N_8120,N_7824,N_7898);
or U8121 (N_8121,N_7939,N_7951);
nor U8122 (N_8122,N_7894,N_7920);
and U8123 (N_8123,N_7891,N_7856);
or U8124 (N_8124,N_7944,N_7821);
and U8125 (N_8125,N_7906,N_7903);
or U8126 (N_8126,N_7935,N_7932);
xor U8127 (N_8127,N_7838,N_7942);
or U8128 (N_8128,N_7886,N_7892);
or U8129 (N_8129,N_7800,N_7976);
or U8130 (N_8130,N_7821,N_7967);
xor U8131 (N_8131,N_7859,N_7902);
xor U8132 (N_8132,N_7990,N_7876);
and U8133 (N_8133,N_7910,N_7898);
xnor U8134 (N_8134,N_7855,N_7816);
and U8135 (N_8135,N_7986,N_7927);
or U8136 (N_8136,N_7995,N_7829);
nor U8137 (N_8137,N_7945,N_7884);
xnor U8138 (N_8138,N_7854,N_7892);
nand U8139 (N_8139,N_7955,N_7933);
nor U8140 (N_8140,N_7942,N_7809);
and U8141 (N_8141,N_7889,N_7909);
nor U8142 (N_8142,N_7813,N_7914);
xor U8143 (N_8143,N_7890,N_7971);
nand U8144 (N_8144,N_7811,N_7935);
or U8145 (N_8145,N_7961,N_7987);
or U8146 (N_8146,N_7901,N_7942);
and U8147 (N_8147,N_7878,N_7967);
and U8148 (N_8148,N_7806,N_7923);
nor U8149 (N_8149,N_7810,N_7832);
nor U8150 (N_8150,N_7836,N_7802);
or U8151 (N_8151,N_7932,N_7980);
nand U8152 (N_8152,N_7909,N_7843);
xor U8153 (N_8153,N_7929,N_7877);
or U8154 (N_8154,N_7949,N_7839);
and U8155 (N_8155,N_7905,N_7820);
and U8156 (N_8156,N_7974,N_7803);
xor U8157 (N_8157,N_7992,N_7823);
or U8158 (N_8158,N_7839,N_7910);
nand U8159 (N_8159,N_7993,N_7960);
nand U8160 (N_8160,N_7873,N_7845);
nand U8161 (N_8161,N_7817,N_7922);
or U8162 (N_8162,N_7981,N_7946);
or U8163 (N_8163,N_7836,N_7807);
and U8164 (N_8164,N_7812,N_7830);
and U8165 (N_8165,N_7901,N_7948);
and U8166 (N_8166,N_7858,N_7890);
xnor U8167 (N_8167,N_7986,N_7878);
nand U8168 (N_8168,N_7962,N_7859);
nor U8169 (N_8169,N_7835,N_7859);
or U8170 (N_8170,N_7817,N_7975);
xor U8171 (N_8171,N_7827,N_7859);
and U8172 (N_8172,N_7819,N_7880);
or U8173 (N_8173,N_7900,N_7973);
nor U8174 (N_8174,N_7938,N_7859);
nor U8175 (N_8175,N_7892,N_7818);
xor U8176 (N_8176,N_7802,N_7817);
and U8177 (N_8177,N_7849,N_7833);
xor U8178 (N_8178,N_7824,N_7909);
nor U8179 (N_8179,N_7915,N_7974);
nand U8180 (N_8180,N_7865,N_7869);
nor U8181 (N_8181,N_7921,N_7929);
and U8182 (N_8182,N_7896,N_7883);
and U8183 (N_8183,N_7991,N_7880);
nor U8184 (N_8184,N_7904,N_7831);
nand U8185 (N_8185,N_7941,N_7876);
nor U8186 (N_8186,N_7805,N_7944);
or U8187 (N_8187,N_7875,N_7992);
or U8188 (N_8188,N_7904,N_7982);
and U8189 (N_8189,N_7889,N_7939);
nor U8190 (N_8190,N_7942,N_7897);
nor U8191 (N_8191,N_7911,N_7890);
nand U8192 (N_8192,N_7919,N_7852);
nand U8193 (N_8193,N_7930,N_7893);
nor U8194 (N_8194,N_7943,N_7972);
nand U8195 (N_8195,N_7852,N_7859);
and U8196 (N_8196,N_7985,N_7970);
xnor U8197 (N_8197,N_7930,N_7812);
nor U8198 (N_8198,N_7900,N_7972);
or U8199 (N_8199,N_7988,N_7925);
or U8200 (N_8200,N_8196,N_8025);
xor U8201 (N_8201,N_8154,N_8180);
nand U8202 (N_8202,N_8173,N_8002);
xnor U8203 (N_8203,N_8089,N_8021);
nand U8204 (N_8204,N_8160,N_8036);
xor U8205 (N_8205,N_8022,N_8100);
nor U8206 (N_8206,N_8014,N_8006);
or U8207 (N_8207,N_8087,N_8043);
xor U8208 (N_8208,N_8137,N_8142);
xor U8209 (N_8209,N_8063,N_8003);
or U8210 (N_8210,N_8148,N_8061);
xor U8211 (N_8211,N_8110,N_8095);
nor U8212 (N_8212,N_8186,N_8123);
or U8213 (N_8213,N_8169,N_8198);
and U8214 (N_8214,N_8053,N_8084);
and U8215 (N_8215,N_8040,N_8105);
nand U8216 (N_8216,N_8023,N_8139);
nor U8217 (N_8217,N_8172,N_8135);
nand U8218 (N_8218,N_8016,N_8039);
and U8219 (N_8219,N_8085,N_8019);
nor U8220 (N_8220,N_8038,N_8018);
or U8221 (N_8221,N_8116,N_8058);
and U8222 (N_8222,N_8109,N_8155);
xor U8223 (N_8223,N_8066,N_8132);
and U8224 (N_8224,N_8140,N_8150);
nand U8225 (N_8225,N_8124,N_8151);
xor U8226 (N_8226,N_8158,N_8190);
and U8227 (N_8227,N_8176,N_8060);
or U8228 (N_8228,N_8091,N_8126);
and U8229 (N_8229,N_8178,N_8080);
xnor U8230 (N_8230,N_8159,N_8162);
or U8231 (N_8231,N_8057,N_8183);
nand U8232 (N_8232,N_8032,N_8076);
or U8233 (N_8233,N_8009,N_8103);
nor U8234 (N_8234,N_8000,N_8088);
and U8235 (N_8235,N_8034,N_8164);
or U8236 (N_8236,N_8111,N_8165);
nor U8237 (N_8237,N_8145,N_8097);
xnor U8238 (N_8238,N_8008,N_8012);
nand U8239 (N_8239,N_8033,N_8055);
and U8240 (N_8240,N_8146,N_8086);
and U8241 (N_8241,N_8144,N_8191);
xnor U8242 (N_8242,N_8072,N_8147);
nand U8243 (N_8243,N_8027,N_8188);
or U8244 (N_8244,N_8028,N_8136);
or U8245 (N_8245,N_8078,N_8031);
or U8246 (N_8246,N_8045,N_8189);
nor U8247 (N_8247,N_8062,N_8079);
and U8248 (N_8248,N_8130,N_8131);
xnor U8249 (N_8249,N_8069,N_8071);
nand U8250 (N_8250,N_8157,N_8052);
and U8251 (N_8251,N_8171,N_8107);
nand U8252 (N_8252,N_8065,N_8106);
nand U8253 (N_8253,N_8120,N_8108);
or U8254 (N_8254,N_8029,N_8153);
and U8255 (N_8255,N_8163,N_8024);
or U8256 (N_8256,N_8129,N_8017);
xor U8257 (N_8257,N_8030,N_8005);
nand U8258 (N_8258,N_8098,N_8112);
nand U8259 (N_8259,N_8068,N_8177);
or U8260 (N_8260,N_8168,N_8101);
or U8261 (N_8261,N_8118,N_8050);
xor U8262 (N_8262,N_8167,N_8149);
or U8263 (N_8263,N_8182,N_8156);
nor U8264 (N_8264,N_8197,N_8195);
or U8265 (N_8265,N_8121,N_8042);
nor U8266 (N_8266,N_8099,N_8187);
xor U8267 (N_8267,N_8161,N_8026);
or U8268 (N_8268,N_8067,N_8073);
nor U8269 (N_8269,N_8138,N_8020);
and U8270 (N_8270,N_8141,N_8170);
xnor U8271 (N_8271,N_8035,N_8115);
xnor U8272 (N_8272,N_8114,N_8127);
xor U8273 (N_8273,N_8046,N_8096);
xnor U8274 (N_8274,N_8102,N_8092);
and U8275 (N_8275,N_8037,N_8064);
nor U8276 (N_8276,N_8051,N_8175);
xor U8277 (N_8277,N_8094,N_8081);
or U8278 (N_8278,N_8125,N_8194);
nor U8279 (N_8279,N_8083,N_8166);
nor U8280 (N_8280,N_8074,N_8119);
or U8281 (N_8281,N_8049,N_8001);
nand U8282 (N_8282,N_8128,N_8192);
nand U8283 (N_8283,N_8059,N_8044);
nand U8284 (N_8284,N_8075,N_8193);
or U8285 (N_8285,N_8184,N_8047);
nor U8286 (N_8286,N_8054,N_8041);
nor U8287 (N_8287,N_8185,N_8174);
nor U8288 (N_8288,N_8122,N_8048);
nand U8289 (N_8289,N_8056,N_8004);
or U8290 (N_8290,N_8007,N_8082);
xor U8291 (N_8291,N_8113,N_8104);
nand U8292 (N_8292,N_8010,N_8077);
nor U8293 (N_8293,N_8093,N_8070);
nor U8294 (N_8294,N_8143,N_8133);
nor U8295 (N_8295,N_8199,N_8090);
xor U8296 (N_8296,N_8179,N_8181);
nand U8297 (N_8297,N_8152,N_8015);
nand U8298 (N_8298,N_8011,N_8134);
nor U8299 (N_8299,N_8013,N_8117);
or U8300 (N_8300,N_8040,N_8163);
nor U8301 (N_8301,N_8093,N_8000);
nor U8302 (N_8302,N_8144,N_8065);
or U8303 (N_8303,N_8051,N_8086);
xnor U8304 (N_8304,N_8024,N_8045);
and U8305 (N_8305,N_8184,N_8131);
nor U8306 (N_8306,N_8009,N_8092);
nand U8307 (N_8307,N_8047,N_8013);
xor U8308 (N_8308,N_8056,N_8053);
and U8309 (N_8309,N_8020,N_8090);
and U8310 (N_8310,N_8020,N_8146);
xor U8311 (N_8311,N_8140,N_8049);
xor U8312 (N_8312,N_8068,N_8176);
xnor U8313 (N_8313,N_8186,N_8172);
xnor U8314 (N_8314,N_8079,N_8030);
nor U8315 (N_8315,N_8150,N_8165);
nand U8316 (N_8316,N_8061,N_8187);
or U8317 (N_8317,N_8146,N_8062);
nand U8318 (N_8318,N_8005,N_8130);
or U8319 (N_8319,N_8127,N_8144);
or U8320 (N_8320,N_8178,N_8171);
nand U8321 (N_8321,N_8020,N_8073);
nand U8322 (N_8322,N_8180,N_8007);
nor U8323 (N_8323,N_8113,N_8016);
xor U8324 (N_8324,N_8078,N_8175);
and U8325 (N_8325,N_8086,N_8041);
nor U8326 (N_8326,N_8037,N_8028);
nor U8327 (N_8327,N_8091,N_8067);
nand U8328 (N_8328,N_8139,N_8063);
nor U8329 (N_8329,N_8022,N_8055);
xor U8330 (N_8330,N_8014,N_8037);
nand U8331 (N_8331,N_8150,N_8130);
nor U8332 (N_8332,N_8176,N_8192);
or U8333 (N_8333,N_8077,N_8155);
nand U8334 (N_8334,N_8099,N_8007);
xor U8335 (N_8335,N_8111,N_8082);
xnor U8336 (N_8336,N_8096,N_8007);
xor U8337 (N_8337,N_8145,N_8116);
nand U8338 (N_8338,N_8084,N_8144);
and U8339 (N_8339,N_8148,N_8044);
or U8340 (N_8340,N_8004,N_8130);
xor U8341 (N_8341,N_8104,N_8043);
nand U8342 (N_8342,N_8145,N_8071);
or U8343 (N_8343,N_8179,N_8169);
xor U8344 (N_8344,N_8146,N_8011);
or U8345 (N_8345,N_8095,N_8019);
or U8346 (N_8346,N_8132,N_8155);
nand U8347 (N_8347,N_8170,N_8127);
xor U8348 (N_8348,N_8058,N_8118);
nand U8349 (N_8349,N_8012,N_8015);
xnor U8350 (N_8350,N_8129,N_8042);
nor U8351 (N_8351,N_8132,N_8168);
and U8352 (N_8352,N_8114,N_8010);
nor U8353 (N_8353,N_8086,N_8037);
nand U8354 (N_8354,N_8012,N_8040);
nand U8355 (N_8355,N_8032,N_8176);
nand U8356 (N_8356,N_8023,N_8021);
xnor U8357 (N_8357,N_8189,N_8106);
nor U8358 (N_8358,N_8082,N_8076);
nand U8359 (N_8359,N_8162,N_8132);
xnor U8360 (N_8360,N_8137,N_8100);
nor U8361 (N_8361,N_8121,N_8055);
nor U8362 (N_8362,N_8149,N_8171);
and U8363 (N_8363,N_8116,N_8127);
xor U8364 (N_8364,N_8023,N_8082);
or U8365 (N_8365,N_8049,N_8071);
and U8366 (N_8366,N_8022,N_8137);
nor U8367 (N_8367,N_8115,N_8140);
xor U8368 (N_8368,N_8037,N_8171);
nor U8369 (N_8369,N_8030,N_8011);
nand U8370 (N_8370,N_8031,N_8024);
nor U8371 (N_8371,N_8152,N_8194);
and U8372 (N_8372,N_8079,N_8174);
nor U8373 (N_8373,N_8005,N_8199);
and U8374 (N_8374,N_8054,N_8046);
nand U8375 (N_8375,N_8068,N_8140);
or U8376 (N_8376,N_8066,N_8128);
nor U8377 (N_8377,N_8034,N_8173);
nor U8378 (N_8378,N_8091,N_8074);
and U8379 (N_8379,N_8068,N_8074);
xor U8380 (N_8380,N_8056,N_8024);
xor U8381 (N_8381,N_8076,N_8045);
nor U8382 (N_8382,N_8011,N_8185);
nand U8383 (N_8383,N_8016,N_8126);
nor U8384 (N_8384,N_8087,N_8188);
xor U8385 (N_8385,N_8167,N_8189);
or U8386 (N_8386,N_8116,N_8192);
nand U8387 (N_8387,N_8084,N_8192);
and U8388 (N_8388,N_8005,N_8174);
and U8389 (N_8389,N_8173,N_8066);
nand U8390 (N_8390,N_8162,N_8046);
xor U8391 (N_8391,N_8186,N_8120);
xor U8392 (N_8392,N_8144,N_8129);
nor U8393 (N_8393,N_8062,N_8139);
xor U8394 (N_8394,N_8014,N_8072);
nor U8395 (N_8395,N_8082,N_8096);
xor U8396 (N_8396,N_8137,N_8023);
and U8397 (N_8397,N_8102,N_8038);
and U8398 (N_8398,N_8104,N_8130);
and U8399 (N_8399,N_8129,N_8154);
and U8400 (N_8400,N_8247,N_8397);
or U8401 (N_8401,N_8269,N_8348);
nor U8402 (N_8402,N_8284,N_8288);
and U8403 (N_8403,N_8390,N_8230);
xor U8404 (N_8404,N_8290,N_8380);
or U8405 (N_8405,N_8398,N_8391);
nand U8406 (N_8406,N_8220,N_8366);
or U8407 (N_8407,N_8212,N_8201);
and U8408 (N_8408,N_8299,N_8250);
nand U8409 (N_8409,N_8297,N_8294);
nor U8410 (N_8410,N_8200,N_8354);
and U8411 (N_8411,N_8218,N_8272);
nor U8412 (N_8412,N_8371,N_8336);
and U8413 (N_8413,N_8375,N_8232);
and U8414 (N_8414,N_8223,N_8275);
or U8415 (N_8415,N_8238,N_8339);
nand U8416 (N_8416,N_8393,N_8304);
or U8417 (N_8417,N_8328,N_8251);
nand U8418 (N_8418,N_8312,N_8327);
or U8419 (N_8419,N_8226,N_8210);
or U8420 (N_8420,N_8314,N_8244);
nand U8421 (N_8421,N_8357,N_8307);
or U8422 (N_8422,N_8236,N_8285);
or U8423 (N_8423,N_8289,N_8319);
nand U8424 (N_8424,N_8264,N_8260);
xor U8425 (N_8425,N_8326,N_8280);
nor U8426 (N_8426,N_8242,N_8266);
and U8427 (N_8427,N_8360,N_8370);
xnor U8428 (N_8428,N_8240,N_8325);
nand U8429 (N_8429,N_8332,N_8346);
or U8430 (N_8430,N_8237,N_8386);
nor U8431 (N_8431,N_8338,N_8355);
or U8432 (N_8432,N_8287,N_8335);
xnor U8433 (N_8433,N_8234,N_8377);
nor U8434 (N_8434,N_8282,N_8270);
or U8435 (N_8435,N_8296,N_8227);
nor U8436 (N_8436,N_8372,N_8235);
or U8437 (N_8437,N_8381,N_8350);
and U8438 (N_8438,N_8363,N_8383);
and U8439 (N_8439,N_8343,N_8208);
nor U8440 (N_8440,N_8376,N_8337);
xnor U8441 (N_8441,N_8379,N_8259);
nor U8442 (N_8442,N_8359,N_8263);
nand U8443 (N_8443,N_8249,N_8274);
nor U8444 (N_8444,N_8229,N_8388);
xor U8445 (N_8445,N_8394,N_8253);
xor U8446 (N_8446,N_8222,N_8203);
and U8447 (N_8447,N_8323,N_8311);
and U8448 (N_8448,N_8301,N_8246);
or U8449 (N_8449,N_8243,N_8308);
xnor U8450 (N_8450,N_8293,N_8356);
and U8451 (N_8451,N_8331,N_8305);
or U8452 (N_8452,N_8310,N_8255);
or U8453 (N_8453,N_8369,N_8216);
and U8454 (N_8454,N_8362,N_8265);
and U8455 (N_8455,N_8329,N_8281);
and U8456 (N_8456,N_8349,N_8277);
and U8457 (N_8457,N_8286,N_8262);
nor U8458 (N_8458,N_8248,N_8302);
xnor U8459 (N_8459,N_8387,N_8291);
and U8460 (N_8460,N_8267,N_8330);
xnor U8461 (N_8461,N_8206,N_8231);
nand U8462 (N_8462,N_8368,N_8258);
nand U8463 (N_8463,N_8384,N_8365);
xor U8464 (N_8464,N_8351,N_8341);
and U8465 (N_8465,N_8217,N_8340);
nor U8466 (N_8466,N_8389,N_8252);
nor U8467 (N_8467,N_8205,N_8345);
and U8468 (N_8468,N_8261,N_8295);
or U8469 (N_8469,N_8306,N_8202);
and U8470 (N_8470,N_8382,N_8333);
or U8471 (N_8471,N_8395,N_8268);
or U8472 (N_8472,N_8298,N_8373);
or U8473 (N_8473,N_8344,N_8211);
xor U8474 (N_8474,N_8317,N_8313);
nand U8475 (N_8475,N_8233,N_8241);
nand U8476 (N_8476,N_8353,N_8322);
and U8477 (N_8477,N_8300,N_8367);
xnor U8478 (N_8478,N_8320,N_8292);
nor U8479 (N_8479,N_8221,N_8224);
and U8480 (N_8480,N_8358,N_8399);
or U8481 (N_8481,N_8257,N_8213);
or U8482 (N_8482,N_8276,N_8385);
xnor U8483 (N_8483,N_8374,N_8342);
and U8484 (N_8484,N_8228,N_8347);
nand U8485 (N_8485,N_8303,N_8309);
nand U8486 (N_8486,N_8209,N_8271);
xor U8487 (N_8487,N_8396,N_8392);
nor U8488 (N_8488,N_8214,N_8279);
nand U8489 (N_8489,N_8256,N_8215);
or U8490 (N_8490,N_8225,N_8318);
or U8491 (N_8491,N_8239,N_8204);
and U8492 (N_8492,N_8324,N_8207);
nand U8493 (N_8493,N_8283,N_8352);
xor U8494 (N_8494,N_8378,N_8254);
xor U8495 (N_8495,N_8219,N_8361);
and U8496 (N_8496,N_8334,N_8316);
nand U8497 (N_8497,N_8321,N_8273);
nand U8498 (N_8498,N_8364,N_8245);
or U8499 (N_8499,N_8278,N_8315);
or U8500 (N_8500,N_8254,N_8312);
and U8501 (N_8501,N_8369,N_8366);
or U8502 (N_8502,N_8237,N_8358);
xnor U8503 (N_8503,N_8334,N_8256);
or U8504 (N_8504,N_8265,N_8245);
xnor U8505 (N_8505,N_8322,N_8340);
and U8506 (N_8506,N_8376,N_8387);
nor U8507 (N_8507,N_8374,N_8307);
nand U8508 (N_8508,N_8318,N_8378);
nor U8509 (N_8509,N_8251,N_8368);
nor U8510 (N_8510,N_8379,N_8374);
xor U8511 (N_8511,N_8319,N_8367);
xor U8512 (N_8512,N_8344,N_8373);
and U8513 (N_8513,N_8367,N_8211);
nor U8514 (N_8514,N_8329,N_8297);
or U8515 (N_8515,N_8347,N_8244);
or U8516 (N_8516,N_8309,N_8370);
nor U8517 (N_8517,N_8319,N_8242);
xor U8518 (N_8518,N_8212,N_8261);
and U8519 (N_8519,N_8249,N_8289);
nor U8520 (N_8520,N_8371,N_8272);
nor U8521 (N_8521,N_8217,N_8341);
nand U8522 (N_8522,N_8228,N_8216);
and U8523 (N_8523,N_8325,N_8309);
and U8524 (N_8524,N_8288,N_8294);
nand U8525 (N_8525,N_8227,N_8349);
nor U8526 (N_8526,N_8375,N_8201);
or U8527 (N_8527,N_8319,N_8379);
nand U8528 (N_8528,N_8362,N_8368);
nand U8529 (N_8529,N_8300,N_8290);
and U8530 (N_8530,N_8387,N_8282);
or U8531 (N_8531,N_8276,N_8263);
nor U8532 (N_8532,N_8235,N_8252);
nor U8533 (N_8533,N_8258,N_8398);
nor U8534 (N_8534,N_8254,N_8250);
nor U8535 (N_8535,N_8232,N_8211);
xor U8536 (N_8536,N_8239,N_8357);
or U8537 (N_8537,N_8371,N_8206);
or U8538 (N_8538,N_8312,N_8274);
nor U8539 (N_8539,N_8302,N_8297);
and U8540 (N_8540,N_8261,N_8368);
nand U8541 (N_8541,N_8308,N_8345);
or U8542 (N_8542,N_8212,N_8384);
and U8543 (N_8543,N_8275,N_8334);
or U8544 (N_8544,N_8283,N_8378);
xnor U8545 (N_8545,N_8355,N_8383);
and U8546 (N_8546,N_8283,N_8364);
nor U8547 (N_8547,N_8260,N_8315);
nand U8548 (N_8548,N_8323,N_8398);
and U8549 (N_8549,N_8376,N_8303);
nor U8550 (N_8550,N_8231,N_8369);
or U8551 (N_8551,N_8278,N_8306);
and U8552 (N_8552,N_8396,N_8357);
or U8553 (N_8553,N_8275,N_8242);
and U8554 (N_8554,N_8328,N_8337);
nand U8555 (N_8555,N_8394,N_8368);
xor U8556 (N_8556,N_8214,N_8363);
or U8557 (N_8557,N_8324,N_8252);
nand U8558 (N_8558,N_8312,N_8361);
nand U8559 (N_8559,N_8320,N_8233);
or U8560 (N_8560,N_8374,N_8237);
nor U8561 (N_8561,N_8394,N_8369);
nor U8562 (N_8562,N_8311,N_8377);
or U8563 (N_8563,N_8256,N_8304);
nor U8564 (N_8564,N_8362,N_8261);
or U8565 (N_8565,N_8394,N_8249);
nor U8566 (N_8566,N_8283,N_8292);
and U8567 (N_8567,N_8357,N_8295);
or U8568 (N_8568,N_8260,N_8299);
xnor U8569 (N_8569,N_8258,N_8286);
nand U8570 (N_8570,N_8378,N_8355);
or U8571 (N_8571,N_8205,N_8341);
xor U8572 (N_8572,N_8307,N_8238);
or U8573 (N_8573,N_8313,N_8201);
nor U8574 (N_8574,N_8386,N_8260);
xor U8575 (N_8575,N_8208,N_8227);
and U8576 (N_8576,N_8341,N_8352);
nor U8577 (N_8577,N_8397,N_8208);
nand U8578 (N_8578,N_8321,N_8293);
or U8579 (N_8579,N_8288,N_8202);
or U8580 (N_8580,N_8315,N_8374);
or U8581 (N_8581,N_8207,N_8200);
nand U8582 (N_8582,N_8352,N_8351);
xor U8583 (N_8583,N_8399,N_8234);
nand U8584 (N_8584,N_8397,N_8388);
and U8585 (N_8585,N_8338,N_8261);
nor U8586 (N_8586,N_8289,N_8232);
nand U8587 (N_8587,N_8233,N_8342);
and U8588 (N_8588,N_8237,N_8367);
and U8589 (N_8589,N_8361,N_8287);
and U8590 (N_8590,N_8394,N_8383);
xnor U8591 (N_8591,N_8243,N_8239);
and U8592 (N_8592,N_8230,N_8296);
and U8593 (N_8593,N_8242,N_8365);
nor U8594 (N_8594,N_8234,N_8205);
or U8595 (N_8595,N_8322,N_8308);
nor U8596 (N_8596,N_8249,N_8365);
nand U8597 (N_8597,N_8301,N_8200);
xnor U8598 (N_8598,N_8256,N_8259);
nor U8599 (N_8599,N_8310,N_8338);
and U8600 (N_8600,N_8567,N_8507);
nand U8601 (N_8601,N_8548,N_8505);
and U8602 (N_8602,N_8572,N_8542);
or U8603 (N_8603,N_8487,N_8556);
and U8604 (N_8604,N_8468,N_8416);
or U8605 (N_8605,N_8521,N_8410);
nand U8606 (N_8606,N_8418,N_8591);
nand U8607 (N_8607,N_8477,N_8497);
or U8608 (N_8608,N_8461,N_8404);
or U8609 (N_8609,N_8547,N_8425);
xor U8610 (N_8610,N_8411,N_8440);
xor U8611 (N_8611,N_8503,N_8500);
xor U8612 (N_8612,N_8463,N_8573);
nor U8613 (N_8613,N_8594,N_8441);
nand U8614 (N_8614,N_8536,N_8589);
or U8615 (N_8615,N_8575,N_8595);
and U8616 (N_8616,N_8563,N_8517);
xor U8617 (N_8617,N_8488,N_8480);
xnor U8618 (N_8618,N_8439,N_8535);
or U8619 (N_8619,N_8454,N_8522);
or U8620 (N_8620,N_8590,N_8415);
xor U8621 (N_8621,N_8466,N_8574);
xnor U8622 (N_8622,N_8495,N_8592);
nor U8623 (N_8623,N_8450,N_8537);
or U8624 (N_8624,N_8509,N_8599);
nor U8625 (N_8625,N_8428,N_8460);
and U8626 (N_8626,N_8456,N_8555);
and U8627 (N_8627,N_8467,N_8593);
or U8628 (N_8628,N_8498,N_8596);
xor U8629 (N_8629,N_8558,N_8557);
and U8630 (N_8630,N_8578,N_8422);
nor U8631 (N_8631,N_8524,N_8502);
xor U8632 (N_8632,N_8570,N_8526);
nor U8633 (N_8633,N_8427,N_8436);
and U8634 (N_8634,N_8409,N_8512);
nor U8635 (N_8635,N_8530,N_8501);
and U8636 (N_8636,N_8519,N_8402);
nor U8637 (N_8637,N_8475,N_8464);
nand U8638 (N_8638,N_8438,N_8479);
nand U8639 (N_8639,N_8420,N_8508);
or U8640 (N_8640,N_8499,N_8518);
nor U8641 (N_8641,N_8474,N_8514);
nand U8642 (N_8642,N_8523,N_8442);
xor U8643 (N_8643,N_8577,N_8545);
nand U8644 (N_8644,N_8485,N_8493);
xnor U8645 (N_8645,N_8412,N_8424);
nor U8646 (N_8646,N_8445,N_8581);
and U8647 (N_8647,N_8433,N_8515);
xnor U8648 (N_8648,N_8403,N_8564);
or U8649 (N_8649,N_8559,N_8587);
or U8650 (N_8650,N_8554,N_8571);
xnor U8651 (N_8651,N_8527,N_8562);
or U8652 (N_8652,N_8486,N_8455);
nor U8653 (N_8653,N_8490,N_8451);
xor U8654 (N_8654,N_8429,N_8452);
xnor U8655 (N_8655,N_8470,N_8588);
nor U8656 (N_8656,N_8489,N_8494);
and U8657 (N_8657,N_8584,N_8435);
nor U8658 (N_8658,N_8506,N_8446);
and U8659 (N_8659,N_8414,N_8560);
nor U8660 (N_8660,N_8525,N_8473);
and U8661 (N_8661,N_8462,N_8413);
xnor U8662 (N_8662,N_8434,N_8417);
xor U8663 (N_8663,N_8476,N_8566);
or U8664 (N_8664,N_8569,N_8437);
and U8665 (N_8665,N_8528,N_8408);
nand U8666 (N_8666,N_8510,N_8449);
nor U8667 (N_8667,N_8576,N_8543);
xor U8668 (N_8668,N_8597,N_8516);
and U8669 (N_8669,N_8544,N_8586);
or U8670 (N_8670,N_8459,N_8419);
nand U8671 (N_8671,N_8580,N_8481);
nor U8672 (N_8672,N_8541,N_8540);
nor U8673 (N_8673,N_8478,N_8453);
xnor U8674 (N_8674,N_8484,N_8400);
nor U8675 (N_8675,N_8407,N_8423);
and U8676 (N_8676,N_8471,N_8447);
xor U8677 (N_8677,N_8483,N_8561);
xnor U8678 (N_8678,N_8458,N_8469);
xor U8679 (N_8679,N_8529,N_8430);
or U8680 (N_8680,N_8465,N_8550);
nand U8681 (N_8681,N_8457,N_8504);
nand U8682 (N_8682,N_8579,N_8539);
nor U8683 (N_8683,N_8496,N_8472);
and U8684 (N_8684,N_8491,N_8582);
or U8685 (N_8685,N_8549,N_8405);
and U8686 (N_8686,N_8533,N_8565);
xor U8687 (N_8687,N_8406,N_8598);
and U8688 (N_8688,N_8511,N_8426);
and U8689 (N_8689,N_8482,N_8546);
nand U8690 (N_8690,N_8583,N_8531);
or U8691 (N_8691,N_8401,N_8534);
nand U8692 (N_8692,N_8492,N_8443);
xnor U8693 (N_8693,N_8553,N_8421);
nand U8694 (N_8694,N_8431,N_8552);
and U8695 (N_8695,N_8448,N_8568);
nor U8696 (N_8696,N_8444,N_8513);
or U8697 (N_8697,N_8532,N_8538);
and U8698 (N_8698,N_8432,N_8551);
xnor U8699 (N_8699,N_8520,N_8585);
xor U8700 (N_8700,N_8462,N_8496);
or U8701 (N_8701,N_8594,N_8507);
nor U8702 (N_8702,N_8567,N_8466);
or U8703 (N_8703,N_8496,N_8453);
nor U8704 (N_8704,N_8598,N_8533);
or U8705 (N_8705,N_8578,N_8552);
nand U8706 (N_8706,N_8572,N_8427);
xor U8707 (N_8707,N_8460,N_8489);
xor U8708 (N_8708,N_8569,N_8473);
nor U8709 (N_8709,N_8536,N_8402);
or U8710 (N_8710,N_8514,N_8425);
nor U8711 (N_8711,N_8464,N_8471);
xnor U8712 (N_8712,N_8498,N_8559);
xnor U8713 (N_8713,N_8483,N_8440);
nand U8714 (N_8714,N_8434,N_8480);
nand U8715 (N_8715,N_8511,N_8578);
nand U8716 (N_8716,N_8483,N_8599);
and U8717 (N_8717,N_8486,N_8566);
and U8718 (N_8718,N_8431,N_8424);
nand U8719 (N_8719,N_8467,N_8478);
and U8720 (N_8720,N_8405,N_8496);
nor U8721 (N_8721,N_8505,N_8568);
and U8722 (N_8722,N_8452,N_8554);
xnor U8723 (N_8723,N_8496,N_8411);
and U8724 (N_8724,N_8574,N_8458);
nand U8725 (N_8725,N_8583,N_8478);
nor U8726 (N_8726,N_8459,N_8452);
or U8727 (N_8727,N_8427,N_8562);
or U8728 (N_8728,N_8512,N_8425);
xnor U8729 (N_8729,N_8491,N_8480);
nor U8730 (N_8730,N_8418,N_8463);
and U8731 (N_8731,N_8595,N_8509);
nor U8732 (N_8732,N_8457,N_8543);
xnor U8733 (N_8733,N_8473,N_8591);
nor U8734 (N_8734,N_8573,N_8581);
xor U8735 (N_8735,N_8494,N_8416);
and U8736 (N_8736,N_8589,N_8498);
and U8737 (N_8737,N_8430,N_8520);
and U8738 (N_8738,N_8583,N_8405);
or U8739 (N_8739,N_8477,N_8464);
xor U8740 (N_8740,N_8554,N_8460);
and U8741 (N_8741,N_8594,N_8545);
or U8742 (N_8742,N_8556,N_8428);
nor U8743 (N_8743,N_8586,N_8581);
nand U8744 (N_8744,N_8417,N_8591);
or U8745 (N_8745,N_8543,N_8495);
xor U8746 (N_8746,N_8438,N_8407);
or U8747 (N_8747,N_8568,N_8518);
xor U8748 (N_8748,N_8589,N_8522);
xor U8749 (N_8749,N_8552,N_8517);
xor U8750 (N_8750,N_8512,N_8584);
nor U8751 (N_8751,N_8571,N_8486);
xnor U8752 (N_8752,N_8411,N_8491);
or U8753 (N_8753,N_8410,N_8535);
nand U8754 (N_8754,N_8533,N_8563);
nor U8755 (N_8755,N_8503,N_8481);
nand U8756 (N_8756,N_8524,N_8456);
xnor U8757 (N_8757,N_8564,N_8473);
or U8758 (N_8758,N_8578,N_8493);
nand U8759 (N_8759,N_8446,N_8436);
xor U8760 (N_8760,N_8499,N_8486);
nor U8761 (N_8761,N_8431,N_8535);
nor U8762 (N_8762,N_8514,N_8548);
nand U8763 (N_8763,N_8454,N_8528);
and U8764 (N_8764,N_8512,N_8498);
or U8765 (N_8765,N_8570,N_8467);
and U8766 (N_8766,N_8421,N_8480);
nor U8767 (N_8767,N_8452,N_8516);
nor U8768 (N_8768,N_8478,N_8505);
nor U8769 (N_8769,N_8479,N_8406);
nand U8770 (N_8770,N_8535,N_8448);
and U8771 (N_8771,N_8517,N_8519);
and U8772 (N_8772,N_8495,N_8590);
xnor U8773 (N_8773,N_8529,N_8566);
and U8774 (N_8774,N_8472,N_8481);
nor U8775 (N_8775,N_8516,N_8509);
or U8776 (N_8776,N_8423,N_8419);
xor U8777 (N_8777,N_8471,N_8579);
nor U8778 (N_8778,N_8481,N_8568);
xor U8779 (N_8779,N_8588,N_8565);
and U8780 (N_8780,N_8427,N_8551);
or U8781 (N_8781,N_8441,N_8414);
xor U8782 (N_8782,N_8542,N_8423);
or U8783 (N_8783,N_8509,N_8420);
nand U8784 (N_8784,N_8593,N_8430);
or U8785 (N_8785,N_8472,N_8416);
xnor U8786 (N_8786,N_8530,N_8419);
and U8787 (N_8787,N_8409,N_8437);
xor U8788 (N_8788,N_8436,N_8561);
nor U8789 (N_8789,N_8553,N_8459);
and U8790 (N_8790,N_8527,N_8575);
nor U8791 (N_8791,N_8529,N_8599);
nor U8792 (N_8792,N_8451,N_8507);
nand U8793 (N_8793,N_8513,N_8450);
or U8794 (N_8794,N_8413,N_8449);
nor U8795 (N_8795,N_8473,N_8587);
nand U8796 (N_8796,N_8461,N_8528);
and U8797 (N_8797,N_8490,N_8582);
nor U8798 (N_8798,N_8528,N_8416);
nand U8799 (N_8799,N_8495,N_8560);
xor U8800 (N_8800,N_8657,N_8621);
nor U8801 (N_8801,N_8706,N_8789);
and U8802 (N_8802,N_8780,N_8645);
or U8803 (N_8803,N_8669,N_8741);
nand U8804 (N_8804,N_8748,N_8757);
or U8805 (N_8805,N_8649,N_8668);
nand U8806 (N_8806,N_8689,N_8790);
or U8807 (N_8807,N_8730,N_8746);
nor U8808 (N_8808,N_8758,N_8788);
or U8809 (N_8809,N_8753,N_8756);
xor U8810 (N_8810,N_8696,N_8615);
or U8811 (N_8811,N_8708,N_8796);
or U8812 (N_8812,N_8760,N_8743);
xor U8813 (N_8813,N_8769,N_8719);
xnor U8814 (N_8814,N_8670,N_8761);
and U8815 (N_8815,N_8784,N_8699);
or U8816 (N_8816,N_8771,N_8609);
xnor U8817 (N_8817,N_8685,N_8713);
nor U8818 (N_8818,N_8722,N_8617);
or U8819 (N_8819,N_8791,N_8750);
xnor U8820 (N_8820,N_8635,N_8684);
xnor U8821 (N_8821,N_8658,N_8785);
nand U8822 (N_8822,N_8659,N_8720);
nand U8823 (N_8823,N_8608,N_8636);
or U8824 (N_8824,N_8717,N_8792);
nor U8825 (N_8825,N_8798,N_8714);
or U8826 (N_8826,N_8775,N_8728);
nor U8827 (N_8827,N_8677,N_8628);
nor U8828 (N_8828,N_8625,N_8783);
and U8829 (N_8829,N_8698,N_8755);
nor U8830 (N_8830,N_8733,N_8622);
and U8831 (N_8831,N_8680,N_8715);
xor U8832 (N_8832,N_8671,N_8744);
nand U8833 (N_8833,N_8793,N_8732);
or U8834 (N_8834,N_8781,N_8778);
xnor U8835 (N_8835,N_8774,N_8773);
or U8836 (N_8836,N_8690,N_8692);
xor U8837 (N_8837,N_8770,N_8694);
and U8838 (N_8838,N_8716,N_8603);
nor U8839 (N_8839,N_8766,N_8644);
or U8840 (N_8840,N_8754,N_8745);
xnor U8841 (N_8841,N_8772,N_8723);
nand U8842 (N_8842,N_8727,N_8633);
xor U8843 (N_8843,N_8620,N_8799);
or U8844 (N_8844,N_8660,N_8638);
and U8845 (N_8845,N_8643,N_8786);
or U8846 (N_8846,N_8678,N_8604);
and U8847 (N_8847,N_8616,N_8724);
xnor U8848 (N_8848,N_8797,N_8777);
and U8849 (N_8849,N_8752,N_8679);
or U8850 (N_8850,N_8665,N_8632);
and U8851 (N_8851,N_8709,N_8647);
and U8852 (N_8852,N_8729,N_8652);
xnor U8853 (N_8853,N_8629,N_8653);
and U8854 (N_8854,N_8641,N_8623);
or U8855 (N_8855,N_8712,N_8639);
and U8856 (N_8856,N_8740,N_8702);
and U8857 (N_8857,N_8686,N_8705);
nand U8858 (N_8858,N_8613,N_8704);
nand U8859 (N_8859,N_8606,N_8640);
nand U8860 (N_8860,N_8612,N_8718);
nand U8861 (N_8861,N_8667,N_8768);
or U8862 (N_8862,N_8666,N_8610);
xnor U8863 (N_8863,N_8675,N_8735);
nor U8864 (N_8864,N_8742,N_8749);
and U8865 (N_8865,N_8600,N_8767);
nand U8866 (N_8866,N_8630,N_8683);
xor U8867 (N_8867,N_8654,N_8765);
nor U8868 (N_8868,N_8751,N_8782);
xor U8869 (N_8869,N_8618,N_8626);
xor U8870 (N_8870,N_8619,N_8726);
or U8871 (N_8871,N_8731,N_8602);
nor U8872 (N_8872,N_8736,N_8721);
or U8873 (N_8873,N_8676,N_8663);
xnor U8874 (N_8874,N_8701,N_8725);
xor U8875 (N_8875,N_8664,N_8651);
nand U8876 (N_8876,N_8738,N_8648);
or U8877 (N_8877,N_8673,N_8764);
nor U8878 (N_8878,N_8697,N_8607);
xnor U8879 (N_8879,N_8688,N_8627);
nand U8880 (N_8880,N_8687,N_8787);
nand U8881 (N_8881,N_8637,N_8703);
nand U8882 (N_8882,N_8650,N_8734);
xnor U8883 (N_8883,N_8776,N_8656);
nor U8884 (N_8884,N_8691,N_8672);
nand U8885 (N_8885,N_8762,N_8759);
or U8886 (N_8886,N_8682,N_8710);
nor U8887 (N_8887,N_8655,N_8601);
and U8888 (N_8888,N_8693,N_8707);
nor U8889 (N_8889,N_8646,N_8763);
nand U8890 (N_8890,N_8794,N_8674);
nand U8891 (N_8891,N_8700,N_8711);
or U8892 (N_8892,N_8695,N_8779);
nor U8893 (N_8893,N_8795,N_8631);
or U8894 (N_8894,N_8642,N_8605);
xor U8895 (N_8895,N_8747,N_8662);
nor U8896 (N_8896,N_8614,N_8681);
xor U8897 (N_8897,N_8611,N_8739);
nor U8898 (N_8898,N_8624,N_8661);
nand U8899 (N_8899,N_8737,N_8634);
or U8900 (N_8900,N_8716,N_8753);
and U8901 (N_8901,N_8747,N_8732);
nand U8902 (N_8902,N_8612,N_8725);
or U8903 (N_8903,N_8672,N_8645);
or U8904 (N_8904,N_8689,N_8664);
and U8905 (N_8905,N_8608,N_8697);
xor U8906 (N_8906,N_8725,N_8711);
and U8907 (N_8907,N_8732,N_8768);
xnor U8908 (N_8908,N_8772,N_8714);
or U8909 (N_8909,N_8674,N_8798);
xor U8910 (N_8910,N_8699,N_8639);
nor U8911 (N_8911,N_8683,N_8695);
or U8912 (N_8912,N_8693,N_8699);
nor U8913 (N_8913,N_8722,N_8607);
xor U8914 (N_8914,N_8671,N_8638);
nor U8915 (N_8915,N_8715,N_8664);
nor U8916 (N_8916,N_8712,N_8641);
xnor U8917 (N_8917,N_8646,N_8666);
nand U8918 (N_8918,N_8793,N_8724);
xnor U8919 (N_8919,N_8654,N_8709);
and U8920 (N_8920,N_8602,N_8725);
xnor U8921 (N_8921,N_8781,N_8664);
and U8922 (N_8922,N_8627,N_8718);
or U8923 (N_8923,N_8786,N_8764);
and U8924 (N_8924,N_8641,N_8637);
and U8925 (N_8925,N_8725,N_8796);
nor U8926 (N_8926,N_8692,N_8700);
xor U8927 (N_8927,N_8671,N_8747);
nand U8928 (N_8928,N_8767,N_8770);
xor U8929 (N_8929,N_8624,N_8628);
nor U8930 (N_8930,N_8613,N_8771);
and U8931 (N_8931,N_8736,N_8678);
and U8932 (N_8932,N_8729,N_8782);
nor U8933 (N_8933,N_8662,N_8721);
nor U8934 (N_8934,N_8640,N_8668);
or U8935 (N_8935,N_8628,N_8745);
nor U8936 (N_8936,N_8702,N_8774);
nor U8937 (N_8937,N_8643,N_8703);
xor U8938 (N_8938,N_8791,N_8655);
and U8939 (N_8939,N_8654,N_8669);
and U8940 (N_8940,N_8625,N_8660);
nor U8941 (N_8941,N_8774,N_8784);
xor U8942 (N_8942,N_8619,N_8613);
and U8943 (N_8943,N_8718,N_8618);
nand U8944 (N_8944,N_8759,N_8611);
nor U8945 (N_8945,N_8706,N_8791);
xor U8946 (N_8946,N_8630,N_8728);
nand U8947 (N_8947,N_8697,N_8719);
nor U8948 (N_8948,N_8655,N_8709);
nand U8949 (N_8949,N_8717,N_8667);
nor U8950 (N_8950,N_8628,N_8672);
and U8951 (N_8951,N_8669,N_8720);
or U8952 (N_8952,N_8679,N_8770);
nor U8953 (N_8953,N_8660,N_8669);
nand U8954 (N_8954,N_8673,N_8729);
nand U8955 (N_8955,N_8643,N_8691);
and U8956 (N_8956,N_8680,N_8692);
or U8957 (N_8957,N_8739,N_8641);
and U8958 (N_8958,N_8716,N_8751);
xnor U8959 (N_8959,N_8610,N_8759);
and U8960 (N_8960,N_8694,N_8711);
or U8961 (N_8961,N_8691,N_8770);
or U8962 (N_8962,N_8798,N_8794);
xor U8963 (N_8963,N_8600,N_8766);
nor U8964 (N_8964,N_8628,N_8728);
or U8965 (N_8965,N_8719,N_8624);
xnor U8966 (N_8966,N_8628,N_8794);
nand U8967 (N_8967,N_8640,N_8756);
xnor U8968 (N_8968,N_8707,N_8715);
or U8969 (N_8969,N_8612,N_8742);
nand U8970 (N_8970,N_8795,N_8681);
nor U8971 (N_8971,N_8653,N_8775);
and U8972 (N_8972,N_8721,N_8618);
nor U8973 (N_8973,N_8734,N_8601);
xnor U8974 (N_8974,N_8681,N_8703);
nand U8975 (N_8975,N_8772,N_8636);
nor U8976 (N_8976,N_8711,N_8669);
xor U8977 (N_8977,N_8755,N_8634);
nor U8978 (N_8978,N_8669,N_8771);
and U8979 (N_8979,N_8648,N_8709);
xor U8980 (N_8980,N_8663,N_8690);
nand U8981 (N_8981,N_8760,N_8645);
nor U8982 (N_8982,N_8626,N_8764);
and U8983 (N_8983,N_8792,N_8636);
nand U8984 (N_8984,N_8610,N_8649);
nand U8985 (N_8985,N_8669,N_8698);
nor U8986 (N_8986,N_8682,N_8696);
nor U8987 (N_8987,N_8715,N_8710);
nand U8988 (N_8988,N_8774,N_8722);
nor U8989 (N_8989,N_8787,N_8671);
nand U8990 (N_8990,N_8735,N_8707);
or U8991 (N_8991,N_8610,N_8706);
and U8992 (N_8992,N_8692,N_8759);
nand U8993 (N_8993,N_8772,N_8786);
nor U8994 (N_8994,N_8687,N_8694);
or U8995 (N_8995,N_8692,N_8729);
nor U8996 (N_8996,N_8661,N_8745);
nand U8997 (N_8997,N_8607,N_8739);
and U8998 (N_8998,N_8603,N_8712);
xor U8999 (N_8999,N_8699,N_8673);
nand U9000 (N_9000,N_8977,N_8876);
nor U9001 (N_9001,N_8873,N_8831);
and U9002 (N_9002,N_8902,N_8928);
xnor U9003 (N_9003,N_8999,N_8868);
nand U9004 (N_9004,N_8909,N_8900);
and U9005 (N_9005,N_8911,N_8810);
and U9006 (N_9006,N_8950,N_8838);
nand U9007 (N_9007,N_8983,N_8933);
or U9008 (N_9008,N_8981,N_8804);
or U9009 (N_9009,N_8997,N_8853);
and U9010 (N_9010,N_8944,N_8937);
xor U9011 (N_9011,N_8920,N_8998);
and U9012 (N_9012,N_8930,N_8863);
and U9013 (N_9013,N_8888,N_8896);
xor U9014 (N_9014,N_8827,N_8962);
xnor U9015 (N_9015,N_8839,N_8803);
or U9016 (N_9016,N_8992,N_8854);
and U9017 (N_9017,N_8882,N_8903);
xor U9018 (N_9018,N_8890,N_8952);
nor U9019 (N_9019,N_8814,N_8975);
or U9020 (N_9020,N_8982,N_8925);
and U9021 (N_9021,N_8832,N_8886);
and U9022 (N_9022,N_8855,N_8851);
and U9023 (N_9023,N_8941,N_8919);
or U9024 (N_9024,N_8864,N_8859);
xnor U9025 (N_9025,N_8893,N_8943);
and U9026 (N_9026,N_8942,N_8852);
and U9027 (N_9027,N_8857,N_8956);
or U9028 (N_9028,N_8967,N_8884);
nand U9029 (N_9029,N_8835,N_8908);
nor U9030 (N_9030,N_8829,N_8817);
nand U9031 (N_9031,N_8812,N_8843);
nand U9032 (N_9032,N_8971,N_8964);
and U9033 (N_9033,N_8877,N_8970);
nand U9034 (N_9034,N_8980,N_8809);
nor U9035 (N_9035,N_8819,N_8833);
nor U9036 (N_9036,N_8880,N_8871);
nand U9037 (N_9037,N_8824,N_8815);
and U9038 (N_9038,N_8988,N_8894);
and U9039 (N_9039,N_8901,N_8828);
nand U9040 (N_9040,N_8953,N_8986);
nand U9041 (N_9041,N_8846,N_8801);
or U9042 (N_9042,N_8913,N_8823);
and U9043 (N_9043,N_8825,N_8939);
or U9044 (N_9044,N_8934,N_8862);
xnor U9045 (N_9045,N_8979,N_8847);
nor U9046 (N_9046,N_8805,N_8822);
nor U9047 (N_9047,N_8938,N_8802);
xnor U9048 (N_9048,N_8905,N_8879);
xor U9049 (N_9049,N_8878,N_8875);
or U9050 (N_9050,N_8960,N_8949);
nor U9051 (N_9051,N_8921,N_8959);
xnor U9052 (N_9052,N_8948,N_8842);
and U9053 (N_9053,N_8897,N_8904);
xnor U9054 (N_9054,N_8808,N_8830);
nand U9055 (N_9055,N_8946,N_8963);
or U9056 (N_9056,N_8929,N_8926);
and U9057 (N_9057,N_8807,N_8881);
or U9058 (N_9058,N_8976,N_8906);
nor U9059 (N_9059,N_8968,N_8818);
nand U9060 (N_9060,N_8860,N_8936);
and U9061 (N_9061,N_8895,N_8958);
or U9062 (N_9062,N_8973,N_8821);
and U9063 (N_9063,N_8816,N_8883);
or U9064 (N_9064,N_8834,N_8995);
nand U9065 (N_9065,N_8907,N_8889);
nor U9066 (N_9066,N_8844,N_8806);
xnor U9067 (N_9067,N_8837,N_8915);
nor U9068 (N_9068,N_8984,N_8899);
or U9069 (N_9069,N_8826,N_8869);
xnor U9070 (N_9070,N_8945,N_8972);
xor U9071 (N_9071,N_8927,N_8951);
and U9072 (N_9072,N_8914,N_8813);
nand U9073 (N_9073,N_8856,N_8916);
or U9074 (N_9074,N_8891,N_8989);
or U9075 (N_9075,N_8800,N_8935);
nor U9076 (N_9076,N_8974,N_8924);
nand U9077 (N_9077,N_8932,N_8965);
xnor U9078 (N_9078,N_8820,N_8993);
nand U9079 (N_9079,N_8858,N_8892);
nor U9080 (N_9080,N_8850,N_8836);
and U9081 (N_9081,N_8861,N_8923);
xnor U9082 (N_9082,N_8845,N_8849);
and U9083 (N_9083,N_8872,N_8867);
nor U9084 (N_9084,N_8931,N_8996);
or U9085 (N_9085,N_8947,N_8848);
nor U9086 (N_9086,N_8887,N_8918);
or U9087 (N_9087,N_8840,N_8811);
xnor U9088 (N_9088,N_8898,N_8966);
xnor U9089 (N_9089,N_8922,N_8985);
xnor U9090 (N_9090,N_8990,N_8910);
nand U9091 (N_9091,N_8841,N_8987);
nor U9092 (N_9092,N_8957,N_8866);
and U9093 (N_9093,N_8885,N_8917);
and U9094 (N_9094,N_8969,N_8874);
nor U9095 (N_9095,N_8994,N_8940);
xor U9096 (N_9096,N_8865,N_8954);
nor U9097 (N_9097,N_8955,N_8978);
or U9098 (N_9098,N_8870,N_8912);
and U9099 (N_9099,N_8961,N_8991);
nand U9100 (N_9100,N_8807,N_8968);
nand U9101 (N_9101,N_8953,N_8878);
and U9102 (N_9102,N_8868,N_8867);
or U9103 (N_9103,N_8929,N_8978);
xnor U9104 (N_9104,N_8924,N_8944);
and U9105 (N_9105,N_8962,N_8980);
xnor U9106 (N_9106,N_8875,N_8833);
xnor U9107 (N_9107,N_8852,N_8802);
xor U9108 (N_9108,N_8953,N_8902);
and U9109 (N_9109,N_8815,N_8954);
or U9110 (N_9110,N_8812,N_8922);
and U9111 (N_9111,N_8909,N_8837);
xnor U9112 (N_9112,N_8864,N_8959);
nor U9113 (N_9113,N_8895,N_8944);
and U9114 (N_9114,N_8887,N_8871);
xor U9115 (N_9115,N_8897,N_8929);
nand U9116 (N_9116,N_8874,N_8831);
xor U9117 (N_9117,N_8888,N_8940);
and U9118 (N_9118,N_8863,N_8957);
xor U9119 (N_9119,N_8919,N_8885);
xor U9120 (N_9120,N_8844,N_8834);
nor U9121 (N_9121,N_8996,N_8861);
nor U9122 (N_9122,N_8975,N_8904);
and U9123 (N_9123,N_8900,N_8904);
nand U9124 (N_9124,N_8830,N_8901);
xor U9125 (N_9125,N_8870,N_8805);
or U9126 (N_9126,N_8842,N_8879);
nand U9127 (N_9127,N_8981,N_8873);
and U9128 (N_9128,N_8994,N_8972);
nand U9129 (N_9129,N_8988,N_8842);
nor U9130 (N_9130,N_8874,N_8959);
xor U9131 (N_9131,N_8894,N_8824);
xor U9132 (N_9132,N_8866,N_8923);
nor U9133 (N_9133,N_8807,N_8805);
or U9134 (N_9134,N_8910,N_8955);
or U9135 (N_9135,N_8965,N_8987);
nand U9136 (N_9136,N_8884,N_8979);
nand U9137 (N_9137,N_8882,N_8825);
xor U9138 (N_9138,N_8867,N_8978);
nand U9139 (N_9139,N_8918,N_8969);
nand U9140 (N_9140,N_8889,N_8955);
nor U9141 (N_9141,N_8878,N_8810);
or U9142 (N_9142,N_8820,N_8918);
nor U9143 (N_9143,N_8948,N_8981);
nand U9144 (N_9144,N_8997,N_8912);
nand U9145 (N_9145,N_8937,N_8995);
nand U9146 (N_9146,N_8811,N_8955);
or U9147 (N_9147,N_8958,N_8843);
nand U9148 (N_9148,N_8815,N_8942);
or U9149 (N_9149,N_8920,N_8874);
xor U9150 (N_9150,N_8964,N_8816);
nor U9151 (N_9151,N_8817,N_8959);
nor U9152 (N_9152,N_8978,N_8962);
and U9153 (N_9153,N_8841,N_8904);
xor U9154 (N_9154,N_8923,N_8989);
nor U9155 (N_9155,N_8841,N_8813);
and U9156 (N_9156,N_8984,N_8810);
nand U9157 (N_9157,N_8910,N_8856);
nor U9158 (N_9158,N_8989,N_8841);
and U9159 (N_9159,N_8847,N_8828);
nand U9160 (N_9160,N_8985,N_8807);
xnor U9161 (N_9161,N_8899,N_8873);
and U9162 (N_9162,N_8915,N_8946);
and U9163 (N_9163,N_8832,N_8978);
and U9164 (N_9164,N_8966,N_8857);
xnor U9165 (N_9165,N_8857,N_8987);
or U9166 (N_9166,N_8874,N_8972);
nor U9167 (N_9167,N_8925,N_8913);
and U9168 (N_9168,N_8835,N_8930);
xnor U9169 (N_9169,N_8865,N_8874);
nor U9170 (N_9170,N_8870,N_8919);
xor U9171 (N_9171,N_8917,N_8875);
nor U9172 (N_9172,N_8993,N_8931);
and U9173 (N_9173,N_8914,N_8883);
nor U9174 (N_9174,N_8924,N_8828);
nand U9175 (N_9175,N_8858,N_8855);
xnor U9176 (N_9176,N_8916,N_8906);
xor U9177 (N_9177,N_8888,N_8827);
nor U9178 (N_9178,N_8892,N_8921);
nand U9179 (N_9179,N_8829,N_8976);
and U9180 (N_9180,N_8887,N_8931);
xor U9181 (N_9181,N_8897,N_8848);
nand U9182 (N_9182,N_8866,N_8906);
and U9183 (N_9183,N_8858,N_8905);
xnor U9184 (N_9184,N_8844,N_8965);
or U9185 (N_9185,N_8853,N_8802);
xnor U9186 (N_9186,N_8823,N_8951);
and U9187 (N_9187,N_8996,N_8969);
or U9188 (N_9188,N_8837,N_8912);
or U9189 (N_9189,N_8847,N_8999);
nor U9190 (N_9190,N_8803,N_8975);
or U9191 (N_9191,N_8909,N_8901);
and U9192 (N_9192,N_8810,N_8821);
xor U9193 (N_9193,N_8802,N_8978);
nand U9194 (N_9194,N_8955,N_8954);
nand U9195 (N_9195,N_8827,N_8996);
nor U9196 (N_9196,N_8847,N_8919);
xnor U9197 (N_9197,N_8897,N_8846);
nor U9198 (N_9198,N_8907,N_8984);
nor U9199 (N_9199,N_8824,N_8874);
nand U9200 (N_9200,N_9019,N_9096);
nand U9201 (N_9201,N_9146,N_9100);
nand U9202 (N_9202,N_9193,N_9067);
or U9203 (N_9203,N_9001,N_9057);
nor U9204 (N_9204,N_9060,N_9179);
or U9205 (N_9205,N_9186,N_9133);
and U9206 (N_9206,N_9029,N_9199);
or U9207 (N_9207,N_9184,N_9104);
nand U9208 (N_9208,N_9031,N_9024);
nor U9209 (N_9209,N_9128,N_9055);
or U9210 (N_9210,N_9190,N_9041);
nor U9211 (N_9211,N_9023,N_9020);
nand U9212 (N_9212,N_9191,N_9078);
or U9213 (N_9213,N_9045,N_9088);
nor U9214 (N_9214,N_9103,N_9097);
nor U9215 (N_9215,N_9108,N_9195);
or U9216 (N_9216,N_9125,N_9132);
and U9217 (N_9217,N_9053,N_9140);
nor U9218 (N_9218,N_9083,N_9012);
nor U9219 (N_9219,N_9052,N_9049);
nand U9220 (N_9220,N_9076,N_9105);
xor U9221 (N_9221,N_9093,N_9173);
or U9222 (N_9222,N_9089,N_9032);
and U9223 (N_9223,N_9009,N_9066);
and U9224 (N_9224,N_9110,N_9004);
nor U9225 (N_9225,N_9056,N_9123);
nor U9226 (N_9226,N_9111,N_9037);
or U9227 (N_9227,N_9065,N_9143);
nand U9228 (N_9228,N_9022,N_9091);
nand U9229 (N_9229,N_9086,N_9137);
and U9230 (N_9230,N_9182,N_9028);
or U9231 (N_9231,N_9003,N_9030);
or U9232 (N_9232,N_9051,N_9021);
or U9233 (N_9233,N_9187,N_9025);
nor U9234 (N_9234,N_9155,N_9099);
nor U9235 (N_9235,N_9172,N_9135);
xnor U9236 (N_9236,N_9177,N_9095);
and U9237 (N_9237,N_9149,N_9035);
xor U9238 (N_9238,N_9157,N_9043);
nor U9239 (N_9239,N_9081,N_9113);
nand U9240 (N_9240,N_9183,N_9080);
nand U9241 (N_9241,N_9114,N_9008);
or U9242 (N_9242,N_9082,N_9117);
nand U9243 (N_9243,N_9197,N_9002);
and U9244 (N_9244,N_9013,N_9185);
xnor U9245 (N_9245,N_9171,N_9121);
and U9246 (N_9246,N_9141,N_9107);
nor U9247 (N_9247,N_9126,N_9077);
and U9248 (N_9248,N_9014,N_9042);
xnor U9249 (N_9249,N_9015,N_9150);
nand U9250 (N_9250,N_9094,N_9112);
xnor U9251 (N_9251,N_9196,N_9147);
and U9252 (N_9252,N_9011,N_9127);
nand U9253 (N_9253,N_9174,N_9169);
nor U9254 (N_9254,N_9178,N_9189);
or U9255 (N_9255,N_9109,N_9124);
nand U9256 (N_9256,N_9070,N_9175);
nand U9257 (N_9257,N_9050,N_9116);
nand U9258 (N_9258,N_9101,N_9079);
nor U9259 (N_9259,N_9153,N_9163);
or U9260 (N_9260,N_9068,N_9168);
xor U9261 (N_9261,N_9069,N_9161);
nand U9262 (N_9262,N_9154,N_9162);
or U9263 (N_9263,N_9152,N_9087);
xnor U9264 (N_9264,N_9194,N_9142);
or U9265 (N_9265,N_9164,N_9148);
and U9266 (N_9266,N_9131,N_9038);
and U9267 (N_9267,N_9016,N_9044);
nand U9268 (N_9268,N_9170,N_9134);
nand U9269 (N_9269,N_9075,N_9064);
nand U9270 (N_9270,N_9129,N_9046);
xnor U9271 (N_9271,N_9092,N_9145);
nand U9272 (N_9272,N_9159,N_9062);
xor U9273 (N_9273,N_9005,N_9118);
xor U9274 (N_9274,N_9084,N_9130);
nor U9275 (N_9275,N_9072,N_9156);
nor U9276 (N_9276,N_9119,N_9166);
xor U9277 (N_9277,N_9176,N_9027);
and U9278 (N_9278,N_9017,N_9054);
and U9279 (N_9279,N_9158,N_9048);
xor U9280 (N_9280,N_9036,N_9165);
xnor U9281 (N_9281,N_9047,N_9139);
nor U9282 (N_9282,N_9120,N_9144);
or U9283 (N_9283,N_9006,N_9063);
nor U9284 (N_9284,N_9007,N_9018);
and U9285 (N_9285,N_9098,N_9026);
nor U9286 (N_9286,N_9192,N_9040);
or U9287 (N_9287,N_9039,N_9160);
xnor U9288 (N_9288,N_9102,N_9034);
and U9289 (N_9289,N_9151,N_9115);
or U9290 (N_9290,N_9033,N_9074);
and U9291 (N_9291,N_9090,N_9106);
and U9292 (N_9292,N_9073,N_9188);
nand U9293 (N_9293,N_9180,N_9138);
nand U9294 (N_9294,N_9058,N_9122);
or U9295 (N_9295,N_9198,N_9059);
or U9296 (N_9296,N_9181,N_9085);
and U9297 (N_9297,N_9071,N_9136);
or U9298 (N_9298,N_9167,N_9000);
or U9299 (N_9299,N_9061,N_9010);
xor U9300 (N_9300,N_9083,N_9107);
nand U9301 (N_9301,N_9057,N_9005);
and U9302 (N_9302,N_9195,N_9155);
nor U9303 (N_9303,N_9007,N_9026);
nor U9304 (N_9304,N_9080,N_9103);
xor U9305 (N_9305,N_9190,N_9104);
or U9306 (N_9306,N_9155,N_9017);
nor U9307 (N_9307,N_9088,N_9060);
and U9308 (N_9308,N_9102,N_9107);
xnor U9309 (N_9309,N_9072,N_9044);
nand U9310 (N_9310,N_9049,N_9082);
xor U9311 (N_9311,N_9042,N_9169);
xor U9312 (N_9312,N_9003,N_9087);
nor U9313 (N_9313,N_9116,N_9158);
xor U9314 (N_9314,N_9167,N_9037);
nand U9315 (N_9315,N_9005,N_9081);
or U9316 (N_9316,N_9145,N_9072);
or U9317 (N_9317,N_9016,N_9092);
xnor U9318 (N_9318,N_9113,N_9046);
and U9319 (N_9319,N_9102,N_9113);
or U9320 (N_9320,N_9088,N_9008);
nor U9321 (N_9321,N_9162,N_9047);
or U9322 (N_9322,N_9059,N_9084);
and U9323 (N_9323,N_9055,N_9190);
nand U9324 (N_9324,N_9039,N_9101);
and U9325 (N_9325,N_9107,N_9137);
and U9326 (N_9326,N_9199,N_9045);
xor U9327 (N_9327,N_9142,N_9044);
xnor U9328 (N_9328,N_9158,N_9025);
nor U9329 (N_9329,N_9157,N_9054);
or U9330 (N_9330,N_9027,N_9191);
nor U9331 (N_9331,N_9121,N_9132);
and U9332 (N_9332,N_9163,N_9167);
or U9333 (N_9333,N_9059,N_9193);
nand U9334 (N_9334,N_9002,N_9070);
and U9335 (N_9335,N_9169,N_9022);
or U9336 (N_9336,N_9176,N_9088);
xnor U9337 (N_9337,N_9166,N_9017);
xnor U9338 (N_9338,N_9086,N_9072);
nor U9339 (N_9339,N_9023,N_9129);
nor U9340 (N_9340,N_9104,N_9019);
nor U9341 (N_9341,N_9072,N_9032);
or U9342 (N_9342,N_9177,N_9044);
nor U9343 (N_9343,N_9121,N_9015);
nor U9344 (N_9344,N_9117,N_9142);
nand U9345 (N_9345,N_9130,N_9147);
xnor U9346 (N_9346,N_9040,N_9025);
xor U9347 (N_9347,N_9009,N_9125);
and U9348 (N_9348,N_9082,N_9059);
or U9349 (N_9349,N_9048,N_9179);
nor U9350 (N_9350,N_9195,N_9175);
nand U9351 (N_9351,N_9009,N_9022);
nor U9352 (N_9352,N_9138,N_9039);
and U9353 (N_9353,N_9157,N_9067);
nor U9354 (N_9354,N_9073,N_9036);
and U9355 (N_9355,N_9033,N_9056);
nor U9356 (N_9356,N_9087,N_9195);
nand U9357 (N_9357,N_9120,N_9104);
nand U9358 (N_9358,N_9116,N_9041);
nor U9359 (N_9359,N_9194,N_9054);
or U9360 (N_9360,N_9043,N_9174);
xor U9361 (N_9361,N_9066,N_9156);
nand U9362 (N_9362,N_9030,N_9177);
xnor U9363 (N_9363,N_9124,N_9069);
or U9364 (N_9364,N_9185,N_9026);
or U9365 (N_9365,N_9053,N_9199);
xor U9366 (N_9366,N_9055,N_9139);
nor U9367 (N_9367,N_9067,N_9044);
or U9368 (N_9368,N_9070,N_9061);
or U9369 (N_9369,N_9108,N_9006);
xor U9370 (N_9370,N_9092,N_9108);
or U9371 (N_9371,N_9040,N_9126);
nand U9372 (N_9372,N_9058,N_9138);
nor U9373 (N_9373,N_9117,N_9194);
nor U9374 (N_9374,N_9167,N_9002);
or U9375 (N_9375,N_9089,N_9071);
xnor U9376 (N_9376,N_9117,N_9163);
xor U9377 (N_9377,N_9161,N_9003);
and U9378 (N_9378,N_9069,N_9048);
and U9379 (N_9379,N_9196,N_9069);
or U9380 (N_9380,N_9198,N_9001);
nand U9381 (N_9381,N_9197,N_9043);
nor U9382 (N_9382,N_9103,N_9160);
and U9383 (N_9383,N_9045,N_9188);
or U9384 (N_9384,N_9160,N_9130);
nor U9385 (N_9385,N_9094,N_9138);
or U9386 (N_9386,N_9123,N_9192);
nand U9387 (N_9387,N_9094,N_9054);
nor U9388 (N_9388,N_9015,N_9165);
nor U9389 (N_9389,N_9158,N_9184);
xnor U9390 (N_9390,N_9175,N_9058);
nor U9391 (N_9391,N_9076,N_9107);
nor U9392 (N_9392,N_9016,N_9109);
nor U9393 (N_9393,N_9068,N_9125);
nand U9394 (N_9394,N_9008,N_9078);
or U9395 (N_9395,N_9102,N_9125);
and U9396 (N_9396,N_9098,N_9080);
xor U9397 (N_9397,N_9011,N_9030);
or U9398 (N_9398,N_9050,N_9082);
and U9399 (N_9399,N_9054,N_9143);
nand U9400 (N_9400,N_9367,N_9324);
nor U9401 (N_9401,N_9313,N_9307);
nor U9402 (N_9402,N_9373,N_9230);
xnor U9403 (N_9403,N_9298,N_9305);
nor U9404 (N_9404,N_9365,N_9258);
or U9405 (N_9405,N_9392,N_9369);
nand U9406 (N_9406,N_9238,N_9317);
or U9407 (N_9407,N_9363,N_9287);
nor U9408 (N_9408,N_9306,N_9393);
xnor U9409 (N_9409,N_9242,N_9286);
and U9410 (N_9410,N_9217,N_9358);
nand U9411 (N_9411,N_9327,N_9297);
or U9412 (N_9412,N_9219,N_9288);
xnor U9413 (N_9413,N_9248,N_9247);
or U9414 (N_9414,N_9376,N_9389);
nor U9415 (N_9415,N_9280,N_9278);
and U9416 (N_9416,N_9385,N_9353);
xnor U9417 (N_9417,N_9379,N_9296);
or U9418 (N_9418,N_9341,N_9319);
nor U9419 (N_9419,N_9315,N_9396);
xor U9420 (N_9420,N_9293,N_9241);
and U9421 (N_9421,N_9218,N_9206);
xnor U9422 (N_9422,N_9209,N_9348);
and U9423 (N_9423,N_9268,N_9277);
nand U9424 (N_9424,N_9370,N_9337);
or U9425 (N_9425,N_9368,N_9282);
nand U9426 (N_9426,N_9361,N_9321);
nand U9427 (N_9427,N_9235,N_9338);
nor U9428 (N_9428,N_9330,N_9260);
and U9429 (N_9429,N_9343,N_9384);
xnor U9430 (N_9430,N_9256,N_9249);
and U9431 (N_9431,N_9284,N_9381);
nand U9432 (N_9432,N_9387,N_9204);
nand U9433 (N_9433,N_9325,N_9394);
xnor U9434 (N_9434,N_9203,N_9303);
and U9435 (N_9435,N_9228,N_9225);
or U9436 (N_9436,N_9372,N_9354);
nor U9437 (N_9437,N_9328,N_9299);
nand U9438 (N_9438,N_9335,N_9388);
nor U9439 (N_9439,N_9243,N_9391);
and U9440 (N_9440,N_9320,N_9221);
or U9441 (N_9441,N_9269,N_9331);
nand U9442 (N_9442,N_9326,N_9347);
xor U9443 (N_9443,N_9255,N_9336);
nor U9444 (N_9444,N_9233,N_9302);
and U9445 (N_9445,N_9213,N_9253);
nor U9446 (N_9446,N_9378,N_9252);
and U9447 (N_9447,N_9291,N_9245);
nand U9448 (N_9448,N_9371,N_9237);
nand U9449 (N_9449,N_9257,N_9356);
nand U9450 (N_9450,N_9267,N_9359);
nand U9451 (N_9451,N_9386,N_9272);
and U9452 (N_9452,N_9236,N_9333);
nor U9453 (N_9453,N_9240,N_9262);
nand U9454 (N_9454,N_9311,N_9322);
xor U9455 (N_9455,N_9263,N_9364);
xnor U9456 (N_9456,N_9366,N_9344);
and U9457 (N_9457,N_9275,N_9292);
xnor U9458 (N_9458,N_9211,N_9300);
nor U9459 (N_9459,N_9232,N_9397);
and U9460 (N_9460,N_9222,N_9316);
or U9461 (N_9461,N_9281,N_9362);
nand U9462 (N_9462,N_9289,N_9398);
or U9463 (N_9463,N_9274,N_9360);
nor U9464 (N_9464,N_9351,N_9227);
and U9465 (N_9465,N_9205,N_9377);
and U9466 (N_9466,N_9314,N_9285);
xnor U9467 (N_9467,N_9208,N_9224);
or U9468 (N_9468,N_9309,N_9216);
and U9469 (N_9469,N_9261,N_9279);
nand U9470 (N_9470,N_9395,N_9270);
and U9471 (N_9471,N_9264,N_9339);
nand U9472 (N_9472,N_9357,N_9271);
or U9473 (N_9473,N_9244,N_9312);
xnor U9474 (N_9474,N_9380,N_9352);
nand U9475 (N_9475,N_9301,N_9201);
or U9476 (N_9476,N_9202,N_9246);
or U9477 (N_9477,N_9346,N_9295);
or U9478 (N_9478,N_9374,N_9283);
and U9479 (N_9479,N_9345,N_9200);
and U9480 (N_9480,N_9323,N_9375);
or U9481 (N_9481,N_9234,N_9332);
nor U9482 (N_9482,N_9214,N_9308);
xor U9483 (N_9483,N_9290,N_9254);
and U9484 (N_9484,N_9355,N_9220);
nand U9485 (N_9485,N_9399,N_9350);
nand U9486 (N_9486,N_9304,N_9212);
xor U9487 (N_9487,N_9340,N_9231);
nand U9488 (N_9488,N_9226,N_9390);
and U9489 (N_9489,N_9273,N_9342);
or U9490 (N_9490,N_9250,N_9251);
nor U9491 (N_9491,N_9259,N_9318);
and U9492 (N_9492,N_9329,N_9229);
and U9493 (N_9493,N_9383,N_9207);
nand U9494 (N_9494,N_9265,N_9294);
xor U9495 (N_9495,N_9310,N_9215);
xnor U9496 (N_9496,N_9266,N_9382);
nor U9497 (N_9497,N_9349,N_9276);
or U9498 (N_9498,N_9334,N_9223);
nand U9499 (N_9499,N_9239,N_9210);
nand U9500 (N_9500,N_9208,N_9341);
and U9501 (N_9501,N_9299,N_9292);
nor U9502 (N_9502,N_9318,N_9308);
xor U9503 (N_9503,N_9205,N_9321);
nand U9504 (N_9504,N_9271,N_9367);
xor U9505 (N_9505,N_9203,N_9258);
or U9506 (N_9506,N_9345,N_9375);
nand U9507 (N_9507,N_9322,N_9273);
nand U9508 (N_9508,N_9396,N_9304);
xnor U9509 (N_9509,N_9221,N_9391);
nor U9510 (N_9510,N_9288,N_9324);
nand U9511 (N_9511,N_9219,N_9222);
nor U9512 (N_9512,N_9273,N_9357);
nand U9513 (N_9513,N_9378,N_9332);
or U9514 (N_9514,N_9395,N_9340);
xor U9515 (N_9515,N_9333,N_9230);
and U9516 (N_9516,N_9368,N_9379);
nor U9517 (N_9517,N_9389,N_9225);
xor U9518 (N_9518,N_9321,N_9391);
and U9519 (N_9519,N_9392,N_9252);
or U9520 (N_9520,N_9367,N_9374);
and U9521 (N_9521,N_9234,N_9372);
nand U9522 (N_9522,N_9338,N_9391);
nor U9523 (N_9523,N_9223,N_9303);
or U9524 (N_9524,N_9337,N_9361);
xor U9525 (N_9525,N_9284,N_9237);
nor U9526 (N_9526,N_9260,N_9371);
nand U9527 (N_9527,N_9261,N_9288);
nand U9528 (N_9528,N_9302,N_9360);
xor U9529 (N_9529,N_9393,N_9240);
or U9530 (N_9530,N_9320,N_9276);
nand U9531 (N_9531,N_9300,N_9282);
nor U9532 (N_9532,N_9210,N_9382);
xor U9533 (N_9533,N_9234,N_9305);
nand U9534 (N_9534,N_9353,N_9382);
xnor U9535 (N_9535,N_9365,N_9288);
nand U9536 (N_9536,N_9211,N_9304);
xor U9537 (N_9537,N_9224,N_9363);
and U9538 (N_9538,N_9276,N_9262);
or U9539 (N_9539,N_9279,N_9374);
xnor U9540 (N_9540,N_9375,N_9231);
or U9541 (N_9541,N_9271,N_9324);
nand U9542 (N_9542,N_9221,N_9214);
and U9543 (N_9543,N_9204,N_9367);
or U9544 (N_9544,N_9328,N_9216);
xnor U9545 (N_9545,N_9354,N_9385);
nand U9546 (N_9546,N_9214,N_9316);
and U9547 (N_9547,N_9304,N_9236);
or U9548 (N_9548,N_9251,N_9287);
and U9549 (N_9549,N_9237,N_9396);
xnor U9550 (N_9550,N_9235,N_9217);
nor U9551 (N_9551,N_9349,N_9269);
nor U9552 (N_9552,N_9295,N_9217);
nand U9553 (N_9553,N_9246,N_9368);
or U9554 (N_9554,N_9361,N_9375);
or U9555 (N_9555,N_9211,N_9219);
nor U9556 (N_9556,N_9314,N_9251);
or U9557 (N_9557,N_9307,N_9382);
nand U9558 (N_9558,N_9241,N_9284);
or U9559 (N_9559,N_9229,N_9351);
xor U9560 (N_9560,N_9262,N_9291);
or U9561 (N_9561,N_9382,N_9321);
nand U9562 (N_9562,N_9319,N_9253);
xnor U9563 (N_9563,N_9377,N_9321);
xor U9564 (N_9564,N_9291,N_9348);
and U9565 (N_9565,N_9288,N_9330);
nor U9566 (N_9566,N_9284,N_9319);
or U9567 (N_9567,N_9254,N_9300);
nand U9568 (N_9568,N_9243,N_9213);
nand U9569 (N_9569,N_9303,N_9215);
nor U9570 (N_9570,N_9231,N_9345);
xor U9571 (N_9571,N_9385,N_9390);
nor U9572 (N_9572,N_9387,N_9243);
nor U9573 (N_9573,N_9368,N_9217);
nand U9574 (N_9574,N_9229,N_9235);
and U9575 (N_9575,N_9386,N_9296);
nand U9576 (N_9576,N_9286,N_9240);
or U9577 (N_9577,N_9209,N_9267);
nand U9578 (N_9578,N_9242,N_9393);
and U9579 (N_9579,N_9238,N_9375);
and U9580 (N_9580,N_9205,N_9360);
nor U9581 (N_9581,N_9368,N_9395);
or U9582 (N_9582,N_9306,N_9289);
xor U9583 (N_9583,N_9265,N_9233);
and U9584 (N_9584,N_9346,N_9238);
nor U9585 (N_9585,N_9270,N_9262);
nand U9586 (N_9586,N_9321,N_9317);
nand U9587 (N_9587,N_9282,N_9366);
xor U9588 (N_9588,N_9353,N_9309);
xor U9589 (N_9589,N_9384,N_9270);
nor U9590 (N_9590,N_9250,N_9278);
and U9591 (N_9591,N_9226,N_9395);
nor U9592 (N_9592,N_9255,N_9263);
nor U9593 (N_9593,N_9364,N_9365);
nand U9594 (N_9594,N_9376,N_9314);
nand U9595 (N_9595,N_9304,N_9397);
and U9596 (N_9596,N_9359,N_9324);
nor U9597 (N_9597,N_9272,N_9223);
nor U9598 (N_9598,N_9395,N_9205);
nor U9599 (N_9599,N_9209,N_9355);
xor U9600 (N_9600,N_9535,N_9485);
nand U9601 (N_9601,N_9484,N_9575);
and U9602 (N_9602,N_9578,N_9415);
nand U9603 (N_9603,N_9489,N_9534);
nor U9604 (N_9604,N_9551,N_9445);
nor U9605 (N_9605,N_9585,N_9492);
and U9606 (N_9606,N_9560,N_9542);
nor U9607 (N_9607,N_9514,N_9550);
or U9608 (N_9608,N_9593,N_9476);
or U9609 (N_9609,N_9523,N_9521);
nand U9610 (N_9610,N_9482,N_9494);
nor U9611 (N_9611,N_9413,N_9419);
nand U9612 (N_9612,N_9519,N_9406);
nor U9613 (N_9613,N_9503,N_9509);
and U9614 (N_9614,N_9487,N_9598);
nand U9615 (N_9615,N_9458,N_9580);
or U9616 (N_9616,N_9414,N_9486);
nand U9617 (N_9617,N_9531,N_9530);
nor U9618 (N_9618,N_9401,N_9451);
and U9619 (N_9619,N_9402,N_9595);
nor U9620 (N_9620,N_9405,N_9525);
and U9621 (N_9621,N_9529,N_9471);
or U9622 (N_9622,N_9495,N_9583);
nor U9623 (N_9623,N_9570,N_9554);
nor U9624 (N_9624,N_9568,N_9411);
xnor U9625 (N_9625,N_9421,N_9460);
nor U9626 (N_9626,N_9581,N_9464);
or U9627 (N_9627,N_9586,N_9475);
or U9628 (N_9628,N_9549,N_9527);
xor U9629 (N_9629,N_9558,N_9592);
nor U9630 (N_9630,N_9505,N_9555);
nor U9631 (N_9631,N_9439,N_9466);
or U9632 (N_9632,N_9434,N_9407);
and U9633 (N_9633,N_9518,N_9517);
nand U9634 (N_9634,N_9540,N_9418);
nor U9635 (N_9635,N_9500,N_9524);
nor U9636 (N_9636,N_9499,N_9467);
nand U9637 (N_9637,N_9403,N_9428);
nor U9638 (N_9638,N_9491,N_9579);
nor U9639 (N_9639,N_9448,N_9459);
nor U9640 (N_9640,N_9571,N_9501);
nor U9641 (N_9641,N_9506,N_9446);
and U9642 (N_9642,N_9450,N_9511);
nand U9643 (N_9643,N_9599,N_9597);
xnor U9644 (N_9644,N_9573,N_9420);
xnor U9645 (N_9645,N_9569,N_9502);
or U9646 (N_9646,N_9539,N_9588);
xor U9647 (N_9647,N_9493,N_9490);
xor U9648 (N_9648,N_9564,N_9438);
nand U9649 (N_9649,N_9456,N_9463);
or U9650 (N_9650,N_9426,N_9548);
and U9651 (N_9651,N_9589,N_9454);
and U9652 (N_9652,N_9477,N_9455);
nand U9653 (N_9653,N_9498,N_9474);
nand U9654 (N_9654,N_9587,N_9512);
or U9655 (N_9655,N_9436,N_9422);
nand U9656 (N_9656,N_9515,N_9537);
nor U9657 (N_9657,N_9430,N_9468);
nor U9658 (N_9658,N_9478,N_9431);
and U9659 (N_9659,N_9507,N_9566);
nand U9660 (N_9660,N_9546,N_9473);
and U9661 (N_9661,N_9556,N_9526);
and U9662 (N_9662,N_9513,N_9433);
or U9663 (N_9663,N_9516,N_9449);
nor U9664 (N_9664,N_9504,N_9469);
nand U9665 (N_9665,N_9409,N_9553);
xnor U9666 (N_9666,N_9404,N_9590);
or U9667 (N_9667,N_9417,N_9472);
nand U9668 (N_9668,N_9481,N_9536);
nor U9669 (N_9669,N_9577,N_9557);
and U9670 (N_9670,N_9510,N_9508);
and U9671 (N_9671,N_9412,N_9522);
nor U9672 (N_9672,N_9462,N_9432);
nor U9673 (N_9673,N_9425,N_9559);
nor U9674 (N_9674,N_9447,N_9457);
and U9675 (N_9675,N_9483,N_9545);
or U9676 (N_9676,N_9572,N_9465);
or U9677 (N_9677,N_9429,N_9461);
nor U9678 (N_9678,N_9441,N_9538);
or U9679 (N_9679,N_9528,N_9565);
or U9680 (N_9680,N_9574,N_9533);
xor U9681 (N_9681,N_9400,N_9443);
nand U9682 (N_9682,N_9563,N_9543);
nand U9683 (N_9683,N_9453,N_9591);
xor U9684 (N_9684,N_9532,N_9427);
nor U9685 (N_9685,N_9435,N_9423);
xnor U9686 (N_9686,N_9408,N_9541);
or U9687 (N_9687,N_9496,N_9488);
nor U9688 (N_9688,N_9424,N_9562);
nand U9689 (N_9689,N_9582,N_9497);
nor U9690 (N_9690,N_9547,N_9596);
or U9691 (N_9691,N_9480,N_9452);
nand U9692 (N_9692,N_9416,N_9594);
xnor U9693 (N_9693,N_9544,N_9479);
xor U9694 (N_9694,N_9567,N_9437);
nor U9695 (N_9695,N_9440,N_9442);
or U9696 (N_9696,N_9561,N_9552);
or U9697 (N_9697,N_9576,N_9520);
nand U9698 (N_9698,N_9410,N_9444);
and U9699 (N_9699,N_9584,N_9470);
and U9700 (N_9700,N_9481,N_9404);
nor U9701 (N_9701,N_9473,N_9448);
and U9702 (N_9702,N_9491,N_9498);
and U9703 (N_9703,N_9442,N_9526);
or U9704 (N_9704,N_9564,N_9453);
and U9705 (N_9705,N_9421,N_9559);
nand U9706 (N_9706,N_9561,N_9520);
or U9707 (N_9707,N_9479,N_9526);
nor U9708 (N_9708,N_9551,N_9537);
and U9709 (N_9709,N_9461,N_9404);
xnor U9710 (N_9710,N_9538,N_9408);
and U9711 (N_9711,N_9427,N_9422);
nand U9712 (N_9712,N_9447,N_9469);
nor U9713 (N_9713,N_9577,N_9564);
and U9714 (N_9714,N_9425,N_9584);
nor U9715 (N_9715,N_9536,N_9483);
nand U9716 (N_9716,N_9506,N_9420);
nor U9717 (N_9717,N_9573,N_9479);
nand U9718 (N_9718,N_9413,N_9578);
xnor U9719 (N_9719,N_9404,N_9579);
or U9720 (N_9720,N_9492,N_9440);
xnor U9721 (N_9721,N_9527,N_9461);
or U9722 (N_9722,N_9466,N_9572);
nor U9723 (N_9723,N_9484,N_9587);
nor U9724 (N_9724,N_9458,N_9523);
xnor U9725 (N_9725,N_9598,N_9472);
nand U9726 (N_9726,N_9478,N_9583);
nor U9727 (N_9727,N_9542,N_9530);
nor U9728 (N_9728,N_9522,N_9529);
or U9729 (N_9729,N_9592,N_9453);
and U9730 (N_9730,N_9500,N_9544);
nand U9731 (N_9731,N_9565,N_9446);
nor U9732 (N_9732,N_9458,N_9448);
nor U9733 (N_9733,N_9597,N_9466);
and U9734 (N_9734,N_9435,N_9458);
xor U9735 (N_9735,N_9527,N_9526);
or U9736 (N_9736,N_9444,N_9570);
or U9737 (N_9737,N_9471,N_9540);
nor U9738 (N_9738,N_9560,N_9577);
and U9739 (N_9739,N_9420,N_9429);
or U9740 (N_9740,N_9440,N_9576);
xnor U9741 (N_9741,N_9519,N_9479);
nor U9742 (N_9742,N_9506,N_9428);
nor U9743 (N_9743,N_9478,N_9539);
xor U9744 (N_9744,N_9478,N_9456);
nor U9745 (N_9745,N_9532,N_9598);
nand U9746 (N_9746,N_9524,N_9565);
nand U9747 (N_9747,N_9434,N_9454);
and U9748 (N_9748,N_9543,N_9437);
nor U9749 (N_9749,N_9425,N_9509);
or U9750 (N_9750,N_9448,N_9502);
nand U9751 (N_9751,N_9599,N_9424);
and U9752 (N_9752,N_9502,N_9535);
nor U9753 (N_9753,N_9599,N_9442);
and U9754 (N_9754,N_9564,N_9520);
nor U9755 (N_9755,N_9569,N_9522);
and U9756 (N_9756,N_9425,N_9547);
nor U9757 (N_9757,N_9592,N_9454);
xnor U9758 (N_9758,N_9494,N_9545);
or U9759 (N_9759,N_9405,N_9461);
xor U9760 (N_9760,N_9486,N_9409);
nor U9761 (N_9761,N_9532,N_9509);
nor U9762 (N_9762,N_9506,N_9411);
nand U9763 (N_9763,N_9521,N_9459);
nand U9764 (N_9764,N_9555,N_9532);
or U9765 (N_9765,N_9512,N_9542);
or U9766 (N_9766,N_9556,N_9485);
and U9767 (N_9767,N_9522,N_9566);
or U9768 (N_9768,N_9442,N_9555);
xor U9769 (N_9769,N_9438,N_9493);
and U9770 (N_9770,N_9485,N_9411);
and U9771 (N_9771,N_9422,N_9505);
nand U9772 (N_9772,N_9573,N_9538);
nand U9773 (N_9773,N_9586,N_9582);
or U9774 (N_9774,N_9506,N_9477);
nand U9775 (N_9775,N_9553,N_9538);
nor U9776 (N_9776,N_9580,N_9503);
xnor U9777 (N_9777,N_9541,N_9589);
and U9778 (N_9778,N_9574,N_9418);
nand U9779 (N_9779,N_9574,N_9445);
nor U9780 (N_9780,N_9585,N_9448);
nand U9781 (N_9781,N_9515,N_9592);
nor U9782 (N_9782,N_9582,N_9442);
nor U9783 (N_9783,N_9549,N_9537);
and U9784 (N_9784,N_9423,N_9490);
xor U9785 (N_9785,N_9516,N_9455);
nor U9786 (N_9786,N_9502,N_9577);
and U9787 (N_9787,N_9481,N_9465);
nand U9788 (N_9788,N_9572,N_9434);
xnor U9789 (N_9789,N_9550,N_9503);
xor U9790 (N_9790,N_9406,N_9573);
nand U9791 (N_9791,N_9546,N_9416);
nor U9792 (N_9792,N_9447,N_9596);
nor U9793 (N_9793,N_9425,N_9430);
and U9794 (N_9794,N_9422,N_9452);
or U9795 (N_9795,N_9521,N_9555);
nor U9796 (N_9796,N_9578,N_9512);
or U9797 (N_9797,N_9521,N_9412);
or U9798 (N_9798,N_9550,N_9421);
xnor U9799 (N_9799,N_9474,N_9496);
or U9800 (N_9800,N_9601,N_9715);
nor U9801 (N_9801,N_9734,N_9748);
or U9802 (N_9802,N_9611,N_9658);
nor U9803 (N_9803,N_9762,N_9775);
xor U9804 (N_9804,N_9758,N_9704);
or U9805 (N_9805,N_9696,N_9780);
or U9806 (N_9806,N_9759,N_9730);
xor U9807 (N_9807,N_9624,N_9673);
xor U9808 (N_9808,N_9798,N_9602);
and U9809 (N_9809,N_9683,N_9689);
xnor U9810 (N_9810,N_9785,N_9667);
xor U9811 (N_9811,N_9700,N_9697);
and U9812 (N_9812,N_9711,N_9732);
nor U9813 (N_9813,N_9681,N_9654);
nand U9814 (N_9814,N_9772,N_9774);
or U9815 (N_9815,N_9605,N_9603);
and U9816 (N_9816,N_9648,N_9692);
nor U9817 (N_9817,N_9642,N_9735);
and U9818 (N_9818,N_9770,N_9706);
and U9819 (N_9819,N_9606,N_9666);
nand U9820 (N_9820,N_9752,N_9663);
nor U9821 (N_9821,N_9795,N_9646);
or U9822 (N_9822,N_9686,N_9768);
nand U9823 (N_9823,N_9764,N_9794);
or U9824 (N_9824,N_9674,N_9699);
or U9825 (N_9825,N_9682,N_9719);
nand U9826 (N_9826,N_9729,N_9799);
and U9827 (N_9827,N_9655,N_9690);
or U9828 (N_9828,N_9652,N_9670);
xor U9829 (N_9829,N_9750,N_9688);
nor U9830 (N_9830,N_9766,N_9657);
or U9831 (N_9831,N_9684,N_9668);
nand U9832 (N_9832,N_9708,N_9733);
nor U9833 (N_9833,N_9713,N_9638);
xnor U9834 (N_9834,N_9662,N_9620);
nand U9835 (N_9835,N_9737,N_9728);
xnor U9836 (N_9836,N_9787,N_9789);
and U9837 (N_9837,N_9660,N_9761);
nor U9838 (N_9838,N_9676,N_9791);
xor U9839 (N_9839,N_9647,N_9619);
nand U9840 (N_9840,N_9705,N_9776);
or U9841 (N_9841,N_9773,N_9765);
or U9842 (N_9842,N_9779,N_9740);
and U9843 (N_9843,N_9747,N_9744);
and U9844 (N_9844,N_9678,N_9788);
xnor U9845 (N_9845,N_9625,N_9783);
xor U9846 (N_9846,N_9640,N_9604);
nor U9847 (N_9847,N_9616,N_9714);
nor U9848 (N_9848,N_9671,N_9639);
xnor U9849 (N_9849,N_9621,N_9736);
and U9850 (N_9850,N_9745,N_9693);
nand U9851 (N_9851,N_9661,N_9623);
or U9852 (N_9852,N_9635,N_9618);
and U9853 (N_9853,N_9701,N_9712);
and U9854 (N_9854,N_9755,N_9687);
nand U9855 (N_9855,N_9796,N_9790);
nor U9856 (N_9856,N_9792,N_9656);
nand U9857 (N_9857,N_9746,N_9626);
xnor U9858 (N_9858,N_9695,N_9716);
nand U9859 (N_9859,N_9782,N_9665);
nand U9860 (N_9860,N_9650,N_9757);
nand U9861 (N_9861,N_9617,N_9710);
and U9862 (N_9862,N_9629,N_9767);
or U9863 (N_9863,N_9723,N_9703);
xnor U9864 (N_9864,N_9784,N_9702);
or U9865 (N_9865,N_9727,N_9709);
nor U9866 (N_9866,N_9786,N_9609);
nor U9867 (N_9867,N_9627,N_9628);
nand U9868 (N_9868,N_9756,N_9610);
nor U9869 (N_9869,N_9653,N_9720);
nor U9870 (N_9870,N_9781,N_9637);
or U9871 (N_9871,N_9726,N_9614);
nand U9872 (N_9872,N_9641,N_9753);
or U9873 (N_9873,N_9622,N_9754);
nor U9874 (N_9874,N_9771,N_9718);
and U9875 (N_9875,N_9607,N_9724);
or U9876 (N_9876,N_9731,N_9707);
and U9877 (N_9877,N_9738,N_9721);
or U9878 (N_9878,N_9651,N_9778);
nor U9879 (N_9879,N_9634,N_9777);
xnor U9880 (N_9880,N_9725,N_9649);
or U9881 (N_9881,N_9760,N_9741);
and U9882 (N_9882,N_9633,N_9717);
or U9883 (N_9883,N_9680,N_9643);
xnor U9884 (N_9884,N_9630,N_9636);
nor U9885 (N_9885,N_9698,N_9675);
xnor U9886 (N_9886,N_9669,N_9608);
xnor U9887 (N_9887,N_9659,N_9797);
nand U9888 (N_9888,N_9632,N_9722);
nor U9889 (N_9889,N_9742,N_9685);
or U9890 (N_9890,N_9739,N_9615);
or U9891 (N_9891,N_9631,N_9644);
and U9892 (N_9892,N_9749,N_9793);
nor U9893 (N_9893,N_9743,N_9672);
xnor U9894 (N_9894,N_9664,N_9694);
nand U9895 (N_9895,N_9769,N_9613);
or U9896 (N_9896,N_9677,N_9679);
or U9897 (N_9897,N_9600,N_9691);
and U9898 (N_9898,N_9612,N_9763);
nand U9899 (N_9899,N_9645,N_9751);
nor U9900 (N_9900,N_9721,N_9697);
or U9901 (N_9901,N_9758,N_9654);
nor U9902 (N_9902,N_9611,N_9716);
xnor U9903 (N_9903,N_9740,N_9785);
and U9904 (N_9904,N_9644,N_9768);
nor U9905 (N_9905,N_9722,N_9624);
or U9906 (N_9906,N_9676,N_9751);
xor U9907 (N_9907,N_9668,N_9729);
and U9908 (N_9908,N_9640,N_9769);
and U9909 (N_9909,N_9608,N_9736);
nor U9910 (N_9910,N_9694,N_9730);
or U9911 (N_9911,N_9701,N_9612);
nand U9912 (N_9912,N_9702,N_9706);
xnor U9913 (N_9913,N_9792,N_9688);
nor U9914 (N_9914,N_9690,N_9685);
xnor U9915 (N_9915,N_9635,N_9705);
nor U9916 (N_9916,N_9742,N_9705);
nand U9917 (N_9917,N_9634,N_9734);
xor U9918 (N_9918,N_9723,N_9798);
and U9919 (N_9919,N_9702,N_9726);
xor U9920 (N_9920,N_9649,N_9774);
nand U9921 (N_9921,N_9693,N_9691);
or U9922 (N_9922,N_9770,N_9707);
or U9923 (N_9923,N_9755,N_9733);
xnor U9924 (N_9924,N_9756,N_9627);
xor U9925 (N_9925,N_9665,N_9623);
nand U9926 (N_9926,N_9660,N_9780);
nand U9927 (N_9927,N_9739,N_9631);
nand U9928 (N_9928,N_9735,N_9757);
xor U9929 (N_9929,N_9726,N_9624);
nand U9930 (N_9930,N_9641,N_9797);
nand U9931 (N_9931,N_9722,N_9681);
nand U9932 (N_9932,N_9618,N_9732);
nor U9933 (N_9933,N_9606,N_9676);
nand U9934 (N_9934,N_9654,N_9776);
and U9935 (N_9935,N_9754,N_9689);
or U9936 (N_9936,N_9695,N_9601);
nand U9937 (N_9937,N_9677,N_9659);
nand U9938 (N_9938,N_9617,N_9765);
and U9939 (N_9939,N_9721,N_9715);
xor U9940 (N_9940,N_9602,N_9687);
nor U9941 (N_9941,N_9667,N_9790);
and U9942 (N_9942,N_9795,N_9719);
xor U9943 (N_9943,N_9620,N_9784);
nand U9944 (N_9944,N_9670,N_9603);
or U9945 (N_9945,N_9658,N_9652);
nand U9946 (N_9946,N_9613,N_9659);
nor U9947 (N_9947,N_9782,N_9697);
xnor U9948 (N_9948,N_9735,N_9745);
nand U9949 (N_9949,N_9778,N_9666);
or U9950 (N_9950,N_9649,N_9689);
nand U9951 (N_9951,N_9755,N_9658);
nand U9952 (N_9952,N_9601,N_9784);
or U9953 (N_9953,N_9684,N_9714);
nand U9954 (N_9954,N_9783,N_9791);
nand U9955 (N_9955,N_9768,N_9790);
nor U9956 (N_9956,N_9691,N_9617);
xor U9957 (N_9957,N_9607,N_9615);
nor U9958 (N_9958,N_9794,N_9627);
or U9959 (N_9959,N_9667,N_9616);
nand U9960 (N_9960,N_9617,N_9656);
xnor U9961 (N_9961,N_9682,N_9744);
nand U9962 (N_9962,N_9786,N_9716);
nand U9963 (N_9963,N_9750,N_9731);
nor U9964 (N_9964,N_9780,N_9611);
nand U9965 (N_9965,N_9798,N_9788);
and U9966 (N_9966,N_9741,N_9774);
nand U9967 (N_9967,N_9698,N_9705);
and U9968 (N_9968,N_9729,N_9779);
or U9969 (N_9969,N_9638,N_9660);
nor U9970 (N_9970,N_9623,N_9736);
nor U9971 (N_9971,N_9683,N_9705);
and U9972 (N_9972,N_9679,N_9663);
and U9973 (N_9973,N_9612,N_9700);
or U9974 (N_9974,N_9663,N_9797);
nor U9975 (N_9975,N_9760,N_9615);
nor U9976 (N_9976,N_9659,N_9748);
or U9977 (N_9977,N_9799,N_9659);
nor U9978 (N_9978,N_9675,N_9717);
xnor U9979 (N_9979,N_9723,N_9685);
nor U9980 (N_9980,N_9651,N_9781);
nor U9981 (N_9981,N_9656,N_9765);
nand U9982 (N_9982,N_9720,N_9630);
nor U9983 (N_9983,N_9655,N_9755);
or U9984 (N_9984,N_9619,N_9606);
xnor U9985 (N_9985,N_9678,N_9680);
and U9986 (N_9986,N_9796,N_9764);
and U9987 (N_9987,N_9735,N_9664);
xor U9988 (N_9988,N_9610,N_9658);
or U9989 (N_9989,N_9621,N_9719);
or U9990 (N_9990,N_9683,N_9743);
or U9991 (N_9991,N_9631,N_9670);
or U9992 (N_9992,N_9629,N_9695);
nor U9993 (N_9993,N_9771,N_9616);
nor U9994 (N_9994,N_9754,N_9664);
and U9995 (N_9995,N_9696,N_9765);
nand U9996 (N_9996,N_9787,N_9684);
xnor U9997 (N_9997,N_9731,N_9783);
xor U9998 (N_9998,N_9604,N_9716);
xnor U9999 (N_9999,N_9790,N_9650);
nor U10000 (N_10000,N_9824,N_9920);
nor U10001 (N_10001,N_9936,N_9997);
or U10002 (N_10002,N_9984,N_9969);
and U10003 (N_10003,N_9926,N_9859);
nor U10004 (N_10004,N_9855,N_9998);
and U10005 (N_10005,N_9891,N_9809);
nor U10006 (N_10006,N_9925,N_9911);
and U10007 (N_10007,N_9933,N_9886);
nand U10008 (N_10008,N_9934,N_9838);
nand U10009 (N_10009,N_9850,N_9975);
and U10010 (N_10010,N_9985,N_9902);
xnor U10011 (N_10011,N_9816,N_9845);
nand U10012 (N_10012,N_9873,N_9822);
and U10013 (N_10013,N_9914,N_9800);
and U10014 (N_10014,N_9875,N_9938);
xnor U10015 (N_10015,N_9930,N_9961);
xnor U10016 (N_10016,N_9804,N_9807);
nor U10017 (N_10017,N_9949,N_9946);
nor U10018 (N_10018,N_9986,N_9959);
nand U10019 (N_10019,N_9993,N_9805);
nor U10020 (N_10020,N_9843,N_9835);
or U10021 (N_10021,N_9977,N_9867);
xor U10022 (N_10022,N_9903,N_9951);
nand U10023 (N_10023,N_9987,N_9839);
xor U10024 (N_10024,N_9806,N_9910);
nor U10025 (N_10025,N_9895,N_9812);
or U10026 (N_10026,N_9917,N_9924);
nand U10027 (N_10027,N_9856,N_9918);
xnor U10028 (N_10028,N_9844,N_9954);
xnor U10029 (N_10029,N_9849,N_9955);
and U10030 (N_10030,N_9865,N_9863);
nor U10031 (N_10031,N_9942,N_9846);
and U10032 (N_10032,N_9966,N_9908);
nor U10033 (N_10033,N_9916,N_9923);
nand U10034 (N_10034,N_9858,N_9825);
nand U10035 (N_10035,N_9929,N_9992);
and U10036 (N_10036,N_9818,N_9853);
xnor U10037 (N_10037,N_9890,N_9906);
or U10038 (N_10038,N_9889,N_9888);
xnor U10039 (N_10039,N_9948,N_9940);
or U10040 (N_10040,N_9877,N_9897);
and U10041 (N_10041,N_9810,N_9848);
nor U10042 (N_10042,N_9995,N_9860);
nor U10043 (N_10043,N_9971,N_9866);
nor U10044 (N_10044,N_9893,N_9999);
and U10045 (N_10045,N_9881,N_9802);
nor U10046 (N_10046,N_9882,N_9935);
or U10047 (N_10047,N_9857,N_9978);
nor U10048 (N_10048,N_9836,N_9862);
xor U10049 (N_10049,N_9973,N_9922);
nor U10050 (N_10050,N_9988,N_9957);
and U10051 (N_10051,N_9967,N_9996);
nor U10052 (N_10052,N_9937,N_9811);
and U10053 (N_10053,N_9814,N_9823);
nor U10054 (N_10054,N_9892,N_9965);
nand U10055 (N_10055,N_9974,N_9960);
nand U10056 (N_10056,N_9912,N_9907);
xnor U10057 (N_10057,N_9833,N_9963);
and U10058 (N_10058,N_9900,N_9980);
xor U10059 (N_10059,N_9831,N_9898);
nand U10060 (N_10060,N_9899,N_9847);
and U10061 (N_10061,N_9880,N_9864);
xnor U10062 (N_10062,N_9945,N_9896);
nand U10063 (N_10063,N_9991,N_9813);
nand U10064 (N_10064,N_9851,N_9837);
nor U10065 (N_10065,N_9979,N_9989);
or U10066 (N_10066,N_9913,N_9905);
nor U10067 (N_10067,N_9976,N_9956);
xnor U10068 (N_10068,N_9808,N_9829);
and U10069 (N_10069,N_9832,N_9801);
nand U10070 (N_10070,N_9964,N_9927);
and U10071 (N_10071,N_9803,N_9874);
and U10072 (N_10072,N_9894,N_9953);
or U10073 (N_10073,N_9981,N_9958);
or U10074 (N_10074,N_9840,N_9878);
nor U10075 (N_10075,N_9854,N_9819);
nand U10076 (N_10076,N_9972,N_9943);
and U10077 (N_10077,N_9915,N_9861);
nand U10078 (N_10078,N_9952,N_9879);
or U10079 (N_10079,N_9950,N_9931);
nand U10080 (N_10080,N_9869,N_9909);
and U10081 (N_10081,N_9939,N_9887);
or U10082 (N_10082,N_9872,N_9968);
nand U10083 (N_10083,N_9830,N_9883);
nand U10084 (N_10084,N_9928,N_9821);
or U10085 (N_10085,N_9884,N_9921);
or U10086 (N_10086,N_9919,N_9941);
nor U10087 (N_10087,N_9815,N_9947);
nand U10088 (N_10088,N_9982,N_9962);
nor U10089 (N_10089,N_9827,N_9868);
nor U10090 (N_10090,N_9841,N_9852);
and U10091 (N_10091,N_9932,N_9834);
or U10092 (N_10092,N_9885,N_9970);
and U10093 (N_10093,N_9826,N_9876);
and U10094 (N_10094,N_9828,N_9983);
nor U10095 (N_10095,N_9871,N_9817);
and U10096 (N_10096,N_9994,N_9990);
nor U10097 (N_10097,N_9944,N_9870);
nor U10098 (N_10098,N_9820,N_9901);
or U10099 (N_10099,N_9904,N_9842);
nand U10100 (N_10100,N_9904,N_9938);
xor U10101 (N_10101,N_9928,N_9936);
xor U10102 (N_10102,N_9896,N_9947);
nand U10103 (N_10103,N_9895,N_9818);
xor U10104 (N_10104,N_9823,N_9992);
xor U10105 (N_10105,N_9917,N_9870);
nand U10106 (N_10106,N_9847,N_9823);
and U10107 (N_10107,N_9881,N_9939);
nand U10108 (N_10108,N_9890,N_9851);
nor U10109 (N_10109,N_9836,N_9800);
and U10110 (N_10110,N_9925,N_9862);
xnor U10111 (N_10111,N_9806,N_9889);
or U10112 (N_10112,N_9815,N_9973);
nand U10113 (N_10113,N_9955,N_9941);
and U10114 (N_10114,N_9998,N_9946);
or U10115 (N_10115,N_9997,N_9886);
nor U10116 (N_10116,N_9903,N_9909);
xor U10117 (N_10117,N_9988,N_9980);
xor U10118 (N_10118,N_9889,N_9923);
and U10119 (N_10119,N_9964,N_9858);
nor U10120 (N_10120,N_9895,N_9800);
or U10121 (N_10121,N_9950,N_9818);
xnor U10122 (N_10122,N_9871,N_9829);
or U10123 (N_10123,N_9825,N_9977);
nor U10124 (N_10124,N_9935,N_9867);
xnor U10125 (N_10125,N_9910,N_9909);
nand U10126 (N_10126,N_9935,N_9995);
nor U10127 (N_10127,N_9901,N_9880);
nand U10128 (N_10128,N_9960,N_9957);
nand U10129 (N_10129,N_9875,N_9821);
nor U10130 (N_10130,N_9867,N_9809);
or U10131 (N_10131,N_9918,N_9909);
nor U10132 (N_10132,N_9996,N_9976);
nor U10133 (N_10133,N_9926,N_9879);
nor U10134 (N_10134,N_9872,N_9907);
nand U10135 (N_10135,N_9924,N_9864);
xnor U10136 (N_10136,N_9942,N_9904);
and U10137 (N_10137,N_9846,N_9870);
xnor U10138 (N_10138,N_9821,N_9939);
nor U10139 (N_10139,N_9911,N_9984);
nor U10140 (N_10140,N_9843,N_9927);
or U10141 (N_10141,N_9933,N_9896);
or U10142 (N_10142,N_9989,N_9906);
xnor U10143 (N_10143,N_9868,N_9858);
or U10144 (N_10144,N_9990,N_9991);
or U10145 (N_10145,N_9954,N_9986);
and U10146 (N_10146,N_9898,N_9805);
xnor U10147 (N_10147,N_9904,N_9968);
nor U10148 (N_10148,N_9915,N_9957);
xor U10149 (N_10149,N_9918,N_9964);
nor U10150 (N_10150,N_9811,N_9833);
nand U10151 (N_10151,N_9862,N_9901);
and U10152 (N_10152,N_9838,N_9859);
and U10153 (N_10153,N_9958,N_9866);
or U10154 (N_10154,N_9863,N_9816);
nand U10155 (N_10155,N_9838,N_9816);
or U10156 (N_10156,N_9912,N_9898);
nor U10157 (N_10157,N_9984,N_9867);
nand U10158 (N_10158,N_9806,N_9884);
and U10159 (N_10159,N_9883,N_9975);
and U10160 (N_10160,N_9861,N_9858);
nand U10161 (N_10161,N_9990,N_9904);
and U10162 (N_10162,N_9858,N_9982);
nand U10163 (N_10163,N_9912,N_9830);
or U10164 (N_10164,N_9873,N_9850);
xnor U10165 (N_10165,N_9913,N_9954);
or U10166 (N_10166,N_9882,N_9851);
or U10167 (N_10167,N_9935,N_9923);
xor U10168 (N_10168,N_9981,N_9830);
nand U10169 (N_10169,N_9975,N_9817);
xnor U10170 (N_10170,N_9812,N_9823);
nor U10171 (N_10171,N_9856,N_9990);
nand U10172 (N_10172,N_9953,N_9911);
and U10173 (N_10173,N_9846,N_9958);
xor U10174 (N_10174,N_9873,N_9892);
xor U10175 (N_10175,N_9983,N_9923);
and U10176 (N_10176,N_9968,N_9925);
or U10177 (N_10177,N_9912,N_9836);
or U10178 (N_10178,N_9866,N_9829);
nor U10179 (N_10179,N_9956,N_9983);
xnor U10180 (N_10180,N_9827,N_9882);
nand U10181 (N_10181,N_9994,N_9960);
and U10182 (N_10182,N_9903,N_9940);
and U10183 (N_10183,N_9940,N_9869);
nor U10184 (N_10184,N_9811,N_9941);
or U10185 (N_10185,N_9833,N_9957);
nand U10186 (N_10186,N_9906,N_9893);
or U10187 (N_10187,N_9973,N_9999);
nor U10188 (N_10188,N_9944,N_9966);
nand U10189 (N_10189,N_9867,N_9947);
nor U10190 (N_10190,N_9973,N_9964);
nand U10191 (N_10191,N_9980,N_9963);
xnor U10192 (N_10192,N_9807,N_9996);
xor U10193 (N_10193,N_9812,N_9822);
xor U10194 (N_10194,N_9971,N_9896);
nand U10195 (N_10195,N_9840,N_9970);
nand U10196 (N_10196,N_9888,N_9919);
and U10197 (N_10197,N_9804,N_9814);
xnor U10198 (N_10198,N_9975,N_9868);
xnor U10199 (N_10199,N_9839,N_9937);
and U10200 (N_10200,N_10174,N_10097);
or U10201 (N_10201,N_10070,N_10060);
and U10202 (N_10202,N_10057,N_10095);
and U10203 (N_10203,N_10107,N_10169);
nor U10204 (N_10204,N_10039,N_10194);
xor U10205 (N_10205,N_10037,N_10019);
or U10206 (N_10206,N_10159,N_10007);
nor U10207 (N_10207,N_10049,N_10038);
or U10208 (N_10208,N_10062,N_10087);
xnor U10209 (N_10209,N_10025,N_10117);
nor U10210 (N_10210,N_10065,N_10138);
or U10211 (N_10211,N_10090,N_10162);
and U10212 (N_10212,N_10118,N_10156);
nor U10213 (N_10213,N_10112,N_10180);
nand U10214 (N_10214,N_10102,N_10066);
and U10215 (N_10215,N_10061,N_10084);
xor U10216 (N_10216,N_10018,N_10101);
nor U10217 (N_10217,N_10130,N_10083);
nand U10218 (N_10218,N_10023,N_10042);
or U10219 (N_10219,N_10050,N_10160);
nor U10220 (N_10220,N_10177,N_10068);
and U10221 (N_10221,N_10073,N_10195);
and U10222 (N_10222,N_10192,N_10085);
nor U10223 (N_10223,N_10030,N_10198);
nor U10224 (N_10224,N_10167,N_10136);
or U10225 (N_10225,N_10149,N_10099);
nand U10226 (N_10226,N_10148,N_10109);
nand U10227 (N_10227,N_10014,N_10092);
or U10228 (N_10228,N_10003,N_10010);
or U10229 (N_10229,N_10029,N_10185);
nand U10230 (N_10230,N_10075,N_10078);
or U10231 (N_10231,N_10187,N_10080);
nand U10232 (N_10232,N_10142,N_10123);
nand U10233 (N_10233,N_10184,N_10013);
or U10234 (N_10234,N_10017,N_10033);
nand U10235 (N_10235,N_10093,N_10100);
or U10236 (N_10236,N_10098,N_10045);
nand U10237 (N_10237,N_10145,N_10076);
nor U10238 (N_10238,N_10058,N_10155);
nand U10239 (N_10239,N_10032,N_10166);
nor U10240 (N_10240,N_10151,N_10119);
xor U10241 (N_10241,N_10041,N_10089);
xor U10242 (N_10242,N_10140,N_10122);
or U10243 (N_10243,N_10196,N_10183);
xnor U10244 (N_10244,N_10163,N_10015);
and U10245 (N_10245,N_10197,N_10081);
xnor U10246 (N_10246,N_10105,N_10168);
nand U10247 (N_10247,N_10114,N_10178);
or U10248 (N_10248,N_10141,N_10082);
and U10249 (N_10249,N_10069,N_10034);
nor U10250 (N_10250,N_10052,N_10026);
xnor U10251 (N_10251,N_10001,N_10129);
xnor U10252 (N_10252,N_10133,N_10027);
nand U10253 (N_10253,N_10055,N_10188);
or U10254 (N_10254,N_10071,N_10153);
or U10255 (N_10255,N_10022,N_10044);
or U10256 (N_10256,N_10046,N_10152);
nor U10257 (N_10257,N_10193,N_10020);
and U10258 (N_10258,N_10189,N_10059);
nor U10259 (N_10259,N_10165,N_10043);
or U10260 (N_10260,N_10000,N_10179);
and U10261 (N_10261,N_10028,N_10008);
and U10262 (N_10262,N_10175,N_10164);
xor U10263 (N_10263,N_10053,N_10063);
and U10264 (N_10264,N_10121,N_10146);
xnor U10265 (N_10265,N_10161,N_10120);
nor U10266 (N_10266,N_10173,N_10124);
nor U10267 (N_10267,N_10147,N_10054);
or U10268 (N_10268,N_10072,N_10012);
nor U10269 (N_10269,N_10077,N_10170);
nor U10270 (N_10270,N_10127,N_10171);
xor U10271 (N_10271,N_10139,N_10048);
nor U10272 (N_10272,N_10005,N_10182);
nand U10273 (N_10273,N_10191,N_10144);
xor U10274 (N_10274,N_10125,N_10016);
xor U10275 (N_10275,N_10096,N_10111);
nor U10276 (N_10276,N_10035,N_10176);
or U10277 (N_10277,N_10051,N_10158);
or U10278 (N_10278,N_10088,N_10132);
or U10279 (N_10279,N_10126,N_10031);
nor U10280 (N_10280,N_10011,N_10067);
nor U10281 (N_10281,N_10004,N_10181);
or U10282 (N_10282,N_10154,N_10172);
nor U10283 (N_10283,N_10157,N_10086);
or U10284 (N_10284,N_10056,N_10199);
and U10285 (N_10285,N_10074,N_10186);
nor U10286 (N_10286,N_10047,N_10091);
xor U10287 (N_10287,N_10108,N_10115);
nor U10288 (N_10288,N_10024,N_10131);
and U10289 (N_10289,N_10104,N_10006);
xnor U10290 (N_10290,N_10190,N_10143);
xor U10291 (N_10291,N_10103,N_10040);
nand U10292 (N_10292,N_10134,N_10110);
xnor U10293 (N_10293,N_10135,N_10137);
nand U10294 (N_10294,N_10150,N_10002);
or U10295 (N_10295,N_10128,N_10106);
or U10296 (N_10296,N_10079,N_10036);
and U10297 (N_10297,N_10021,N_10116);
nand U10298 (N_10298,N_10064,N_10113);
nand U10299 (N_10299,N_10009,N_10094);
xor U10300 (N_10300,N_10165,N_10134);
nor U10301 (N_10301,N_10143,N_10007);
and U10302 (N_10302,N_10007,N_10161);
nor U10303 (N_10303,N_10089,N_10055);
and U10304 (N_10304,N_10070,N_10019);
nand U10305 (N_10305,N_10052,N_10056);
and U10306 (N_10306,N_10181,N_10092);
and U10307 (N_10307,N_10107,N_10139);
nor U10308 (N_10308,N_10110,N_10126);
or U10309 (N_10309,N_10024,N_10190);
or U10310 (N_10310,N_10131,N_10039);
or U10311 (N_10311,N_10106,N_10187);
and U10312 (N_10312,N_10078,N_10074);
xor U10313 (N_10313,N_10116,N_10096);
nor U10314 (N_10314,N_10151,N_10118);
and U10315 (N_10315,N_10043,N_10134);
or U10316 (N_10316,N_10016,N_10060);
nand U10317 (N_10317,N_10188,N_10079);
nand U10318 (N_10318,N_10085,N_10170);
xor U10319 (N_10319,N_10120,N_10051);
nor U10320 (N_10320,N_10147,N_10169);
and U10321 (N_10321,N_10178,N_10152);
nand U10322 (N_10322,N_10127,N_10097);
and U10323 (N_10323,N_10006,N_10164);
xnor U10324 (N_10324,N_10136,N_10084);
nor U10325 (N_10325,N_10138,N_10197);
xor U10326 (N_10326,N_10034,N_10041);
and U10327 (N_10327,N_10114,N_10176);
nand U10328 (N_10328,N_10180,N_10123);
and U10329 (N_10329,N_10053,N_10193);
or U10330 (N_10330,N_10047,N_10193);
xnor U10331 (N_10331,N_10041,N_10046);
xnor U10332 (N_10332,N_10153,N_10128);
xor U10333 (N_10333,N_10142,N_10121);
xnor U10334 (N_10334,N_10130,N_10100);
xor U10335 (N_10335,N_10164,N_10011);
nand U10336 (N_10336,N_10164,N_10182);
and U10337 (N_10337,N_10169,N_10180);
and U10338 (N_10338,N_10105,N_10032);
nand U10339 (N_10339,N_10029,N_10174);
nand U10340 (N_10340,N_10196,N_10094);
xnor U10341 (N_10341,N_10091,N_10027);
nor U10342 (N_10342,N_10165,N_10051);
nand U10343 (N_10343,N_10056,N_10030);
nand U10344 (N_10344,N_10057,N_10053);
nand U10345 (N_10345,N_10159,N_10056);
or U10346 (N_10346,N_10066,N_10039);
nor U10347 (N_10347,N_10162,N_10169);
nand U10348 (N_10348,N_10068,N_10034);
and U10349 (N_10349,N_10046,N_10134);
or U10350 (N_10350,N_10181,N_10030);
xnor U10351 (N_10351,N_10117,N_10187);
nand U10352 (N_10352,N_10085,N_10181);
nor U10353 (N_10353,N_10017,N_10043);
xor U10354 (N_10354,N_10098,N_10022);
and U10355 (N_10355,N_10109,N_10115);
xor U10356 (N_10356,N_10073,N_10190);
and U10357 (N_10357,N_10099,N_10154);
nand U10358 (N_10358,N_10014,N_10159);
or U10359 (N_10359,N_10009,N_10085);
nor U10360 (N_10360,N_10117,N_10182);
nand U10361 (N_10361,N_10118,N_10024);
or U10362 (N_10362,N_10047,N_10015);
or U10363 (N_10363,N_10088,N_10041);
nand U10364 (N_10364,N_10154,N_10130);
nor U10365 (N_10365,N_10174,N_10131);
and U10366 (N_10366,N_10168,N_10110);
nand U10367 (N_10367,N_10120,N_10052);
and U10368 (N_10368,N_10165,N_10186);
or U10369 (N_10369,N_10011,N_10152);
nand U10370 (N_10370,N_10108,N_10189);
nand U10371 (N_10371,N_10175,N_10103);
xor U10372 (N_10372,N_10050,N_10137);
and U10373 (N_10373,N_10106,N_10185);
and U10374 (N_10374,N_10040,N_10116);
nand U10375 (N_10375,N_10151,N_10156);
and U10376 (N_10376,N_10129,N_10053);
nand U10377 (N_10377,N_10002,N_10139);
xor U10378 (N_10378,N_10075,N_10108);
and U10379 (N_10379,N_10087,N_10078);
or U10380 (N_10380,N_10122,N_10123);
or U10381 (N_10381,N_10053,N_10103);
nor U10382 (N_10382,N_10186,N_10169);
and U10383 (N_10383,N_10144,N_10038);
nor U10384 (N_10384,N_10119,N_10027);
or U10385 (N_10385,N_10003,N_10017);
xor U10386 (N_10386,N_10096,N_10002);
nand U10387 (N_10387,N_10052,N_10034);
and U10388 (N_10388,N_10003,N_10189);
nand U10389 (N_10389,N_10149,N_10185);
nor U10390 (N_10390,N_10115,N_10028);
or U10391 (N_10391,N_10069,N_10117);
nand U10392 (N_10392,N_10184,N_10149);
or U10393 (N_10393,N_10116,N_10183);
nand U10394 (N_10394,N_10070,N_10043);
nand U10395 (N_10395,N_10131,N_10075);
or U10396 (N_10396,N_10174,N_10178);
and U10397 (N_10397,N_10031,N_10101);
xor U10398 (N_10398,N_10010,N_10094);
nor U10399 (N_10399,N_10196,N_10014);
xor U10400 (N_10400,N_10234,N_10245);
xnor U10401 (N_10401,N_10376,N_10200);
nand U10402 (N_10402,N_10276,N_10322);
xor U10403 (N_10403,N_10394,N_10243);
nor U10404 (N_10404,N_10248,N_10347);
or U10405 (N_10405,N_10207,N_10360);
and U10406 (N_10406,N_10355,N_10235);
or U10407 (N_10407,N_10203,N_10379);
nand U10408 (N_10408,N_10268,N_10382);
xnor U10409 (N_10409,N_10393,N_10367);
nor U10410 (N_10410,N_10217,N_10252);
nand U10411 (N_10411,N_10221,N_10265);
xnor U10412 (N_10412,N_10392,N_10363);
nand U10413 (N_10413,N_10277,N_10375);
xnor U10414 (N_10414,N_10333,N_10242);
and U10415 (N_10415,N_10377,N_10349);
nand U10416 (N_10416,N_10292,N_10261);
xor U10417 (N_10417,N_10301,N_10285);
and U10418 (N_10418,N_10315,N_10353);
xnor U10419 (N_10419,N_10259,N_10237);
xor U10420 (N_10420,N_10205,N_10345);
nor U10421 (N_10421,N_10212,N_10346);
and U10422 (N_10422,N_10358,N_10303);
or U10423 (N_10423,N_10283,N_10220);
nand U10424 (N_10424,N_10371,N_10256);
xnor U10425 (N_10425,N_10238,N_10378);
and U10426 (N_10426,N_10330,N_10362);
nor U10427 (N_10427,N_10291,N_10325);
nor U10428 (N_10428,N_10269,N_10339);
nor U10429 (N_10429,N_10227,N_10289);
and U10430 (N_10430,N_10372,N_10228);
nor U10431 (N_10431,N_10241,N_10391);
xor U10432 (N_10432,N_10273,N_10249);
or U10433 (N_10433,N_10232,N_10388);
nand U10434 (N_10434,N_10326,N_10262);
or U10435 (N_10435,N_10264,N_10223);
nand U10436 (N_10436,N_10387,N_10306);
or U10437 (N_10437,N_10260,N_10370);
nor U10438 (N_10438,N_10397,N_10302);
xnor U10439 (N_10439,N_10216,N_10318);
or U10440 (N_10440,N_10218,N_10300);
and U10441 (N_10441,N_10298,N_10255);
nor U10442 (N_10442,N_10356,N_10284);
or U10443 (N_10443,N_10328,N_10295);
or U10444 (N_10444,N_10229,N_10253);
and U10445 (N_10445,N_10386,N_10314);
nand U10446 (N_10446,N_10321,N_10398);
or U10447 (N_10447,N_10257,N_10389);
xor U10448 (N_10448,N_10309,N_10350);
or U10449 (N_10449,N_10365,N_10226);
nand U10450 (N_10450,N_10396,N_10399);
xnor U10451 (N_10451,N_10266,N_10219);
nor U10452 (N_10452,N_10236,N_10327);
nand U10453 (N_10453,N_10373,N_10383);
and U10454 (N_10454,N_10351,N_10240);
nor U10455 (N_10455,N_10213,N_10204);
and U10456 (N_10456,N_10305,N_10280);
nand U10457 (N_10457,N_10274,N_10317);
or U10458 (N_10458,N_10211,N_10381);
nor U10459 (N_10459,N_10352,N_10310);
or U10460 (N_10460,N_10384,N_10331);
or U10461 (N_10461,N_10320,N_10354);
nor U10462 (N_10462,N_10272,N_10335);
and U10463 (N_10463,N_10319,N_10225);
or U10464 (N_10464,N_10290,N_10294);
and U10465 (N_10465,N_10281,N_10369);
xor U10466 (N_10466,N_10230,N_10222);
nor U10467 (N_10467,N_10390,N_10364);
and U10468 (N_10468,N_10224,N_10316);
and U10469 (N_10469,N_10296,N_10201);
xnor U10470 (N_10470,N_10214,N_10250);
nand U10471 (N_10471,N_10374,N_10247);
and U10472 (N_10472,N_10395,N_10340);
xnor U10473 (N_10473,N_10282,N_10278);
xnor U10474 (N_10474,N_10323,N_10293);
and U10475 (N_10475,N_10202,N_10279);
xor U10476 (N_10476,N_10359,N_10368);
xor U10477 (N_10477,N_10267,N_10297);
or U10478 (N_10478,N_10246,N_10304);
or U10479 (N_10479,N_10338,N_10244);
and U10480 (N_10480,N_10271,N_10357);
nor U10481 (N_10481,N_10343,N_10215);
nor U10482 (N_10482,N_10348,N_10329);
xnor U10483 (N_10483,N_10233,N_10312);
and U10484 (N_10484,N_10210,N_10311);
nor U10485 (N_10485,N_10275,N_10336);
nor U10486 (N_10486,N_10263,N_10286);
nand U10487 (N_10487,N_10344,N_10270);
and U10488 (N_10488,N_10385,N_10366);
nor U10489 (N_10489,N_10206,N_10254);
nand U10490 (N_10490,N_10334,N_10342);
or U10491 (N_10491,N_10208,N_10361);
or U10492 (N_10492,N_10239,N_10324);
and U10493 (N_10493,N_10258,N_10307);
or U10494 (N_10494,N_10313,N_10380);
or U10495 (N_10495,N_10287,N_10308);
and U10496 (N_10496,N_10341,N_10332);
nor U10497 (N_10497,N_10231,N_10209);
or U10498 (N_10498,N_10299,N_10337);
nand U10499 (N_10499,N_10288,N_10251);
and U10500 (N_10500,N_10312,N_10236);
or U10501 (N_10501,N_10314,N_10252);
or U10502 (N_10502,N_10360,N_10292);
xnor U10503 (N_10503,N_10332,N_10388);
or U10504 (N_10504,N_10378,N_10363);
and U10505 (N_10505,N_10301,N_10219);
nor U10506 (N_10506,N_10218,N_10318);
and U10507 (N_10507,N_10319,N_10239);
or U10508 (N_10508,N_10225,N_10284);
nand U10509 (N_10509,N_10362,N_10369);
or U10510 (N_10510,N_10298,N_10346);
nand U10511 (N_10511,N_10302,N_10308);
and U10512 (N_10512,N_10235,N_10206);
nor U10513 (N_10513,N_10274,N_10226);
nor U10514 (N_10514,N_10397,N_10394);
nor U10515 (N_10515,N_10333,N_10311);
and U10516 (N_10516,N_10362,N_10274);
xor U10517 (N_10517,N_10240,N_10328);
nand U10518 (N_10518,N_10266,N_10296);
and U10519 (N_10519,N_10277,N_10256);
xnor U10520 (N_10520,N_10213,N_10242);
nand U10521 (N_10521,N_10370,N_10237);
nor U10522 (N_10522,N_10261,N_10399);
xnor U10523 (N_10523,N_10258,N_10321);
xor U10524 (N_10524,N_10213,N_10343);
nor U10525 (N_10525,N_10319,N_10259);
xnor U10526 (N_10526,N_10355,N_10253);
nor U10527 (N_10527,N_10351,N_10236);
and U10528 (N_10528,N_10245,N_10214);
or U10529 (N_10529,N_10340,N_10210);
nor U10530 (N_10530,N_10208,N_10266);
nand U10531 (N_10531,N_10228,N_10391);
xor U10532 (N_10532,N_10296,N_10352);
or U10533 (N_10533,N_10217,N_10376);
xor U10534 (N_10534,N_10366,N_10375);
nor U10535 (N_10535,N_10256,N_10241);
or U10536 (N_10536,N_10307,N_10369);
nand U10537 (N_10537,N_10206,N_10213);
nand U10538 (N_10538,N_10339,N_10371);
nand U10539 (N_10539,N_10311,N_10397);
nand U10540 (N_10540,N_10296,N_10318);
nor U10541 (N_10541,N_10222,N_10301);
nor U10542 (N_10542,N_10392,N_10288);
nand U10543 (N_10543,N_10262,N_10380);
nand U10544 (N_10544,N_10278,N_10399);
nor U10545 (N_10545,N_10285,N_10281);
and U10546 (N_10546,N_10221,N_10301);
xor U10547 (N_10547,N_10251,N_10299);
xor U10548 (N_10548,N_10371,N_10338);
and U10549 (N_10549,N_10285,N_10278);
or U10550 (N_10550,N_10333,N_10347);
and U10551 (N_10551,N_10334,N_10271);
or U10552 (N_10552,N_10277,N_10212);
or U10553 (N_10553,N_10344,N_10262);
or U10554 (N_10554,N_10245,N_10297);
and U10555 (N_10555,N_10337,N_10350);
xnor U10556 (N_10556,N_10227,N_10229);
and U10557 (N_10557,N_10377,N_10229);
xnor U10558 (N_10558,N_10222,N_10217);
nor U10559 (N_10559,N_10379,N_10220);
or U10560 (N_10560,N_10291,N_10311);
nand U10561 (N_10561,N_10238,N_10353);
nand U10562 (N_10562,N_10228,N_10313);
or U10563 (N_10563,N_10272,N_10277);
or U10564 (N_10564,N_10255,N_10355);
and U10565 (N_10565,N_10309,N_10334);
or U10566 (N_10566,N_10229,N_10311);
nor U10567 (N_10567,N_10271,N_10279);
nor U10568 (N_10568,N_10295,N_10264);
nor U10569 (N_10569,N_10227,N_10359);
nor U10570 (N_10570,N_10263,N_10352);
nand U10571 (N_10571,N_10215,N_10305);
and U10572 (N_10572,N_10313,N_10252);
nor U10573 (N_10573,N_10340,N_10257);
nor U10574 (N_10574,N_10368,N_10214);
nand U10575 (N_10575,N_10303,N_10376);
and U10576 (N_10576,N_10274,N_10254);
nand U10577 (N_10577,N_10263,N_10239);
and U10578 (N_10578,N_10233,N_10252);
nand U10579 (N_10579,N_10279,N_10366);
or U10580 (N_10580,N_10293,N_10259);
nor U10581 (N_10581,N_10366,N_10322);
or U10582 (N_10582,N_10257,N_10309);
nor U10583 (N_10583,N_10271,N_10346);
xor U10584 (N_10584,N_10238,N_10300);
nor U10585 (N_10585,N_10323,N_10246);
and U10586 (N_10586,N_10280,N_10360);
or U10587 (N_10587,N_10251,N_10244);
xor U10588 (N_10588,N_10375,N_10361);
and U10589 (N_10589,N_10213,N_10351);
and U10590 (N_10590,N_10267,N_10374);
and U10591 (N_10591,N_10214,N_10311);
or U10592 (N_10592,N_10349,N_10289);
nor U10593 (N_10593,N_10297,N_10246);
and U10594 (N_10594,N_10323,N_10229);
nand U10595 (N_10595,N_10332,N_10204);
nor U10596 (N_10596,N_10356,N_10338);
or U10597 (N_10597,N_10251,N_10381);
xnor U10598 (N_10598,N_10273,N_10372);
xnor U10599 (N_10599,N_10365,N_10249);
or U10600 (N_10600,N_10594,N_10401);
nor U10601 (N_10601,N_10406,N_10539);
or U10602 (N_10602,N_10413,N_10417);
or U10603 (N_10603,N_10469,N_10433);
nand U10604 (N_10604,N_10421,N_10548);
and U10605 (N_10605,N_10590,N_10573);
nand U10606 (N_10606,N_10557,N_10400);
nor U10607 (N_10607,N_10476,N_10513);
xnor U10608 (N_10608,N_10564,N_10482);
nor U10609 (N_10609,N_10595,N_10427);
and U10610 (N_10610,N_10428,N_10467);
or U10611 (N_10611,N_10546,N_10487);
or U10612 (N_10612,N_10544,N_10515);
nor U10613 (N_10613,N_10575,N_10506);
or U10614 (N_10614,N_10446,N_10424);
and U10615 (N_10615,N_10423,N_10472);
or U10616 (N_10616,N_10597,N_10471);
nand U10617 (N_10617,N_10484,N_10567);
and U10618 (N_10618,N_10504,N_10415);
xor U10619 (N_10619,N_10583,N_10524);
and U10620 (N_10620,N_10519,N_10462);
and U10621 (N_10621,N_10532,N_10402);
nand U10622 (N_10622,N_10509,N_10456);
or U10623 (N_10623,N_10577,N_10412);
xor U10624 (N_10624,N_10522,N_10550);
nand U10625 (N_10625,N_10481,N_10449);
or U10626 (N_10626,N_10414,N_10501);
nor U10627 (N_10627,N_10475,N_10470);
xor U10628 (N_10628,N_10422,N_10478);
xnor U10629 (N_10629,N_10457,N_10510);
nor U10630 (N_10630,N_10559,N_10518);
xor U10631 (N_10631,N_10444,N_10570);
or U10632 (N_10632,N_10486,N_10566);
or U10633 (N_10633,N_10453,N_10502);
or U10634 (N_10634,N_10445,N_10463);
xor U10635 (N_10635,N_10585,N_10419);
or U10636 (N_10636,N_10547,N_10571);
and U10637 (N_10637,N_10578,N_10512);
nor U10638 (N_10638,N_10541,N_10526);
and U10639 (N_10639,N_10454,N_10480);
or U10640 (N_10640,N_10439,N_10536);
xnor U10641 (N_10641,N_10551,N_10507);
and U10642 (N_10642,N_10552,N_10591);
or U10643 (N_10643,N_10485,N_10474);
xor U10644 (N_10644,N_10572,N_10561);
xnor U10645 (N_10645,N_10473,N_10530);
or U10646 (N_10646,N_10404,N_10516);
nand U10647 (N_10647,N_10436,N_10587);
and U10648 (N_10648,N_10465,N_10574);
and U10649 (N_10649,N_10488,N_10576);
or U10650 (N_10650,N_10535,N_10565);
or U10651 (N_10651,N_10599,N_10430);
xor U10652 (N_10652,N_10549,N_10553);
nand U10653 (N_10653,N_10517,N_10496);
xnor U10654 (N_10654,N_10443,N_10477);
xor U10655 (N_10655,N_10468,N_10581);
and U10656 (N_10656,N_10556,N_10407);
and U10657 (N_10657,N_10568,N_10503);
or U10658 (N_10658,N_10435,N_10540);
nor U10659 (N_10659,N_10460,N_10589);
and U10660 (N_10660,N_10409,N_10533);
nor U10661 (N_10661,N_10429,N_10560);
and U10662 (N_10662,N_10442,N_10563);
and U10663 (N_10663,N_10529,N_10447);
nor U10664 (N_10664,N_10431,N_10514);
xnor U10665 (N_10665,N_10531,N_10493);
or U10666 (N_10666,N_10494,N_10542);
nand U10667 (N_10667,N_10466,N_10579);
xnor U10668 (N_10668,N_10558,N_10592);
and U10669 (N_10669,N_10543,N_10491);
or U10670 (N_10670,N_10489,N_10438);
nand U10671 (N_10671,N_10410,N_10459);
xor U10672 (N_10672,N_10452,N_10520);
and U10673 (N_10673,N_10495,N_10434);
xnor U10674 (N_10674,N_10437,N_10555);
nand U10675 (N_10675,N_10416,N_10426);
nand U10676 (N_10676,N_10498,N_10461);
or U10677 (N_10677,N_10420,N_10479);
nor U10678 (N_10678,N_10569,N_10483);
and U10679 (N_10679,N_10508,N_10492);
nor U10680 (N_10680,N_10440,N_10584);
nand U10681 (N_10681,N_10450,N_10458);
nand U10682 (N_10682,N_10562,N_10405);
and U10683 (N_10683,N_10545,N_10527);
and U10684 (N_10684,N_10528,N_10497);
nand U10685 (N_10685,N_10455,N_10588);
nor U10686 (N_10686,N_10500,N_10582);
xnor U10687 (N_10687,N_10523,N_10525);
or U10688 (N_10688,N_10554,N_10403);
or U10689 (N_10689,N_10441,N_10586);
nand U10690 (N_10690,N_10432,N_10418);
nand U10691 (N_10691,N_10521,N_10499);
or U10692 (N_10692,N_10511,N_10538);
or U10693 (N_10693,N_10411,N_10408);
nand U10694 (N_10694,N_10596,N_10490);
and U10695 (N_10695,N_10593,N_10425);
xnor U10696 (N_10696,N_10451,N_10598);
xnor U10697 (N_10697,N_10580,N_10534);
xnor U10698 (N_10698,N_10505,N_10464);
xor U10699 (N_10699,N_10537,N_10448);
nand U10700 (N_10700,N_10496,N_10572);
xor U10701 (N_10701,N_10540,N_10567);
nor U10702 (N_10702,N_10451,N_10570);
or U10703 (N_10703,N_10562,N_10589);
nor U10704 (N_10704,N_10471,N_10489);
and U10705 (N_10705,N_10587,N_10427);
and U10706 (N_10706,N_10443,N_10486);
xnor U10707 (N_10707,N_10479,N_10553);
nand U10708 (N_10708,N_10528,N_10545);
nand U10709 (N_10709,N_10416,N_10583);
or U10710 (N_10710,N_10539,N_10494);
and U10711 (N_10711,N_10442,N_10571);
xnor U10712 (N_10712,N_10571,N_10469);
nand U10713 (N_10713,N_10427,N_10512);
or U10714 (N_10714,N_10574,N_10415);
xor U10715 (N_10715,N_10475,N_10457);
nand U10716 (N_10716,N_10568,N_10579);
and U10717 (N_10717,N_10464,N_10515);
or U10718 (N_10718,N_10546,N_10499);
and U10719 (N_10719,N_10520,N_10439);
nor U10720 (N_10720,N_10437,N_10535);
nand U10721 (N_10721,N_10582,N_10416);
and U10722 (N_10722,N_10436,N_10475);
nand U10723 (N_10723,N_10477,N_10561);
nand U10724 (N_10724,N_10538,N_10473);
nand U10725 (N_10725,N_10403,N_10552);
xor U10726 (N_10726,N_10519,N_10529);
xor U10727 (N_10727,N_10515,N_10563);
or U10728 (N_10728,N_10526,N_10511);
nand U10729 (N_10729,N_10501,N_10523);
or U10730 (N_10730,N_10416,N_10553);
nor U10731 (N_10731,N_10573,N_10574);
nor U10732 (N_10732,N_10582,N_10523);
nor U10733 (N_10733,N_10408,N_10544);
and U10734 (N_10734,N_10405,N_10542);
nand U10735 (N_10735,N_10502,N_10429);
nand U10736 (N_10736,N_10513,N_10481);
nor U10737 (N_10737,N_10409,N_10540);
nand U10738 (N_10738,N_10516,N_10483);
xor U10739 (N_10739,N_10444,N_10584);
nand U10740 (N_10740,N_10506,N_10412);
nor U10741 (N_10741,N_10549,N_10416);
or U10742 (N_10742,N_10401,N_10425);
or U10743 (N_10743,N_10599,N_10539);
nor U10744 (N_10744,N_10507,N_10522);
or U10745 (N_10745,N_10566,N_10437);
or U10746 (N_10746,N_10532,N_10441);
xor U10747 (N_10747,N_10463,N_10509);
xnor U10748 (N_10748,N_10484,N_10415);
nor U10749 (N_10749,N_10426,N_10518);
or U10750 (N_10750,N_10597,N_10479);
or U10751 (N_10751,N_10528,N_10513);
nor U10752 (N_10752,N_10541,N_10423);
nand U10753 (N_10753,N_10427,N_10470);
and U10754 (N_10754,N_10496,N_10523);
nor U10755 (N_10755,N_10454,N_10443);
and U10756 (N_10756,N_10476,N_10439);
or U10757 (N_10757,N_10443,N_10452);
nand U10758 (N_10758,N_10574,N_10476);
or U10759 (N_10759,N_10528,N_10457);
or U10760 (N_10760,N_10505,N_10578);
nand U10761 (N_10761,N_10403,N_10426);
nand U10762 (N_10762,N_10520,N_10567);
xor U10763 (N_10763,N_10401,N_10491);
and U10764 (N_10764,N_10471,N_10590);
nor U10765 (N_10765,N_10565,N_10567);
xor U10766 (N_10766,N_10554,N_10585);
or U10767 (N_10767,N_10405,N_10508);
nor U10768 (N_10768,N_10428,N_10430);
and U10769 (N_10769,N_10421,N_10422);
nand U10770 (N_10770,N_10521,N_10442);
and U10771 (N_10771,N_10509,N_10419);
xor U10772 (N_10772,N_10443,N_10458);
xor U10773 (N_10773,N_10492,N_10570);
nor U10774 (N_10774,N_10445,N_10440);
xnor U10775 (N_10775,N_10427,N_10454);
and U10776 (N_10776,N_10541,N_10420);
nand U10777 (N_10777,N_10431,N_10568);
and U10778 (N_10778,N_10459,N_10408);
nor U10779 (N_10779,N_10554,N_10488);
nand U10780 (N_10780,N_10533,N_10582);
and U10781 (N_10781,N_10493,N_10565);
xor U10782 (N_10782,N_10401,N_10417);
nor U10783 (N_10783,N_10539,N_10592);
or U10784 (N_10784,N_10548,N_10504);
nand U10785 (N_10785,N_10528,N_10558);
and U10786 (N_10786,N_10474,N_10483);
nand U10787 (N_10787,N_10424,N_10431);
nor U10788 (N_10788,N_10490,N_10582);
xnor U10789 (N_10789,N_10484,N_10586);
xnor U10790 (N_10790,N_10573,N_10497);
xnor U10791 (N_10791,N_10506,N_10461);
and U10792 (N_10792,N_10431,N_10502);
xnor U10793 (N_10793,N_10586,N_10407);
or U10794 (N_10794,N_10477,N_10598);
xor U10795 (N_10795,N_10514,N_10547);
or U10796 (N_10796,N_10525,N_10579);
and U10797 (N_10797,N_10593,N_10438);
and U10798 (N_10798,N_10540,N_10467);
nor U10799 (N_10799,N_10422,N_10511);
or U10800 (N_10800,N_10617,N_10722);
or U10801 (N_10801,N_10669,N_10672);
and U10802 (N_10802,N_10680,N_10618);
xor U10803 (N_10803,N_10629,N_10797);
nand U10804 (N_10804,N_10671,N_10741);
or U10805 (N_10805,N_10723,N_10656);
xor U10806 (N_10806,N_10696,N_10645);
nor U10807 (N_10807,N_10615,N_10790);
xor U10808 (N_10808,N_10730,N_10627);
nand U10809 (N_10809,N_10699,N_10609);
and U10810 (N_10810,N_10694,N_10710);
and U10811 (N_10811,N_10632,N_10726);
xor U10812 (N_10812,N_10626,N_10714);
nand U10813 (N_10813,N_10707,N_10700);
and U10814 (N_10814,N_10716,N_10762);
nor U10815 (N_10815,N_10650,N_10796);
or U10816 (N_10816,N_10621,N_10701);
xnor U10817 (N_10817,N_10674,N_10789);
nand U10818 (N_10818,N_10668,N_10743);
nor U10819 (N_10819,N_10685,N_10660);
nand U10820 (N_10820,N_10739,N_10642);
nor U10821 (N_10821,N_10654,N_10677);
or U10822 (N_10822,N_10745,N_10765);
or U10823 (N_10823,N_10653,N_10784);
xnor U10824 (N_10824,N_10690,N_10795);
nand U10825 (N_10825,N_10753,N_10704);
nor U10826 (N_10826,N_10759,N_10610);
nor U10827 (N_10827,N_10778,N_10736);
xor U10828 (N_10828,N_10623,N_10752);
and U10829 (N_10829,N_10738,N_10768);
and U10830 (N_10830,N_10773,N_10604);
or U10831 (N_10831,N_10608,N_10721);
or U10832 (N_10832,N_10639,N_10683);
nand U10833 (N_10833,N_10785,N_10719);
and U10834 (N_10834,N_10729,N_10709);
nand U10835 (N_10835,N_10662,N_10692);
nor U10836 (N_10836,N_10625,N_10611);
xnor U10837 (N_10837,N_10687,N_10786);
xnor U10838 (N_10838,N_10655,N_10792);
nand U10839 (N_10839,N_10775,N_10757);
xnor U10840 (N_10840,N_10652,N_10619);
xnor U10841 (N_10841,N_10770,N_10640);
and U10842 (N_10842,N_10600,N_10737);
xnor U10843 (N_10843,N_10670,N_10760);
nand U10844 (N_10844,N_10673,N_10788);
and U10845 (N_10845,N_10798,N_10733);
and U10846 (N_10846,N_10676,N_10746);
xnor U10847 (N_10847,N_10780,N_10612);
nand U10848 (N_10848,N_10658,N_10606);
xnor U10849 (N_10849,N_10706,N_10666);
xnor U10850 (N_10850,N_10659,N_10742);
nand U10851 (N_10851,N_10767,N_10637);
and U10852 (N_10852,N_10764,N_10607);
and U10853 (N_10853,N_10631,N_10732);
xor U10854 (N_10854,N_10689,N_10712);
xnor U10855 (N_10855,N_10682,N_10684);
or U10856 (N_10856,N_10636,N_10693);
nand U10857 (N_10857,N_10601,N_10643);
and U10858 (N_10858,N_10794,N_10667);
nand U10859 (N_10859,N_10755,N_10624);
or U10860 (N_10860,N_10657,N_10748);
or U10861 (N_10861,N_10782,N_10695);
and U10862 (N_10862,N_10720,N_10781);
or U10863 (N_10863,N_10605,N_10776);
xnor U10864 (N_10864,N_10756,N_10681);
xor U10865 (N_10865,N_10679,N_10661);
or U10866 (N_10866,N_10638,N_10711);
xor U10867 (N_10867,N_10686,N_10634);
xor U10868 (N_10868,N_10774,N_10761);
and U10869 (N_10869,N_10705,N_10630);
and U10870 (N_10870,N_10688,N_10675);
or U10871 (N_10871,N_10791,N_10787);
xnor U10872 (N_10872,N_10799,N_10648);
and U10873 (N_10873,N_10703,N_10702);
and U10874 (N_10874,N_10664,N_10633);
or U10875 (N_10875,N_10717,N_10735);
and U10876 (N_10876,N_10644,N_10725);
xnor U10877 (N_10877,N_10763,N_10731);
xor U10878 (N_10878,N_10678,N_10744);
xnor U10879 (N_10879,N_10647,N_10758);
nand U10880 (N_10880,N_10779,N_10740);
and U10881 (N_10881,N_10620,N_10777);
and U10882 (N_10882,N_10665,N_10747);
nand U10883 (N_10883,N_10635,N_10641);
nand U10884 (N_10884,N_10691,N_10628);
nor U10885 (N_10885,N_10771,N_10754);
nand U10886 (N_10886,N_10622,N_10651);
nor U10887 (N_10887,N_10783,N_10649);
nand U10888 (N_10888,N_10769,N_10616);
nand U10889 (N_10889,N_10715,N_10728);
and U10890 (N_10890,N_10734,N_10793);
nand U10891 (N_10891,N_10602,N_10613);
nor U10892 (N_10892,N_10614,N_10727);
xnor U10893 (N_10893,N_10718,N_10772);
nor U10894 (N_10894,N_10697,N_10698);
or U10895 (N_10895,N_10646,N_10663);
and U10896 (N_10896,N_10713,N_10603);
nand U10897 (N_10897,N_10750,N_10766);
or U10898 (N_10898,N_10751,N_10724);
xor U10899 (N_10899,N_10708,N_10749);
or U10900 (N_10900,N_10757,N_10712);
xor U10901 (N_10901,N_10746,N_10768);
nand U10902 (N_10902,N_10733,N_10642);
or U10903 (N_10903,N_10757,N_10648);
or U10904 (N_10904,N_10693,N_10677);
nand U10905 (N_10905,N_10675,N_10642);
xor U10906 (N_10906,N_10662,N_10771);
and U10907 (N_10907,N_10790,N_10631);
nor U10908 (N_10908,N_10663,N_10747);
and U10909 (N_10909,N_10751,N_10693);
or U10910 (N_10910,N_10732,N_10782);
or U10911 (N_10911,N_10683,N_10621);
xnor U10912 (N_10912,N_10608,N_10753);
nor U10913 (N_10913,N_10642,N_10748);
xnor U10914 (N_10914,N_10792,N_10780);
xnor U10915 (N_10915,N_10701,N_10727);
nand U10916 (N_10916,N_10756,N_10745);
or U10917 (N_10917,N_10703,N_10643);
nand U10918 (N_10918,N_10742,N_10740);
nand U10919 (N_10919,N_10621,N_10758);
and U10920 (N_10920,N_10667,N_10697);
nor U10921 (N_10921,N_10713,N_10740);
and U10922 (N_10922,N_10752,N_10602);
and U10923 (N_10923,N_10611,N_10708);
or U10924 (N_10924,N_10702,N_10636);
and U10925 (N_10925,N_10703,N_10688);
nor U10926 (N_10926,N_10679,N_10757);
and U10927 (N_10927,N_10688,N_10701);
nor U10928 (N_10928,N_10605,N_10751);
or U10929 (N_10929,N_10643,N_10709);
or U10930 (N_10930,N_10713,N_10687);
xnor U10931 (N_10931,N_10726,N_10730);
and U10932 (N_10932,N_10718,N_10657);
xor U10933 (N_10933,N_10665,N_10789);
nor U10934 (N_10934,N_10617,N_10659);
nand U10935 (N_10935,N_10705,N_10780);
nand U10936 (N_10936,N_10798,N_10653);
nand U10937 (N_10937,N_10691,N_10777);
xnor U10938 (N_10938,N_10741,N_10678);
nand U10939 (N_10939,N_10639,N_10641);
and U10940 (N_10940,N_10687,N_10794);
xnor U10941 (N_10941,N_10613,N_10620);
xnor U10942 (N_10942,N_10740,N_10796);
and U10943 (N_10943,N_10614,N_10782);
and U10944 (N_10944,N_10636,N_10712);
and U10945 (N_10945,N_10631,N_10741);
xor U10946 (N_10946,N_10611,N_10725);
nor U10947 (N_10947,N_10696,N_10622);
and U10948 (N_10948,N_10754,N_10642);
xor U10949 (N_10949,N_10747,N_10780);
xnor U10950 (N_10950,N_10758,N_10602);
or U10951 (N_10951,N_10674,N_10659);
or U10952 (N_10952,N_10657,N_10615);
and U10953 (N_10953,N_10652,N_10717);
and U10954 (N_10954,N_10663,N_10714);
or U10955 (N_10955,N_10683,N_10668);
nand U10956 (N_10956,N_10748,N_10611);
and U10957 (N_10957,N_10765,N_10657);
and U10958 (N_10958,N_10729,N_10619);
nor U10959 (N_10959,N_10660,N_10691);
nand U10960 (N_10960,N_10680,N_10737);
nor U10961 (N_10961,N_10618,N_10655);
and U10962 (N_10962,N_10679,N_10654);
nand U10963 (N_10963,N_10740,N_10738);
and U10964 (N_10964,N_10778,N_10662);
or U10965 (N_10965,N_10631,N_10701);
xnor U10966 (N_10966,N_10731,N_10746);
nor U10967 (N_10967,N_10696,N_10771);
or U10968 (N_10968,N_10628,N_10617);
xor U10969 (N_10969,N_10729,N_10679);
nand U10970 (N_10970,N_10655,N_10627);
nor U10971 (N_10971,N_10707,N_10668);
and U10972 (N_10972,N_10771,N_10692);
nor U10973 (N_10973,N_10644,N_10722);
nand U10974 (N_10974,N_10738,N_10794);
and U10975 (N_10975,N_10759,N_10717);
and U10976 (N_10976,N_10670,N_10654);
xnor U10977 (N_10977,N_10638,N_10641);
or U10978 (N_10978,N_10602,N_10673);
and U10979 (N_10979,N_10702,N_10676);
xor U10980 (N_10980,N_10604,N_10779);
or U10981 (N_10981,N_10789,N_10664);
xor U10982 (N_10982,N_10628,N_10636);
and U10983 (N_10983,N_10662,N_10720);
nand U10984 (N_10984,N_10604,N_10608);
nor U10985 (N_10985,N_10683,N_10782);
nor U10986 (N_10986,N_10743,N_10788);
or U10987 (N_10987,N_10738,N_10790);
nor U10988 (N_10988,N_10674,N_10714);
and U10989 (N_10989,N_10742,N_10642);
or U10990 (N_10990,N_10728,N_10756);
nand U10991 (N_10991,N_10761,N_10619);
or U10992 (N_10992,N_10642,N_10718);
and U10993 (N_10993,N_10759,N_10779);
xor U10994 (N_10994,N_10780,N_10646);
nor U10995 (N_10995,N_10777,N_10680);
and U10996 (N_10996,N_10646,N_10671);
and U10997 (N_10997,N_10631,N_10672);
nor U10998 (N_10998,N_10679,N_10687);
xor U10999 (N_10999,N_10771,N_10641);
or U11000 (N_11000,N_10922,N_10864);
or U11001 (N_11001,N_10872,N_10917);
xnor U11002 (N_11002,N_10983,N_10833);
nand U11003 (N_11003,N_10956,N_10957);
nor U11004 (N_11004,N_10986,N_10952);
or U11005 (N_11005,N_10846,N_10978);
and U11006 (N_11006,N_10891,N_10859);
or U11007 (N_11007,N_10822,N_10892);
or U11008 (N_11008,N_10874,N_10897);
nor U11009 (N_11009,N_10987,N_10849);
or U11010 (N_11010,N_10933,N_10930);
or U11011 (N_11011,N_10816,N_10903);
and U11012 (N_11012,N_10838,N_10860);
and U11013 (N_11013,N_10946,N_10958);
and U11014 (N_11014,N_10841,N_10847);
and U11015 (N_11015,N_10994,N_10951);
nand U11016 (N_11016,N_10955,N_10904);
nand U11017 (N_11017,N_10887,N_10858);
and U11018 (N_11018,N_10916,N_10975);
nand U11019 (N_11019,N_10912,N_10837);
nand U11020 (N_11020,N_10880,N_10932);
nor U11021 (N_11021,N_10959,N_10905);
or U11022 (N_11022,N_10811,N_10909);
nor U11023 (N_11023,N_10857,N_10876);
and U11024 (N_11024,N_10999,N_10913);
xnor U11025 (N_11025,N_10843,N_10800);
xnor U11026 (N_11026,N_10801,N_10856);
and U11027 (N_11027,N_10873,N_10942);
nor U11028 (N_11028,N_10899,N_10971);
or U11029 (N_11029,N_10940,N_10921);
xor U11030 (N_11030,N_10862,N_10883);
or U11031 (N_11031,N_10855,N_10911);
or U11032 (N_11032,N_10980,N_10947);
and U11033 (N_11033,N_10949,N_10884);
xnor U11034 (N_11034,N_10981,N_10906);
xnor U11035 (N_11035,N_10818,N_10854);
xnor U11036 (N_11036,N_10902,N_10826);
nor U11037 (N_11037,N_10842,N_10937);
or U11038 (N_11038,N_10961,N_10962);
xor U11039 (N_11039,N_10945,N_10870);
xnor U11040 (N_11040,N_10943,N_10893);
or U11041 (N_11041,N_10821,N_10819);
or U11042 (N_11042,N_10886,N_10964);
and U11043 (N_11043,N_10820,N_10993);
and U11044 (N_11044,N_10813,N_10831);
nand U11045 (N_11045,N_10806,N_10944);
nand U11046 (N_11046,N_10900,N_10827);
and U11047 (N_11047,N_10895,N_10882);
nor U11048 (N_11048,N_10966,N_10844);
nor U11049 (N_11049,N_10866,N_10823);
and U11050 (N_11050,N_10936,N_10901);
nand U11051 (N_11051,N_10894,N_10918);
xor U11052 (N_11052,N_10852,N_10889);
or U11053 (N_11053,N_10914,N_10969);
nor U11054 (N_11054,N_10929,N_10853);
and U11055 (N_11055,N_10878,N_10840);
nand U11056 (N_11056,N_10898,N_10881);
and U11057 (N_11057,N_10834,N_10809);
nand U11058 (N_11058,N_10803,N_10997);
or U11059 (N_11059,N_10845,N_10808);
or U11060 (N_11060,N_10863,N_10968);
nor U11061 (N_11061,N_10954,N_10976);
and U11062 (N_11062,N_10972,N_10877);
or U11063 (N_11063,N_10825,N_10868);
or U11064 (N_11064,N_10817,N_10979);
or U11065 (N_11065,N_10850,N_10805);
and U11066 (N_11066,N_10867,N_10991);
nand U11067 (N_11067,N_10888,N_10998);
xnor U11068 (N_11068,N_10875,N_10848);
nor U11069 (N_11069,N_10814,N_10824);
nand U11070 (N_11070,N_10920,N_10829);
and U11071 (N_11071,N_10938,N_10965);
xor U11072 (N_11072,N_10995,N_10941);
or U11073 (N_11073,N_10931,N_10832);
nand U11074 (N_11074,N_10984,N_10908);
and U11075 (N_11075,N_10835,N_10926);
nand U11076 (N_11076,N_10915,N_10896);
xnor U11077 (N_11077,N_10974,N_10963);
nor U11078 (N_11078,N_10970,N_10925);
nand U11079 (N_11079,N_10934,N_10927);
and U11080 (N_11080,N_10990,N_10815);
or U11081 (N_11081,N_10907,N_10928);
and U11082 (N_11082,N_10967,N_10935);
nand U11083 (N_11083,N_10953,N_10923);
nor U11084 (N_11084,N_10973,N_10977);
xor U11085 (N_11085,N_10890,N_10950);
xor U11086 (N_11086,N_10851,N_10948);
nor U11087 (N_11087,N_10992,N_10989);
and U11088 (N_11088,N_10960,N_10871);
or U11089 (N_11089,N_10865,N_10996);
and U11090 (N_11090,N_10939,N_10879);
nor U11091 (N_11091,N_10812,N_10828);
xnor U11092 (N_11092,N_10830,N_10807);
nand U11093 (N_11093,N_10919,N_10924);
xnor U11094 (N_11094,N_10836,N_10810);
and U11095 (N_11095,N_10861,N_10988);
and U11096 (N_11096,N_10802,N_10839);
and U11097 (N_11097,N_10885,N_10869);
nor U11098 (N_11098,N_10982,N_10985);
xnor U11099 (N_11099,N_10804,N_10910);
or U11100 (N_11100,N_10930,N_10924);
and U11101 (N_11101,N_10871,N_10991);
nor U11102 (N_11102,N_10941,N_10971);
and U11103 (N_11103,N_10957,N_10912);
or U11104 (N_11104,N_10910,N_10969);
nor U11105 (N_11105,N_10950,N_10835);
nand U11106 (N_11106,N_10941,N_10936);
xnor U11107 (N_11107,N_10965,N_10881);
nor U11108 (N_11108,N_10867,N_10944);
nor U11109 (N_11109,N_10870,N_10995);
xor U11110 (N_11110,N_10963,N_10968);
nand U11111 (N_11111,N_10874,N_10961);
and U11112 (N_11112,N_10875,N_10977);
nor U11113 (N_11113,N_10994,N_10933);
nor U11114 (N_11114,N_10915,N_10870);
nand U11115 (N_11115,N_10891,N_10835);
xor U11116 (N_11116,N_10934,N_10861);
nor U11117 (N_11117,N_10879,N_10890);
nor U11118 (N_11118,N_10814,N_10918);
xnor U11119 (N_11119,N_10869,N_10925);
xor U11120 (N_11120,N_10801,N_10844);
xor U11121 (N_11121,N_10883,N_10984);
nor U11122 (N_11122,N_10917,N_10950);
xnor U11123 (N_11123,N_10935,N_10800);
nand U11124 (N_11124,N_10950,N_10901);
or U11125 (N_11125,N_10926,N_10848);
or U11126 (N_11126,N_10939,N_10933);
xnor U11127 (N_11127,N_10931,N_10921);
nor U11128 (N_11128,N_10823,N_10872);
nor U11129 (N_11129,N_10897,N_10947);
and U11130 (N_11130,N_10825,N_10998);
xnor U11131 (N_11131,N_10996,N_10886);
and U11132 (N_11132,N_10872,N_10801);
and U11133 (N_11133,N_10848,N_10898);
nand U11134 (N_11134,N_10994,N_10941);
nand U11135 (N_11135,N_10977,N_10905);
nor U11136 (N_11136,N_10831,N_10991);
nand U11137 (N_11137,N_10974,N_10975);
and U11138 (N_11138,N_10816,N_10930);
nand U11139 (N_11139,N_10992,N_10963);
and U11140 (N_11140,N_10889,N_10815);
nor U11141 (N_11141,N_10973,N_10884);
nor U11142 (N_11142,N_10886,N_10992);
nor U11143 (N_11143,N_10926,N_10981);
nand U11144 (N_11144,N_10888,N_10875);
and U11145 (N_11145,N_10814,N_10941);
nand U11146 (N_11146,N_10919,N_10830);
and U11147 (N_11147,N_10862,N_10918);
and U11148 (N_11148,N_10923,N_10938);
nand U11149 (N_11149,N_10961,N_10857);
and U11150 (N_11150,N_10844,N_10806);
nand U11151 (N_11151,N_10926,N_10803);
nand U11152 (N_11152,N_10943,N_10901);
xor U11153 (N_11153,N_10958,N_10878);
nor U11154 (N_11154,N_10869,N_10862);
nand U11155 (N_11155,N_10943,N_10942);
or U11156 (N_11156,N_10813,N_10958);
xnor U11157 (N_11157,N_10805,N_10942);
or U11158 (N_11158,N_10977,N_10923);
nor U11159 (N_11159,N_10908,N_10904);
nor U11160 (N_11160,N_10831,N_10959);
or U11161 (N_11161,N_10894,N_10857);
or U11162 (N_11162,N_10938,N_10830);
or U11163 (N_11163,N_10880,N_10813);
nand U11164 (N_11164,N_10871,N_10813);
and U11165 (N_11165,N_10967,N_10870);
or U11166 (N_11166,N_10876,N_10819);
or U11167 (N_11167,N_10871,N_10976);
nor U11168 (N_11168,N_10918,N_10954);
nand U11169 (N_11169,N_10818,N_10919);
and U11170 (N_11170,N_10913,N_10893);
or U11171 (N_11171,N_10854,N_10916);
xnor U11172 (N_11172,N_10855,N_10931);
nor U11173 (N_11173,N_10915,N_10997);
xnor U11174 (N_11174,N_10886,N_10831);
nor U11175 (N_11175,N_10854,N_10883);
xor U11176 (N_11176,N_10995,N_10948);
xor U11177 (N_11177,N_10971,N_10983);
and U11178 (N_11178,N_10848,N_10906);
nand U11179 (N_11179,N_10815,N_10818);
or U11180 (N_11180,N_10831,N_10805);
or U11181 (N_11181,N_10948,N_10955);
or U11182 (N_11182,N_10944,N_10949);
xnor U11183 (N_11183,N_10862,N_10853);
or U11184 (N_11184,N_10914,N_10827);
and U11185 (N_11185,N_10905,N_10989);
and U11186 (N_11186,N_10931,N_10901);
nand U11187 (N_11187,N_10820,N_10912);
nand U11188 (N_11188,N_10890,N_10839);
nor U11189 (N_11189,N_10840,N_10841);
and U11190 (N_11190,N_10913,N_10806);
nand U11191 (N_11191,N_10989,N_10971);
xor U11192 (N_11192,N_10898,N_10973);
xnor U11193 (N_11193,N_10844,N_10949);
and U11194 (N_11194,N_10965,N_10993);
or U11195 (N_11195,N_10897,N_10948);
and U11196 (N_11196,N_10875,N_10981);
nand U11197 (N_11197,N_10957,N_10907);
or U11198 (N_11198,N_10920,N_10994);
xor U11199 (N_11199,N_10857,N_10924);
and U11200 (N_11200,N_11080,N_11073);
or U11201 (N_11201,N_11039,N_11170);
xnor U11202 (N_11202,N_11146,N_11103);
and U11203 (N_11203,N_11153,N_11044);
xnor U11204 (N_11204,N_11158,N_11054);
xnor U11205 (N_11205,N_11114,N_11083);
xnor U11206 (N_11206,N_11183,N_11070);
nor U11207 (N_11207,N_11067,N_11042);
nor U11208 (N_11208,N_11018,N_11078);
nor U11209 (N_11209,N_11087,N_11189);
or U11210 (N_11210,N_11156,N_11137);
and U11211 (N_11211,N_11021,N_11141);
xor U11212 (N_11212,N_11108,N_11188);
nand U11213 (N_11213,N_11035,N_11048);
and U11214 (N_11214,N_11192,N_11079);
xor U11215 (N_11215,N_11016,N_11033);
or U11216 (N_11216,N_11012,N_11068);
xnor U11217 (N_11217,N_11050,N_11123);
nand U11218 (N_11218,N_11071,N_11027);
or U11219 (N_11219,N_11008,N_11149);
and U11220 (N_11220,N_11164,N_11166);
nor U11221 (N_11221,N_11101,N_11106);
nand U11222 (N_11222,N_11161,N_11095);
nand U11223 (N_11223,N_11090,N_11117);
or U11224 (N_11224,N_11126,N_11125);
nand U11225 (N_11225,N_11124,N_11185);
nor U11226 (N_11226,N_11029,N_11081);
nand U11227 (N_11227,N_11005,N_11194);
and U11228 (N_11228,N_11020,N_11074);
nor U11229 (N_11229,N_11198,N_11134);
nor U11230 (N_11230,N_11061,N_11131);
nor U11231 (N_11231,N_11136,N_11017);
and U11232 (N_11232,N_11168,N_11142);
and U11233 (N_11233,N_11178,N_11115);
xor U11234 (N_11234,N_11129,N_11046);
or U11235 (N_11235,N_11197,N_11152);
nand U11236 (N_11236,N_11196,N_11034);
or U11237 (N_11237,N_11147,N_11037);
and U11238 (N_11238,N_11144,N_11069);
xor U11239 (N_11239,N_11043,N_11065);
or U11240 (N_11240,N_11132,N_11036);
and U11241 (N_11241,N_11025,N_11000);
and U11242 (N_11242,N_11075,N_11176);
xnor U11243 (N_11243,N_11055,N_11066);
xor U11244 (N_11244,N_11002,N_11118);
and U11245 (N_11245,N_11171,N_11187);
nor U11246 (N_11246,N_11006,N_11127);
xor U11247 (N_11247,N_11133,N_11184);
nor U11248 (N_11248,N_11135,N_11096);
or U11249 (N_11249,N_11140,N_11177);
or U11250 (N_11250,N_11179,N_11102);
or U11251 (N_11251,N_11077,N_11122);
xor U11252 (N_11252,N_11173,N_11191);
nand U11253 (N_11253,N_11180,N_11195);
xnor U11254 (N_11254,N_11172,N_11120);
or U11255 (N_11255,N_11084,N_11104);
nor U11256 (N_11256,N_11182,N_11064);
xor U11257 (N_11257,N_11009,N_11091);
nand U11258 (N_11258,N_11139,N_11190);
or U11259 (N_11259,N_11072,N_11150);
nor U11260 (N_11260,N_11162,N_11024);
and U11261 (N_11261,N_11003,N_11053);
or U11262 (N_11262,N_11110,N_11099);
xor U11263 (N_11263,N_11022,N_11093);
nand U11264 (N_11264,N_11119,N_11098);
and U11265 (N_11265,N_11011,N_11138);
or U11266 (N_11266,N_11026,N_11089);
and U11267 (N_11267,N_11100,N_11051);
and U11268 (N_11268,N_11057,N_11023);
nor U11269 (N_11269,N_11130,N_11169);
or U11270 (N_11270,N_11014,N_11094);
and U11271 (N_11271,N_11097,N_11085);
xnor U11272 (N_11272,N_11128,N_11088);
nor U11273 (N_11273,N_11052,N_11181);
nor U11274 (N_11274,N_11186,N_11047);
xor U11275 (N_11275,N_11121,N_11111);
and U11276 (N_11276,N_11030,N_11159);
xor U11277 (N_11277,N_11040,N_11060);
and U11278 (N_11278,N_11063,N_11157);
xor U11279 (N_11279,N_11007,N_11148);
xnor U11280 (N_11280,N_11160,N_11059);
nand U11281 (N_11281,N_11032,N_11193);
nor U11282 (N_11282,N_11151,N_11105);
or U11283 (N_11283,N_11154,N_11001);
xnor U11284 (N_11284,N_11143,N_11086);
or U11285 (N_11285,N_11109,N_11165);
nor U11286 (N_11286,N_11107,N_11028);
and U11287 (N_11287,N_11045,N_11041);
and U11288 (N_11288,N_11013,N_11155);
xor U11289 (N_11289,N_11058,N_11163);
xor U11290 (N_11290,N_11116,N_11175);
or U11291 (N_11291,N_11167,N_11031);
nor U11292 (N_11292,N_11199,N_11145);
or U11293 (N_11293,N_11174,N_11076);
nor U11294 (N_11294,N_11015,N_11019);
and U11295 (N_11295,N_11049,N_11092);
nor U11296 (N_11296,N_11056,N_11113);
xnor U11297 (N_11297,N_11010,N_11082);
nor U11298 (N_11298,N_11062,N_11038);
xnor U11299 (N_11299,N_11004,N_11112);
or U11300 (N_11300,N_11005,N_11160);
nand U11301 (N_11301,N_11174,N_11080);
and U11302 (N_11302,N_11178,N_11059);
nand U11303 (N_11303,N_11170,N_11117);
and U11304 (N_11304,N_11017,N_11081);
and U11305 (N_11305,N_11107,N_11058);
nand U11306 (N_11306,N_11137,N_11033);
nand U11307 (N_11307,N_11093,N_11145);
nor U11308 (N_11308,N_11153,N_11117);
nor U11309 (N_11309,N_11026,N_11071);
or U11310 (N_11310,N_11144,N_11044);
xnor U11311 (N_11311,N_11022,N_11173);
nor U11312 (N_11312,N_11024,N_11106);
nor U11313 (N_11313,N_11115,N_11124);
xnor U11314 (N_11314,N_11041,N_11178);
and U11315 (N_11315,N_11114,N_11167);
or U11316 (N_11316,N_11016,N_11138);
xnor U11317 (N_11317,N_11016,N_11195);
or U11318 (N_11318,N_11155,N_11051);
xnor U11319 (N_11319,N_11144,N_11145);
nand U11320 (N_11320,N_11035,N_11058);
nand U11321 (N_11321,N_11013,N_11004);
nand U11322 (N_11322,N_11048,N_11158);
nor U11323 (N_11323,N_11101,N_11107);
nand U11324 (N_11324,N_11103,N_11056);
nor U11325 (N_11325,N_11161,N_11100);
nor U11326 (N_11326,N_11112,N_11037);
xnor U11327 (N_11327,N_11007,N_11159);
and U11328 (N_11328,N_11062,N_11015);
xor U11329 (N_11329,N_11122,N_11135);
and U11330 (N_11330,N_11112,N_11109);
nand U11331 (N_11331,N_11110,N_11194);
xor U11332 (N_11332,N_11151,N_11076);
or U11333 (N_11333,N_11176,N_11109);
nand U11334 (N_11334,N_11171,N_11075);
or U11335 (N_11335,N_11060,N_11086);
xnor U11336 (N_11336,N_11181,N_11191);
and U11337 (N_11337,N_11063,N_11027);
nor U11338 (N_11338,N_11069,N_11021);
or U11339 (N_11339,N_11083,N_11130);
nor U11340 (N_11340,N_11033,N_11038);
xnor U11341 (N_11341,N_11168,N_11162);
nor U11342 (N_11342,N_11068,N_11121);
or U11343 (N_11343,N_11134,N_11132);
nor U11344 (N_11344,N_11134,N_11031);
or U11345 (N_11345,N_11068,N_11170);
or U11346 (N_11346,N_11167,N_11123);
xnor U11347 (N_11347,N_11110,N_11151);
and U11348 (N_11348,N_11054,N_11021);
nand U11349 (N_11349,N_11110,N_11162);
nand U11350 (N_11350,N_11108,N_11027);
or U11351 (N_11351,N_11097,N_11189);
nand U11352 (N_11352,N_11072,N_11184);
nand U11353 (N_11353,N_11145,N_11198);
nor U11354 (N_11354,N_11133,N_11031);
nand U11355 (N_11355,N_11123,N_11152);
nor U11356 (N_11356,N_11104,N_11139);
or U11357 (N_11357,N_11182,N_11046);
nor U11358 (N_11358,N_11051,N_11045);
nand U11359 (N_11359,N_11006,N_11190);
nor U11360 (N_11360,N_11184,N_11193);
or U11361 (N_11361,N_11048,N_11083);
xor U11362 (N_11362,N_11154,N_11083);
or U11363 (N_11363,N_11112,N_11036);
xor U11364 (N_11364,N_11064,N_11047);
nor U11365 (N_11365,N_11002,N_11061);
or U11366 (N_11366,N_11022,N_11016);
nor U11367 (N_11367,N_11010,N_11169);
and U11368 (N_11368,N_11011,N_11149);
xnor U11369 (N_11369,N_11155,N_11076);
or U11370 (N_11370,N_11073,N_11095);
or U11371 (N_11371,N_11171,N_11161);
nor U11372 (N_11372,N_11107,N_11071);
xor U11373 (N_11373,N_11074,N_11097);
and U11374 (N_11374,N_11113,N_11101);
nand U11375 (N_11375,N_11121,N_11171);
xor U11376 (N_11376,N_11024,N_11127);
nand U11377 (N_11377,N_11166,N_11049);
and U11378 (N_11378,N_11007,N_11145);
and U11379 (N_11379,N_11174,N_11041);
nor U11380 (N_11380,N_11032,N_11194);
nand U11381 (N_11381,N_11077,N_11052);
or U11382 (N_11382,N_11063,N_11141);
nand U11383 (N_11383,N_11004,N_11105);
and U11384 (N_11384,N_11126,N_11026);
nand U11385 (N_11385,N_11002,N_11020);
and U11386 (N_11386,N_11134,N_11051);
nand U11387 (N_11387,N_11184,N_11100);
or U11388 (N_11388,N_11177,N_11006);
nor U11389 (N_11389,N_11179,N_11063);
nor U11390 (N_11390,N_11172,N_11135);
nor U11391 (N_11391,N_11006,N_11102);
or U11392 (N_11392,N_11046,N_11089);
nand U11393 (N_11393,N_11145,N_11077);
or U11394 (N_11394,N_11140,N_11175);
nand U11395 (N_11395,N_11092,N_11030);
nand U11396 (N_11396,N_11038,N_11092);
or U11397 (N_11397,N_11139,N_11188);
nor U11398 (N_11398,N_11129,N_11058);
nor U11399 (N_11399,N_11044,N_11100);
nand U11400 (N_11400,N_11348,N_11307);
nand U11401 (N_11401,N_11395,N_11247);
and U11402 (N_11402,N_11363,N_11210);
nor U11403 (N_11403,N_11254,N_11213);
or U11404 (N_11404,N_11231,N_11337);
nor U11405 (N_11405,N_11344,N_11301);
and U11406 (N_11406,N_11245,N_11288);
nor U11407 (N_11407,N_11379,N_11282);
xor U11408 (N_11408,N_11291,N_11203);
nor U11409 (N_11409,N_11243,N_11289);
or U11410 (N_11410,N_11236,N_11300);
xor U11411 (N_11411,N_11393,N_11362);
or U11412 (N_11412,N_11330,N_11322);
nand U11413 (N_11413,N_11294,N_11341);
nand U11414 (N_11414,N_11279,N_11336);
and U11415 (N_11415,N_11372,N_11350);
and U11416 (N_11416,N_11234,N_11218);
xnor U11417 (N_11417,N_11229,N_11293);
and U11418 (N_11418,N_11326,N_11351);
and U11419 (N_11419,N_11373,N_11280);
and U11420 (N_11420,N_11318,N_11207);
xnor U11421 (N_11421,N_11285,N_11325);
xor U11422 (N_11422,N_11276,N_11292);
xor U11423 (N_11423,N_11262,N_11334);
xnor U11424 (N_11424,N_11239,N_11246);
nor U11425 (N_11425,N_11274,N_11304);
and U11426 (N_11426,N_11399,N_11319);
or U11427 (N_11427,N_11343,N_11267);
xor U11428 (N_11428,N_11224,N_11258);
and U11429 (N_11429,N_11365,N_11283);
and U11430 (N_11430,N_11320,N_11250);
nand U11431 (N_11431,N_11238,N_11369);
or U11432 (N_11432,N_11358,N_11278);
xor U11433 (N_11433,N_11205,N_11221);
nand U11434 (N_11434,N_11271,N_11244);
nor U11435 (N_11435,N_11375,N_11345);
nor U11436 (N_11436,N_11323,N_11390);
xor U11437 (N_11437,N_11383,N_11310);
nor U11438 (N_11438,N_11255,N_11387);
or U11439 (N_11439,N_11211,N_11315);
xor U11440 (N_11440,N_11397,N_11321);
nor U11441 (N_11441,N_11302,N_11342);
xnor U11442 (N_11442,N_11316,N_11331);
or U11443 (N_11443,N_11273,N_11256);
or U11444 (N_11444,N_11349,N_11378);
nand U11445 (N_11445,N_11312,N_11268);
xnor U11446 (N_11446,N_11392,N_11306);
nand U11447 (N_11447,N_11233,N_11385);
nand U11448 (N_11448,N_11257,N_11261);
or U11449 (N_11449,N_11277,N_11396);
or U11450 (N_11450,N_11388,N_11217);
nor U11451 (N_11451,N_11311,N_11209);
nor U11452 (N_11452,N_11297,N_11249);
xnor U11453 (N_11453,N_11225,N_11296);
and U11454 (N_11454,N_11340,N_11228);
nand U11455 (N_11455,N_11286,N_11281);
and U11456 (N_11456,N_11335,N_11241);
nor U11457 (N_11457,N_11370,N_11204);
and U11458 (N_11458,N_11364,N_11398);
xor U11459 (N_11459,N_11368,N_11366);
nor U11460 (N_11460,N_11347,N_11308);
nor U11461 (N_11461,N_11248,N_11382);
xnor U11462 (N_11462,N_11381,N_11242);
or U11463 (N_11463,N_11299,N_11371);
nor U11464 (N_11464,N_11360,N_11214);
or U11465 (N_11465,N_11327,N_11324);
nand U11466 (N_11466,N_11376,N_11338);
or U11467 (N_11467,N_11266,N_11226);
and U11468 (N_11468,N_11269,N_11235);
nor U11469 (N_11469,N_11284,N_11377);
nor U11470 (N_11470,N_11252,N_11290);
or U11471 (N_11471,N_11295,N_11206);
nand U11472 (N_11472,N_11275,N_11272);
nor U11473 (N_11473,N_11216,N_11201);
nand U11474 (N_11474,N_11339,N_11309);
nand U11475 (N_11475,N_11305,N_11263);
xor U11476 (N_11476,N_11223,N_11361);
nand U11477 (N_11477,N_11367,N_11313);
and U11478 (N_11478,N_11394,N_11317);
or U11479 (N_11479,N_11329,N_11219);
xnor U11480 (N_11480,N_11208,N_11240);
nand U11481 (N_11481,N_11380,N_11202);
or U11482 (N_11482,N_11215,N_11353);
xnor U11483 (N_11483,N_11356,N_11303);
nor U11484 (N_11484,N_11260,N_11384);
or U11485 (N_11485,N_11270,N_11332);
nor U11486 (N_11486,N_11265,N_11346);
nor U11487 (N_11487,N_11251,N_11359);
nor U11488 (N_11488,N_11389,N_11230);
nor U11489 (N_11489,N_11259,N_11212);
nand U11490 (N_11490,N_11374,N_11287);
or U11491 (N_11491,N_11352,N_11328);
xnor U11492 (N_11492,N_11333,N_11264);
xor U11493 (N_11493,N_11355,N_11314);
xnor U11494 (N_11494,N_11200,N_11391);
xnor U11495 (N_11495,N_11237,N_11298);
nor U11496 (N_11496,N_11232,N_11357);
or U11497 (N_11497,N_11227,N_11220);
and U11498 (N_11498,N_11354,N_11222);
or U11499 (N_11499,N_11386,N_11253);
nor U11500 (N_11500,N_11227,N_11277);
xnor U11501 (N_11501,N_11365,N_11281);
or U11502 (N_11502,N_11321,N_11389);
nor U11503 (N_11503,N_11361,N_11325);
and U11504 (N_11504,N_11385,N_11377);
and U11505 (N_11505,N_11274,N_11207);
or U11506 (N_11506,N_11216,N_11207);
xor U11507 (N_11507,N_11366,N_11321);
or U11508 (N_11508,N_11232,N_11361);
and U11509 (N_11509,N_11364,N_11240);
xnor U11510 (N_11510,N_11239,N_11356);
or U11511 (N_11511,N_11264,N_11226);
nor U11512 (N_11512,N_11268,N_11218);
nor U11513 (N_11513,N_11289,N_11288);
nor U11514 (N_11514,N_11293,N_11245);
or U11515 (N_11515,N_11241,N_11260);
xor U11516 (N_11516,N_11392,N_11225);
nand U11517 (N_11517,N_11352,N_11295);
nand U11518 (N_11518,N_11386,N_11269);
nor U11519 (N_11519,N_11353,N_11327);
nor U11520 (N_11520,N_11381,N_11247);
and U11521 (N_11521,N_11399,N_11395);
nor U11522 (N_11522,N_11326,N_11346);
and U11523 (N_11523,N_11208,N_11360);
or U11524 (N_11524,N_11303,N_11379);
xor U11525 (N_11525,N_11332,N_11336);
nor U11526 (N_11526,N_11357,N_11231);
nor U11527 (N_11527,N_11353,N_11392);
nor U11528 (N_11528,N_11231,N_11232);
or U11529 (N_11529,N_11356,N_11207);
or U11530 (N_11530,N_11337,N_11323);
nand U11531 (N_11531,N_11355,N_11207);
nor U11532 (N_11532,N_11365,N_11367);
or U11533 (N_11533,N_11359,N_11353);
xnor U11534 (N_11534,N_11275,N_11240);
nor U11535 (N_11535,N_11353,N_11214);
nand U11536 (N_11536,N_11220,N_11267);
nor U11537 (N_11537,N_11375,N_11378);
xor U11538 (N_11538,N_11229,N_11334);
or U11539 (N_11539,N_11298,N_11395);
or U11540 (N_11540,N_11310,N_11273);
and U11541 (N_11541,N_11355,N_11230);
xor U11542 (N_11542,N_11337,N_11211);
xnor U11543 (N_11543,N_11337,N_11311);
xnor U11544 (N_11544,N_11262,N_11364);
and U11545 (N_11545,N_11306,N_11211);
or U11546 (N_11546,N_11350,N_11247);
or U11547 (N_11547,N_11369,N_11226);
or U11548 (N_11548,N_11350,N_11235);
or U11549 (N_11549,N_11386,N_11306);
nor U11550 (N_11550,N_11261,N_11265);
and U11551 (N_11551,N_11250,N_11330);
or U11552 (N_11552,N_11250,N_11298);
and U11553 (N_11553,N_11382,N_11291);
and U11554 (N_11554,N_11245,N_11300);
or U11555 (N_11555,N_11270,N_11296);
or U11556 (N_11556,N_11388,N_11246);
nand U11557 (N_11557,N_11294,N_11228);
nand U11558 (N_11558,N_11244,N_11318);
and U11559 (N_11559,N_11378,N_11353);
and U11560 (N_11560,N_11205,N_11278);
and U11561 (N_11561,N_11295,N_11343);
xnor U11562 (N_11562,N_11299,N_11353);
xnor U11563 (N_11563,N_11380,N_11310);
xnor U11564 (N_11564,N_11311,N_11376);
nand U11565 (N_11565,N_11393,N_11246);
xor U11566 (N_11566,N_11212,N_11242);
or U11567 (N_11567,N_11384,N_11215);
and U11568 (N_11568,N_11266,N_11345);
and U11569 (N_11569,N_11348,N_11326);
nor U11570 (N_11570,N_11311,N_11314);
and U11571 (N_11571,N_11233,N_11398);
nor U11572 (N_11572,N_11266,N_11309);
or U11573 (N_11573,N_11316,N_11283);
or U11574 (N_11574,N_11203,N_11339);
or U11575 (N_11575,N_11290,N_11291);
nand U11576 (N_11576,N_11317,N_11327);
and U11577 (N_11577,N_11249,N_11336);
nor U11578 (N_11578,N_11239,N_11269);
and U11579 (N_11579,N_11251,N_11349);
nor U11580 (N_11580,N_11340,N_11265);
nor U11581 (N_11581,N_11272,N_11373);
nor U11582 (N_11582,N_11262,N_11345);
and U11583 (N_11583,N_11309,N_11249);
nor U11584 (N_11584,N_11331,N_11368);
or U11585 (N_11585,N_11390,N_11228);
xnor U11586 (N_11586,N_11205,N_11327);
or U11587 (N_11587,N_11376,N_11382);
nand U11588 (N_11588,N_11253,N_11255);
xor U11589 (N_11589,N_11296,N_11272);
xor U11590 (N_11590,N_11243,N_11325);
or U11591 (N_11591,N_11331,N_11273);
or U11592 (N_11592,N_11382,N_11300);
xor U11593 (N_11593,N_11380,N_11231);
nand U11594 (N_11594,N_11207,N_11283);
xor U11595 (N_11595,N_11317,N_11218);
nor U11596 (N_11596,N_11382,N_11318);
and U11597 (N_11597,N_11290,N_11399);
or U11598 (N_11598,N_11261,N_11287);
xor U11599 (N_11599,N_11253,N_11338);
and U11600 (N_11600,N_11467,N_11496);
and U11601 (N_11601,N_11538,N_11477);
and U11602 (N_11602,N_11573,N_11508);
nand U11603 (N_11603,N_11544,N_11562);
nand U11604 (N_11604,N_11570,N_11531);
nand U11605 (N_11605,N_11439,N_11561);
nand U11606 (N_11606,N_11501,N_11539);
nor U11607 (N_11607,N_11493,N_11429);
and U11608 (N_11608,N_11553,N_11437);
nor U11609 (N_11609,N_11524,N_11404);
nor U11610 (N_11610,N_11590,N_11465);
nor U11611 (N_11611,N_11489,N_11475);
or U11612 (N_11612,N_11588,N_11441);
or U11613 (N_11613,N_11457,N_11476);
nand U11614 (N_11614,N_11438,N_11547);
xor U11615 (N_11615,N_11402,N_11462);
xnor U11616 (N_11616,N_11479,N_11537);
and U11617 (N_11617,N_11409,N_11517);
xnor U11618 (N_11618,N_11578,N_11579);
xnor U11619 (N_11619,N_11571,N_11411);
xor U11620 (N_11620,N_11415,N_11400);
or U11621 (N_11621,N_11416,N_11559);
nor U11622 (N_11622,N_11473,N_11596);
nand U11623 (N_11623,N_11463,N_11581);
nor U11624 (N_11624,N_11526,N_11456);
xor U11625 (N_11625,N_11563,N_11480);
nand U11626 (N_11626,N_11403,N_11490);
nor U11627 (N_11627,N_11474,N_11454);
nand U11628 (N_11628,N_11512,N_11527);
xor U11629 (N_11629,N_11426,N_11583);
nor U11630 (N_11630,N_11491,N_11565);
nand U11631 (N_11631,N_11460,N_11428);
or U11632 (N_11632,N_11558,N_11498);
and U11633 (N_11633,N_11497,N_11525);
nand U11634 (N_11634,N_11468,N_11481);
or U11635 (N_11635,N_11566,N_11568);
nand U11636 (N_11636,N_11423,N_11500);
nor U11637 (N_11637,N_11452,N_11422);
xor U11638 (N_11638,N_11433,N_11458);
nand U11639 (N_11639,N_11587,N_11495);
nor U11640 (N_11640,N_11412,N_11413);
and U11641 (N_11641,N_11552,N_11466);
and U11642 (N_11642,N_11407,N_11599);
or U11643 (N_11643,N_11431,N_11430);
xnor U11644 (N_11644,N_11436,N_11488);
nor U11645 (N_11645,N_11516,N_11446);
nand U11646 (N_11646,N_11520,N_11405);
and U11647 (N_11647,N_11542,N_11471);
xnor U11648 (N_11648,N_11515,N_11591);
nand U11649 (N_11649,N_11518,N_11469);
xor U11650 (N_11650,N_11546,N_11556);
or U11651 (N_11651,N_11507,N_11574);
and U11652 (N_11652,N_11521,N_11577);
or U11653 (N_11653,N_11464,N_11504);
and U11654 (N_11654,N_11549,N_11576);
nand U11655 (N_11655,N_11593,N_11505);
nand U11656 (N_11656,N_11519,N_11470);
nand U11657 (N_11657,N_11408,N_11486);
nor U11658 (N_11658,N_11483,N_11580);
nor U11659 (N_11659,N_11447,N_11595);
and U11660 (N_11660,N_11472,N_11543);
xor U11661 (N_11661,N_11503,N_11540);
nor U11662 (N_11662,N_11410,N_11592);
xor U11663 (N_11663,N_11586,N_11582);
and U11664 (N_11664,N_11510,N_11449);
nand U11665 (N_11665,N_11494,N_11557);
and U11666 (N_11666,N_11487,N_11424);
or U11667 (N_11667,N_11522,N_11451);
and U11668 (N_11668,N_11584,N_11535);
or U11669 (N_11669,N_11594,N_11482);
nor U11670 (N_11670,N_11461,N_11529);
xor U11671 (N_11671,N_11567,N_11511);
and U11672 (N_11672,N_11548,N_11550);
and U11673 (N_11673,N_11509,N_11598);
nand U11674 (N_11674,N_11414,N_11506);
nor U11675 (N_11675,N_11545,N_11406);
and U11676 (N_11676,N_11432,N_11523);
nor U11677 (N_11677,N_11585,N_11421);
or U11678 (N_11678,N_11445,N_11569);
and U11679 (N_11679,N_11575,N_11541);
or U11680 (N_11680,N_11555,N_11533);
nor U11681 (N_11681,N_11418,N_11443);
nand U11682 (N_11682,N_11453,N_11532);
nor U11683 (N_11683,N_11513,N_11442);
xnor U11684 (N_11684,N_11551,N_11589);
xor U11685 (N_11685,N_11440,N_11530);
nor U11686 (N_11686,N_11420,N_11572);
xnor U11687 (N_11687,N_11560,N_11478);
nor U11688 (N_11688,N_11554,N_11435);
and U11689 (N_11689,N_11401,N_11502);
or U11690 (N_11690,N_11564,N_11528);
xnor U11691 (N_11691,N_11434,N_11499);
nor U11692 (N_11692,N_11597,N_11450);
nand U11693 (N_11693,N_11536,N_11417);
or U11694 (N_11694,N_11534,N_11492);
and U11695 (N_11695,N_11425,N_11514);
xor U11696 (N_11696,N_11427,N_11444);
nor U11697 (N_11697,N_11485,N_11459);
nand U11698 (N_11698,N_11419,N_11484);
xor U11699 (N_11699,N_11455,N_11448);
xor U11700 (N_11700,N_11462,N_11555);
nand U11701 (N_11701,N_11596,N_11447);
and U11702 (N_11702,N_11518,N_11478);
or U11703 (N_11703,N_11518,N_11579);
or U11704 (N_11704,N_11522,N_11595);
nand U11705 (N_11705,N_11488,N_11562);
xor U11706 (N_11706,N_11578,N_11415);
xor U11707 (N_11707,N_11517,N_11542);
and U11708 (N_11708,N_11498,N_11490);
nand U11709 (N_11709,N_11437,N_11463);
nand U11710 (N_11710,N_11568,N_11579);
or U11711 (N_11711,N_11577,N_11535);
or U11712 (N_11712,N_11577,N_11424);
and U11713 (N_11713,N_11553,N_11506);
nor U11714 (N_11714,N_11516,N_11543);
and U11715 (N_11715,N_11403,N_11492);
nand U11716 (N_11716,N_11429,N_11454);
and U11717 (N_11717,N_11525,N_11540);
nand U11718 (N_11718,N_11532,N_11550);
xnor U11719 (N_11719,N_11400,N_11451);
xor U11720 (N_11720,N_11582,N_11513);
xor U11721 (N_11721,N_11471,N_11547);
and U11722 (N_11722,N_11506,N_11453);
nand U11723 (N_11723,N_11561,N_11521);
nor U11724 (N_11724,N_11426,N_11511);
xor U11725 (N_11725,N_11470,N_11509);
nor U11726 (N_11726,N_11547,N_11475);
xor U11727 (N_11727,N_11538,N_11555);
xnor U11728 (N_11728,N_11567,N_11480);
xnor U11729 (N_11729,N_11599,N_11513);
xor U11730 (N_11730,N_11504,N_11463);
and U11731 (N_11731,N_11413,N_11411);
nor U11732 (N_11732,N_11434,N_11462);
xnor U11733 (N_11733,N_11419,N_11503);
nor U11734 (N_11734,N_11428,N_11586);
nand U11735 (N_11735,N_11460,N_11484);
and U11736 (N_11736,N_11432,N_11581);
or U11737 (N_11737,N_11521,N_11535);
xor U11738 (N_11738,N_11521,N_11416);
and U11739 (N_11739,N_11429,N_11517);
or U11740 (N_11740,N_11467,N_11502);
xnor U11741 (N_11741,N_11527,N_11479);
xnor U11742 (N_11742,N_11452,N_11527);
xnor U11743 (N_11743,N_11501,N_11400);
nand U11744 (N_11744,N_11519,N_11513);
nor U11745 (N_11745,N_11512,N_11428);
and U11746 (N_11746,N_11429,N_11489);
or U11747 (N_11747,N_11468,N_11466);
nor U11748 (N_11748,N_11400,N_11583);
nand U11749 (N_11749,N_11462,N_11534);
xnor U11750 (N_11750,N_11543,N_11523);
nor U11751 (N_11751,N_11504,N_11569);
and U11752 (N_11752,N_11574,N_11409);
xnor U11753 (N_11753,N_11538,N_11458);
nand U11754 (N_11754,N_11453,N_11543);
nand U11755 (N_11755,N_11548,N_11523);
nand U11756 (N_11756,N_11503,N_11597);
or U11757 (N_11757,N_11434,N_11410);
nor U11758 (N_11758,N_11456,N_11477);
xnor U11759 (N_11759,N_11572,N_11495);
nand U11760 (N_11760,N_11492,N_11564);
or U11761 (N_11761,N_11574,N_11510);
xnor U11762 (N_11762,N_11539,N_11484);
or U11763 (N_11763,N_11592,N_11531);
and U11764 (N_11764,N_11482,N_11522);
or U11765 (N_11765,N_11566,N_11401);
xor U11766 (N_11766,N_11409,N_11500);
nand U11767 (N_11767,N_11451,N_11574);
or U11768 (N_11768,N_11458,N_11568);
nor U11769 (N_11769,N_11520,N_11489);
or U11770 (N_11770,N_11578,N_11484);
nor U11771 (N_11771,N_11459,N_11553);
and U11772 (N_11772,N_11536,N_11432);
or U11773 (N_11773,N_11498,N_11517);
and U11774 (N_11774,N_11515,N_11472);
nand U11775 (N_11775,N_11536,N_11555);
and U11776 (N_11776,N_11464,N_11596);
nand U11777 (N_11777,N_11576,N_11592);
or U11778 (N_11778,N_11459,N_11435);
xnor U11779 (N_11779,N_11418,N_11413);
xnor U11780 (N_11780,N_11541,N_11587);
or U11781 (N_11781,N_11585,N_11560);
or U11782 (N_11782,N_11595,N_11557);
nor U11783 (N_11783,N_11492,N_11567);
and U11784 (N_11784,N_11475,N_11578);
nand U11785 (N_11785,N_11455,N_11493);
or U11786 (N_11786,N_11416,N_11567);
xnor U11787 (N_11787,N_11455,N_11472);
xor U11788 (N_11788,N_11517,N_11422);
nand U11789 (N_11789,N_11556,N_11415);
and U11790 (N_11790,N_11455,N_11505);
nor U11791 (N_11791,N_11422,N_11473);
nor U11792 (N_11792,N_11556,N_11460);
or U11793 (N_11793,N_11448,N_11597);
and U11794 (N_11794,N_11526,N_11572);
nor U11795 (N_11795,N_11483,N_11539);
or U11796 (N_11796,N_11530,N_11420);
or U11797 (N_11797,N_11544,N_11522);
xor U11798 (N_11798,N_11455,N_11443);
nor U11799 (N_11799,N_11441,N_11409);
and U11800 (N_11800,N_11727,N_11771);
and U11801 (N_11801,N_11655,N_11627);
xor U11802 (N_11802,N_11671,N_11620);
xor U11803 (N_11803,N_11795,N_11675);
and U11804 (N_11804,N_11613,N_11626);
nand U11805 (N_11805,N_11633,N_11789);
and U11806 (N_11806,N_11700,N_11780);
nand U11807 (N_11807,N_11615,N_11657);
xor U11808 (N_11808,N_11720,N_11665);
xor U11809 (N_11809,N_11604,N_11723);
nor U11810 (N_11810,N_11611,N_11709);
xor U11811 (N_11811,N_11725,N_11710);
xnor U11812 (N_11812,N_11691,N_11798);
xor U11813 (N_11813,N_11608,N_11659);
xnor U11814 (N_11814,N_11638,N_11707);
or U11815 (N_11815,N_11740,N_11708);
nor U11816 (N_11816,N_11678,N_11742);
nor U11817 (N_11817,N_11670,N_11612);
and U11818 (N_11818,N_11667,N_11622);
xnor U11819 (N_11819,N_11746,N_11763);
or U11820 (N_11820,N_11760,N_11761);
xnor U11821 (N_11821,N_11651,N_11792);
or U11822 (N_11822,N_11787,N_11619);
nor U11823 (N_11823,N_11684,N_11734);
nor U11824 (N_11824,N_11751,N_11722);
or U11825 (N_11825,N_11628,N_11681);
nor U11826 (N_11826,N_11730,N_11753);
nor U11827 (N_11827,N_11766,N_11649);
nor U11828 (N_11828,N_11768,N_11656);
nand U11829 (N_11829,N_11685,N_11729);
nand U11830 (N_11830,N_11756,N_11762);
nand U11831 (N_11831,N_11704,N_11791);
xnor U11832 (N_11832,N_11703,N_11648);
and U11833 (N_11833,N_11603,N_11694);
nor U11834 (N_11834,N_11717,N_11646);
and U11835 (N_11835,N_11636,N_11785);
nand U11836 (N_11836,N_11640,N_11706);
or U11837 (N_11837,N_11643,N_11774);
and U11838 (N_11838,N_11769,N_11669);
xnor U11839 (N_11839,N_11793,N_11645);
nand U11840 (N_11840,N_11777,N_11772);
nand U11841 (N_11841,N_11737,N_11690);
nor U11842 (N_11842,N_11759,N_11617);
and U11843 (N_11843,N_11660,N_11765);
or U11844 (N_11844,N_11702,N_11750);
nor U11845 (N_11845,N_11697,N_11739);
and U11846 (N_11846,N_11757,N_11668);
xnor U11847 (N_11847,N_11610,N_11716);
and U11848 (N_11848,N_11754,N_11601);
and U11849 (N_11849,N_11719,N_11618);
and U11850 (N_11850,N_11712,N_11693);
and U11851 (N_11851,N_11755,N_11606);
nand U11852 (N_11852,N_11621,N_11688);
nand U11853 (N_11853,N_11600,N_11650);
nor U11854 (N_11854,N_11713,N_11642);
nor U11855 (N_11855,N_11796,N_11732);
nor U11856 (N_11856,N_11682,N_11733);
xnor U11857 (N_11857,N_11758,N_11749);
nand U11858 (N_11858,N_11797,N_11687);
nor U11859 (N_11859,N_11711,N_11647);
and U11860 (N_11860,N_11614,N_11724);
or U11861 (N_11861,N_11705,N_11699);
nor U11862 (N_11862,N_11653,N_11654);
or U11863 (N_11863,N_11767,N_11676);
xnor U11864 (N_11864,N_11752,N_11764);
nand U11865 (N_11865,N_11673,N_11698);
nor U11866 (N_11866,N_11663,N_11701);
nor U11867 (N_11867,N_11661,N_11728);
nand U11868 (N_11868,N_11624,N_11686);
nor U11869 (N_11869,N_11639,N_11794);
nor U11870 (N_11870,N_11743,N_11788);
and U11871 (N_11871,N_11662,N_11784);
nand U11872 (N_11872,N_11629,N_11731);
xor U11873 (N_11873,N_11747,N_11634);
nand U11874 (N_11874,N_11602,N_11770);
or U11875 (N_11875,N_11666,N_11605);
nor U11876 (N_11876,N_11721,N_11736);
xnor U11877 (N_11877,N_11741,N_11695);
nand U11878 (N_11878,N_11745,N_11748);
xnor U11879 (N_11879,N_11738,N_11609);
or U11880 (N_11880,N_11683,N_11637);
and U11881 (N_11881,N_11631,N_11689);
nand U11882 (N_11882,N_11632,N_11718);
and U11883 (N_11883,N_11692,N_11607);
or U11884 (N_11884,N_11625,N_11744);
or U11885 (N_11885,N_11714,N_11781);
or U11886 (N_11886,N_11779,N_11635);
nor U11887 (N_11887,N_11790,N_11644);
nor U11888 (N_11888,N_11658,N_11786);
or U11889 (N_11889,N_11775,N_11623);
xnor U11890 (N_11890,N_11773,N_11677);
nor U11891 (N_11891,N_11696,N_11616);
xor U11892 (N_11892,N_11664,N_11776);
nor U11893 (N_11893,N_11735,N_11630);
or U11894 (N_11894,N_11652,N_11674);
or U11895 (N_11895,N_11641,N_11726);
or U11896 (N_11896,N_11783,N_11782);
nand U11897 (N_11897,N_11778,N_11679);
or U11898 (N_11898,N_11680,N_11715);
nor U11899 (N_11899,N_11672,N_11799);
xor U11900 (N_11900,N_11656,N_11649);
nor U11901 (N_11901,N_11651,N_11752);
or U11902 (N_11902,N_11653,N_11603);
nor U11903 (N_11903,N_11706,N_11629);
or U11904 (N_11904,N_11704,N_11620);
nor U11905 (N_11905,N_11633,N_11750);
and U11906 (N_11906,N_11705,N_11749);
or U11907 (N_11907,N_11761,N_11735);
nand U11908 (N_11908,N_11661,N_11704);
xnor U11909 (N_11909,N_11756,N_11728);
xor U11910 (N_11910,N_11697,N_11616);
and U11911 (N_11911,N_11726,N_11609);
and U11912 (N_11912,N_11788,N_11701);
nand U11913 (N_11913,N_11768,N_11795);
or U11914 (N_11914,N_11649,N_11622);
nand U11915 (N_11915,N_11786,N_11748);
and U11916 (N_11916,N_11609,N_11787);
nor U11917 (N_11917,N_11688,N_11619);
and U11918 (N_11918,N_11657,N_11677);
or U11919 (N_11919,N_11754,N_11731);
and U11920 (N_11920,N_11735,N_11657);
nor U11921 (N_11921,N_11693,N_11700);
nand U11922 (N_11922,N_11608,N_11689);
nor U11923 (N_11923,N_11725,N_11643);
xnor U11924 (N_11924,N_11775,N_11765);
nor U11925 (N_11925,N_11625,N_11642);
or U11926 (N_11926,N_11632,N_11767);
or U11927 (N_11927,N_11630,N_11792);
and U11928 (N_11928,N_11688,N_11702);
or U11929 (N_11929,N_11730,N_11774);
nand U11930 (N_11930,N_11729,N_11762);
xor U11931 (N_11931,N_11759,N_11796);
xor U11932 (N_11932,N_11793,N_11792);
nand U11933 (N_11933,N_11787,N_11732);
nor U11934 (N_11934,N_11740,N_11687);
or U11935 (N_11935,N_11775,N_11794);
nand U11936 (N_11936,N_11711,N_11627);
nor U11937 (N_11937,N_11793,N_11739);
and U11938 (N_11938,N_11632,N_11704);
xnor U11939 (N_11939,N_11610,N_11693);
nor U11940 (N_11940,N_11651,N_11646);
nand U11941 (N_11941,N_11666,N_11610);
nor U11942 (N_11942,N_11629,N_11762);
and U11943 (N_11943,N_11683,N_11793);
nor U11944 (N_11944,N_11763,N_11672);
nand U11945 (N_11945,N_11794,N_11606);
and U11946 (N_11946,N_11601,N_11795);
nand U11947 (N_11947,N_11775,N_11700);
or U11948 (N_11948,N_11626,N_11715);
or U11949 (N_11949,N_11722,N_11617);
and U11950 (N_11950,N_11771,N_11728);
xnor U11951 (N_11951,N_11799,N_11753);
nor U11952 (N_11952,N_11615,N_11740);
nand U11953 (N_11953,N_11766,N_11632);
nand U11954 (N_11954,N_11692,N_11699);
and U11955 (N_11955,N_11605,N_11753);
or U11956 (N_11956,N_11720,N_11755);
nor U11957 (N_11957,N_11659,N_11686);
nand U11958 (N_11958,N_11752,N_11796);
or U11959 (N_11959,N_11623,N_11798);
or U11960 (N_11960,N_11729,N_11653);
or U11961 (N_11961,N_11691,N_11632);
xor U11962 (N_11962,N_11644,N_11793);
and U11963 (N_11963,N_11706,N_11736);
or U11964 (N_11964,N_11609,N_11661);
nand U11965 (N_11965,N_11778,N_11628);
or U11966 (N_11966,N_11717,N_11723);
or U11967 (N_11967,N_11767,N_11639);
xor U11968 (N_11968,N_11621,N_11794);
and U11969 (N_11969,N_11796,N_11717);
nor U11970 (N_11970,N_11760,N_11669);
or U11971 (N_11971,N_11662,N_11722);
nand U11972 (N_11972,N_11720,N_11630);
and U11973 (N_11973,N_11689,N_11624);
and U11974 (N_11974,N_11605,N_11641);
and U11975 (N_11975,N_11768,N_11788);
or U11976 (N_11976,N_11709,N_11627);
xnor U11977 (N_11977,N_11637,N_11634);
and U11978 (N_11978,N_11783,N_11725);
nor U11979 (N_11979,N_11743,N_11602);
or U11980 (N_11980,N_11708,N_11771);
nand U11981 (N_11981,N_11763,N_11709);
xnor U11982 (N_11982,N_11787,N_11630);
or U11983 (N_11983,N_11710,N_11715);
or U11984 (N_11984,N_11737,N_11756);
xnor U11985 (N_11985,N_11796,N_11626);
nor U11986 (N_11986,N_11618,N_11602);
nand U11987 (N_11987,N_11731,N_11626);
nand U11988 (N_11988,N_11728,N_11785);
xnor U11989 (N_11989,N_11787,N_11686);
xnor U11990 (N_11990,N_11643,N_11775);
xnor U11991 (N_11991,N_11672,N_11655);
nand U11992 (N_11992,N_11767,N_11624);
xnor U11993 (N_11993,N_11714,N_11678);
xor U11994 (N_11994,N_11665,N_11785);
xor U11995 (N_11995,N_11739,N_11789);
nand U11996 (N_11996,N_11636,N_11633);
and U11997 (N_11997,N_11638,N_11672);
or U11998 (N_11998,N_11736,N_11771);
xor U11999 (N_11999,N_11662,N_11768);
xor U12000 (N_12000,N_11868,N_11971);
nor U12001 (N_12001,N_11934,N_11851);
or U12002 (N_12002,N_11828,N_11817);
or U12003 (N_12003,N_11973,N_11922);
nor U12004 (N_12004,N_11967,N_11872);
nor U12005 (N_12005,N_11949,N_11824);
nand U12006 (N_12006,N_11902,N_11923);
and U12007 (N_12007,N_11816,N_11829);
or U12008 (N_12008,N_11867,N_11838);
and U12009 (N_12009,N_11890,N_11980);
and U12010 (N_12010,N_11880,N_11858);
xor U12011 (N_12011,N_11871,N_11970);
nand U12012 (N_12012,N_11881,N_11836);
and U12013 (N_12013,N_11945,N_11944);
xnor U12014 (N_12014,N_11981,N_11908);
nor U12015 (N_12015,N_11834,N_11889);
xnor U12016 (N_12016,N_11946,N_11958);
and U12017 (N_12017,N_11900,N_11933);
nor U12018 (N_12018,N_11942,N_11917);
nor U12019 (N_12019,N_11972,N_11940);
nand U12020 (N_12020,N_11879,N_11861);
xnor U12021 (N_12021,N_11840,N_11921);
and U12022 (N_12022,N_11991,N_11926);
or U12023 (N_12023,N_11911,N_11813);
and U12024 (N_12024,N_11863,N_11935);
and U12025 (N_12025,N_11976,N_11957);
and U12026 (N_12026,N_11882,N_11826);
and U12027 (N_12027,N_11894,N_11930);
nand U12028 (N_12028,N_11956,N_11906);
or U12029 (N_12029,N_11801,N_11918);
nand U12030 (N_12030,N_11877,N_11909);
xor U12031 (N_12031,N_11805,N_11939);
or U12032 (N_12032,N_11975,N_11857);
nor U12033 (N_12033,N_11913,N_11999);
or U12034 (N_12034,N_11866,N_11915);
or U12035 (N_12035,N_11994,N_11819);
xor U12036 (N_12036,N_11842,N_11837);
and U12037 (N_12037,N_11962,N_11883);
and U12038 (N_12038,N_11878,N_11959);
and U12039 (N_12039,N_11827,N_11961);
xnor U12040 (N_12040,N_11841,N_11952);
xor U12041 (N_12041,N_11924,N_11986);
nor U12042 (N_12042,N_11941,N_11912);
or U12043 (N_12043,N_11993,N_11870);
nand U12044 (N_12044,N_11804,N_11873);
and U12045 (N_12045,N_11865,N_11964);
nand U12046 (N_12046,N_11891,N_11965);
xnor U12047 (N_12047,N_11850,N_11974);
xnor U12048 (N_12048,N_11925,N_11963);
nand U12049 (N_12049,N_11953,N_11920);
and U12050 (N_12050,N_11807,N_11904);
or U12051 (N_12051,N_11950,N_11888);
nor U12052 (N_12052,N_11914,N_11886);
nand U12053 (N_12053,N_11892,N_11899);
and U12054 (N_12054,N_11853,N_11839);
nor U12055 (N_12055,N_11802,N_11947);
nand U12056 (N_12056,N_11910,N_11860);
xnor U12057 (N_12057,N_11822,N_11955);
xor U12058 (N_12058,N_11985,N_11916);
and U12059 (N_12059,N_11896,N_11927);
xor U12060 (N_12060,N_11905,N_11898);
nand U12061 (N_12061,N_11897,N_11808);
nand U12062 (N_12062,N_11830,N_11951);
or U12063 (N_12063,N_11854,N_11814);
xnor U12064 (N_12064,N_11876,N_11997);
nand U12065 (N_12065,N_11812,N_11928);
or U12066 (N_12066,N_11978,N_11845);
xnor U12067 (N_12067,N_11979,N_11869);
and U12068 (N_12068,N_11983,N_11843);
and U12069 (N_12069,N_11938,N_11966);
or U12070 (N_12070,N_11864,N_11844);
or U12071 (N_12071,N_11856,N_11989);
and U12072 (N_12072,N_11874,N_11936);
and U12073 (N_12073,N_11875,N_11847);
or U12074 (N_12074,N_11806,N_11982);
xnor U12075 (N_12075,N_11893,N_11821);
nor U12076 (N_12076,N_11948,N_11996);
nand U12077 (N_12077,N_11992,N_11884);
xnor U12078 (N_12078,N_11818,N_11852);
xnor U12079 (N_12079,N_11895,N_11803);
xor U12080 (N_12080,N_11815,N_11835);
nor U12081 (N_12081,N_11937,N_11987);
nor U12082 (N_12082,N_11998,N_11988);
nor U12083 (N_12083,N_11820,N_11990);
xnor U12084 (N_12084,N_11929,N_11907);
nor U12085 (N_12085,N_11919,N_11885);
or U12086 (N_12086,N_11977,N_11800);
nand U12087 (N_12087,N_11846,N_11832);
and U12088 (N_12088,N_11825,N_11811);
nand U12089 (N_12089,N_11901,N_11831);
and U12090 (N_12090,N_11931,N_11862);
nor U12091 (N_12091,N_11968,N_11960);
or U12092 (N_12092,N_11855,N_11859);
or U12093 (N_12093,N_11995,N_11848);
and U12094 (N_12094,N_11809,N_11833);
nand U12095 (N_12095,N_11849,N_11984);
xnor U12096 (N_12096,N_11943,N_11969);
nor U12097 (N_12097,N_11810,N_11903);
xor U12098 (N_12098,N_11887,N_11823);
or U12099 (N_12099,N_11932,N_11954);
xnor U12100 (N_12100,N_11892,N_11875);
xor U12101 (N_12101,N_11851,N_11891);
xnor U12102 (N_12102,N_11965,N_11937);
nand U12103 (N_12103,N_11900,N_11881);
and U12104 (N_12104,N_11915,N_11958);
nor U12105 (N_12105,N_11811,N_11833);
and U12106 (N_12106,N_11814,N_11951);
nand U12107 (N_12107,N_11817,N_11936);
xnor U12108 (N_12108,N_11911,N_11987);
and U12109 (N_12109,N_11801,N_11929);
nor U12110 (N_12110,N_11959,N_11802);
nor U12111 (N_12111,N_11966,N_11939);
or U12112 (N_12112,N_11817,N_11860);
xor U12113 (N_12113,N_11922,N_11961);
xnor U12114 (N_12114,N_11986,N_11962);
nand U12115 (N_12115,N_11819,N_11962);
or U12116 (N_12116,N_11926,N_11833);
and U12117 (N_12117,N_11811,N_11952);
and U12118 (N_12118,N_11989,N_11863);
nand U12119 (N_12119,N_11977,N_11938);
and U12120 (N_12120,N_11906,N_11937);
xnor U12121 (N_12121,N_11978,N_11828);
xnor U12122 (N_12122,N_11928,N_11862);
nand U12123 (N_12123,N_11978,N_11836);
and U12124 (N_12124,N_11994,N_11979);
nor U12125 (N_12125,N_11859,N_11958);
xnor U12126 (N_12126,N_11807,N_11931);
xnor U12127 (N_12127,N_11956,N_11948);
or U12128 (N_12128,N_11962,N_11890);
xor U12129 (N_12129,N_11918,N_11852);
nor U12130 (N_12130,N_11934,N_11820);
and U12131 (N_12131,N_11902,N_11872);
nor U12132 (N_12132,N_11966,N_11948);
and U12133 (N_12133,N_11903,N_11866);
and U12134 (N_12134,N_11931,N_11996);
or U12135 (N_12135,N_11963,N_11954);
or U12136 (N_12136,N_11870,N_11856);
nand U12137 (N_12137,N_11957,N_11869);
nand U12138 (N_12138,N_11927,N_11989);
nor U12139 (N_12139,N_11975,N_11865);
or U12140 (N_12140,N_11853,N_11855);
and U12141 (N_12141,N_11872,N_11880);
nor U12142 (N_12142,N_11834,N_11975);
and U12143 (N_12143,N_11801,N_11856);
or U12144 (N_12144,N_11870,N_11992);
or U12145 (N_12145,N_11911,N_11867);
nor U12146 (N_12146,N_11825,N_11917);
nand U12147 (N_12147,N_11801,N_11992);
xnor U12148 (N_12148,N_11836,N_11988);
and U12149 (N_12149,N_11928,N_11808);
or U12150 (N_12150,N_11928,N_11996);
and U12151 (N_12151,N_11924,N_11922);
nor U12152 (N_12152,N_11893,N_11968);
xor U12153 (N_12153,N_11958,N_11868);
or U12154 (N_12154,N_11897,N_11932);
nand U12155 (N_12155,N_11941,N_11889);
and U12156 (N_12156,N_11942,N_11842);
nor U12157 (N_12157,N_11927,N_11895);
nor U12158 (N_12158,N_11997,N_11924);
nor U12159 (N_12159,N_11998,N_11847);
nand U12160 (N_12160,N_11883,N_11907);
xnor U12161 (N_12161,N_11941,N_11848);
and U12162 (N_12162,N_11937,N_11857);
nor U12163 (N_12163,N_11943,N_11830);
nor U12164 (N_12164,N_11854,N_11865);
and U12165 (N_12165,N_11956,N_11844);
or U12166 (N_12166,N_11826,N_11995);
or U12167 (N_12167,N_11919,N_11871);
nor U12168 (N_12168,N_11863,N_11943);
nor U12169 (N_12169,N_11841,N_11806);
xnor U12170 (N_12170,N_11828,N_11884);
nand U12171 (N_12171,N_11951,N_11802);
xnor U12172 (N_12172,N_11873,N_11999);
and U12173 (N_12173,N_11975,N_11875);
and U12174 (N_12174,N_11813,N_11933);
xnor U12175 (N_12175,N_11958,N_11990);
nand U12176 (N_12176,N_11861,N_11823);
or U12177 (N_12177,N_11910,N_11999);
xnor U12178 (N_12178,N_11888,N_11899);
nor U12179 (N_12179,N_11805,N_11811);
xor U12180 (N_12180,N_11930,N_11992);
nand U12181 (N_12181,N_11821,N_11881);
nand U12182 (N_12182,N_11812,N_11967);
and U12183 (N_12183,N_11833,N_11976);
nand U12184 (N_12184,N_11999,N_11979);
nand U12185 (N_12185,N_11844,N_11940);
nand U12186 (N_12186,N_11895,N_11869);
and U12187 (N_12187,N_11881,N_11898);
nor U12188 (N_12188,N_11863,N_11900);
xnor U12189 (N_12189,N_11878,N_11991);
xor U12190 (N_12190,N_11923,N_11994);
nand U12191 (N_12191,N_11820,N_11871);
nor U12192 (N_12192,N_11928,N_11921);
nor U12193 (N_12193,N_11835,N_11964);
and U12194 (N_12194,N_11845,N_11889);
nor U12195 (N_12195,N_11904,N_11924);
and U12196 (N_12196,N_11959,N_11833);
nand U12197 (N_12197,N_11907,N_11997);
and U12198 (N_12198,N_11815,N_11912);
nor U12199 (N_12199,N_11840,N_11987);
and U12200 (N_12200,N_12059,N_12074);
or U12201 (N_12201,N_12139,N_12101);
xor U12202 (N_12202,N_12012,N_12007);
or U12203 (N_12203,N_12022,N_12154);
nor U12204 (N_12204,N_12041,N_12026);
nor U12205 (N_12205,N_12085,N_12162);
xnor U12206 (N_12206,N_12056,N_12018);
and U12207 (N_12207,N_12153,N_12109);
and U12208 (N_12208,N_12047,N_12040);
nor U12209 (N_12209,N_12163,N_12098);
nor U12210 (N_12210,N_12055,N_12020);
xnor U12211 (N_12211,N_12156,N_12144);
nand U12212 (N_12212,N_12019,N_12130);
or U12213 (N_12213,N_12196,N_12184);
or U12214 (N_12214,N_12028,N_12011);
nand U12215 (N_12215,N_12160,N_12181);
xnor U12216 (N_12216,N_12077,N_12089);
nor U12217 (N_12217,N_12037,N_12029);
nor U12218 (N_12218,N_12158,N_12097);
or U12219 (N_12219,N_12152,N_12024);
xor U12220 (N_12220,N_12048,N_12043);
and U12221 (N_12221,N_12188,N_12119);
and U12222 (N_12222,N_12164,N_12129);
and U12223 (N_12223,N_12106,N_12067);
xnor U12224 (N_12224,N_12151,N_12114);
nor U12225 (N_12225,N_12082,N_12124);
and U12226 (N_12226,N_12166,N_12103);
and U12227 (N_12227,N_12083,N_12030);
nor U12228 (N_12228,N_12023,N_12049);
and U12229 (N_12229,N_12009,N_12167);
nor U12230 (N_12230,N_12081,N_12071);
and U12231 (N_12231,N_12112,N_12033);
xnor U12232 (N_12232,N_12175,N_12195);
xor U12233 (N_12233,N_12168,N_12079);
nor U12234 (N_12234,N_12118,N_12187);
nand U12235 (N_12235,N_12004,N_12185);
or U12236 (N_12236,N_12027,N_12104);
and U12237 (N_12237,N_12178,N_12174);
or U12238 (N_12238,N_12076,N_12150);
nand U12239 (N_12239,N_12005,N_12183);
xor U12240 (N_12240,N_12051,N_12165);
or U12241 (N_12241,N_12138,N_12013);
nor U12242 (N_12242,N_12179,N_12133);
xor U12243 (N_12243,N_12094,N_12099);
nand U12244 (N_12244,N_12084,N_12032);
nor U12245 (N_12245,N_12053,N_12116);
and U12246 (N_12246,N_12131,N_12042);
and U12247 (N_12247,N_12021,N_12111);
nor U12248 (N_12248,N_12039,N_12147);
nand U12249 (N_12249,N_12014,N_12117);
nand U12250 (N_12250,N_12031,N_12108);
xnor U12251 (N_12251,N_12177,N_12189);
nor U12252 (N_12252,N_12115,N_12045);
nand U12253 (N_12253,N_12171,N_12137);
and U12254 (N_12254,N_12170,N_12073);
and U12255 (N_12255,N_12063,N_12090);
xor U12256 (N_12256,N_12182,N_12044);
or U12257 (N_12257,N_12062,N_12015);
xnor U12258 (N_12258,N_12198,N_12002);
nand U12259 (N_12259,N_12052,N_12105);
and U12260 (N_12260,N_12149,N_12001);
nor U12261 (N_12261,N_12126,N_12122);
nand U12262 (N_12262,N_12161,N_12064);
nand U12263 (N_12263,N_12121,N_12110);
nor U12264 (N_12264,N_12003,N_12113);
and U12265 (N_12265,N_12006,N_12038);
nand U12266 (N_12266,N_12008,N_12025);
or U12267 (N_12267,N_12146,N_12036);
nand U12268 (N_12268,N_12078,N_12066);
nor U12269 (N_12269,N_12148,N_12194);
nand U12270 (N_12270,N_12191,N_12125);
or U12271 (N_12271,N_12155,N_12128);
and U12272 (N_12272,N_12157,N_12199);
or U12273 (N_12273,N_12169,N_12050);
or U12274 (N_12274,N_12143,N_12069);
nor U12275 (N_12275,N_12134,N_12061);
nor U12276 (N_12276,N_12080,N_12140);
nand U12277 (N_12277,N_12186,N_12075);
and U12278 (N_12278,N_12096,N_12034);
xor U12279 (N_12279,N_12123,N_12159);
and U12280 (N_12280,N_12070,N_12135);
xor U12281 (N_12281,N_12132,N_12010);
and U12282 (N_12282,N_12142,N_12093);
nand U12283 (N_12283,N_12173,N_12046);
nor U12284 (N_12284,N_12060,N_12176);
and U12285 (N_12285,N_12057,N_12087);
xnor U12286 (N_12286,N_12172,N_12102);
and U12287 (N_12287,N_12072,N_12192);
or U12288 (N_12288,N_12068,N_12193);
nand U12289 (N_12289,N_12017,N_12000);
or U12290 (N_12290,N_12091,N_12127);
and U12291 (N_12291,N_12095,N_12065);
and U12292 (N_12292,N_12120,N_12107);
xor U12293 (N_12293,N_12141,N_12180);
and U12294 (N_12294,N_12016,N_12190);
nand U12295 (N_12295,N_12088,N_12100);
or U12296 (N_12296,N_12035,N_12197);
xnor U12297 (N_12297,N_12092,N_12136);
nand U12298 (N_12298,N_12086,N_12145);
nor U12299 (N_12299,N_12054,N_12058);
or U12300 (N_12300,N_12110,N_12016);
or U12301 (N_12301,N_12095,N_12064);
nand U12302 (N_12302,N_12138,N_12146);
or U12303 (N_12303,N_12128,N_12160);
xnor U12304 (N_12304,N_12044,N_12009);
and U12305 (N_12305,N_12147,N_12082);
or U12306 (N_12306,N_12194,N_12032);
xor U12307 (N_12307,N_12149,N_12126);
and U12308 (N_12308,N_12020,N_12009);
xor U12309 (N_12309,N_12122,N_12119);
nand U12310 (N_12310,N_12012,N_12143);
xor U12311 (N_12311,N_12095,N_12108);
xnor U12312 (N_12312,N_12087,N_12193);
nor U12313 (N_12313,N_12087,N_12040);
xor U12314 (N_12314,N_12189,N_12102);
and U12315 (N_12315,N_12050,N_12036);
and U12316 (N_12316,N_12102,N_12005);
nand U12317 (N_12317,N_12046,N_12084);
nor U12318 (N_12318,N_12101,N_12024);
and U12319 (N_12319,N_12094,N_12102);
xor U12320 (N_12320,N_12127,N_12107);
and U12321 (N_12321,N_12056,N_12093);
and U12322 (N_12322,N_12183,N_12009);
nor U12323 (N_12323,N_12139,N_12070);
nand U12324 (N_12324,N_12133,N_12131);
nor U12325 (N_12325,N_12008,N_12173);
nand U12326 (N_12326,N_12034,N_12041);
and U12327 (N_12327,N_12184,N_12034);
and U12328 (N_12328,N_12146,N_12085);
nor U12329 (N_12329,N_12103,N_12146);
or U12330 (N_12330,N_12059,N_12099);
xor U12331 (N_12331,N_12139,N_12103);
nor U12332 (N_12332,N_12192,N_12074);
and U12333 (N_12333,N_12043,N_12183);
nor U12334 (N_12334,N_12118,N_12086);
nand U12335 (N_12335,N_12001,N_12137);
or U12336 (N_12336,N_12142,N_12099);
and U12337 (N_12337,N_12065,N_12043);
xnor U12338 (N_12338,N_12063,N_12052);
and U12339 (N_12339,N_12144,N_12167);
nor U12340 (N_12340,N_12027,N_12011);
xor U12341 (N_12341,N_12073,N_12150);
nand U12342 (N_12342,N_12074,N_12108);
nand U12343 (N_12343,N_12025,N_12190);
nand U12344 (N_12344,N_12105,N_12088);
and U12345 (N_12345,N_12175,N_12129);
or U12346 (N_12346,N_12192,N_12152);
or U12347 (N_12347,N_12007,N_12130);
nand U12348 (N_12348,N_12139,N_12175);
or U12349 (N_12349,N_12079,N_12184);
or U12350 (N_12350,N_12140,N_12090);
or U12351 (N_12351,N_12028,N_12097);
nor U12352 (N_12352,N_12108,N_12092);
nor U12353 (N_12353,N_12071,N_12185);
xor U12354 (N_12354,N_12140,N_12028);
and U12355 (N_12355,N_12156,N_12038);
xor U12356 (N_12356,N_12021,N_12011);
xnor U12357 (N_12357,N_12118,N_12167);
nand U12358 (N_12358,N_12014,N_12157);
nand U12359 (N_12359,N_12194,N_12083);
and U12360 (N_12360,N_12043,N_12109);
nor U12361 (N_12361,N_12007,N_12027);
nor U12362 (N_12362,N_12165,N_12038);
xor U12363 (N_12363,N_12195,N_12032);
nand U12364 (N_12364,N_12047,N_12025);
nor U12365 (N_12365,N_12185,N_12079);
or U12366 (N_12366,N_12034,N_12121);
xnor U12367 (N_12367,N_12112,N_12119);
nor U12368 (N_12368,N_12047,N_12046);
and U12369 (N_12369,N_12029,N_12186);
nor U12370 (N_12370,N_12147,N_12136);
nor U12371 (N_12371,N_12079,N_12044);
xnor U12372 (N_12372,N_12051,N_12008);
xor U12373 (N_12373,N_12089,N_12131);
xor U12374 (N_12374,N_12063,N_12100);
xor U12375 (N_12375,N_12175,N_12120);
and U12376 (N_12376,N_12181,N_12050);
or U12377 (N_12377,N_12161,N_12092);
nor U12378 (N_12378,N_12085,N_12062);
and U12379 (N_12379,N_12195,N_12005);
xor U12380 (N_12380,N_12004,N_12155);
or U12381 (N_12381,N_12040,N_12025);
or U12382 (N_12382,N_12091,N_12001);
and U12383 (N_12383,N_12158,N_12195);
and U12384 (N_12384,N_12075,N_12178);
and U12385 (N_12385,N_12058,N_12002);
nor U12386 (N_12386,N_12078,N_12068);
or U12387 (N_12387,N_12075,N_12152);
xnor U12388 (N_12388,N_12158,N_12009);
nor U12389 (N_12389,N_12158,N_12059);
nand U12390 (N_12390,N_12171,N_12166);
xor U12391 (N_12391,N_12076,N_12173);
and U12392 (N_12392,N_12179,N_12129);
and U12393 (N_12393,N_12090,N_12007);
xnor U12394 (N_12394,N_12063,N_12165);
or U12395 (N_12395,N_12143,N_12059);
and U12396 (N_12396,N_12062,N_12170);
nand U12397 (N_12397,N_12161,N_12164);
and U12398 (N_12398,N_12186,N_12080);
nor U12399 (N_12399,N_12180,N_12167);
and U12400 (N_12400,N_12245,N_12331);
nor U12401 (N_12401,N_12201,N_12215);
xnor U12402 (N_12402,N_12225,N_12309);
and U12403 (N_12403,N_12365,N_12207);
xor U12404 (N_12404,N_12205,N_12249);
nor U12405 (N_12405,N_12327,N_12264);
or U12406 (N_12406,N_12366,N_12325);
and U12407 (N_12407,N_12210,N_12300);
and U12408 (N_12408,N_12364,N_12328);
or U12409 (N_12409,N_12208,N_12272);
nand U12410 (N_12410,N_12346,N_12335);
nand U12411 (N_12411,N_12209,N_12311);
or U12412 (N_12412,N_12271,N_12336);
nor U12413 (N_12413,N_12242,N_12200);
xor U12414 (N_12414,N_12342,N_12322);
and U12415 (N_12415,N_12216,N_12397);
nor U12416 (N_12416,N_12305,N_12258);
nand U12417 (N_12417,N_12363,N_12256);
nor U12418 (N_12418,N_12308,N_12387);
nand U12419 (N_12419,N_12385,N_12319);
nand U12420 (N_12420,N_12394,N_12218);
and U12421 (N_12421,N_12266,N_12273);
nand U12422 (N_12422,N_12312,N_12375);
xnor U12423 (N_12423,N_12368,N_12381);
or U12424 (N_12424,N_12285,N_12231);
nor U12425 (N_12425,N_12203,N_12310);
nand U12426 (N_12426,N_12339,N_12223);
xnor U12427 (N_12427,N_12276,N_12265);
nand U12428 (N_12428,N_12283,N_12240);
nand U12429 (N_12429,N_12262,N_12350);
and U12430 (N_12430,N_12376,N_12287);
nand U12431 (N_12431,N_12292,N_12221);
and U12432 (N_12432,N_12332,N_12263);
nor U12433 (N_12433,N_12257,N_12280);
nor U12434 (N_12434,N_12211,N_12357);
nand U12435 (N_12435,N_12279,N_12326);
nand U12436 (N_12436,N_12274,N_12302);
xnor U12437 (N_12437,N_12399,N_12323);
and U12438 (N_12438,N_12226,N_12389);
nand U12439 (N_12439,N_12284,N_12396);
or U12440 (N_12440,N_12252,N_12289);
or U12441 (N_12441,N_12286,N_12269);
and U12442 (N_12442,N_12329,N_12253);
nand U12443 (N_12443,N_12373,N_12372);
and U12444 (N_12444,N_12202,N_12369);
xor U12445 (N_12445,N_12377,N_12237);
nand U12446 (N_12446,N_12290,N_12298);
xnor U12447 (N_12447,N_12371,N_12227);
nor U12448 (N_12448,N_12352,N_12359);
xor U12449 (N_12449,N_12299,N_12247);
nor U12450 (N_12450,N_12212,N_12214);
or U12451 (N_12451,N_12244,N_12259);
nand U12452 (N_12452,N_12206,N_12246);
nor U12453 (N_12453,N_12267,N_12341);
nor U12454 (N_12454,N_12294,N_12293);
nand U12455 (N_12455,N_12224,N_12243);
nand U12456 (N_12456,N_12250,N_12313);
and U12457 (N_12457,N_12234,N_12238);
nor U12458 (N_12458,N_12384,N_12354);
xnor U12459 (N_12459,N_12334,N_12383);
nor U12460 (N_12460,N_12282,N_12229);
or U12461 (N_12461,N_12348,N_12261);
and U12462 (N_12462,N_12378,N_12318);
nor U12463 (N_12463,N_12296,N_12340);
nor U12464 (N_12464,N_12230,N_12317);
nor U12465 (N_12465,N_12297,N_12367);
and U12466 (N_12466,N_12316,N_12379);
nand U12467 (N_12467,N_12232,N_12248);
nor U12468 (N_12468,N_12291,N_12338);
xor U12469 (N_12469,N_12344,N_12356);
xnor U12470 (N_12470,N_12220,N_12374);
nand U12471 (N_12471,N_12347,N_12260);
and U12472 (N_12472,N_12382,N_12315);
nand U12473 (N_12473,N_12255,N_12270);
xor U12474 (N_12474,N_12337,N_12391);
xor U12475 (N_12475,N_12380,N_12254);
nand U12476 (N_12476,N_12239,N_12393);
nand U12477 (N_12477,N_12295,N_12390);
nor U12478 (N_12478,N_12204,N_12388);
nand U12479 (N_12479,N_12361,N_12358);
and U12480 (N_12480,N_12303,N_12343);
nor U12481 (N_12481,N_12281,N_12321);
or U12482 (N_12482,N_12301,N_12333);
nand U12483 (N_12483,N_12324,N_12213);
nand U12484 (N_12484,N_12222,N_12219);
nor U12485 (N_12485,N_12320,N_12355);
xnor U12486 (N_12486,N_12351,N_12349);
nor U12487 (N_12487,N_12370,N_12228);
nor U12488 (N_12488,N_12392,N_12275);
or U12489 (N_12489,N_12236,N_12330);
nand U12490 (N_12490,N_12398,N_12360);
xnor U12491 (N_12491,N_12235,N_12386);
nor U12492 (N_12492,N_12306,N_12233);
xnor U12493 (N_12493,N_12345,N_12241);
xnor U12494 (N_12494,N_12251,N_12395);
and U12495 (N_12495,N_12278,N_12277);
and U12496 (N_12496,N_12362,N_12314);
nor U12497 (N_12497,N_12217,N_12307);
nor U12498 (N_12498,N_12353,N_12288);
and U12499 (N_12499,N_12304,N_12268);
xnor U12500 (N_12500,N_12269,N_12313);
or U12501 (N_12501,N_12298,N_12221);
nand U12502 (N_12502,N_12284,N_12269);
xnor U12503 (N_12503,N_12280,N_12307);
or U12504 (N_12504,N_12234,N_12258);
nand U12505 (N_12505,N_12262,N_12219);
or U12506 (N_12506,N_12306,N_12216);
and U12507 (N_12507,N_12248,N_12284);
or U12508 (N_12508,N_12256,N_12203);
nand U12509 (N_12509,N_12251,N_12264);
and U12510 (N_12510,N_12309,N_12218);
nor U12511 (N_12511,N_12287,N_12280);
and U12512 (N_12512,N_12314,N_12207);
nor U12513 (N_12513,N_12388,N_12301);
and U12514 (N_12514,N_12343,N_12364);
and U12515 (N_12515,N_12384,N_12342);
or U12516 (N_12516,N_12224,N_12259);
or U12517 (N_12517,N_12251,N_12324);
or U12518 (N_12518,N_12269,N_12216);
and U12519 (N_12519,N_12203,N_12279);
xor U12520 (N_12520,N_12359,N_12260);
xnor U12521 (N_12521,N_12254,N_12318);
and U12522 (N_12522,N_12292,N_12201);
nand U12523 (N_12523,N_12239,N_12313);
and U12524 (N_12524,N_12380,N_12224);
xor U12525 (N_12525,N_12235,N_12273);
xor U12526 (N_12526,N_12398,N_12240);
and U12527 (N_12527,N_12251,N_12389);
nor U12528 (N_12528,N_12238,N_12372);
and U12529 (N_12529,N_12230,N_12395);
or U12530 (N_12530,N_12311,N_12304);
and U12531 (N_12531,N_12203,N_12295);
nor U12532 (N_12532,N_12358,N_12362);
or U12533 (N_12533,N_12325,N_12232);
or U12534 (N_12534,N_12286,N_12313);
xnor U12535 (N_12535,N_12336,N_12209);
or U12536 (N_12536,N_12213,N_12229);
xor U12537 (N_12537,N_12396,N_12202);
nand U12538 (N_12538,N_12381,N_12288);
nand U12539 (N_12539,N_12351,N_12328);
nor U12540 (N_12540,N_12371,N_12319);
nand U12541 (N_12541,N_12390,N_12207);
nand U12542 (N_12542,N_12226,N_12356);
xnor U12543 (N_12543,N_12357,N_12309);
and U12544 (N_12544,N_12333,N_12201);
nor U12545 (N_12545,N_12328,N_12292);
and U12546 (N_12546,N_12335,N_12333);
nor U12547 (N_12547,N_12348,N_12343);
or U12548 (N_12548,N_12392,N_12328);
nor U12549 (N_12549,N_12327,N_12237);
nand U12550 (N_12550,N_12305,N_12364);
nand U12551 (N_12551,N_12225,N_12365);
or U12552 (N_12552,N_12275,N_12205);
and U12553 (N_12553,N_12312,N_12333);
and U12554 (N_12554,N_12265,N_12249);
xnor U12555 (N_12555,N_12323,N_12250);
nand U12556 (N_12556,N_12257,N_12330);
xor U12557 (N_12557,N_12366,N_12228);
xnor U12558 (N_12558,N_12206,N_12242);
nor U12559 (N_12559,N_12327,N_12236);
and U12560 (N_12560,N_12359,N_12385);
nor U12561 (N_12561,N_12244,N_12391);
nor U12562 (N_12562,N_12319,N_12225);
or U12563 (N_12563,N_12235,N_12239);
xnor U12564 (N_12564,N_12249,N_12337);
xor U12565 (N_12565,N_12303,N_12216);
xnor U12566 (N_12566,N_12249,N_12262);
nor U12567 (N_12567,N_12209,N_12264);
nand U12568 (N_12568,N_12217,N_12206);
xnor U12569 (N_12569,N_12332,N_12208);
or U12570 (N_12570,N_12216,N_12348);
or U12571 (N_12571,N_12341,N_12357);
nand U12572 (N_12572,N_12289,N_12383);
and U12573 (N_12573,N_12317,N_12377);
or U12574 (N_12574,N_12219,N_12306);
or U12575 (N_12575,N_12360,N_12390);
nand U12576 (N_12576,N_12200,N_12366);
nand U12577 (N_12577,N_12200,N_12373);
xnor U12578 (N_12578,N_12214,N_12312);
nor U12579 (N_12579,N_12222,N_12304);
xor U12580 (N_12580,N_12276,N_12365);
and U12581 (N_12581,N_12368,N_12222);
and U12582 (N_12582,N_12279,N_12388);
or U12583 (N_12583,N_12243,N_12394);
xor U12584 (N_12584,N_12283,N_12320);
nor U12585 (N_12585,N_12304,N_12271);
nor U12586 (N_12586,N_12320,N_12243);
xor U12587 (N_12587,N_12278,N_12221);
or U12588 (N_12588,N_12246,N_12247);
nand U12589 (N_12589,N_12288,N_12342);
nand U12590 (N_12590,N_12224,N_12365);
or U12591 (N_12591,N_12350,N_12385);
nand U12592 (N_12592,N_12285,N_12355);
or U12593 (N_12593,N_12307,N_12250);
and U12594 (N_12594,N_12223,N_12294);
xor U12595 (N_12595,N_12341,N_12287);
or U12596 (N_12596,N_12272,N_12299);
nor U12597 (N_12597,N_12232,N_12366);
or U12598 (N_12598,N_12313,N_12263);
and U12599 (N_12599,N_12213,N_12273);
or U12600 (N_12600,N_12445,N_12491);
xor U12601 (N_12601,N_12431,N_12588);
and U12602 (N_12602,N_12406,N_12553);
nand U12603 (N_12603,N_12470,N_12451);
nand U12604 (N_12604,N_12434,N_12484);
and U12605 (N_12605,N_12453,N_12595);
and U12606 (N_12606,N_12450,N_12401);
nand U12607 (N_12607,N_12419,N_12459);
or U12608 (N_12608,N_12418,N_12527);
and U12609 (N_12609,N_12426,N_12481);
xnor U12610 (N_12610,N_12587,N_12545);
nor U12611 (N_12611,N_12467,N_12578);
nand U12612 (N_12612,N_12540,N_12511);
and U12613 (N_12613,N_12579,N_12519);
or U12614 (N_12614,N_12506,N_12437);
nor U12615 (N_12615,N_12425,N_12525);
nand U12616 (N_12616,N_12454,N_12576);
nand U12617 (N_12617,N_12599,N_12490);
or U12618 (N_12618,N_12513,N_12552);
xor U12619 (N_12619,N_12492,N_12403);
xor U12620 (N_12620,N_12410,N_12427);
nor U12621 (N_12621,N_12569,N_12543);
nor U12622 (N_12622,N_12440,N_12478);
and U12623 (N_12623,N_12452,N_12412);
nor U12624 (N_12624,N_12479,N_12496);
nand U12625 (N_12625,N_12449,N_12574);
xnor U12626 (N_12626,N_12529,N_12524);
or U12627 (N_12627,N_12458,N_12423);
nand U12628 (N_12628,N_12542,N_12477);
nor U12629 (N_12629,N_12499,N_12518);
and U12630 (N_12630,N_12420,N_12556);
nor U12631 (N_12631,N_12590,N_12494);
nor U12632 (N_12632,N_12544,N_12593);
nand U12633 (N_12633,N_12554,N_12582);
and U12634 (N_12634,N_12560,N_12537);
nor U12635 (N_12635,N_12523,N_12501);
nor U12636 (N_12636,N_12476,N_12417);
and U12637 (N_12637,N_12514,N_12487);
xnor U12638 (N_12638,N_12432,N_12485);
nor U12639 (N_12639,N_12448,N_12565);
and U12640 (N_12640,N_12473,N_12500);
and U12641 (N_12641,N_12571,N_12515);
and U12642 (N_12642,N_12480,N_12598);
and U12643 (N_12643,N_12555,N_12503);
and U12644 (N_12644,N_12568,N_12522);
nand U12645 (N_12645,N_12517,N_12455);
xnor U12646 (N_12646,N_12497,N_12549);
and U12647 (N_12647,N_12559,N_12584);
or U12648 (N_12648,N_12446,N_12483);
xor U12649 (N_12649,N_12520,N_12502);
nor U12650 (N_12650,N_12586,N_12474);
nand U12651 (N_12651,N_12441,N_12585);
and U12652 (N_12652,N_12566,N_12488);
xnor U12653 (N_12653,N_12468,N_12534);
and U12654 (N_12654,N_12541,N_12589);
or U12655 (N_12655,N_12548,N_12409);
nand U12656 (N_12656,N_12411,N_12413);
nand U12657 (N_12657,N_12443,N_12498);
nand U12658 (N_12658,N_12428,N_12505);
nand U12659 (N_12659,N_12464,N_12504);
nor U12660 (N_12660,N_12563,N_12557);
xor U12661 (N_12661,N_12561,N_12422);
nand U12662 (N_12662,N_12550,N_12430);
nand U12663 (N_12663,N_12564,N_12546);
nand U12664 (N_12664,N_12439,N_12509);
xor U12665 (N_12665,N_12402,N_12526);
xor U12666 (N_12666,N_12472,N_12530);
and U12667 (N_12667,N_12400,N_12482);
xor U12668 (N_12668,N_12442,N_12562);
nand U12669 (N_12669,N_12528,N_12575);
or U12670 (N_12670,N_12572,N_12493);
nand U12671 (N_12671,N_12536,N_12516);
xor U12672 (N_12672,N_12407,N_12465);
xnor U12673 (N_12673,N_12508,N_12456);
xnor U12674 (N_12674,N_12533,N_12594);
and U12675 (N_12675,N_12444,N_12404);
xnor U12676 (N_12676,N_12436,N_12551);
nor U12677 (N_12677,N_12495,N_12583);
xor U12678 (N_12678,N_12521,N_12424);
or U12679 (N_12679,N_12447,N_12421);
xor U12680 (N_12680,N_12457,N_12475);
xor U12681 (N_12681,N_12538,N_12577);
xnor U12682 (N_12682,N_12558,N_12580);
or U12683 (N_12683,N_12462,N_12429);
and U12684 (N_12684,N_12414,N_12573);
xor U12685 (N_12685,N_12460,N_12512);
xor U12686 (N_12686,N_12415,N_12489);
or U12687 (N_12687,N_12581,N_12507);
and U12688 (N_12688,N_12597,N_12461);
and U12689 (N_12689,N_12463,N_12510);
or U12690 (N_12690,N_12547,N_12532);
and U12691 (N_12691,N_12405,N_12469);
xnor U12692 (N_12692,N_12471,N_12435);
or U12693 (N_12693,N_12592,N_12570);
nor U12694 (N_12694,N_12535,N_12591);
nand U12695 (N_12695,N_12596,N_12408);
xor U12696 (N_12696,N_12486,N_12416);
nand U12697 (N_12697,N_12438,N_12466);
nor U12698 (N_12698,N_12539,N_12433);
nand U12699 (N_12699,N_12531,N_12567);
and U12700 (N_12700,N_12498,N_12510);
xor U12701 (N_12701,N_12481,N_12463);
or U12702 (N_12702,N_12581,N_12497);
nor U12703 (N_12703,N_12595,N_12429);
nand U12704 (N_12704,N_12582,N_12558);
nand U12705 (N_12705,N_12558,N_12576);
and U12706 (N_12706,N_12526,N_12587);
nand U12707 (N_12707,N_12540,N_12468);
nand U12708 (N_12708,N_12440,N_12521);
or U12709 (N_12709,N_12497,N_12559);
xor U12710 (N_12710,N_12461,N_12575);
and U12711 (N_12711,N_12461,N_12583);
and U12712 (N_12712,N_12518,N_12402);
nor U12713 (N_12713,N_12539,N_12412);
or U12714 (N_12714,N_12462,N_12599);
nor U12715 (N_12715,N_12444,N_12591);
nor U12716 (N_12716,N_12432,N_12560);
and U12717 (N_12717,N_12420,N_12408);
or U12718 (N_12718,N_12575,N_12400);
or U12719 (N_12719,N_12538,N_12442);
or U12720 (N_12720,N_12573,N_12593);
nor U12721 (N_12721,N_12500,N_12567);
nand U12722 (N_12722,N_12401,N_12595);
and U12723 (N_12723,N_12533,N_12504);
or U12724 (N_12724,N_12524,N_12417);
nor U12725 (N_12725,N_12420,N_12487);
nor U12726 (N_12726,N_12560,N_12455);
xnor U12727 (N_12727,N_12465,N_12416);
nor U12728 (N_12728,N_12537,N_12535);
nand U12729 (N_12729,N_12428,N_12410);
nor U12730 (N_12730,N_12486,N_12499);
or U12731 (N_12731,N_12449,N_12496);
nor U12732 (N_12732,N_12568,N_12407);
xor U12733 (N_12733,N_12427,N_12595);
nor U12734 (N_12734,N_12570,N_12412);
xnor U12735 (N_12735,N_12524,N_12535);
nand U12736 (N_12736,N_12441,N_12511);
or U12737 (N_12737,N_12449,N_12471);
nor U12738 (N_12738,N_12516,N_12546);
nand U12739 (N_12739,N_12598,N_12594);
nor U12740 (N_12740,N_12415,N_12468);
xor U12741 (N_12741,N_12599,N_12504);
and U12742 (N_12742,N_12598,N_12429);
or U12743 (N_12743,N_12534,N_12531);
nor U12744 (N_12744,N_12414,N_12566);
and U12745 (N_12745,N_12455,N_12569);
nor U12746 (N_12746,N_12556,N_12407);
nand U12747 (N_12747,N_12589,N_12402);
xor U12748 (N_12748,N_12551,N_12460);
xnor U12749 (N_12749,N_12509,N_12584);
nor U12750 (N_12750,N_12526,N_12501);
xnor U12751 (N_12751,N_12575,N_12510);
xor U12752 (N_12752,N_12503,N_12496);
and U12753 (N_12753,N_12483,N_12565);
xnor U12754 (N_12754,N_12565,N_12464);
and U12755 (N_12755,N_12528,N_12563);
nand U12756 (N_12756,N_12450,N_12517);
and U12757 (N_12757,N_12417,N_12585);
and U12758 (N_12758,N_12542,N_12573);
or U12759 (N_12759,N_12598,N_12557);
nor U12760 (N_12760,N_12472,N_12446);
and U12761 (N_12761,N_12565,N_12525);
and U12762 (N_12762,N_12548,N_12584);
nand U12763 (N_12763,N_12480,N_12503);
or U12764 (N_12764,N_12565,N_12561);
xor U12765 (N_12765,N_12447,N_12430);
or U12766 (N_12766,N_12448,N_12415);
and U12767 (N_12767,N_12525,N_12589);
nor U12768 (N_12768,N_12580,N_12438);
or U12769 (N_12769,N_12474,N_12456);
and U12770 (N_12770,N_12545,N_12407);
and U12771 (N_12771,N_12422,N_12577);
xor U12772 (N_12772,N_12516,N_12504);
nand U12773 (N_12773,N_12516,N_12482);
or U12774 (N_12774,N_12582,N_12501);
or U12775 (N_12775,N_12411,N_12435);
and U12776 (N_12776,N_12422,N_12510);
and U12777 (N_12777,N_12492,N_12491);
nand U12778 (N_12778,N_12565,N_12470);
nand U12779 (N_12779,N_12429,N_12504);
nor U12780 (N_12780,N_12564,N_12599);
and U12781 (N_12781,N_12493,N_12587);
nor U12782 (N_12782,N_12486,N_12502);
and U12783 (N_12783,N_12462,N_12588);
xnor U12784 (N_12784,N_12494,N_12564);
nor U12785 (N_12785,N_12410,N_12435);
nor U12786 (N_12786,N_12424,N_12466);
or U12787 (N_12787,N_12486,N_12497);
and U12788 (N_12788,N_12448,N_12471);
xor U12789 (N_12789,N_12438,N_12552);
and U12790 (N_12790,N_12530,N_12425);
and U12791 (N_12791,N_12418,N_12405);
and U12792 (N_12792,N_12548,N_12528);
nor U12793 (N_12793,N_12475,N_12512);
or U12794 (N_12794,N_12410,N_12485);
nand U12795 (N_12795,N_12500,N_12466);
nor U12796 (N_12796,N_12407,N_12460);
xnor U12797 (N_12797,N_12509,N_12576);
nand U12798 (N_12798,N_12498,N_12446);
xor U12799 (N_12799,N_12544,N_12577);
or U12800 (N_12800,N_12723,N_12731);
nand U12801 (N_12801,N_12611,N_12734);
nor U12802 (N_12802,N_12621,N_12602);
xor U12803 (N_12803,N_12631,N_12725);
or U12804 (N_12804,N_12746,N_12653);
or U12805 (N_12805,N_12622,N_12702);
xor U12806 (N_12806,N_12788,N_12641);
xor U12807 (N_12807,N_12697,N_12669);
xor U12808 (N_12808,N_12608,N_12676);
xnor U12809 (N_12809,N_12728,N_12696);
nand U12810 (N_12810,N_12717,N_12714);
or U12811 (N_12811,N_12713,N_12614);
or U12812 (N_12812,N_12703,N_12662);
nand U12813 (N_12813,N_12786,N_12638);
and U12814 (N_12814,N_12644,N_12687);
nor U12815 (N_12815,N_12666,N_12749);
nand U12816 (N_12816,N_12757,N_12642);
and U12817 (N_12817,N_12795,N_12707);
or U12818 (N_12818,N_12724,N_12754);
nand U12819 (N_12819,N_12793,N_12693);
xor U12820 (N_12820,N_12718,N_12605);
and U12821 (N_12821,N_12668,N_12737);
xor U12822 (N_12822,N_12615,N_12701);
nand U12823 (N_12823,N_12628,N_12719);
and U12824 (N_12824,N_12655,N_12623);
nor U12825 (N_12825,N_12705,N_12775);
nor U12826 (N_12826,N_12685,N_12625);
nor U12827 (N_12827,N_12679,N_12726);
and U12828 (N_12828,N_12667,N_12601);
nand U12829 (N_12829,N_12681,N_12698);
xnor U12830 (N_12830,N_12646,N_12633);
xnor U12831 (N_12831,N_12750,N_12771);
nand U12832 (N_12832,N_12721,N_12764);
and U12833 (N_12833,N_12634,N_12678);
nor U12834 (N_12834,N_12799,N_12770);
nor U12835 (N_12835,N_12682,N_12767);
xor U12836 (N_12836,N_12629,N_12619);
nand U12837 (N_12837,N_12677,N_12773);
and U12838 (N_12838,N_12607,N_12643);
nand U12839 (N_12839,N_12792,N_12658);
nand U12840 (N_12840,N_12732,N_12798);
nor U12841 (N_12841,N_12675,N_12782);
nand U12842 (N_12842,N_12691,N_12797);
nand U12843 (N_12843,N_12672,N_12654);
nand U12844 (N_12844,N_12722,N_12657);
nor U12845 (N_12845,N_12626,N_12783);
nand U12846 (N_12846,N_12747,N_12661);
and U12847 (N_12847,N_12694,N_12704);
nor U12848 (N_12848,N_12651,N_12688);
or U12849 (N_12849,N_12711,N_12743);
xnor U12850 (N_12850,N_12755,N_12680);
and U12851 (N_12851,N_12710,N_12742);
and U12852 (N_12852,N_12778,N_12618);
or U12853 (N_12853,N_12700,N_12789);
nor U12854 (N_12854,N_12761,N_12659);
xnor U12855 (N_12855,N_12744,N_12616);
or U12856 (N_12856,N_12781,N_12727);
nand U12857 (N_12857,N_12785,N_12612);
nor U12858 (N_12858,N_12787,N_12709);
xnor U12859 (N_12859,N_12752,N_12738);
nor U12860 (N_12860,N_12766,N_12630);
and U12861 (N_12861,N_12600,N_12617);
nor U12862 (N_12862,N_12636,N_12620);
nand U12863 (N_12863,N_12663,N_12748);
or U12864 (N_12864,N_12650,N_12673);
xor U12865 (N_12865,N_12674,N_12791);
xor U12866 (N_12866,N_12706,N_12699);
nor U12867 (N_12867,N_12664,N_12606);
nor U12868 (N_12868,N_12649,N_12686);
nand U12869 (N_12869,N_12796,N_12739);
nand U12870 (N_12870,N_12647,N_12768);
and U12871 (N_12871,N_12652,N_12776);
nand U12872 (N_12872,N_12604,N_12695);
xor U12873 (N_12873,N_12640,N_12689);
and U12874 (N_12874,N_12715,N_12656);
xor U12875 (N_12875,N_12756,N_12741);
nand U12876 (N_12876,N_12683,N_12627);
or U12877 (N_12877,N_12730,N_12690);
or U12878 (N_12878,N_12692,N_12779);
and U12879 (N_12879,N_12684,N_12758);
xor U12880 (N_12880,N_12736,N_12774);
nand U12881 (N_12881,N_12753,N_12784);
nor U12882 (N_12882,N_12632,N_12765);
or U12883 (N_12883,N_12762,N_12603);
nand U12884 (N_12884,N_12790,N_12780);
or U12885 (N_12885,N_12639,N_12609);
and U12886 (N_12886,N_12624,N_12645);
xor U12887 (N_12887,N_12708,N_12751);
or U12888 (N_12888,N_12745,N_12716);
or U12889 (N_12889,N_12740,N_12763);
or U12890 (N_12890,N_12665,N_12637);
xor U12891 (N_12891,N_12648,N_12735);
and U12892 (N_12892,N_12733,N_12769);
nor U12893 (N_12893,N_12777,N_12794);
and U12894 (N_12894,N_12772,N_12729);
nand U12895 (N_12895,N_12671,N_12720);
and U12896 (N_12896,N_12610,N_12613);
nand U12897 (N_12897,N_12759,N_12760);
and U12898 (N_12898,N_12712,N_12670);
nand U12899 (N_12899,N_12635,N_12660);
nor U12900 (N_12900,N_12620,N_12779);
and U12901 (N_12901,N_12627,N_12757);
and U12902 (N_12902,N_12654,N_12605);
nand U12903 (N_12903,N_12657,N_12750);
nor U12904 (N_12904,N_12650,N_12692);
and U12905 (N_12905,N_12652,N_12602);
and U12906 (N_12906,N_12643,N_12788);
nor U12907 (N_12907,N_12723,N_12616);
nor U12908 (N_12908,N_12793,N_12607);
or U12909 (N_12909,N_12621,N_12760);
nand U12910 (N_12910,N_12732,N_12600);
nor U12911 (N_12911,N_12786,N_12763);
xor U12912 (N_12912,N_12788,N_12733);
nor U12913 (N_12913,N_12682,N_12688);
nor U12914 (N_12914,N_12636,N_12655);
or U12915 (N_12915,N_12658,N_12671);
xnor U12916 (N_12916,N_12712,N_12766);
nand U12917 (N_12917,N_12742,N_12781);
nor U12918 (N_12918,N_12645,N_12786);
or U12919 (N_12919,N_12675,N_12686);
nand U12920 (N_12920,N_12628,N_12641);
nor U12921 (N_12921,N_12755,N_12773);
nor U12922 (N_12922,N_12704,N_12691);
and U12923 (N_12923,N_12793,N_12712);
nor U12924 (N_12924,N_12765,N_12607);
xnor U12925 (N_12925,N_12695,N_12780);
or U12926 (N_12926,N_12732,N_12651);
and U12927 (N_12927,N_12755,N_12694);
nor U12928 (N_12928,N_12626,N_12647);
xor U12929 (N_12929,N_12602,N_12689);
nand U12930 (N_12930,N_12696,N_12642);
xor U12931 (N_12931,N_12708,N_12684);
nand U12932 (N_12932,N_12764,N_12684);
nor U12933 (N_12933,N_12616,N_12699);
xnor U12934 (N_12934,N_12656,N_12600);
or U12935 (N_12935,N_12668,N_12700);
xnor U12936 (N_12936,N_12718,N_12708);
and U12937 (N_12937,N_12694,N_12647);
xnor U12938 (N_12938,N_12621,N_12665);
or U12939 (N_12939,N_12771,N_12783);
xnor U12940 (N_12940,N_12774,N_12746);
or U12941 (N_12941,N_12756,N_12789);
or U12942 (N_12942,N_12775,N_12747);
xor U12943 (N_12943,N_12682,N_12787);
nor U12944 (N_12944,N_12610,N_12790);
and U12945 (N_12945,N_12765,N_12610);
and U12946 (N_12946,N_12767,N_12786);
nand U12947 (N_12947,N_12692,N_12609);
nand U12948 (N_12948,N_12610,N_12660);
or U12949 (N_12949,N_12759,N_12634);
or U12950 (N_12950,N_12711,N_12616);
xnor U12951 (N_12951,N_12657,N_12735);
or U12952 (N_12952,N_12615,N_12610);
nand U12953 (N_12953,N_12611,N_12787);
or U12954 (N_12954,N_12602,N_12693);
xnor U12955 (N_12955,N_12649,N_12652);
or U12956 (N_12956,N_12684,N_12608);
nand U12957 (N_12957,N_12770,N_12649);
xor U12958 (N_12958,N_12630,N_12613);
and U12959 (N_12959,N_12739,N_12617);
and U12960 (N_12960,N_12753,N_12620);
xor U12961 (N_12961,N_12710,N_12711);
and U12962 (N_12962,N_12759,N_12701);
nor U12963 (N_12963,N_12792,N_12743);
or U12964 (N_12964,N_12703,N_12637);
and U12965 (N_12965,N_12756,N_12753);
and U12966 (N_12966,N_12785,N_12744);
xor U12967 (N_12967,N_12663,N_12775);
or U12968 (N_12968,N_12742,N_12663);
nand U12969 (N_12969,N_12729,N_12604);
xor U12970 (N_12970,N_12782,N_12628);
nand U12971 (N_12971,N_12703,N_12791);
nor U12972 (N_12972,N_12656,N_12687);
nand U12973 (N_12973,N_12658,N_12761);
or U12974 (N_12974,N_12771,N_12649);
xnor U12975 (N_12975,N_12760,N_12756);
and U12976 (N_12976,N_12617,N_12650);
nor U12977 (N_12977,N_12697,N_12642);
nand U12978 (N_12978,N_12759,N_12763);
xnor U12979 (N_12979,N_12616,N_12784);
nor U12980 (N_12980,N_12676,N_12745);
nor U12981 (N_12981,N_12713,N_12695);
nand U12982 (N_12982,N_12703,N_12649);
or U12983 (N_12983,N_12725,N_12765);
xnor U12984 (N_12984,N_12682,N_12732);
nand U12985 (N_12985,N_12603,N_12770);
or U12986 (N_12986,N_12652,N_12625);
or U12987 (N_12987,N_12794,N_12678);
nor U12988 (N_12988,N_12727,N_12768);
and U12989 (N_12989,N_12645,N_12670);
nand U12990 (N_12990,N_12738,N_12724);
nand U12991 (N_12991,N_12633,N_12746);
xor U12992 (N_12992,N_12607,N_12741);
and U12993 (N_12993,N_12767,N_12712);
nor U12994 (N_12994,N_12618,N_12781);
and U12995 (N_12995,N_12772,N_12662);
nor U12996 (N_12996,N_12708,N_12769);
and U12997 (N_12997,N_12771,N_12627);
and U12998 (N_12998,N_12770,N_12768);
or U12999 (N_12999,N_12678,N_12706);
nand U13000 (N_13000,N_12802,N_12900);
xor U13001 (N_13001,N_12948,N_12924);
xnor U13002 (N_13002,N_12945,N_12861);
or U13003 (N_13003,N_12801,N_12984);
nor U13004 (N_13004,N_12963,N_12850);
and U13005 (N_13005,N_12846,N_12864);
nand U13006 (N_13006,N_12830,N_12936);
nand U13007 (N_13007,N_12999,N_12839);
nand U13008 (N_13008,N_12889,N_12987);
or U13009 (N_13009,N_12813,N_12940);
or U13010 (N_13010,N_12968,N_12949);
and U13011 (N_13011,N_12904,N_12928);
nand U13012 (N_13012,N_12894,N_12881);
or U13013 (N_13013,N_12821,N_12962);
xor U13014 (N_13014,N_12932,N_12970);
xnor U13015 (N_13015,N_12847,N_12921);
and U13016 (N_13016,N_12982,N_12837);
xor U13017 (N_13017,N_12833,N_12874);
nor U13018 (N_13018,N_12906,N_12989);
or U13019 (N_13019,N_12840,N_12927);
nand U13020 (N_13020,N_12937,N_12981);
or U13021 (N_13021,N_12951,N_12955);
xnor U13022 (N_13022,N_12865,N_12965);
xor U13023 (N_13023,N_12986,N_12854);
and U13024 (N_13024,N_12966,N_12944);
nand U13025 (N_13025,N_12871,N_12817);
and U13026 (N_13026,N_12895,N_12980);
and U13027 (N_13027,N_12994,N_12979);
nor U13028 (N_13028,N_12803,N_12903);
and U13029 (N_13029,N_12931,N_12993);
xnor U13030 (N_13030,N_12905,N_12884);
nand U13031 (N_13031,N_12841,N_12880);
or U13032 (N_13032,N_12976,N_12914);
or U13033 (N_13033,N_12814,N_12831);
nand U13034 (N_13034,N_12818,N_12899);
nand U13035 (N_13035,N_12909,N_12959);
xnor U13036 (N_13036,N_12870,N_12848);
nor U13037 (N_13037,N_12923,N_12810);
or U13038 (N_13038,N_12898,N_12812);
and U13039 (N_13039,N_12827,N_12912);
and U13040 (N_13040,N_12882,N_12893);
or U13041 (N_13041,N_12890,N_12964);
and U13042 (N_13042,N_12942,N_12954);
nor U13043 (N_13043,N_12869,N_12855);
xnor U13044 (N_13044,N_12907,N_12852);
nand U13045 (N_13045,N_12971,N_12834);
nor U13046 (N_13046,N_12851,N_12910);
or U13047 (N_13047,N_12943,N_12958);
nor U13048 (N_13048,N_12888,N_12997);
or U13049 (N_13049,N_12857,N_12856);
and U13050 (N_13050,N_12991,N_12918);
nor U13051 (N_13051,N_12967,N_12908);
nor U13052 (N_13052,N_12866,N_12800);
and U13053 (N_13053,N_12974,N_12863);
or U13054 (N_13054,N_12878,N_12862);
nor U13055 (N_13055,N_12952,N_12879);
nand U13056 (N_13056,N_12915,N_12825);
and U13057 (N_13057,N_12956,N_12824);
nand U13058 (N_13058,N_12875,N_12992);
nor U13059 (N_13059,N_12805,N_12977);
or U13060 (N_13060,N_12872,N_12985);
or U13061 (N_13061,N_12816,N_12933);
nand U13062 (N_13062,N_12925,N_12960);
and U13063 (N_13063,N_12941,N_12867);
xor U13064 (N_13064,N_12828,N_12930);
xnor U13065 (N_13065,N_12804,N_12807);
and U13066 (N_13066,N_12806,N_12946);
or U13067 (N_13067,N_12990,N_12896);
nand U13068 (N_13068,N_12916,N_12988);
nand U13069 (N_13069,N_12835,N_12913);
xnor U13070 (N_13070,N_12820,N_12919);
nand U13071 (N_13071,N_12996,N_12836);
xor U13072 (N_13072,N_12838,N_12885);
and U13073 (N_13073,N_12808,N_12973);
or U13074 (N_13074,N_12823,N_12975);
and U13075 (N_13075,N_12926,N_12858);
nand U13076 (N_13076,N_12883,N_12972);
and U13077 (N_13077,N_12902,N_12859);
or U13078 (N_13078,N_12920,N_12876);
nand U13079 (N_13079,N_12845,N_12950);
nand U13080 (N_13080,N_12938,N_12843);
nor U13081 (N_13081,N_12917,N_12998);
or U13082 (N_13082,N_12868,N_12901);
or U13083 (N_13083,N_12873,N_12829);
nand U13084 (N_13084,N_12886,N_12891);
or U13085 (N_13085,N_12819,N_12983);
xor U13086 (N_13086,N_12877,N_12978);
xor U13087 (N_13087,N_12832,N_12969);
or U13088 (N_13088,N_12809,N_12934);
nor U13089 (N_13089,N_12844,N_12935);
and U13090 (N_13090,N_12961,N_12815);
xor U13091 (N_13091,N_12957,N_12860);
or U13092 (N_13092,N_12953,N_12811);
nor U13093 (N_13093,N_12842,N_12826);
or U13094 (N_13094,N_12849,N_12995);
nand U13095 (N_13095,N_12939,N_12929);
and U13096 (N_13096,N_12897,N_12892);
xnor U13097 (N_13097,N_12911,N_12947);
or U13098 (N_13098,N_12822,N_12853);
nand U13099 (N_13099,N_12887,N_12922);
nor U13100 (N_13100,N_12990,N_12963);
nor U13101 (N_13101,N_12866,N_12902);
nand U13102 (N_13102,N_12972,N_12807);
nor U13103 (N_13103,N_12826,N_12986);
or U13104 (N_13104,N_12920,N_12865);
nand U13105 (N_13105,N_12921,N_12990);
and U13106 (N_13106,N_12939,N_12936);
and U13107 (N_13107,N_12888,N_12835);
or U13108 (N_13108,N_12942,N_12828);
and U13109 (N_13109,N_12949,N_12827);
or U13110 (N_13110,N_12812,N_12867);
or U13111 (N_13111,N_12901,N_12974);
xnor U13112 (N_13112,N_12905,N_12971);
nor U13113 (N_13113,N_12992,N_12823);
and U13114 (N_13114,N_12872,N_12890);
nor U13115 (N_13115,N_12824,N_12930);
nor U13116 (N_13116,N_12965,N_12847);
nor U13117 (N_13117,N_12893,N_12811);
nor U13118 (N_13118,N_12936,N_12880);
or U13119 (N_13119,N_12985,N_12995);
nor U13120 (N_13120,N_12950,N_12850);
xnor U13121 (N_13121,N_12851,N_12953);
nor U13122 (N_13122,N_12938,N_12900);
nor U13123 (N_13123,N_12862,N_12894);
xor U13124 (N_13124,N_12960,N_12985);
or U13125 (N_13125,N_12817,N_12897);
or U13126 (N_13126,N_12863,N_12840);
xor U13127 (N_13127,N_12948,N_12957);
xnor U13128 (N_13128,N_12842,N_12914);
nor U13129 (N_13129,N_12925,N_12846);
nand U13130 (N_13130,N_12913,N_12916);
or U13131 (N_13131,N_12925,N_12902);
and U13132 (N_13132,N_12869,N_12922);
nor U13133 (N_13133,N_12823,N_12811);
nand U13134 (N_13134,N_12836,N_12905);
and U13135 (N_13135,N_12942,N_12931);
nor U13136 (N_13136,N_12818,N_12838);
and U13137 (N_13137,N_12836,N_12918);
and U13138 (N_13138,N_12849,N_12814);
and U13139 (N_13139,N_12863,N_12928);
or U13140 (N_13140,N_12816,N_12945);
nor U13141 (N_13141,N_12993,N_12990);
and U13142 (N_13142,N_12880,N_12866);
and U13143 (N_13143,N_12889,N_12993);
xnor U13144 (N_13144,N_12960,N_12900);
or U13145 (N_13145,N_12805,N_12995);
or U13146 (N_13146,N_12976,N_12990);
xor U13147 (N_13147,N_12919,N_12823);
xor U13148 (N_13148,N_12816,N_12806);
xnor U13149 (N_13149,N_12921,N_12872);
xor U13150 (N_13150,N_12925,N_12888);
nor U13151 (N_13151,N_12809,N_12879);
and U13152 (N_13152,N_12832,N_12928);
xnor U13153 (N_13153,N_12877,N_12916);
xnor U13154 (N_13154,N_12851,N_12860);
and U13155 (N_13155,N_12885,N_12969);
and U13156 (N_13156,N_12819,N_12934);
and U13157 (N_13157,N_12956,N_12952);
nor U13158 (N_13158,N_12845,N_12826);
nor U13159 (N_13159,N_12927,N_12900);
nor U13160 (N_13160,N_12911,N_12837);
nor U13161 (N_13161,N_12954,N_12841);
or U13162 (N_13162,N_12962,N_12894);
xnor U13163 (N_13163,N_12873,N_12887);
nand U13164 (N_13164,N_12883,N_12869);
or U13165 (N_13165,N_12984,N_12864);
or U13166 (N_13166,N_12849,N_12874);
xor U13167 (N_13167,N_12841,N_12846);
nand U13168 (N_13168,N_12939,N_12963);
and U13169 (N_13169,N_12809,N_12914);
or U13170 (N_13170,N_12827,N_12927);
or U13171 (N_13171,N_12886,N_12963);
and U13172 (N_13172,N_12966,N_12942);
and U13173 (N_13173,N_12893,N_12828);
or U13174 (N_13174,N_12941,N_12944);
and U13175 (N_13175,N_12903,N_12967);
and U13176 (N_13176,N_12981,N_12917);
nand U13177 (N_13177,N_12850,N_12827);
or U13178 (N_13178,N_12991,N_12922);
nor U13179 (N_13179,N_12954,N_12833);
and U13180 (N_13180,N_12949,N_12932);
nand U13181 (N_13181,N_12832,N_12914);
and U13182 (N_13182,N_12825,N_12867);
nor U13183 (N_13183,N_12904,N_12850);
nor U13184 (N_13184,N_12954,N_12945);
nor U13185 (N_13185,N_12945,N_12911);
xnor U13186 (N_13186,N_12909,N_12925);
nand U13187 (N_13187,N_12887,N_12812);
or U13188 (N_13188,N_12997,N_12836);
nand U13189 (N_13189,N_12949,N_12972);
nand U13190 (N_13190,N_12995,N_12892);
nand U13191 (N_13191,N_12889,N_12947);
xnor U13192 (N_13192,N_12848,N_12920);
nand U13193 (N_13193,N_12837,N_12913);
or U13194 (N_13194,N_12932,N_12901);
xnor U13195 (N_13195,N_12853,N_12924);
or U13196 (N_13196,N_12922,N_12820);
nor U13197 (N_13197,N_12864,N_12895);
nand U13198 (N_13198,N_12905,N_12805);
nand U13199 (N_13199,N_12981,N_12956);
or U13200 (N_13200,N_13035,N_13016);
xnor U13201 (N_13201,N_13183,N_13112);
or U13202 (N_13202,N_13146,N_13103);
nor U13203 (N_13203,N_13111,N_13050);
nand U13204 (N_13204,N_13110,N_13039);
and U13205 (N_13205,N_13005,N_13190);
nand U13206 (N_13206,N_13121,N_13140);
nand U13207 (N_13207,N_13045,N_13062);
nand U13208 (N_13208,N_13082,N_13093);
nor U13209 (N_13209,N_13067,N_13132);
nor U13210 (N_13210,N_13078,N_13088);
nor U13211 (N_13211,N_13085,N_13114);
xnor U13212 (N_13212,N_13027,N_13047);
and U13213 (N_13213,N_13194,N_13100);
nor U13214 (N_13214,N_13177,N_13053);
nand U13215 (N_13215,N_13126,N_13063);
nand U13216 (N_13216,N_13116,N_13097);
xnor U13217 (N_13217,N_13007,N_13059);
and U13218 (N_13218,N_13124,N_13134);
or U13219 (N_13219,N_13105,N_13170);
and U13220 (N_13220,N_13084,N_13172);
nand U13221 (N_13221,N_13196,N_13028);
and U13222 (N_13222,N_13163,N_13167);
and U13223 (N_13223,N_13139,N_13023);
or U13224 (N_13224,N_13098,N_13025);
or U13225 (N_13225,N_13021,N_13069);
and U13226 (N_13226,N_13024,N_13101);
and U13227 (N_13227,N_13015,N_13109);
and U13228 (N_13228,N_13041,N_13072);
xnor U13229 (N_13229,N_13030,N_13185);
nor U13230 (N_13230,N_13008,N_13153);
xor U13231 (N_13231,N_13157,N_13179);
and U13232 (N_13232,N_13147,N_13189);
nand U13233 (N_13233,N_13150,N_13131);
nand U13234 (N_13234,N_13042,N_13149);
xnor U13235 (N_13235,N_13145,N_13113);
nand U13236 (N_13236,N_13026,N_13010);
xor U13237 (N_13237,N_13086,N_13187);
xnor U13238 (N_13238,N_13182,N_13119);
nor U13239 (N_13239,N_13193,N_13123);
nor U13240 (N_13240,N_13044,N_13032);
and U13241 (N_13241,N_13058,N_13003);
and U13242 (N_13242,N_13091,N_13161);
or U13243 (N_13243,N_13095,N_13006);
and U13244 (N_13244,N_13165,N_13138);
nand U13245 (N_13245,N_13137,N_13004);
nand U13246 (N_13246,N_13195,N_13087);
xor U13247 (N_13247,N_13019,N_13043);
or U13248 (N_13248,N_13074,N_13128);
nand U13249 (N_13249,N_13160,N_13040);
and U13250 (N_13250,N_13038,N_13135);
nor U13251 (N_13251,N_13031,N_13054);
and U13252 (N_13252,N_13155,N_13186);
nor U13253 (N_13253,N_13188,N_13048);
nand U13254 (N_13254,N_13017,N_13120);
xnor U13255 (N_13255,N_13061,N_13029);
nor U13256 (N_13256,N_13060,N_13133);
xor U13257 (N_13257,N_13130,N_13020);
nand U13258 (N_13258,N_13051,N_13118);
nand U13259 (N_13259,N_13037,N_13141);
and U13260 (N_13260,N_13168,N_13056);
or U13261 (N_13261,N_13081,N_13011);
nor U13262 (N_13262,N_13129,N_13181);
nand U13263 (N_13263,N_13154,N_13075);
nand U13264 (N_13264,N_13012,N_13174);
and U13265 (N_13265,N_13180,N_13106);
nor U13266 (N_13266,N_13178,N_13073);
xor U13267 (N_13267,N_13175,N_13159);
or U13268 (N_13268,N_13104,N_13117);
xor U13269 (N_13269,N_13001,N_13136);
and U13270 (N_13270,N_13192,N_13068);
nand U13271 (N_13271,N_13191,N_13049);
and U13272 (N_13272,N_13142,N_13052);
and U13273 (N_13273,N_13171,N_13036);
and U13274 (N_13274,N_13018,N_13080);
nor U13275 (N_13275,N_13013,N_13057);
nor U13276 (N_13276,N_13034,N_13083);
and U13277 (N_13277,N_13144,N_13071);
nand U13278 (N_13278,N_13046,N_13122);
nor U13279 (N_13279,N_13127,N_13102);
nand U13280 (N_13280,N_13151,N_13108);
or U13281 (N_13281,N_13089,N_13158);
or U13282 (N_13282,N_13197,N_13164);
nand U13283 (N_13283,N_13094,N_13066);
or U13284 (N_13284,N_13156,N_13000);
xnor U13285 (N_13285,N_13064,N_13143);
and U13286 (N_13286,N_13166,N_13090);
nand U13287 (N_13287,N_13002,N_13099);
and U13288 (N_13288,N_13199,N_13107);
xor U13289 (N_13289,N_13033,N_13198);
or U13290 (N_13290,N_13070,N_13152);
nor U13291 (N_13291,N_13125,N_13092);
and U13292 (N_13292,N_13009,N_13014);
and U13293 (N_13293,N_13184,N_13115);
nor U13294 (N_13294,N_13022,N_13173);
and U13295 (N_13295,N_13076,N_13096);
or U13296 (N_13296,N_13162,N_13169);
nor U13297 (N_13297,N_13148,N_13079);
nand U13298 (N_13298,N_13055,N_13065);
or U13299 (N_13299,N_13176,N_13077);
nand U13300 (N_13300,N_13045,N_13143);
and U13301 (N_13301,N_13071,N_13067);
and U13302 (N_13302,N_13195,N_13041);
nand U13303 (N_13303,N_13161,N_13159);
xnor U13304 (N_13304,N_13177,N_13109);
or U13305 (N_13305,N_13070,N_13081);
nor U13306 (N_13306,N_13139,N_13123);
nor U13307 (N_13307,N_13174,N_13014);
xnor U13308 (N_13308,N_13055,N_13048);
nand U13309 (N_13309,N_13037,N_13100);
xor U13310 (N_13310,N_13170,N_13169);
or U13311 (N_13311,N_13125,N_13011);
or U13312 (N_13312,N_13163,N_13070);
xor U13313 (N_13313,N_13051,N_13187);
or U13314 (N_13314,N_13088,N_13174);
xor U13315 (N_13315,N_13145,N_13185);
xnor U13316 (N_13316,N_13007,N_13003);
nor U13317 (N_13317,N_13065,N_13032);
or U13318 (N_13318,N_13041,N_13099);
or U13319 (N_13319,N_13046,N_13169);
xnor U13320 (N_13320,N_13153,N_13096);
nand U13321 (N_13321,N_13084,N_13157);
nand U13322 (N_13322,N_13193,N_13081);
nand U13323 (N_13323,N_13068,N_13029);
nand U13324 (N_13324,N_13062,N_13190);
xor U13325 (N_13325,N_13035,N_13155);
nor U13326 (N_13326,N_13133,N_13055);
nand U13327 (N_13327,N_13036,N_13044);
or U13328 (N_13328,N_13014,N_13052);
or U13329 (N_13329,N_13106,N_13123);
nand U13330 (N_13330,N_13063,N_13107);
and U13331 (N_13331,N_13155,N_13015);
xnor U13332 (N_13332,N_13041,N_13118);
xnor U13333 (N_13333,N_13187,N_13098);
and U13334 (N_13334,N_13068,N_13144);
nor U13335 (N_13335,N_13010,N_13099);
xor U13336 (N_13336,N_13189,N_13000);
nand U13337 (N_13337,N_13095,N_13112);
nand U13338 (N_13338,N_13042,N_13099);
xnor U13339 (N_13339,N_13119,N_13173);
and U13340 (N_13340,N_13072,N_13025);
nor U13341 (N_13341,N_13095,N_13044);
nand U13342 (N_13342,N_13138,N_13175);
and U13343 (N_13343,N_13024,N_13141);
xor U13344 (N_13344,N_13031,N_13014);
xor U13345 (N_13345,N_13077,N_13108);
xnor U13346 (N_13346,N_13028,N_13159);
nor U13347 (N_13347,N_13198,N_13128);
xor U13348 (N_13348,N_13057,N_13113);
xor U13349 (N_13349,N_13050,N_13156);
nand U13350 (N_13350,N_13080,N_13016);
nand U13351 (N_13351,N_13130,N_13184);
xor U13352 (N_13352,N_13121,N_13182);
nand U13353 (N_13353,N_13099,N_13184);
xor U13354 (N_13354,N_13022,N_13053);
or U13355 (N_13355,N_13059,N_13129);
or U13356 (N_13356,N_13075,N_13199);
nor U13357 (N_13357,N_13095,N_13165);
nor U13358 (N_13358,N_13151,N_13179);
xnor U13359 (N_13359,N_13180,N_13130);
or U13360 (N_13360,N_13176,N_13144);
and U13361 (N_13361,N_13102,N_13181);
and U13362 (N_13362,N_13151,N_13089);
and U13363 (N_13363,N_13037,N_13079);
nand U13364 (N_13364,N_13101,N_13121);
nor U13365 (N_13365,N_13095,N_13069);
nor U13366 (N_13366,N_13056,N_13164);
nand U13367 (N_13367,N_13046,N_13114);
nor U13368 (N_13368,N_13004,N_13112);
xor U13369 (N_13369,N_13108,N_13184);
and U13370 (N_13370,N_13034,N_13147);
nor U13371 (N_13371,N_13046,N_13193);
and U13372 (N_13372,N_13107,N_13100);
and U13373 (N_13373,N_13053,N_13125);
nand U13374 (N_13374,N_13098,N_13185);
and U13375 (N_13375,N_13085,N_13108);
or U13376 (N_13376,N_13072,N_13010);
nand U13377 (N_13377,N_13180,N_13137);
or U13378 (N_13378,N_13119,N_13133);
and U13379 (N_13379,N_13154,N_13008);
nand U13380 (N_13380,N_13066,N_13003);
nand U13381 (N_13381,N_13174,N_13001);
nand U13382 (N_13382,N_13055,N_13167);
nor U13383 (N_13383,N_13189,N_13035);
and U13384 (N_13384,N_13128,N_13092);
and U13385 (N_13385,N_13106,N_13081);
xnor U13386 (N_13386,N_13198,N_13175);
or U13387 (N_13387,N_13150,N_13176);
and U13388 (N_13388,N_13086,N_13070);
nand U13389 (N_13389,N_13063,N_13088);
nor U13390 (N_13390,N_13152,N_13012);
and U13391 (N_13391,N_13130,N_13012);
or U13392 (N_13392,N_13027,N_13004);
xor U13393 (N_13393,N_13178,N_13083);
and U13394 (N_13394,N_13004,N_13106);
and U13395 (N_13395,N_13194,N_13169);
nand U13396 (N_13396,N_13084,N_13183);
and U13397 (N_13397,N_13151,N_13090);
or U13398 (N_13398,N_13112,N_13042);
xnor U13399 (N_13399,N_13104,N_13165);
or U13400 (N_13400,N_13228,N_13239);
and U13401 (N_13401,N_13246,N_13309);
nand U13402 (N_13402,N_13291,N_13379);
nand U13403 (N_13403,N_13330,N_13249);
nand U13404 (N_13404,N_13332,N_13337);
or U13405 (N_13405,N_13203,N_13304);
and U13406 (N_13406,N_13320,N_13248);
nor U13407 (N_13407,N_13279,N_13206);
or U13408 (N_13408,N_13307,N_13321);
xnor U13409 (N_13409,N_13384,N_13289);
nor U13410 (N_13410,N_13334,N_13361);
or U13411 (N_13411,N_13333,N_13331);
or U13412 (N_13412,N_13340,N_13273);
nand U13413 (N_13413,N_13244,N_13299);
nor U13414 (N_13414,N_13323,N_13342);
nand U13415 (N_13415,N_13281,N_13378);
nor U13416 (N_13416,N_13201,N_13255);
and U13417 (N_13417,N_13352,N_13267);
or U13418 (N_13418,N_13297,N_13218);
xnor U13419 (N_13419,N_13236,N_13354);
or U13420 (N_13420,N_13283,N_13350);
or U13421 (N_13421,N_13393,N_13305);
or U13422 (N_13422,N_13369,N_13306);
nand U13423 (N_13423,N_13371,N_13329);
and U13424 (N_13424,N_13314,N_13359);
xnor U13425 (N_13425,N_13274,N_13343);
nand U13426 (N_13426,N_13229,N_13312);
and U13427 (N_13427,N_13292,N_13336);
and U13428 (N_13428,N_13214,N_13260);
xor U13429 (N_13429,N_13245,N_13385);
nor U13430 (N_13430,N_13327,N_13285);
nand U13431 (N_13431,N_13240,N_13375);
nand U13432 (N_13432,N_13395,N_13315);
and U13433 (N_13433,N_13205,N_13286);
nor U13434 (N_13434,N_13319,N_13234);
nor U13435 (N_13435,N_13364,N_13287);
xor U13436 (N_13436,N_13313,N_13377);
and U13437 (N_13437,N_13356,N_13316);
nor U13438 (N_13438,N_13294,N_13200);
xnor U13439 (N_13439,N_13250,N_13380);
nand U13440 (N_13440,N_13272,N_13398);
and U13441 (N_13441,N_13269,N_13222);
xor U13442 (N_13442,N_13310,N_13278);
nor U13443 (N_13443,N_13325,N_13341);
or U13444 (N_13444,N_13210,N_13280);
and U13445 (N_13445,N_13302,N_13216);
xnor U13446 (N_13446,N_13295,N_13373);
or U13447 (N_13447,N_13290,N_13296);
or U13448 (N_13448,N_13238,N_13293);
xnor U13449 (N_13449,N_13300,N_13265);
xnor U13450 (N_13450,N_13202,N_13360);
nand U13451 (N_13451,N_13243,N_13207);
xor U13452 (N_13452,N_13376,N_13318);
nand U13453 (N_13453,N_13220,N_13317);
nand U13454 (N_13454,N_13308,N_13247);
nand U13455 (N_13455,N_13284,N_13212);
or U13456 (N_13456,N_13399,N_13204);
xnor U13457 (N_13457,N_13357,N_13221);
nor U13458 (N_13458,N_13224,N_13230);
and U13459 (N_13459,N_13282,N_13226);
nand U13460 (N_13460,N_13382,N_13338);
nand U13461 (N_13461,N_13368,N_13241);
and U13462 (N_13462,N_13301,N_13339);
nand U13463 (N_13463,N_13253,N_13387);
nor U13464 (N_13464,N_13367,N_13219);
nor U13465 (N_13465,N_13366,N_13383);
xor U13466 (N_13466,N_13237,N_13355);
or U13467 (N_13467,N_13345,N_13326);
xor U13468 (N_13468,N_13266,N_13348);
nand U13469 (N_13469,N_13217,N_13235);
and U13470 (N_13470,N_13363,N_13381);
nor U13471 (N_13471,N_13372,N_13365);
nor U13472 (N_13472,N_13394,N_13215);
nor U13473 (N_13473,N_13227,N_13258);
and U13474 (N_13474,N_13391,N_13257);
nor U13475 (N_13475,N_13389,N_13263);
and U13476 (N_13476,N_13390,N_13264);
and U13477 (N_13477,N_13259,N_13358);
and U13478 (N_13478,N_13209,N_13271);
nand U13479 (N_13479,N_13277,N_13392);
nor U13480 (N_13480,N_13349,N_13335);
and U13481 (N_13481,N_13353,N_13256);
and U13482 (N_13482,N_13397,N_13362);
or U13483 (N_13483,N_13254,N_13346);
nor U13484 (N_13484,N_13303,N_13396);
nor U13485 (N_13485,N_13324,N_13233);
nand U13486 (N_13486,N_13242,N_13213);
and U13487 (N_13487,N_13261,N_13223);
nand U13488 (N_13488,N_13344,N_13328);
or U13489 (N_13489,N_13374,N_13386);
or U13490 (N_13490,N_13288,N_13275);
nand U13491 (N_13491,N_13211,N_13370);
xor U13492 (N_13492,N_13232,N_13298);
nand U13493 (N_13493,N_13270,N_13311);
xor U13494 (N_13494,N_13231,N_13322);
xnor U13495 (N_13495,N_13351,N_13388);
nor U13496 (N_13496,N_13268,N_13208);
nand U13497 (N_13497,N_13347,N_13252);
nor U13498 (N_13498,N_13225,N_13276);
xnor U13499 (N_13499,N_13251,N_13262);
nor U13500 (N_13500,N_13264,N_13248);
nor U13501 (N_13501,N_13251,N_13331);
nor U13502 (N_13502,N_13310,N_13358);
nor U13503 (N_13503,N_13290,N_13249);
and U13504 (N_13504,N_13360,N_13356);
xnor U13505 (N_13505,N_13296,N_13240);
and U13506 (N_13506,N_13332,N_13338);
and U13507 (N_13507,N_13339,N_13377);
nor U13508 (N_13508,N_13289,N_13254);
nor U13509 (N_13509,N_13230,N_13259);
nor U13510 (N_13510,N_13343,N_13341);
nand U13511 (N_13511,N_13269,N_13388);
xnor U13512 (N_13512,N_13368,N_13305);
nand U13513 (N_13513,N_13308,N_13281);
xnor U13514 (N_13514,N_13362,N_13231);
xor U13515 (N_13515,N_13217,N_13215);
nor U13516 (N_13516,N_13280,N_13204);
nor U13517 (N_13517,N_13249,N_13321);
nor U13518 (N_13518,N_13255,N_13230);
xnor U13519 (N_13519,N_13261,N_13205);
or U13520 (N_13520,N_13302,N_13268);
xor U13521 (N_13521,N_13243,N_13307);
xnor U13522 (N_13522,N_13234,N_13278);
xnor U13523 (N_13523,N_13298,N_13363);
nor U13524 (N_13524,N_13396,N_13223);
nor U13525 (N_13525,N_13272,N_13254);
or U13526 (N_13526,N_13374,N_13349);
or U13527 (N_13527,N_13337,N_13312);
and U13528 (N_13528,N_13356,N_13202);
nand U13529 (N_13529,N_13259,N_13204);
or U13530 (N_13530,N_13291,N_13382);
nand U13531 (N_13531,N_13362,N_13250);
or U13532 (N_13532,N_13359,N_13306);
xor U13533 (N_13533,N_13225,N_13272);
and U13534 (N_13534,N_13291,N_13376);
or U13535 (N_13535,N_13358,N_13327);
nand U13536 (N_13536,N_13363,N_13399);
nand U13537 (N_13537,N_13333,N_13327);
nor U13538 (N_13538,N_13321,N_13326);
or U13539 (N_13539,N_13264,N_13350);
nor U13540 (N_13540,N_13354,N_13233);
or U13541 (N_13541,N_13225,N_13368);
xor U13542 (N_13542,N_13266,N_13260);
and U13543 (N_13543,N_13205,N_13397);
or U13544 (N_13544,N_13386,N_13311);
nor U13545 (N_13545,N_13281,N_13264);
and U13546 (N_13546,N_13294,N_13375);
or U13547 (N_13547,N_13322,N_13378);
and U13548 (N_13548,N_13242,N_13356);
nand U13549 (N_13549,N_13324,N_13303);
nor U13550 (N_13550,N_13244,N_13274);
or U13551 (N_13551,N_13383,N_13368);
or U13552 (N_13552,N_13393,N_13303);
and U13553 (N_13553,N_13396,N_13354);
or U13554 (N_13554,N_13323,N_13252);
nand U13555 (N_13555,N_13296,N_13334);
nor U13556 (N_13556,N_13319,N_13392);
nor U13557 (N_13557,N_13271,N_13230);
or U13558 (N_13558,N_13284,N_13394);
nand U13559 (N_13559,N_13325,N_13324);
or U13560 (N_13560,N_13258,N_13224);
and U13561 (N_13561,N_13224,N_13317);
or U13562 (N_13562,N_13307,N_13266);
nor U13563 (N_13563,N_13369,N_13344);
nor U13564 (N_13564,N_13291,N_13398);
xor U13565 (N_13565,N_13205,N_13276);
xnor U13566 (N_13566,N_13314,N_13237);
and U13567 (N_13567,N_13224,N_13228);
nor U13568 (N_13568,N_13206,N_13337);
nand U13569 (N_13569,N_13322,N_13350);
nor U13570 (N_13570,N_13333,N_13225);
and U13571 (N_13571,N_13268,N_13355);
nand U13572 (N_13572,N_13318,N_13345);
nand U13573 (N_13573,N_13232,N_13397);
xor U13574 (N_13574,N_13264,N_13340);
or U13575 (N_13575,N_13258,N_13252);
xor U13576 (N_13576,N_13378,N_13346);
and U13577 (N_13577,N_13356,N_13255);
nand U13578 (N_13578,N_13361,N_13217);
nand U13579 (N_13579,N_13279,N_13229);
nor U13580 (N_13580,N_13297,N_13311);
nor U13581 (N_13581,N_13208,N_13236);
nand U13582 (N_13582,N_13331,N_13212);
nor U13583 (N_13583,N_13232,N_13367);
nor U13584 (N_13584,N_13322,N_13288);
or U13585 (N_13585,N_13302,N_13322);
nor U13586 (N_13586,N_13282,N_13304);
nor U13587 (N_13587,N_13287,N_13252);
nor U13588 (N_13588,N_13217,N_13335);
and U13589 (N_13589,N_13232,N_13347);
or U13590 (N_13590,N_13328,N_13257);
and U13591 (N_13591,N_13290,N_13303);
and U13592 (N_13592,N_13216,N_13305);
nor U13593 (N_13593,N_13206,N_13320);
nand U13594 (N_13594,N_13349,N_13259);
and U13595 (N_13595,N_13382,N_13355);
nor U13596 (N_13596,N_13276,N_13338);
xnor U13597 (N_13597,N_13277,N_13343);
or U13598 (N_13598,N_13212,N_13316);
or U13599 (N_13599,N_13237,N_13223);
and U13600 (N_13600,N_13462,N_13472);
or U13601 (N_13601,N_13498,N_13434);
xnor U13602 (N_13602,N_13427,N_13523);
xor U13603 (N_13603,N_13587,N_13517);
and U13604 (N_13604,N_13405,N_13572);
xnor U13605 (N_13605,N_13482,N_13538);
and U13606 (N_13606,N_13481,N_13526);
or U13607 (N_13607,N_13590,N_13442);
nand U13608 (N_13608,N_13420,N_13402);
and U13609 (N_13609,N_13528,N_13458);
nor U13610 (N_13610,N_13595,N_13545);
or U13611 (N_13611,N_13469,N_13484);
and U13612 (N_13612,N_13423,N_13502);
xor U13613 (N_13613,N_13553,N_13443);
and U13614 (N_13614,N_13499,N_13519);
nor U13615 (N_13615,N_13480,N_13552);
xor U13616 (N_13616,N_13513,N_13586);
nand U13617 (N_13617,N_13429,N_13467);
nand U13618 (N_13618,N_13589,N_13470);
nand U13619 (N_13619,N_13493,N_13403);
and U13620 (N_13620,N_13419,N_13475);
nand U13621 (N_13621,N_13500,N_13566);
nor U13622 (N_13622,N_13464,N_13497);
xor U13623 (N_13623,N_13571,N_13578);
and U13624 (N_13624,N_13501,N_13400);
nand U13625 (N_13625,N_13486,N_13478);
nand U13626 (N_13626,N_13577,N_13559);
nand U13627 (N_13627,N_13431,N_13556);
nand U13628 (N_13628,N_13522,N_13585);
and U13629 (N_13629,N_13495,N_13460);
and U13630 (N_13630,N_13409,N_13448);
nor U13631 (N_13631,N_13598,N_13451);
or U13632 (N_13632,N_13562,N_13537);
xor U13633 (N_13633,N_13567,N_13547);
and U13634 (N_13634,N_13592,N_13539);
or U13635 (N_13635,N_13490,N_13516);
xnor U13636 (N_13636,N_13555,N_13591);
or U13637 (N_13637,N_13540,N_13452);
or U13638 (N_13638,N_13548,N_13574);
and U13639 (N_13639,N_13441,N_13444);
xor U13640 (N_13640,N_13426,N_13487);
nor U13641 (N_13641,N_13542,N_13473);
xor U13642 (N_13642,N_13477,N_13508);
xor U13643 (N_13643,N_13581,N_13417);
or U13644 (N_13644,N_13465,N_13468);
nor U13645 (N_13645,N_13558,N_13489);
or U13646 (N_13646,N_13597,N_13525);
nand U13647 (N_13647,N_13579,N_13410);
nand U13648 (N_13648,N_13575,N_13549);
xnor U13649 (N_13649,N_13536,N_13492);
or U13650 (N_13650,N_13424,N_13569);
nor U13651 (N_13651,N_13433,N_13425);
nor U13652 (N_13652,N_13401,N_13404);
or U13653 (N_13653,N_13599,N_13584);
xor U13654 (N_13654,N_13514,N_13412);
xnor U13655 (N_13655,N_13479,N_13494);
nand U13656 (N_13656,N_13518,N_13594);
or U13657 (N_13657,N_13456,N_13532);
or U13658 (N_13658,N_13459,N_13439);
xnor U13659 (N_13659,N_13413,N_13580);
and U13660 (N_13660,N_13560,N_13557);
or U13661 (N_13661,N_13507,N_13406);
nor U13662 (N_13662,N_13440,N_13534);
xor U13663 (N_13663,N_13438,N_13471);
and U13664 (N_13664,N_13568,N_13411);
and U13665 (N_13665,N_13466,N_13582);
or U13666 (N_13666,N_13563,N_13415);
xor U13667 (N_13667,N_13504,N_13445);
nand U13668 (N_13668,N_13461,N_13463);
and U13669 (N_13669,N_13488,N_13449);
or U13670 (N_13670,N_13550,N_13446);
xnor U13671 (N_13671,N_13483,N_13455);
nand U13672 (N_13672,N_13533,N_13437);
and U13673 (N_13673,N_13509,N_13551);
xnor U13674 (N_13674,N_13512,N_13503);
nand U13675 (N_13675,N_13447,N_13596);
and U13676 (N_13676,N_13529,N_13521);
nand U13677 (N_13677,N_13476,N_13408);
or U13678 (N_13678,N_13583,N_13546);
xor U13679 (N_13679,N_13506,N_13418);
xor U13680 (N_13680,N_13421,N_13531);
nor U13681 (N_13681,N_13511,N_13570);
nor U13682 (N_13682,N_13430,N_13544);
and U13683 (N_13683,N_13474,N_13496);
and U13684 (N_13684,N_13593,N_13454);
nor U13685 (N_13685,N_13524,N_13414);
nor U13686 (N_13686,N_13564,N_13565);
and U13687 (N_13687,N_13527,N_13457);
nor U13688 (N_13688,N_13407,N_13561);
and U13689 (N_13689,N_13428,N_13515);
xor U13690 (N_13690,N_13535,N_13588);
xnor U13691 (N_13691,N_13416,N_13510);
xor U13692 (N_13692,N_13573,N_13450);
nor U13693 (N_13693,N_13505,N_13422);
or U13694 (N_13694,N_13520,N_13576);
nand U13695 (N_13695,N_13436,N_13541);
nand U13696 (N_13696,N_13435,N_13543);
nand U13697 (N_13697,N_13491,N_13453);
nand U13698 (N_13698,N_13485,N_13530);
nand U13699 (N_13699,N_13554,N_13432);
nand U13700 (N_13700,N_13417,N_13430);
or U13701 (N_13701,N_13507,N_13525);
or U13702 (N_13702,N_13436,N_13424);
or U13703 (N_13703,N_13433,N_13448);
or U13704 (N_13704,N_13471,N_13430);
nand U13705 (N_13705,N_13550,N_13564);
nor U13706 (N_13706,N_13411,N_13483);
and U13707 (N_13707,N_13571,N_13502);
and U13708 (N_13708,N_13509,N_13595);
or U13709 (N_13709,N_13554,N_13513);
nand U13710 (N_13710,N_13529,N_13551);
xor U13711 (N_13711,N_13524,N_13518);
xnor U13712 (N_13712,N_13469,N_13414);
or U13713 (N_13713,N_13516,N_13419);
or U13714 (N_13714,N_13597,N_13524);
and U13715 (N_13715,N_13477,N_13571);
and U13716 (N_13716,N_13400,N_13575);
xnor U13717 (N_13717,N_13446,N_13441);
or U13718 (N_13718,N_13531,N_13597);
or U13719 (N_13719,N_13487,N_13534);
and U13720 (N_13720,N_13571,N_13543);
and U13721 (N_13721,N_13571,N_13450);
xor U13722 (N_13722,N_13446,N_13574);
nor U13723 (N_13723,N_13445,N_13474);
or U13724 (N_13724,N_13513,N_13597);
nor U13725 (N_13725,N_13431,N_13563);
nand U13726 (N_13726,N_13536,N_13451);
xor U13727 (N_13727,N_13517,N_13554);
xnor U13728 (N_13728,N_13449,N_13404);
nor U13729 (N_13729,N_13446,N_13557);
nand U13730 (N_13730,N_13513,N_13524);
nand U13731 (N_13731,N_13559,N_13468);
nand U13732 (N_13732,N_13478,N_13451);
or U13733 (N_13733,N_13478,N_13530);
or U13734 (N_13734,N_13412,N_13436);
or U13735 (N_13735,N_13551,N_13517);
and U13736 (N_13736,N_13434,N_13530);
xor U13737 (N_13737,N_13493,N_13489);
nor U13738 (N_13738,N_13438,N_13491);
or U13739 (N_13739,N_13555,N_13589);
and U13740 (N_13740,N_13487,N_13520);
xor U13741 (N_13741,N_13553,N_13573);
and U13742 (N_13742,N_13412,N_13545);
nor U13743 (N_13743,N_13455,N_13402);
nor U13744 (N_13744,N_13484,N_13569);
nor U13745 (N_13745,N_13400,N_13430);
or U13746 (N_13746,N_13553,N_13476);
nand U13747 (N_13747,N_13432,N_13413);
or U13748 (N_13748,N_13483,N_13555);
nor U13749 (N_13749,N_13561,N_13494);
xor U13750 (N_13750,N_13588,N_13521);
nand U13751 (N_13751,N_13430,N_13408);
nor U13752 (N_13752,N_13588,N_13412);
xnor U13753 (N_13753,N_13452,N_13480);
nor U13754 (N_13754,N_13482,N_13465);
nand U13755 (N_13755,N_13542,N_13459);
or U13756 (N_13756,N_13448,N_13545);
and U13757 (N_13757,N_13498,N_13532);
nor U13758 (N_13758,N_13450,N_13559);
xnor U13759 (N_13759,N_13516,N_13472);
or U13760 (N_13760,N_13446,N_13502);
xor U13761 (N_13761,N_13568,N_13466);
and U13762 (N_13762,N_13572,N_13590);
and U13763 (N_13763,N_13461,N_13552);
and U13764 (N_13764,N_13406,N_13407);
nor U13765 (N_13765,N_13502,N_13543);
xor U13766 (N_13766,N_13438,N_13413);
nand U13767 (N_13767,N_13484,N_13548);
and U13768 (N_13768,N_13543,N_13494);
nand U13769 (N_13769,N_13579,N_13550);
and U13770 (N_13770,N_13536,N_13522);
nor U13771 (N_13771,N_13538,N_13572);
nand U13772 (N_13772,N_13519,N_13584);
nor U13773 (N_13773,N_13449,N_13458);
xnor U13774 (N_13774,N_13577,N_13519);
nand U13775 (N_13775,N_13429,N_13468);
xor U13776 (N_13776,N_13590,N_13402);
and U13777 (N_13777,N_13584,N_13514);
xnor U13778 (N_13778,N_13428,N_13568);
and U13779 (N_13779,N_13563,N_13487);
xnor U13780 (N_13780,N_13435,N_13493);
nor U13781 (N_13781,N_13525,N_13476);
nor U13782 (N_13782,N_13469,N_13514);
xor U13783 (N_13783,N_13574,N_13424);
nor U13784 (N_13784,N_13406,N_13514);
nand U13785 (N_13785,N_13444,N_13583);
nand U13786 (N_13786,N_13475,N_13444);
nand U13787 (N_13787,N_13464,N_13588);
or U13788 (N_13788,N_13558,N_13447);
and U13789 (N_13789,N_13571,N_13559);
and U13790 (N_13790,N_13588,N_13458);
nand U13791 (N_13791,N_13505,N_13487);
and U13792 (N_13792,N_13489,N_13479);
and U13793 (N_13793,N_13595,N_13598);
nor U13794 (N_13794,N_13548,N_13528);
nand U13795 (N_13795,N_13484,N_13468);
and U13796 (N_13796,N_13599,N_13509);
nor U13797 (N_13797,N_13575,N_13529);
and U13798 (N_13798,N_13400,N_13595);
nand U13799 (N_13799,N_13509,N_13593);
or U13800 (N_13800,N_13717,N_13625);
or U13801 (N_13801,N_13653,N_13737);
nor U13802 (N_13802,N_13630,N_13643);
or U13803 (N_13803,N_13740,N_13718);
and U13804 (N_13804,N_13699,N_13770);
xor U13805 (N_13805,N_13602,N_13750);
nand U13806 (N_13806,N_13725,N_13670);
nor U13807 (N_13807,N_13722,N_13700);
nand U13808 (N_13808,N_13655,N_13787);
and U13809 (N_13809,N_13771,N_13743);
or U13810 (N_13810,N_13615,N_13617);
or U13811 (N_13811,N_13603,N_13776);
xnor U13812 (N_13812,N_13632,N_13606);
nand U13813 (N_13813,N_13792,N_13605);
nand U13814 (N_13814,N_13600,N_13634);
and U13815 (N_13815,N_13721,N_13692);
or U13816 (N_13816,N_13616,N_13646);
or U13817 (N_13817,N_13611,N_13618);
nand U13818 (N_13818,N_13635,N_13773);
xor U13819 (N_13819,N_13642,N_13759);
nor U13820 (N_13820,N_13620,N_13755);
and U13821 (N_13821,N_13720,N_13652);
xnor U13822 (N_13822,N_13724,N_13681);
xnor U13823 (N_13823,N_13650,N_13629);
or U13824 (N_13824,N_13664,N_13744);
or U13825 (N_13825,N_13685,N_13715);
xor U13826 (N_13826,N_13628,N_13785);
and U13827 (N_13827,N_13768,N_13799);
and U13828 (N_13828,N_13788,N_13619);
nand U13829 (N_13829,N_13735,N_13703);
xor U13830 (N_13830,N_13648,N_13601);
or U13831 (N_13831,N_13647,N_13779);
nand U13832 (N_13832,N_13610,N_13623);
and U13833 (N_13833,N_13797,N_13730);
xnor U13834 (N_13834,N_13680,N_13775);
xor U13835 (N_13835,N_13752,N_13665);
nor U13836 (N_13836,N_13783,N_13733);
nor U13837 (N_13837,N_13649,N_13687);
xnor U13838 (N_13838,N_13660,N_13696);
nor U13839 (N_13839,N_13753,N_13702);
or U13840 (N_13840,N_13636,N_13672);
and U13841 (N_13841,N_13645,N_13719);
or U13842 (N_13842,N_13693,N_13608);
nor U13843 (N_13843,N_13641,N_13777);
and U13844 (N_13844,N_13637,N_13612);
nor U13845 (N_13845,N_13661,N_13690);
xor U13846 (N_13846,N_13677,N_13631);
nor U13847 (N_13847,N_13626,N_13604);
or U13848 (N_13848,N_13711,N_13644);
nand U13849 (N_13849,N_13746,N_13607);
nand U13850 (N_13850,N_13682,N_13749);
or U13851 (N_13851,N_13688,N_13684);
and U13852 (N_13852,N_13723,N_13669);
nand U13853 (N_13853,N_13728,N_13657);
xnor U13854 (N_13854,N_13760,N_13784);
and U13855 (N_13855,N_13621,N_13751);
and U13856 (N_13856,N_13736,N_13676);
nor U13857 (N_13857,N_13763,N_13698);
nand U13858 (N_13858,N_13782,N_13683);
nand U13859 (N_13859,N_13747,N_13795);
and U13860 (N_13860,N_13761,N_13614);
and U13861 (N_13861,N_13691,N_13732);
or U13862 (N_13862,N_13673,N_13624);
and U13863 (N_13863,N_13609,N_13695);
xnor U13864 (N_13864,N_13796,N_13706);
nand U13865 (N_13865,N_13769,N_13686);
xor U13866 (N_13866,N_13671,N_13668);
nand U13867 (N_13867,N_13716,N_13758);
or U13868 (N_13868,N_13790,N_13662);
xnor U13869 (N_13869,N_13633,N_13767);
nand U13870 (N_13870,N_13638,N_13748);
xor U13871 (N_13871,N_13663,N_13741);
nor U13872 (N_13872,N_13780,N_13651);
and U13873 (N_13873,N_13734,N_13764);
nor U13874 (N_13874,N_13708,N_13731);
and U13875 (N_13875,N_13674,N_13778);
nor U13876 (N_13876,N_13710,N_13622);
nor U13877 (N_13877,N_13754,N_13772);
nand U13878 (N_13878,N_13738,N_13656);
xor U13879 (N_13879,N_13667,N_13781);
or U13880 (N_13880,N_13639,N_13697);
or U13881 (N_13881,N_13679,N_13745);
and U13882 (N_13882,N_13659,N_13705);
nand U13883 (N_13883,N_13627,N_13678);
nor U13884 (N_13884,N_13712,N_13713);
or U13885 (N_13885,N_13704,N_13786);
nor U13886 (N_13886,N_13726,N_13765);
nand U13887 (N_13887,N_13701,N_13727);
or U13888 (N_13888,N_13729,N_13757);
or U13889 (N_13889,N_13709,N_13742);
or U13890 (N_13890,N_13640,N_13658);
or U13891 (N_13891,N_13794,N_13675);
or U13892 (N_13892,N_13694,N_13789);
nand U13893 (N_13893,N_13762,N_13793);
nor U13894 (N_13894,N_13791,N_13756);
and U13895 (N_13895,N_13689,N_13739);
nor U13896 (N_13896,N_13766,N_13774);
or U13897 (N_13897,N_13707,N_13613);
xor U13898 (N_13898,N_13666,N_13798);
and U13899 (N_13899,N_13714,N_13654);
or U13900 (N_13900,N_13610,N_13675);
nand U13901 (N_13901,N_13761,N_13634);
xnor U13902 (N_13902,N_13788,N_13705);
nand U13903 (N_13903,N_13716,N_13664);
or U13904 (N_13904,N_13731,N_13728);
xor U13905 (N_13905,N_13678,N_13637);
or U13906 (N_13906,N_13666,N_13605);
nand U13907 (N_13907,N_13678,N_13705);
nor U13908 (N_13908,N_13623,N_13693);
nand U13909 (N_13909,N_13621,N_13778);
or U13910 (N_13910,N_13784,N_13798);
and U13911 (N_13911,N_13605,N_13641);
nand U13912 (N_13912,N_13619,N_13729);
xnor U13913 (N_13913,N_13651,N_13663);
nor U13914 (N_13914,N_13680,N_13665);
xor U13915 (N_13915,N_13781,N_13743);
xnor U13916 (N_13916,N_13642,N_13623);
xor U13917 (N_13917,N_13698,N_13749);
xor U13918 (N_13918,N_13612,N_13628);
nor U13919 (N_13919,N_13647,N_13790);
nand U13920 (N_13920,N_13741,N_13611);
nor U13921 (N_13921,N_13733,N_13700);
xnor U13922 (N_13922,N_13746,N_13656);
nand U13923 (N_13923,N_13657,N_13704);
nor U13924 (N_13924,N_13780,N_13689);
or U13925 (N_13925,N_13602,N_13680);
or U13926 (N_13926,N_13612,N_13693);
xnor U13927 (N_13927,N_13674,N_13668);
nor U13928 (N_13928,N_13709,N_13776);
nand U13929 (N_13929,N_13615,N_13603);
and U13930 (N_13930,N_13777,N_13697);
nand U13931 (N_13931,N_13690,N_13784);
nor U13932 (N_13932,N_13624,N_13687);
or U13933 (N_13933,N_13687,N_13627);
or U13934 (N_13934,N_13750,N_13660);
nor U13935 (N_13935,N_13708,N_13779);
nor U13936 (N_13936,N_13680,N_13723);
xnor U13937 (N_13937,N_13700,N_13784);
nand U13938 (N_13938,N_13712,N_13714);
nor U13939 (N_13939,N_13728,N_13664);
or U13940 (N_13940,N_13639,N_13751);
nor U13941 (N_13941,N_13663,N_13739);
and U13942 (N_13942,N_13683,N_13753);
nand U13943 (N_13943,N_13668,N_13788);
nand U13944 (N_13944,N_13719,N_13690);
nand U13945 (N_13945,N_13702,N_13751);
nand U13946 (N_13946,N_13791,N_13684);
nand U13947 (N_13947,N_13763,N_13778);
nor U13948 (N_13948,N_13705,N_13628);
nor U13949 (N_13949,N_13697,N_13629);
and U13950 (N_13950,N_13708,N_13739);
nor U13951 (N_13951,N_13644,N_13710);
and U13952 (N_13952,N_13735,N_13604);
nor U13953 (N_13953,N_13623,N_13753);
and U13954 (N_13954,N_13685,N_13710);
nor U13955 (N_13955,N_13678,N_13602);
and U13956 (N_13956,N_13723,N_13697);
nor U13957 (N_13957,N_13652,N_13756);
nor U13958 (N_13958,N_13761,N_13788);
nand U13959 (N_13959,N_13768,N_13634);
xor U13960 (N_13960,N_13660,N_13732);
nor U13961 (N_13961,N_13781,N_13735);
nor U13962 (N_13962,N_13689,N_13604);
xnor U13963 (N_13963,N_13641,N_13797);
or U13964 (N_13964,N_13633,N_13766);
xnor U13965 (N_13965,N_13681,N_13798);
nand U13966 (N_13966,N_13671,N_13636);
nor U13967 (N_13967,N_13649,N_13699);
xor U13968 (N_13968,N_13666,N_13682);
xor U13969 (N_13969,N_13788,N_13650);
and U13970 (N_13970,N_13624,N_13778);
nand U13971 (N_13971,N_13668,N_13713);
nor U13972 (N_13972,N_13764,N_13759);
nand U13973 (N_13973,N_13763,N_13659);
nor U13974 (N_13974,N_13685,N_13687);
xnor U13975 (N_13975,N_13756,N_13650);
nor U13976 (N_13976,N_13724,N_13605);
xor U13977 (N_13977,N_13705,N_13734);
nand U13978 (N_13978,N_13606,N_13659);
nand U13979 (N_13979,N_13637,N_13751);
and U13980 (N_13980,N_13617,N_13752);
and U13981 (N_13981,N_13623,N_13734);
and U13982 (N_13982,N_13694,N_13710);
and U13983 (N_13983,N_13780,N_13756);
and U13984 (N_13984,N_13608,N_13741);
or U13985 (N_13985,N_13700,N_13695);
nor U13986 (N_13986,N_13647,N_13747);
nand U13987 (N_13987,N_13739,N_13678);
or U13988 (N_13988,N_13629,N_13646);
nor U13989 (N_13989,N_13767,N_13786);
and U13990 (N_13990,N_13675,N_13630);
xor U13991 (N_13991,N_13637,N_13775);
and U13992 (N_13992,N_13747,N_13727);
nand U13993 (N_13993,N_13725,N_13612);
nand U13994 (N_13994,N_13724,N_13705);
nor U13995 (N_13995,N_13732,N_13635);
nor U13996 (N_13996,N_13774,N_13664);
nand U13997 (N_13997,N_13736,N_13649);
nor U13998 (N_13998,N_13695,N_13744);
or U13999 (N_13999,N_13628,N_13650);
nor U14000 (N_14000,N_13884,N_13921);
and U14001 (N_14001,N_13870,N_13915);
nor U14002 (N_14002,N_13866,N_13999);
or U14003 (N_14003,N_13904,N_13907);
or U14004 (N_14004,N_13824,N_13983);
xnor U14005 (N_14005,N_13997,N_13965);
or U14006 (N_14006,N_13917,N_13889);
or U14007 (N_14007,N_13931,N_13814);
nand U14008 (N_14008,N_13908,N_13918);
nor U14009 (N_14009,N_13985,N_13869);
xor U14010 (N_14010,N_13909,N_13805);
nor U14011 (N_14011,N_13945,N_13966);
xnor U14012 (N_14012,N_13850,N_13820);
nand U14013 (N_14013,N_13925,N_13877);
and U14014 (N_14014,N_13808,N_13880);
nor U14015 (N_14015,N_13988,N_13943);
xnor U14016 (N_14016,N_13937,N_13922);
nand U14017 (N_14017,N_13950,N_13926);
nand U14018 (N_14018,N_13991,N_13848);
xor U14019 (N_14019,N_13989,N_13829);
nor U14020 (N_14020,N_13971,N_13847);
and U14021 (N_14021,N_13845,N_13809);
xnor U14022 (N_14022,N_13895,N_13978);
nand U14023 (N_14023,N_13894,N_13810);
xor U14024 (N_14024,N_13876,N_13896);
nand U14025 (N_14025,N_13942,N_13812);
xor U14026 (N_14026,N_13963,N_13835);
nand U14027 (N_14027,N_13928,N_13984);
nand U14028 (N_14028,N_13929,N_13952);
xnor U14029 (N_14029,N_13864,N_13806);
nand U14030 (N_14030,N_13944,N_13886);
xnor U14031 (N_14031,N_13927,N_13957);
or U14032 (N_14032,N_13879,N_13953);
or U14033 (N_14033,N_13804,N_13939);
xor U14034 (N_14034,N_13843,N_13856);
or U14035 (N_14035,N_13972,N_13802);
or U14036 (N_14036,N_13818,N_13958);
xnor U14037 (N_14037,N_13852,N_13967);
nand U14038 (N_14038,N_13891,N_13867);
and U14039 (N_14039,N_13977,N_13872);
nand U14040 (N_14040,N_13893,N_13949);
xnor U14041 (N_14041,N_13849,N_13823);
or U14042 (N_14042,N_13834,N_13962);
nand U14043 (N_14043,N_13955,N_13956);
nand U14044 (N_14044,N_13998,N_13913);
xor U14045 (N_14045,N_13844,N_13923);
xor U14046 (N_14046,N_13946,N_13853);
and U14047 (N_14047,N_13947,N_13873);
nand U14048 (N_14048,N_13826,N_13800);
xor U14049 (N_14049,N_13881,N_13861);
nor U14050 (N_14050,N_13885,N_13898);
nor U14051 (N_14051,N_13875,N_13865);
xor U14052 (N_14052,N_13961,N_13831);
nor U14053 (N_14053,N_13816,N_13906);
or U14054 (N_14054,N_13839,N_13980);
or U14055 (N_14055,N_13897,N_13903);
nand U14056 (N_14056,N_13899,N_13951);
xnor U14057 (N_14057,N_13924,N_13874);
xor U14058 (N_14058,N_13887,N_13973);
nand U14059 (N_14059,N_13836,N_13854);
nand U14060 (N_14060,N_13914,N_13832);
nor U14061 (N_14061,N_13828,N_13916);
xnor U14062 (N_14062,N_13868,N_13933);
nand U14063 (N_14063,N_13911,N_13871);
or U14064 (N_14064,N_13968,N_13846);
nor U14065 (N_14065,N_13910,N_13859);
nand U14066 (N_14066,N_13930,N_13993);
xor U14067 (N_14067,N_13982,N_13841);
and U14068 (N_14068,N_13935,N_13815);
nor U14069 (N_14069,N_13981,N_13919);
nand U14070 (N_14070,N_13940,N_13964);
or U14071 (N_14071,N_13905,N_13838);
xor U14072 (N_14072,N_13822,N_13948);
nor U14073 (N_14073,N_13842,N_13979);
and U14074 (N_14074,N_13862,N_13996);
nor U14075 (N_14075,N_13860,N_13901);
nand U14076 (N_14076,N_13890,N_13830);
and U14077 (N_14077,N_13851,N_13882);
xor U14078 (N_14078,N_13994,N_13819);
and U14079 (N_14079,N_13986,N_13932);
or U14080 (N_14080,N_13878,N_13813);
xnor U14081 (N_14081,N_13920,N_13987);
nor U14082 (N_14082,N_13938,N_13954);
nor U14083 (N_14083,N_13833,N_13960);
xnor U14084 (N_14084,N_13827,N_13888);
nand U14085 (N_14085,N_13941,N_13934);
or U14086 (N_14086,N_13840,N_13990);
or U14087 (N_14087,N_13821,N_13975);
or U14088 (N_14088,N_13936,N_13976);
xnor U14089 (N_14089,N_13825,N_13807);
nand U14090 (N_14090,N_13855,N_13969);
and U14091 (N_14091,N_13857,N_13858);
and U14092 (N_14092,N_13995,N_13974);
nor U14093 (N_14093,N_13892,N_13900);
nor U14094 (N_14094,N_13992,N_13970);
nor U14095 (N_14095,N_13959,N_13863);
xor U14096 (N_14096,N_13811,N_13837);
xnor U14097 (N_14097,N_13912,N_13803);
or U14098 (N_14098,N_13801,N_13883);
xor U14099 (N_14099,N_13817,N_13902);
nor U14100 (N_14100,N_13984,N_13833);
nor U14101 (N_14101,N_13999,N_13891);
or U14102 (N_14102,N_13949,N_13901);
xnor U14103 (N_14103,N_13830,N_13852);
nor U14104 (N_14104,N_13969,N_13900);
nor U14105 (N_14105,N_13833,N_13835);
and U14106 (N_14106,N_13928,N_13927);
nor U14107 (N_14107,N_13951,N_13921);
and U14108 (N_14108,N_13803,N_13883);
nor U14109 (N_14109,N_13945,N_13982);
nor U14110 (N_14110,N_13887,N_13953);
xnor U14111 (N_14111,N_13905,N_13987);
or U14112 (N_14112,N_13802,N_13890);
nand U14113 (N_14113,N_13913,N_13906);
nand U14114 (N_14114,N_13834,N_13976);
nor U14115 (N_14115,N_13870,N_13897);
xor U14116 (N_14116,N_13969,N_13886);
and U14117 (N_14117,N_13983,N_13931);
xor U14118 (N_14118,N_13869,N_13804);
nor U14119 (N_14119,N_13971,N_13950);
and U14120 (N_14120,N_13844,N_13852);
xor U14121 (N_14121,N_13892,N_13861);
or U14122 (N_14122,N_13992,N_13987);
or U14123 (N_14123,N_13959,N_13938);
nor U14124 (N_14124,N_13975,N_13865);
nand U14125 (N_14125,N_13856,N_13999);
or U14126 (N_14126,N_13918,N_13890);
nand U14127 (N_14127,N_13847,N_13833);
nor U14128 (N_14128,N_13837,N_13812);
nor U14129 (N_14129,N_13938,N_13845);
nor U14130 (N_14130,N_13868,N_13802);
or U14131 (N_14131,N_13925,N_13894);
and U14132 (N_14132,N_13868,N_13991);
nor U14133 (N_14133,N_13891,N_13893);
nor U14134 (N_14134,N_13968,N_13969);
xnor U14135 (N_14135,N_13987,N_13933);
nand U14136 (N_14136,N_13985,N_13880);
nand U14137 (N_14137,N_13943,N_13877);
nor U14138 (N_14138,N_13993,N_13851);
nand U14139 (N_14139,N_13948,N_13983);
and U14140 (N_14140,N_13902,N_13920);
or U14141 (N_14141,N_13841,N_13804);
or U14142 (N_14142,N_13918,N_13895);
xor U14143 (N_14143,N_13801,N_13843);
nor U14144 (N_14144,N_13886,N_13804);
nor U14145 (N_14145,N_13844,N_13884);
nor U14146 (N_14146,N_13851,N_13964);
and U14147 (N_14147,N_13995,N_13939);
nor U14148 (N_14148,N_13823,N_13899);
nand U14149 (N_14149,N_13854,N_13873);
or U14150 (N_14150,N_13850,N_13871);
xor U14151 (N_14151,N_13980,N_13957);
and U14152 (N_14152,N_13835,N_13918);
nor U14153 (N_14153,N_13892,N_13867);
nand U14154 (N_14154,N_13964,N_13899);
nand U14155 (N_14155,N_13851,N_13802);
nand U14156 (N_14156,N_13937,N_13889);
xnor U14157 (N_14157,N_13824,N_13969);
nor U14158 (N_14158,N_13871,N_13987);
nor U14159 (N_14159,N_13880,N_13943);
nor U14160 (N_14160,N_13833,N_13804);
xnor U14161 (N_14161,N_13856,N_13971);
and U14162 (N_14162,N_13836,N_13991);
xnor U14163 (N_14163,N_13928,N_13925);
nand U14164 (N_14164,N_13945,N_13991);
nor U14165 (N_14165,N_13986,N_13921);
xnor U14166 (N_14166,N_13836,N_13862);
xnor U14167 (N_14167,N_13810,N_13888);
nor U14168 (N_14168,N_13808,N_13989);
nand U14169 (N_14169,N_13847,N_13899);
or U14170 (N_14170,N_13845,N_13891);
nand U14171 (N_14171,N_13897,N_13834);
nor U14172 (N_14172,N_13883,N_13946);
and U14173 (N_14173,N_13872,N_13899);
or U14174 (N_14174,N_13980,N_13842);
or U14175 (N_14175,N_13968,N_13879);
xor U14176 (N_14176,N_13850,N_13869);
nor U14177 (N_14177,N_13860,N_13985);
xnor U14178 (N_14178,N_13831,N_13829);
or U14179 (N_14179,N_13897,N_13985);
nand U14180 (N_14180,N_13850,N_13930);
xor U14181 (N_14181,N_13826,N_13879);
or U14182 (N_14182,N_13944,N_13898);
and U14183 (N_14183,N_13973,N_13952);
nand U14184 (N_14184,N_13845,N_13823);
or U14185 (N_14185,N_13825,N_13895);
nand U14186 (N_14186,N_13907,N_13998);
and U14187 (N_14187,N_13986,N_13819);
and U14188 (N_14188,N_13858,N_13925);
or U14189 (N_14189,N_13966,N_13920);
nor U14190 (N_14190,N_13867,N_13979);
or U14191 (N_14191,N_13980,N_13891);
nand U14192 (N_14192,N_13818,N_13893);
nor U14193 (N_14193,N_13943,N_13974);
nand U14194 (N_14194,N_13943,N_13808);
or U14195 (N_14195,N_13889,N_13819);
nand U14196 (N_14196,N_13832,N_13906);
xor U14197 (N_14197,N_13809,N_13952);
nor U14198 (N_14198,N_13813,N_13873);
nand U14199 (N_14199,N_13895,N_13955);
and U14200 (N_14200,N_14101,N_14057);
nor U14201 (N_14201,N_14027,N_14130);
nand U14202 (N_14202,N_14131,N_14105);
nand U14203 (N_14203,N_14189,N_14030);
or U14204 (N_14204,N_14185,N_14049);
xor U14205 (N_14205,N_14113,N_14160);
nand U14206 (N_14206,N_14088,N_14174);
or U14207 (N_14207,N_14079,N_14043);
or U14208 (N_14208,N_14186,N_14070);
or U14209 (N_14209,N_14072,N_14129);
or U14210 (N_14210,N_14055,N_14000);
and U14211 (N_14211,N_14173,N_14059);
xnor U14212 (N_14212,N_14022,N_14050);
nand U14213 (N_14213,N_14077,N_14047);
or U14214 (N_14214,N_14006,N_14074);
or U14215 (N_14215,N_14081,N_14182);
nor U14216 (N_14216,N_14147,N_14175);
nand U14217 (N_14217,N_14149,N_14142);
nand U14218 (N_14218,N_14075,N_14112);
or U14219 (N_14219,N_14126,N_14107);
xor U14220 (N_14220,N_14051,N_14148);
nand U14221 (N_14221,N_14120,N_14013);
nand U14222 (N_14222,N_14183,N_14082);
or U14223 (N_14223,N_14090,N_14080);
xnor U14224 (N_14224,N_14008,N_14170);
and U14225 (N_14225,N_14018,N_14195);
nand U14226 (N_14226,N_14196,N_14181);
or U14227 (N_14227,N_14172,N_14024);
or U14228 (N_14228,N_14119,N_14128);
or U14229 (N_14229,N_14188,N_14110);
nor U14230 (N_14230,N_14028,N_14062);
or U14231 (N_14231,N_14092,N_14121);
and U14232 (N_14232,N_14056,N_14089);
and U14233 (N_14233,N_14083,N_14033);
xor U14234 (N_14234,N_14073,N_14031);
and U14235 (N_14235,N_14199,N_14054);
nand U14236 (N_14236,N_14168,N_14011);
xnor U14237 (N_14237,N_14178,N_14005);
nand U14238 (N_14238,N_14171,N_14094);
nand U14239 (N_14239,N_14015,N_14058);
or U14240 (N_14240,N_14026,N_14097);
xor U14241 (N_14241,N_14103,N_14091);
nor U14242 (N_14242,N_14125,N_14066);
xnor U14243 (N_14243,N_14020,N_14150);
and U14244 (N_14244,N_14136,N_14108);
or U14245 (N_14245,N_14085,N_14095);
nor U14246 (N_14246,N_14102,N_14084);
nor U14247 (N_14247,N_14025,N_14064);
nor U14248 (N_14248,N_14063,N_14179);
nor U14249 (N_14249,N_14021,N_14145);
nand U14250 (N_14250,N_14190,N_14096);
nor U14251 (N_14251,N_14001,N_14193);
nand U14252 (N_14252,N_14019,N_14122);
and U14253 (N_14253,N_14032,N_14042);
nor U14254 (N_14254,N_14109,N_14146);
nor U14255 (N_14255,N_14127,N_14071);
and U14256 (N_14256,N_14036,N_14065);
and U14257 (N_14257,N_14176,N_14144);
xor U14258 (N_14258,N_14093,N_14117);
nor U14259 (N_14259,N_14163,N_14133);
nor U14260 (N_14260,N_14053,N_14039);
or U14261 (N_14261,N_14154,N_14157);
nor U14262 (N_14262,N_14029,N_14135);
and U14263 (N_14263,N_14158,N_14007);
xnor U14264 (N_14264,N_14106,N_14187);
xnor U14265 (N_14265,N_14184,N_14132);
and U14266 (N_14266,N_14139,N_14061);
and U14267 (N_14267,N_14035,N_14010);
nor U14268 (N_14268,N_14044,N_14004);
and U14269 (N_14269,N_14152,N_14155);
nor U14270 (N_14270,N_14137,N_14164);
nand U14271 (N_14271,N_14040,N_14014);
nor U14272 (N_14272,N_14098,N_14076);
and U14273 (N_14273,N_14177,N_14017);
nor U14274 (N_14274,N_14140,N_14115);
nand U14275 (N_14275,N_14104,N_14041);
nand U14276 (N_14276,N_14161,N_14099);
nor U14277 (N_14277,N_14009,N_14169);
and U14278 (N_14278,N_14111,N_14034);
nand U14279 (N_14279,N_14141,N_14123);
nand U14280 (N_14280,N_14012,N_14198);
and U14281 (N_14281,N_14023,N_14060);
nor U14282 (N_14282,N_14143,N_14067);
xor U14283 (N_14283,N_14086,N_14191);
and U14284 (N_14284,N_14052,N_14046);
and U14285 (N_14285,N_14087,N_14003);
and U14286 (N_14286,N_14165,N_14194);
xnor U14287 (N_14287,N_14138,N_14069);
and U14288 (N_14288,N_14068,N_14153);
nor U14289 (N_14289,N_14197,N_14038);
nand U14290 (N_14290,N_14037,N_14045);
or U14291 (N_14291,N_14192,N_14162);
xor U14292 (N_14292,N_14156,N_14124);
nand U14293 (N_14293,N_14078,N_14159);
or U14294 (N_14294,N_14166,N_14016);
nand U14295 (N_14295,N_14180,N_14134);
and U14296 (N_14296,N_14048,N_14100);
or U14297 (N_14297,N_14116,N_14114);
or U14298 (N_14298,N_14167,N_14151);
xnor U14299 (N_14299,N_14118,N_14002);
nand U14300 (N_14300,N_14002,N_14159);
and U14301 (N_14301,N_14140,N_14028);
and U14302 (N_14302,N_14008,N_14019);
xor U14303 (N_14303,N_14042,N_14198);
or U14304 (N_14304,N_14153,N_14075);
and U14305 (N_14305,N_14022,N_14190);
xor U14306 (N_14306,N_14157,N_14064);
or U14307 (N_14307,N_14005,N_14057);
xor U14308 (N_14308,N_14095,N_14014);
or U14309 (N_14309,N_14099,N_14085);
or U14310 (N_14310,N_14149,N_14132);
nand U14311 (N_14311,N_14165,N_14098);
and U14312 (N_14312,N_14191,N_14154);
xnor U14313 (N_14313,N_14028,N_14068);
or U14314 (N_14314,N_14100,N_14199);
or U14315 (N_14315,N_14048,N_14181);
xnor U14316 (N_14316,N_14130,N_14065);
nand U14317 (N_14317,N_14194,N_14199);
nor U14318 (N_14318,N_14140,N_14045);
xnor U14319 (N_14319,N_14070,N_14046);
and U14320 (N_14320,N_14160,N_14102);
and U14321 (N_14321,N_14025,N_14008);
nor U14322 (N_14322,N_14044,N_14079);
or U14323 (N_14323,N_14056,N_14127);
xnor U14324 (N_14324,N_14162,N_14197);
nor U14325 (N_14325,N_14057,N_14043);
or U14326 (N_14326,N_14031,N_14181);
xor U14327 (N_14327,N_14001,N_14035);
or U14328 (N_14328,N_14028,N_14135);
xnor U14329 (N_14329,N_14163,N_14192);
and U14330 (N_14330,N_14188,N_14011);
and U14331 (N_14331,N_14076,N_14087);
or U14332 (N_14332,N_14008,N_14029);
nor U14333 (N_14333,N_14091,N_14031);
nor U14334 (N_14334,N_14083,N_14029);
or U14335 (N_14335,N_14113,N_14072);
nor U14336 (N_14336,N_14031,N_14069);
and U14337 (N_14337,N_14007,N_14142);
or U14338 (N_14338,N_14077,N_14190);
nand U14339 (N_14339,N_14034,N_14126);
nand U14340 (N_14340,N_14191,N_14005);
nor U14341 (N_14341,N_14067,N_14173);
and U14342 (N_14342,N_14178,N_14140);
or U14343 (N_14343,N_14107,N_14102);
or U14344 (N_14344,N_14163,N_14121);
nand U14345 (N_14345,N_14142,N_14138);
nand U14346 (N_14346,N_14189,N_14123);
and U14347 (N_14347,N_14010,N_14079);
nor U14348 (N_14348,N_14177,N_14014);
and U14349 (N_14349,N_14114,N_14168);
or U14350 (N_14350,N_14119,N_14191);
or U14351 (N_14351,N_14138,N_14171);
or U14352 (N_14352,N_14112,N_14110);
nor U14353 (N_14353,N_14041,N_14063);
xor U14354 (N_14354,N_14176,N_14187);
or U14355 (N_14355,N_14140,N_14074);
or U14356 (N_14356,N_14169,N_14095);
nand U14357 (N_14357,N_14145,N_14059);
xnor U14358 (N_14358,N_14160,N_14078);
nand U14359 (N_14359,N_14100,N_14000);
or U14360 (N_14360,N_14011,N_14085);
or U14361 (N_14361,N_14059,N_14194);
or U14362 (N_14362,N_14111,N_14007);
xnor U14363 (N_14363,N_14129,N_14150);
nor U14364 (N_14364,N_14139,N_14174);
or U14365 (N_14365,N_14070,N_14001);
and U14366 (N_14366,N_14018,N_14033);
and U14367 (N_14367,N_14011,N_14047);
and U14368 (N_14368,N_14114,N_14130);
nor U14369 (N_14369,N_14174,N_14011);
or U14370 (N_14370,N_14188,N_14006);
or U14371 (N_14371,N_14195,N_14050);
or U14372 (N_14372,N_14183,N_14147);
nand U14373 (N_14373,N_14152,N_14039);
and U14374 (N_14374,N_14074,N_14069);
xor U14375 (N_14375,N_14162,N_14010);
nor U14376 (N_14376,N_14022,N_14117);
or U14377 (N_14377,N_14031,N_14085);
nand U14378 (N_14378,N_14015,N_14166);
nor U14379 (N_14379,N_14142,N_14136);
and U14380 (N_14380,N_14090,N_14062);
and U14381 (N_14381,N_14027,N_14187);
nand U14382 (N_14382,N_14149,N_14126);
or U14383 (N_14383,N_14096,N_14023);
nor U14384 (N_14384,N_14077,N_14188);
nor U14385 (N_14385,N_14041,N_14197);
and U14386 (N_14386,N_14183,N_14102);
nor U14387 (N_14387,N_14067,N_14115);
xor U14388 (N_14388,N_14082,N_14092);
nor U14389 (N_14389,N_14045,N_14195);
xnor U14390 (N_14390,N_14198,N_14091);
nor U14391 (N_14391,N_14195,N_14160);
nor U14392 (N_14392,N_14119,N_14018);
or U14393 (N_14393,N_14094,N_14135);
nand U14394 (N_14394,N_14132,N_14075);
or U14395 (N_14395,N_14086,N_14008);
xor U14396 (N_14396,N_14042,N_14011);
and U14397 (N_14397,N_14014,N_14021);
nor U14398 (N_14398,N_14080,N_14184);
nand U14399 (N_14399,N_14176,N_14131);
or U14400 (N_14400,N_14363,N_14374);
and U14401 (N_14401,N_14218,N_14256);
xnor U14402 (N_14402,N_14319,N_14392);
nand U14403 (N_14403,N_14236,N_14230);
and U14404 (N_14404,N_14239,N_14235);
and U14405 (N_14405,N_14377,N_14204);
and U14406 (N_14406,N_14330,N_14340);
and U14407 (N_14407,N_14353,N_14397);
xnor U14408 (N_14408,N_14238,N_14313);
xor U14409 (N_14409,N_14315,N_14344);
xor U14410 (N_14410,N_14399,N_14263);
xnor U14411 (N_14411,N_14387,N_14247);
and U14412 (N_14412,N_14314,N_14208);
xnor U14413 (N_14413,N_14336,N_14282);
xnor U14414 (N_14414,N_14381,N_14250);
or U14415 (N_14415,N_14356,N_14398);
nand U14416 (N_14416,N_14354,N_14249);
or U14417 (N_14417,N_14335,N_14373);
and U14418 (N_14418,N_14268,N_14292);
and U14419 (N_14419,N_14357,N_14346);
or U14420 (N_14420,N_14287,N_14270);
nor U14421 (N_14421,N_14364,N_14216);
or U14422 (N_14422,N_14224,N_14355);
or U14423 (N_14423,N_14371,N_14306);
or U14424 (N_14424,N_14237,N_14280);
nor U14425 (N_14425,N_14205,N_14207);
and U14426 (N_14426,N_14322,N_14394);
or U14427 (N_14427,N_14307,N_14283);
nand U14428 (N_14428,N_14244,N_14200);
or U14429 (N_14429,N_14290,N_14385);
and U14430 (N_14430,N_14327,N_14217);
xnor U14431 (N_14431,N_14255,N_14240);
nor U14432 (N_14432,N_14302,N_14380);
or U14433 (N_14433,N_14226,N_14360);
xor U14434 (N_14434,N_14286,N_14301);
and U14435 (N_14435,N_14316,N_14219);
nand U14436 (N_14436,N_14288,N_14349);
and U14437 (N_14437,N_14276,N_14289);
and U14438 (N_14438,N_14333,N_14367);
and U14439 (N_14439,N_14227,N_14246);
xnor U14440 (N_14440,N_14245,N_14345);
nand U14441 (N_14441,N_14383,N_14368);
nand U14442 (N_14442,N_14296,N_14273);
and U14443 (N_14443,N_14221,N_14309);
and U14444 (N_14444,N_14391,N_14232);
xnor U14445 (N_14445,N_14274,N_14329);
nor U14446 (N_14446,N_14262,N_14293);
xnor U14447 (N_14447,N_14229,N_14211);
nor U14448 (N_14448,N_14341,N_14261);
nor U14449 (N_14449,N_14212,N_14384);
xor U14450 (N_14450,N_14201,N_14390);
nor U14451 (N_14451,N_14325,N_14334);
xnor U14452 (N_14452,N_14365,N_14254);
nand U14453 (N_14453,N_14303,N_14359);
nor U14454 (N_14454,N_14332,N_14362);
nand U14455 (N_14455,N_14267,N_14304);
xor U14456 (N_14456,N_14366,N_14311);
and U14457 (N_14457,N_14310,N_14395);
xnor U14458 (N_14458,N_14266,N_14358);
nor U14459 (N_14459,N_14203,N_14231);
nor U14460 (N_14460,N_14281,N_14251);
and U14461 (N_14461,N_14347,N_14298);
or U14462 (N_14462,N_14284,N_14258);
xor U14463 (N_14463,N_14378,N_14294);
and U14464 (N_14464,N_14202,N_14372);
xnor U14465 (N_14465,N_14389,N_14342);
nor U14466 (N_14466,N_14337,N_14352);
nor U14467 (N_14467,N_14388,N_14265);
nand U14468 (N_14468,N_14339,N_14343);
nand U14469 (N_14469,N_14318,N_14259);
or U14470 (N_14470,N_14328,N_14321);
and U14471 (N_14471,N_14348,N_14233);
and U14472 (N_14472,N_14376,N_14285);
or U14473 (N_14473,N_14350,N_14210);
and U14474 (N_14474,N_14279,N_14297);
nand U14475 (N_14475,N_14243,N_14248);
nor U14476 (N_14476,N_14338,N_14312);
nor U14477 (N_14477,N_14241,N_14379);
xor U14478 (N_14478,N_14222,N_14257);
nand U14479 (N_14479,N_14295,N_14351);
xor U14480 (N_14480,N_14393,N_14382);
and U14481 (N_14481,N_14275,N_14278);
and U14482 (N_14482,N_14223,N_14213);
nand U14483 (N_14483,N_14323,N_14300);
or U14484 (N_14484,N_14271,N_14228);
nand U14485 (N_14485,N_14206,N_14260);
and U14486 (N_14486,N_14269,N_14326);
nand U14487 (N_14487,N_14291,N_14209);
or U14488 (N_14488,N_14299,N_14277);
and U14489 (N_14489,N_14324,N_14375);
nor U14490 (N_14490,N_14214,N_14215);
xnor U14491 (N_14491,N_14234,N_14369);
and U14492 (N_14492,N_14253,N_14242);
or U14493 (N_14493,N_14272,N_14220);
xor U14494 (N_14494,N_14305,N_14386);
xor U14495 (N_14495,N_14320,N_14370);
and U14496 (N_14496,N_14331,N_14396);
xnor U14497 (N_14497,N_14252,N_14317);
and U14498 (N_14498,N_14361,N_14264);
xor U14499 (N_14499,N_14225,N_14308);
nand U14500 (N_14500,N_14292,N_14326);
or U14501 (N_14501,N_14368,N_14340);
nand U14502 (N_14502,N_14209,N_14395);
xor U14503 (N_14503,N_14393,N_14322);
and U14504 (N_14504,N_14370,N_14246);
nand U14505 (N_14505,N_14370,N_14257);
or U14506 (N_14506,N_14299,N_14252);
and U14507 (N_14507,N_14294,N_14346);
xor U14508 (N_14508,N_14344,N_14223);
nand U14509 (N_14509,N_14263,N_14314);
nor U14510 (N_14510,N_14311,N_14388);
xor U14511 (N_14511,N_14331,N_14259);
nand U14512 (N_14512,N_14352,N_14327);
xnor U14513 (N_14513,N_14262,N_14382);
nor U14514 (N_14514,N_14361,N_14367);
or U14515 (N_14515,N_14202,N_14307);
or U14516 (N_14516,N_14269,N_14241);
nand U14517 (N_14517,N_14240,N_14262);
or U14518 (N_14518,N_14260,N_14328);
or U14519 (N_14519,N_14262,N_14288);
nor U14520 (N_14520,N_14201,N_14356);
xor U14521 (N_14521,N_14322,N_14317);
nand U14522 (N_14522,N_14351,N_14335);
or U14523 (N_14523,N_14332,N_14338);
xnor U14524 (N_14524,N_14261,N_14339);
nand U14525 (N_14525,N_14278,N_14376);
nand U14526 (N_14526,N_14369,N_14275);
nor U14527 (N_14527,N_14204,N_14205);
nand U14528 (N_14528,N_14227,N_14221);
or U14529 (N_14529,N_14347,N_14399);
and U14530 (N_14530,N_14337,N_14305);
nand U14531 (N_14531,N_14323,N_14243);
and U14532 (N_14532,N_14344,N_14300);
nor U14533 (N_14533,N_14343,N_14294);
or U14534 (N_14534,N_14210,N_14235);
xor U14535 (N_14535,N_14314,N_14254);
and U14536 (N_14536,N_14367,N_14302);
xor U14537 (N_14537,N_14342,N_14396);
or U14538 (N_14538,N_14397,N_14278);
and U14539 (N_14539,N_14203,N_14200);
or U14540 (N_14540,N_14301,N_14357);
nor U14541 (N_14541,N_14213,N_14217);
and U14542 (N_14542,N_14397,N_14310);
nand U14543 (N_14543,N_14375,N_14289);
nor U14544 (N_14544,N_14233,N_14291);
nand U14545 (N_14545,N_14250,N_14308);
xor U14546 (N_14546,N_14386,N_14344);
and U14547 (N_14547,N_14262,N_14257);
and U14548 (N_14548,N_14253,N_14310);
and U14549 (N_14549,N_14271,N_14327);
nor U14550 (N_14550,N_14287,N_14258);
xor U14551 (N_14551,N_14375,N_14292);
nand U14552 (N_14552,N_14333,N_14288);
nand U14553 (N_14553,N_14202,N_14366);
or U14554 (N_14554,N_14336,N_14234);
and U14555 (N_14555,N_14240,N_14366);
nand U14556 (N_14556,N_14286,N_14219);
nor U14557 (N_14557,N_14285,N_14234);
nand U14558 (N_14558,N_14277,N_14261);
nand U14559 (N_14559,N_14242,N_14270);
nand U14560 (N_14560,N_14232,N_14241);
or U14561 (N_14561,N_14264,N_14287);
nor U14562 (N_14562,N_14370,N_14262);
or U14563 (N_14563,N_14310,N_14360);
and U14564 (N_14564,N_14368,N_14246);
nand U14565 (N_14565,N_14303,N_14232);
nand U14566 (N_14566,N_14233,N_14260);
or U14567 (N_14567,N_14373,N_14314);
or U14568 (N_14568,N_14374,N_14364);
or U14569 (N_14569,N_14214,N_14372);
xnor U14570 (N_14570,N_14215,N_14357);
nor U14571 (N_14571,N_14286,N_14343);
nor U14572 (N_14572,N_14378,N_14280);
xnor U14573 (N_14573,N_14284,N_14315);
xnor U14574 (N_14574,N_14329,N_14213);
and U14575 (N_14575,N_14288,N_14247);
xnor U14576 (N_14576,N_14238,N_14396);
nand U14577 (N_14577,N_14227,N_14352);
or U14578 (N_14578,N_14356,N_14271);
nand U14579 (N_14579,N_14220,N_14369);
nor U14580 (N_14580,N_14367,N_14282);
nand U14581 (N_14581,N_14302,N_14262);
xor U14582 (N_14582,N_14396,N_14336);
or U14583 (N_14583,N_14371,N_14240);
nor U14584 (N_14584,N_14270,N_14379);
or U14585 (N_14585,N_14230,N_14352);
nand U14586 (N_14586,N_14267,N_14328);
xnor U14587 (N_14587,N_14279,N_14324);
nand U14588 (N_14588,N_14206,N_14227);
nand U14589 (N_14589,N_14210,N_14272);
and U14590 (N_14590,N_14363,N_14253);
or U14591 (N_14591,N_14235,N_14230);
nor U14592 (N_14592,N_14304,N_14294);
nand U14593 (N_14593,N_14240,N_14345);
nor U14594 (N_14594,N_14394,N_14251);
and U14595 (N_14595,N_14312,N_14360);
and U14596 (N_14596,N_14376,N_14293);
nand U14597 (N_14597,N_14207,N_14297);
nand U14598 (N_14598,N_14324,N_14202);
or U14599 (N_14599,N_14335,N_14296);
and U14600 (N_14600,N_14581,N_14449);
nor U14601 (N_14601,N_14415,N_14572);
and U14602 (N_14602,N_14493,N_14448);
nor U14603 (N_14603,N_14435,N_14516);
nor U14604 (N_14604,N_14541,N_14528);
and U14605 (N_14605,N_14504,N_14416);
and U14606 (N_14606,N_14468,N_14540);
nand U14607 (N_14607,N_14485,N_14433);
and U14608 (N_14608,N_14563,N_14530);
and U14609 (N_14609,N_14569,N_14513);
and U14610 (N_14610,N_14555,N_14546);
and U14611 (N_14611,N_14525,N_14437);
or U14612 (N_14612,N_14580,N_14432);
nor U14613 (N_14613,N_14514,N_14599);
nor U14614 (N_14614,N_14512,N_14529);
nand U14615 (N_14615,N_14508,N_14548);
nor U14616 (N_14616,N_14428,N_14550);
and U14617 (N_14617,N_14488,N_14421);
nor U14618 (N_14618,N_14413,N_14480);
or U14619 (N_14619,N_14526,N_14477);
nor U14620 (N_14620,N_14545,N_14559);
nor U14621 (N_14621,N_14596,N_14463);
xnor U14622 (N_14622,N_14562,N_14492);
and U14623 (N_14623,N_14411,N_14589);
nand U14624 (N_14624,N_14462,N_14498);
nor U14625 (N_14625,N_14558,N_14429);
and U14626 (N_14626,N_14439,N_14460);
nand U14627 (N_14627,N_14466,N_14533);
nand U14628 (N_14628,N_14431,N_14497);
nor U14629 (N_14629,N_14487,N_14471);
xnor U14630 (N_14630,N_14509,N_14424);
and U14631 (N_14631,N_14543,N_14406);
xor U14632 (N_14632,N_14592,N_14505);
nand U14633 (N_14633,N_14531,N_14567);
nor U14634 (N_14634,N_14453,N_14475);
or U14635 (N_14635,N_14451,N_14486);
nor U14636 (N_14636,N_14455,N_14409);
nor U14637 (N_14637,N_14425,N_14419);
or U14638 (N_14638,N_14444,N_14427);
nand U14639 (N_14639,N_14483,N_14459);
or U14640 (N_14640,N_14420,N_14539);
xnor U14641 (N_14641,N_14408,N_14423);
and U14642 (N_14642,N_14561,N_14405);
or U14643 (N_14643,N_14454,N_14554);
nor U14644 (N_14644,N_14410,N_14422);
nand U14645 (N_14645,N_14467,N_14591);
or U14646 (N_14646,N_14584,N_14538);
nand U14647 (N_14647,N_14520,N_14574);
or U14648 (N_14648,N_14403,N_14490);
nor U14649 (N_14649,N_14519,N_14418);
and U14650 (N_14650,N_14524,N_14579);
or U14651 (N_14651,N_14565,N_14577);
or U14652 (N_14652,N_14401,N_14452);
nand U14653 (N_14653,N_14560,N_14489);
xor U14654 (N_14654,N_14400,N_14445);
nor U14655 (N_14655,N_14583,N_14501);
xor U14656 (N_14656,N_14442,N_14491);
nand U14657 (N_14657,N_14597,N_14476);
and U14658 (N_14658,N_14570,N_14465);
nor U14659 (N_14659,N_14495,N_14456);
and U14660 (N_14660,N_14590,N_14535);
or U14661 (N_14661,N_14523,N_14564);
xor U14662 (N_14662,N_14515,N_14537);
nor U14663 (N_14663,N_14496,N_14447);
or U14664 (N_14664,N_14521,N_14500);
xor U14665 (N_14665,N_14441,N_14549);
nor U14666 (N_14666,N_14553,N_14474);
or U14667 (N_14667,N_14458,N_14473);
xor U14668 (N_14668,N_14438,N_14430);
and U14669 (N_14669,N_14557,N_14440);
nand U14670 (N_14670,N_14547,N_14478);
nand U14671 (N_14671,N_14407,N_14417);
or U14672 (N_14672,N_14556,N_14494);
and U14673 (N_14673,N_14595,N_14510);
nand U14674 (N_14674,N_14536,N_14522);
and U14675 (N_14675,N_14594,N_14542);
nand U14676 (N_14676,N_14552,N_14436);
nor U14677 (N_14677,N_14585,N_14470);
nor U14678 (N_14678,N_14566,N_14434);
nand U14679 (N_14679,N_14481,N_14527);
nand U14680 (N_14680,N_14587,N_14503);
nand U14681 (N_14681,N_14464,N_14502);
or U14682 (N_14682,N_14532,N_14457);
xnor U14683 (N_14683,N_14404,N_14443);
and U14684 (N_14684,N_14588,N_14582);
nor U14685 (N_14685,N_14472,N_14575);
and U14686 (N_14686,N_14551,N_14412);
nor U14687 (N_14687,N_14414,N_14576);
or U14688 (N_14688,N_14479,N_14598);
xnor U14689 (N_14689,N_14507,N_14426);
xor U14690 (N_14690,N_14518,N_14402);
nand U14691 (N_14691,N_14482,N_14450);
nand U14692 (N_14692,N_14573,N_14593);
and U14693 (N_14693,N_14511,N_14484);
and U14694 (N_14694,N_14571,N_14446);
nand U14695 (N_14695,N_14499,N_14544);
nor U14696 (N_14696,N_14578,N_14534);
or U14697 (N_14697,N_14586,N_14517);
or U14698 (N_14698,N_14461,N_14469);
nand U14699 (N_14699,N_14506,N_14568);
and U14700 (N_14700,N_14441,N_14404);
nand U14701 (N_14701,N_14560,N_14592);
nand U14702 (N_14702,N_14517,N_14541);
xor U14703 (N_14703,N_14401,N_14522);
nor U14704 (N_14704,N_14480,N_14592);
and U14705 (N_14705,N_14461,N_14517);
nand U14706 (N_14706,N_14537,N_14470);
nor U14707 (N_14707,N_14429,N_14516);
or U14708 (N_14708,N_14496,N_14493);
xor U14709 (N_14709,N_14444,N_14454);
and U14710 (N_14710,N_14497,N_14562);
nand U14711 (N_14711,N_14587,N_14572);
xnor U14712 (N_14712,N_14566,N_14432);
xnor U14713 (N_14713,N_14512,N_14410);
nand U14714 (N_14714,N_14427,N_14459);
and U14715 (N_14715,N_14529,N_14412);
nand U14716 (N_14716,N_14590,N_14464);
and U14717 (N_14717,N_14429,N_14441);
or U14718 (N_14718,N_14445,N_14570);
or U14719 (N_14719,N_14503,N_14588);
nand U14720 (N_14720,N_14582,N_14543);
or U14721 (N_14721,N_14532,N_14514);
nand U14722 (N_14722,N_14510,N_14431);
nand U14723 (N_14723,N_14536,N_14417);
and U14724 (N_14724,N_14520,N_14582);
or U14725 (N_14725,N_14422,N_14460);
and U14726 (N_14726,N_14480,N_14445);
or U14727 (N_14727,N_14524,N_14441);
or U14728 (N_14728,N_14484,N_14532);
nand U14729 (N_14729,N_14403,N_14563);
nor U14730 (N_14730,N_14460,N_14538);
nor U14731 (N_14731,N_14450,N_14400);
nor U14732 (N_14732,N_14547,N_14559);
nor U14733 (N_14733,N_14512,N_14587);
nor U14734 (N_14734,N_14532,N_14493);
or U14735 (N_14735,N_14500,N_14407);
or U14736 (N_14736,N_14493,N_14521);
xor U14737 (N_14737,N_14425,N_14402);
nand U14738 (N_14738,N_14536,N_14535);
and U14739 (N_14739,N_14474,N_14455);
xnor U14740 (N_14740,N_14586,N_14467);
xor U14741 (N_14741,N_14569,N_14473);
xor U14742 (N_14742,N_14550,N_14421);
nor U14743 (N_14743,N_14426,N_14562);
and U14744 (N_14744,N_14430,N_14475);
or U14745 (N_14745,N_14521,N_14581);
xor U14746 (N_14746,N_14499,N_14482);
xor U14747 (N_14747,N_14563,N_14542);
xnor U14748 (N_14748,N_14542,N_14592);
nand U14749 (N_14749,N_14545,N_14556);
xnor U14750 (N_14750,N_14409,N_14457);
nor U14751 (N_14751,N_14593,N_14449);
nand U14752 (N_14752,N_14513,N_14505);
nor U14753 (N_14753,N_14565,N_14535);
and U14754 (N_14754,N_14439,N_14518);
xor U14755 (N_14755,N_14521,N_14588);
nand U14756 (N_14756,N_14405,N_14500);
or U14757 (N_14757,N_14517,N_14464);
nand U14758 (N_14758,N_14450,N_14491);
nand U14759 (N_14759,N_14439,N_14446);
nor U14760 (N_14760,N_14516,N_14534);
nor U14761 (N_14761,N_14515,N_14492);
and U14762 (N_14762,N_14482,N_14438);
or U14763 (N_14763,N_14453,N_14581);
and U14764 (N_14764,N_14556,N_14422);
nand U14765 (N_14765,N_14512,N_14455);
nor U14766 (N_14766,N_14582,N_14537);
or U14767 (N_14767,N_14471,N_14543);
or U14768 (N_14768,N_14599,N_14468);
or U14769 (N_14769,N_14550,N_14548);
or U14770 (N_14770,N_14454,N_14502);
nand U14771 (N_14771,N_14428,N_14544);
nand U14772 (N_14772,N_14585,N_14464);
or U14773 (N_14773,N_14517,N_14488);
xor U14774 (N_14774,N_14425,N_14531);
nand U14775 (N_14775,N_14572,N_14523);
or U14776 (N_14776,N_14407,N_14411);
or U14777 (N_14777,N_14430,N_14405);
or U14778 (N_14778,N_14539,N_14402);
and U14779 (N_14779,N_14416,N_14524);
nor U14780 (N_14780,N_14512,N_14428);
xnor U14781 (N_14781,N_14448,N_14545);
xor U14782 (N_14782,N_14501,N_14513);
and U14783 (N_14783,N_14409,N_14410);
or U14784 (N_14784,N_14444,N_14505);
xnor U14785 (N_14785,N_14424,N_14531);
nor U14786 (N_14786,N_14489,N_14583);
and U14787 (N_14787,N_14501,N_14530);
nor U14788 (N_14788,N_14564,N_14555);
nor U14789 (N_14789,N_14589,N_14453);
nand U14790 (N_14790,N_14479,N_14562);
nand U14791 (N_14791,N_14433,N_14462);
and U14792 (N_14792,N_14458,N_14419);
and U14793 (N_14793,N_14402,N_14432);
nor U14794 (N_14794,N_14560,N_14580);
nor U14795 (N_14795,N_14516,N_14577);
and U14796 (N_14796,N_14410,N_14587);
and U14797 (N_14797,N_14460,N_14468);
and U14798 (N_14798,N_14487,N_14534);
nor U14799 (N_14799,N_14431,N_14436);
nand U14800 (N_14800,N_14675,N_14734);
or U14801 (N_14801,N_14720,N_14617);
xnor U14802 (N_14802,N_14666,N_14779);
nor U14803 (N_14803,N_14798,N_14750);
nor U14804 (N_14804,N_14611,N_14748);
nor U14805 (N_14805,N_14607,N_14702);
or U14806 (N_14806,N_14629,N_14655);
xnor U14807 (N_14807,N_14739,N_14648);
or U14808 (N_14808,N_14696,N_14662);
nand U14809 (N_14809,N_14704,N_14766);
nor U14810 (N_14810,N_14612,N_14642);
or U14811 (N_14811,N_14692,N_14621);
nand U14812 (N_14812,N_14600,N_14682);
and U14813 (N_14813,N_14697,N_14773);
nor U14814 (N_14814,N_14610,N_14619);
nor U14815 (N_14815,N_14679,N_14640);
and U14816 (N_14816,N_14756,N_14703);
nor U14817 (N_14817,N_14691,N_14622);
or U14818 (N_14818,N_14695,N_14745);
and U14819 (N_14819,N_14794,N_14693);
and U14820 (N_14820,N_14762,N_14632);
nand U14821 (N_14821,N_14705,N_14661);
and U14822 (N_14822,N_14780,N_14646);
and U14823 (N_14823,N_14764,N_14669);
xor U14824 (N_14824,N_14625,N_14627);
nand U14825 (N_14825,N_14608,N_14711);
and U14826 (N_14826,N_14736,N_14652);
nor U14827 (N_14827,N_14623,N_14647);
nand U14828 (N_14828,N_14659,N_14616);
nor U14829 (N_14829,N_14728,N_14656);
and U14830 (N_14830,N_14641,N_14624);
nand U14831 (N_14831,N_14778,N_14664);
nand U14832 (N_14832,N_14602,N_14751);
or U14833 (N_14833,N_14781,N_14665);
nand U14834 (N_14834,N_14742,N_14615);
xnor U14835 (N_14835,N_14609,N_14788);
nand U14836 (N_14836,N_14799,N_14789);
xor U14837 (N_14837,N_14644,N_14613);
and U14838 (N_14838,N_14713,N_14604);
and U14839 (N_14839,N_14730,N_14735);
and U14840 (N_14840,N_14790,N_14716);
or U14841 (N_14841,N_14688,N_14714);
xor U14842 (N_14842,N_14694,N_14686);
and U14843 (N_14843,N_14606,N_14658);
nor U14844 (N_14844,N_14732,N_14700);
xor U14845 (N_14845,N_14796,N_14729);
or U14846 (N_14846,N_14784,N_14752);
or U14847 (N_14847,N_14620,N_14701);
and U14848 (N_14848,N_14667,N_14718);
or U14849 (N_14849,N_14723,N_14689);
or U14850 (N_14850,N_14654,N_14746);
xnor U14851 (N_14851,N_14630,N_14601);
and U14852 (N_14852,N_14634,N_14676);
nand U14853 (N_14853,N_14782,N_14614);
nor U14854 (N_14854,N_14708,N_14671);
and U14855 (N_14855,N_14638,N_14677);
xor U14856 (N_14856,N_14740,N_14761);
nor U14857 (N_14857,N_14709,N_14681);
nor U14858 (N_14858,N_14722,N_14772);
or U14859 (N_14859,N_14719,N_14637);
nor U14860 (N_14860,N_14793,N_14618);
nor U14861 (N_14861,N_14791,N_14738);
nand U14862 (N_14862,N_14605,N_14721);
nor U14863 (N_14863,N_14660,N_14639);
xor U14864 (N_14864,N_14792,N_14707);
xnor U14865 (N_14865,N_14643,N_14771);
nor U14866 (N_14866,N_14754,N_14651);
xor U14867 (N_14867,N_14770,N_14724);
and U14868 (N_14868,N_14767,N_14777);
nand U14869 (N_14869,N_14657,N_14685);
nand U14870 (N_14870,N_14673,N_14741);
xor U14871 (N_14871,N_14635,N_14795);
xor U14872 (N_14872,N_14710,N_14717);
nand U14873 (N_14873,N_14786,N_14749);
and U14874 (N_14874,N_14757,N_14760);
xor U14875 (N_14875,N_14733,N_14747);
nor U14876 (N_14876,N_14712,N_14765);
or U14877 (N_14877,N_14668,N_14725);
or U14878 (N_14878,N_14768,N_14680);
xor U14879 (N_14879,N_14753,N_14649);
or U14880 (N_14880,N_14672,N_14678);
nor U14881 (N_14881,N_14785,N_14653);
xnor U14882 (N_14882,N_14628,N_14763);
xnor U14883 (N_14883,N_14687,N_14726);
nor U14884 (N_14884,N_14769,N_14699);
or U14885 (N_14885,N_14737,N_14797);
or U14886 (N_14886,N_14758,N_14603);
and U14887 (N_14887,N_14706,N_14633);
or U14888 (N_14888,N_14755,N_14759);
or U14889 (N_14889,N_14775,N_14684);
or U14890 (N_14890,N_14663,N_14727);
nor U14891 (N_14891,N_14744,N_14698);
nor U14892 (N_14892,N_14670,N_14645);
xnor U14893 (N_14893,N_14774,N_14743);
and U14894 (N_14894,N_14650,N_14690);
and U14895 (N_14895,N_14715,N_14787);
and U14896 (N_14896,N_14783,N_14674);
and U14897 (N_14897,N_14626,N_14683);
or U14898 (N_14898,N_14631,N_14636);
and U14899 (N_14899,N_14731,N_14776);
nand U14900 (N_14900,N_14736,N_14681);
and U14901 (N_14901,N_14604,N_14654);
xnor U14902 (N_14902,N_14683,N_14763);
nor U14903 (N_14903,N_14629,N_14700);
nor U14904 (N_14904,N_14754,N_14778);
and U14905 (N_14905,N_14641,N_14726);
xnor U14906 (N_14906,N_14653,N_14678);
or U14907 (N_14907,N_14778,N_14766);
nand U14908 (N_14908,N_14700,N_14677);
and U14909 (N_14909,N_14705,N_14749);
or U14910 (N_14910,N_14729,N_14782);
nand U14911 (N_14911,N_14623,N_14702);
and U14912 (N_14912,N_14735,N_14714);
or U14913 (N_14913,N_14754,N_14660);
xor U14914 (N_14914,N_14631,N_14737);
or U14915 (N_14915,N_14746,N_14607);
and U14916 (N_14916,N_14686,N_14642);
nor U14917 (N_14917,N_14669,N_14711);
xnor U14918 (N_14918,N_14653,N_14731);
xor U14919 (N_14919,N_14652,N_14761);
nand U14920 (N_14920,N_14688,N_14605);
nor U14921 (N_14921,N_14775,N_14771);
nand U14922 (N_14922,N_14730,N_14749);
or U14923 (N_14923,N_14684,N_14725);
xor U14924 (N_14924,N_14763,N_14693);
or U14925 (N_14925,N_14714,N_14680);
nand U14926 (N_14926,N_14790,N_14623);
or U14927 (N_14927,N_14712,N_14714);
or U14928 (N_14928,N_14694,N_14630);
nor U14929 (N_14929,N_14777,N_14606);
and U14930 (N_14930,N_14695,N_14731);
nand U14931 (N_14931,N_14772,N_14625);
xor U14932 (N_14932,N_14752,N_14638);
nor U14933 (N_14933,N_14795,N_14743);
nand U14934 (N_14934,N_14646,N_14698);
xnor U14935 (N_14935,N_14662,N_14789);
or U14936 (N_14936,N_14691,N_14740);
and U14937 (N_14937,N_14792,N_14696);
or U14938 (N_14938,N_14734,N_14682);
and U14939 (N_14939,N_14692,N_14712);
xnor U14940 (N_14940,N_14728,N_14755);
and U14941 (N_14941,N_14604,N_14787);
xor U14942 (N_14942,N_14738,N_14601);
xnor U14943 (N_14943,N_14630,N_14729);
and U14944 (N_14944,N_14769,N_14702);
nand U14945 (N_14945,N_14748,N_14601);
and U14946 (N_14946,N_14720,N_14636);
or U14947 (N_14947,N_14687,N_14716);
xnor U14948 (N_14948,N_14622,N_14652);
nand U14949 (N_14949,N_14704,N_14771);
or U14950 (N_14950,N_14766,N_14659);
nor U14951 (N_14951,N_14736,N_14695);
nor U14952 (N_14952,N_14677,N_14748);
or U14953 (N_14953,N_14652,N_14673);
nand U14954 (N_14954,N_14636,N_14799);
nand U14955 (N_14955,N_14645,N_14736);
or U14956 (N_14956,N_14723,N_14690);
xnor U14957 (N_14957,N_14637,N_14636);
or U14958 (N_14958,N_14792,N_14636);
or U14959 (N_14959,N_14606,N_14650);
nand U14960 (N_14960,N_14668,N_14757);
nor U14961 (N_14961,N_14724,N_14709);
or U14962 (N_14962,N_14795,N_14633);
nor U14963 (N_14963,N_14777,N_14798);
or U14964 (N_14964,N_14670,N_14602);
nor U14965 (N_14965,N_14654,N_14665);
or U14966 (N_14966,N_14657,N_14637);
nor U14967 (N_14967,N_14657,N_14742);
or U14968 (N_14968,N_14775,N_14720);
nand U14969 (N_14969,N_14666,N_14760);
nand U14970 (N_14970,N_14602,N_14690);
nand U14971 (N_14971,N_14775,N_14659);
nor U14972 (N_14972,N_14755,N_14618);
nand U14973 (N_14973,N_14626,N_14731);
xor U14974 (N_14974,N_14791,N_14774);
nand U14975 (N_14975,N_14796,N_14626);
nor U14976 (N_14976,N_14685,N_14677);
nor U14977 (N_14977,N_14783,N_14772);
or U14978 (N_14978,N_14729,N_14775);
and U14979 (N_14979,N_14684,N_14628);
nor U14980 (N_14980,N_14628,N_14710);
nand U14981 (N_14981,N_14614,N_14646);
nor U14982 (N_14982,N_14705,N_14649);
nand U14983 (N_14983,N_14697,N_14661);
nor U14984 (N_14984,N_14662,N_14726);
xor U14985 (N_14985,N_14671,N_14674);
xnor U14986 (N_14986,N_14774,N_14635);
xor U14987 (N_14987,N_14701,N_14708);
nor U14988 (N_14988,N_14770,N_14700);
or U14989 (N_14989,N_14669,N_14729);
nor U14990 (N_14990,N_14783,N_14604);
and U14991 (N_14991,N_14761,N_14690);
xnor U14992 (N_14992,N_14651,N_14793);
or U14993 (N_14993,N_14603,N_14648);
or U14994 (N_14994,N_14723,N_14777);
nor U14995 (N_14995,N_14744,N_14752);
nand U14996 (N_14996,N_14676,N_14798);
nand U14997 (N_14997,N_14708,N_14694);
nand U14998 (N_14998,N_14732,N_14659);
or U14999 (N_14999,N_14704,N_14765);
and U15000 (N_15000,N_14970,N_14875);
or U15001 (N_15001,N_14919,N_14924);
nor U15002 (N_15002,N_14960,N_14990);
and U15003 (N_15003,N_14951,N_14905);
or U15004 (N_15004,N_14849,N_14822);
or U15005 (N_15005,N_14836,N_14915);
or U15006 (N_15006,N_14814,N_14938);
nor U15007 (N_15007,N_14807,N_14856);
nor U15008 (N_15008,N_14884,N_14879);
xnor U15009 (N_15009,N_14817,N_14940);
and U15010 (N_15010,N_14899,N_14941);
and U15011 (N_15011,N_14843,N_14949);
or U15012 (N_15012,N_14844,N_14857);
xnor U15013 (N_15013,N_14885,N_14812);
xnor U15014 (N_15014,N_14911,N_14937);
or U15015 (N_15015,N_14991,N_14962);
and U15016 (N_15016,N_14922,N_14883);
or U15017 (N_15017,N_14867,N_14815);
nor U15018 (N_15018,N_14926,N_14823);
nand U15019 (N_15019,N_14892,N_14876);
nor U15020 (N_15020,N_14918,N_14805);
and U15021 (N_15021,N_14818,N_14808);
or U15022 (N_15022,N_14933,N_14983);
and U15023 (N_15023,N_14816,N_14925);
xnor U15024 (N_15024,N_14907,N_14861);
and U15025 (N_15025,N_14846,N_14819);
nand U15026 (N_15026,N_14985,N_14889);
and U15027 (N_15027,N_14838,N_14860);
and U15028 (N_15028,N_14967,N_14989);
nor U15029 (N_15029,N_14801,N_14864);
nor U15030 (N_15030,N_14984,N_14897);
and U15031 (N_15031,N_14996,N_14971);
xor U15032 (N_15032,N_14909,N_14802);
or U15033 (N_15033,N_14961,N_14908);
xor U15034 (N_15034,N_14906,N_14871);
and U15035 (N_15035,N_14901,N_14946);
and U15036 (N_15036,N_14923,N_14969);
nand U15037 (N_15037,N_14835,N_14800);
and U15038 (N_15038,N_14904,N_14998);
xnor U15039 (N_15039,N_14981,N_14834);
xor U15040 (N_15040,N_14929,N_14854);
and U15041 (N_15041,N_14886,N_14995);
nand U15042 (N_15042,N_14903,N_14881);
nor U15043 (N_15043,N_14913,N_14890);
xnor U15044 (N_15044,N_14898,N_14964);
nor U15045 (N_15045,N_14865,N_14963);
and U15046 (N_15046,N_14955,N_14832);
nand U15047 (N_15047,N_14927,N_14806);
xnor U15048 (N_15048,N_14988,N_14979);
nand U15049 (N_15049,N_14982,N_14966);
nand U15050 (N_15050,N_14975,N_14945);
or U15051 (N_15051,N_14896,N_14976);
or U15052 (N_15052,N_14870,N_14978);
or U15053 (N_15053,N_14921,N_14873);
nor U15054 (N_15054,N_14891,N_14887);
xnor U15055 (N_15055,N_14845,N_14831);
nand U15056 (N_15056,N_14930,N_14895);
xor U15057 (N_15057,N_14934,N_14830);
xnor U15058 (N_15058,N_14841,N_14882);
nand U15059 (N_15059,N_14855,N_14850);
xnor U15060 (N_15060,N_14993,N_14847);
xnor U15061 (N_15061,N_14920,N_14944);
nand U15062 (N_15062,N_14912,N_14974);
xnor U15063 (N_15063,N_14936,N_14900);
nand U15064 (N_15064,N_14986,N_14910);
nand U15065 (N_15065,N_14957,N_14977);
or U15066 (N_15066,N_14863,N_14821);
xnor U15067 (N_15067,N_14953,N_14869);
or U15068 (N_15068,N_14943,N_14948);
xor U15069 (N_15069,N_14853,N_14858);
or U15070 (N_15070,N_14968,N_14932);
nand U15071 (N_15071,N_14917,N_14874);
and U15072 (N_15072,N_14833,N_14868);
and U15073 (N_15073,N_14880,N_14973);
nor U15074 (N_15074,N_14827,N_14987);
nor U15075 (N_15075,N_14828,N_14992);
nand U15076 (N_15076,N_14931,N_14826);
or U15077 (N_15077,N_14840,N_14839);
nand U15078 (N_15078,N_14820,N_14994);
nand U15079 (N_15079,N_14959,N_14939);
or U15080 (N_15080,N_14866,N_14888);
nor U15081 (N_15081,N_14804,N_14972);
nand U15082 (N_15082,N_14999,N_14935);
or U15083 (N_15083,N_14859,N_14997);
and U15084 (N_15084,N_14851,N_14829);
nor U15085 (N_15085,N_14902,N_14810);
nor U15086 (N_15086,N_14947,N_14862);
xnor U15087 (N_15087,N_14980,N_14824);
xor U15088 (N_15088,N_14956,N_14914);
and U15089 (N_15089,N_14848,N_14842);
or U15090 (N_15090,N_14852,N_14965);
or U15091 (N_15091,N_14878,N_14893);
nand U15092 (N_15092,N_14877,N_14952);
or U15093 (N_15093,N_14928,N_14894);
nand U15094 (N_15094,N_14837,N_14958);
xor U15095 (N_15095,N_14825,N_14803);
nor U15096 (N_15096,N_14950,N_14872);
and U15097 (N_15097,N_14954,N_14942);
xor U15098 (N_15098,N_14916,N_14809);
or U15099 (N_15099,N_14811,N_14813);
or U15100 (N_15100,N_14883,N_14808);
or U15101 (N_15101,N_14851,N_14974);
xor U15102 (N_15102,N_14984,N_14945);
or U15103 (N_15103,N_14812,N_14837);
or U15104 (N_15104,N_14862,N_14941);
and U15105 (N_15105,N_14851,N_14883);
or U15106 (N_15106,N_14884,N_14920);
or U15107 (N_15107,N_14807,N_14903);
xnor U15108 (N_15108,N_14953,N_14957);
nor U15109 (N_15109,N_14906,N_14945);
xnor U15110 (N_15110,N_14824,N_14957);
or U15111 (N_15111,N_14964,N_14886);
xnor U15112 (N_15112,N_14914,N_14837);
nor U15113 (N_15113,N_14837,N_14963);
and U15114 (N_15114,N_14958,N_14829);
or U15115 (N_15115,N_14806,N_14856);
xnor U15116 (N_15116,N_14981,N_14836);
nor U15117 (N_15117,N_14923,N_14964);
nor U15118 (N_15118,N_14856,N_14879);
nor U15119 (N_15119,N_14889,N_14982);
nand U15120 (N_15120,N_14968,N_14915);
or U15121 (N_15121,N_14924,N_14884);
and U15122 (N_15122,N_14801,N_14806);
and U15123 (N_15123,N_14857,N_14992);
xnor U15124 (N_15124,N_14837,N_14956);
xnor U15125 (N_15125,N_14822,N_14805);
nor U15126 (N_15126,N_14860,N_14894);
and U15127 (N_15127,N_14832,N_14951);
nor U15128 (N_15128,N_14976,N_14972);
nand U15129 (N_15129,N_14837,N_14885);
and U15130 (N_15130,N_14985,N_14865);
xnor U15131 (N_15131,N_14958,N_14818);
and U15132 (N_15132,N_14972,N_14823);
and U15133 (N_15133,N_14949,N_14811);
and U15134 (N_15134,N_14938,N_14855);
and U15135 (N_15135,N_14952,N_14987);
or U15136 (N_15136,N_14925,N_14959);
and U15137 (N_15137,N_14959,N_14879);
xnor U15138 (N_15138,N_14824,N_14863);
and U15139 (N_15139,N_14895,N_14905);
and U15140 (N_15140,N_14989,N_14902);
and U15141 (N_15141,N_14932,N_14916);
or U15142 (N_15142,N_14852,N_14925);
and U15143 (N_15143,N_14883,N_14809);
nor U15144 (N_15144,N_14889,N_14958);
nand U15145 (N_15145,N_14830,N_14881);
and U15146 (N_15146,N_14876,N_14883);
or U15147 (N_15147,N_14943,N_14854);
xnor U15148 (N_15148,N_14864,N_14932);
nor U15149 (N_15149,N_14928,N_14908);
and U15150 (N_15150,N_14950,N_14832);
nand U15151 (N_15151,N_14902,N_14832);
nand U15152 (N_15152,N_14998,N_14886);
nand U15153 (N_15153,N_14890,N_14927);
nand U15154 (N_15154,N_14913,N_14915);
nand U15155 (N_15155,N_14885,N_14934);
and U15156 (N_15156,N_14922,N_14967);
and U15157 (N_15157,N_14842,N_14901);
nor U15158 (N_15158,N_14802,N_14918);
or U15159 (N_15159,N_14923,N_14845);
and U15160 (N_15160,N_14939,N_14811);
or U15161 (N_15161,N_14992,N_14878);
nand U15162 (N_15162,N_14891,N_14966);
and U15163 (N_15163,N_14993,N_14859);
or U15164 (N_15164,N_14823,N_14800);
or U15165 (N_15165,N_14801,N_14971);
nor U15166 (N_15166,N_14955,N_14880);
or U15167 (N_15167,N_14987,N_14851);
and U15168 (N_15168,N_14833,N_14888);
or U15169 (N_15169,N_14910,N_14808);
nand U15170 (N_15170,N_14893,N_14864);
and U15171 (N_15171,N_14830,N_14993);
or U15172 (N_15172,N_14886,N_14979);
and U15173 (N_15173,N_14954,N_14986);
xnor U15174 (N_15174,N_14898,N_14860);
nor U15175 (N_15175,N_14817,N_14827);
nor U15176 (N_15176,N_14897,N_14989);
or U15177 (N_15177,N_14866,N_14845);
or U15178 (N_15178,N_14883,N_14934);
nand U15179 (N_15179,N_14806,N_14886);
and U15180 (N_15180,N_14984,N_14823);
nor U15181 (N_15181,N_14870,N_14810);
xor U15182 (N_15182,N_14896,N_14986);
nor U15183 (N_15183,N_14910,N_14871);
nand U15184 (N_15184,N_14985,N_14952);
nor U15185 (N_15185,N_14897,N_14831);
and U15186 (N_15186,N_14865,N_14889);
nand U15187 (N_15187,N_14935,N_14998);
or U15188 (N_15188,N_14923,N_14892);
nor U15189 (N_15189,N_14985,N_14937);
and U15190 (N_15190,N_14954,N_14812);
or U15191 (N_15191,N_14909,N_14926);
or U15192 (N_15192,N_14813,N_14901);
or U15193 (N_15193,N_14908,N_14863);
and U15194 (N_15194,N_14834,N_14963);
nor U15195 (N_15195,N_14914,N_14939);
nor U15196 (N_15196,N_14927,N_14947);
and U15197 (N_15197,N_14824,N_14943);
and U15198 (N_15198,N_14846,N_14965);
xnor U15199 (N_15199,N_14840,N_14826);
or U15200 (N_15200,N_15008,N_15111);
nand U15201 (N_15201,N_15045,N_15186);
nand U15202 (N_15202,N_15050,N_15141);
nand U15203 (N_15203,N_15166,N_15167);
nor U15204 (N_15204,N_15177,N_15022);
and U15205 (N_15205,N_15089,N_15007);
nand U15206 (N_15206,N_15105,N_15189);
and U15207 (N_15207,N_15194,N_15010);
nand U15208 (N_15208,N_15055,N_15054);
nand U15209 (N_15209,N_15187,N_15199);
or U15210 (N_15210,N_15058,N_15128);
or U15211 (N_15211,N_15002,N_15121);
and U15212 (N_15212,N_15075,N_15068);
xor U15213 (N_15213,N_15140,N_15033);
xnor U15214 (N_15214,N_15072,N_15184);
nand U15215 (N_15215,N_15195,N_15154);
or U15216 (N_15216,N_15173,N_15013);
nand U15217 (N_15217,N_15197,N_15172);
xor U15218 (N_15218,N_15133,N_15135);
and U15219 (N_15219,N_15061,N_15087);
nor U15220 (N_15220,N_15136,N_15034);
or U15221 (N_15221,N_15159,N_15000);
and U15222 (N_15222,N_15139,N_15145);
xor U15223 (N_15223,N_15042,N_15095);
or U15224 (N_15224,N_15081,N_15106);
nand U15225 (N_15225,N_15104,N_15052);
nand U15226 (N_15226,N_15162,N_15014);
nor U15227 (N_15227,N_15191,N_15150);
and U15228 (N_15228,N_15188,N_15181);
or U15229 (N_15229,N_15192,N_15078);
or U15230 (N_15230,N_15093,N_15005);
xnor U15231 (N_15231,N_15153,N_15158);
nor U15232 (N_15232,N_15018,N_15049);
or U15233 (N_15233,N_15028,N_15067);
and U15234 (N_15234,N_15100,N_15143);
xor U15235 (N_15235,N_15174,N_15063);
nor U15236 (N_15236,N_15099,N_15023);
xnor U15237 (N_15237,N_15124,N_15085);
nor U15238 (N_15238,N_15009,N_15073);
xor U15239 (N_15239,N_15171,N_15156);
nand U15240 (N_15240,N_15151,N_15129);
nand U15241 (N_15241,N_15064,N_15101);
and U15242 (N_15242,N_15137,N_15126);
nor U15243 (N_15243,N_15122,N_15047);
and U15244 (N_15244,N_15032,N_15107);
or U15245 (N_15245,N_15098,N_15112);
xor U15246 (N_15246,N_15190,N_15036);
and U15247 (N_15247,N_15040,N_15020);
or U15248 (N_15248,N_15138,N_15025);
nor U15249 (N_15249,N_15026,N_15070);
nand U15250 (N_15250,N_15071,N_15037);
nand U15251 (N_15251,N_15127,N_15060);
or U15252 (N_15252,N_15169,N_15092);
xor U15253 (N_15253,N_15051,N_15001);
or U15254 (N_15254,N_15146,N_15094);
and U15255 (N_15255,N_15003,N_15134);
and U15256 (N_15256,N_15065,N_15086);
or U15257 (N_15257,N_15066,N_15027);
nand U15258 (N_15258,N_15059,N_15091);
nor U15259 (N_15259,N_15115,N_15168);
or U15260 (N_15260,N_15142,N_15165);
xor U15261 (N_15261,N_15083,N_15119);
or U15262 (N_15262,N_15043,N_15102);
nor U15263 (N_15263,N_15179,N_15148);
nor U15264 (N_15264,N_15015,N_15017);
or U15265 (N_15265,N_15113,N_15196);
xnor U15266 (N_15266,N_15021,N_15031);
nand U15267 (N_15267,N_15012,N_15030);
and U15268 (N_15268,N_15057,N_15110);
nor U15269 (N_15269,N_15097,N_15046);
xnor U15270 (N_15270,N_15116,N_15123);
xnor U15271 (N_15271,N_15118,N_15004);
nor U15272 (N_15272,N_15198,N_15080);
nor U15273 (N_15273,N_15062,N_15011);
xor U15274 (N_15274,N_15164,N_15006);
nand U15275 (N_15275,N_15048,N_15125);
or U15276 (N_15276,N_15175,N_15163);
nor U15277 (N_15277,N_15024,N_15131);
or U15278 (N_15278,N_15157,N_15117);
xnor U15279 (N_15279,N_15155,N_15096);
nand U15280 (N_15280,N_15180,N_15182);
nor U15281 (N_15281,N_15039,N_15147);
xor U15282 (N_15282,N_15074,N_15035);
xnor U15283 (N_15283,N_15056,N_15016);
and U15284 (N_15284,N_15041,N_15090);
or U15285 (N_15285,N_15193,N_15103);
nor U15286 (N_15286,N_15019,N_15170);
nand U15287 (N_15287,N_15120,N_15082);
and U15288 (N_15288,N_15029,N_15160);
nor U15289 (N_15289,N_15044,N_15077);
nand U15290 (N_15290,N_15144,N_15076);
nor U15291 (N_15291,N_15149,N_15114);
xnor U15292 (N_15292,N_15038,N_15178);
or U15293 (N_15293,N_15084,N_15069);
and U15294 (N_15294,N_15161,N_15053);
nand U15295 (N_15295,N_15109,N_15130);
xor U15296 (N_15296,N_15079,N_15183);
xnor U15297 (N_15297,N_15176,N_15185);
nor U15298 (N_15298,N_15088,N_15108);
xor U15299 (N_15299,N_15132,N_15152);
or U15300 (N_15300,N_15039,N_15096);
or U15301 (N_15301,N_15005,N_15022);
or U15302 (N_15302,N_15017,N_15115);
xor U15303 (N_15303,N_15106,N_15118);
nand U15304 (N_15304,N_15187,N_15044);
and U15305 (N_15305,N_15166,N_15159);
nor U15306 (N_15306,N_15152,N_15079);
nand U15307 (N_15307,N_15104,N_15004);
nand U15308 (N_15308,N_15102,N_15080);
and U15309 (N_15309,N_15013,N_15006);
or U15310 (N_15310,N_15119,N_15012);
and U15311 (N_15311,N_15131,N_15102);
xnor U15312 (N_15312,N_15102,N_15181);
xnor U15313 (N_15313,N_15096,N_15067);
xnor U15314 (N_15314,N_15025,N_15060);
xor U15315 (N_15315,N_15188,N_15159);
nand U15316 (N_15316,N_15166,N_15076);
xnor U15317 (N_15317,N_15092,N_15166);
nand U15318 (N_15318,N_15049,N_15167);
nor U15319 (N_15319,N_15063,N_15026);
nand U15320 (N_15320,N_15063,N_15173);
and U15321 (N_15321,N_15016,N_15001);
nor U15322 (N_15322,N_15058,N_15071);
and U15323 (N_15323,N_15175,N_15135);
nand U15324 (N_15324,N_15006,N_15128);
or U15325 (N_15325,N_15103,N_15009);
xnor U15326 (N_15326,N_15037,N_15166);
and U15327 (N_15327,N_15066,N_15187);
and U15328 (N_15328,N_15096,N_15083);
nor U15329 (N_15329,N_15183,N_15056);
or U15330 (N_15330,N_15138,N_15060);
and U15331 (N_15331,N_15029,N_15163);
or U15332 (N_15332,N_15047,N_15077);
nor U15333 (N_15333,N_15030,N_15081);
xor U15334 (N_15334,N_15084,N_15081);
nand U15335 (N_15335,N_15142,N_15110);
nor U15336 (N_15336,N_15009,N_15195);
and U15337 (N_15337,N_15183,N_15099);
or U15338 (N_15338,N_15107,N_15112);
or U15339 (N_15339,N_15002,N_15077);
or U15340 (N_15340,N_15146,N_15111);
nor U15341 (N_15341,N_15133,N_15128);
nor U15342 (N_15342,N_15126,N_15185);
and U15343 (N_15343,N_15066,N_15164);
nor U15344 (N_15344,N_15086,N_15150);
nand U15345 (N_15345,N_15053,N_15122);
and U15346 (N_15346,N_15188,N_15176);
and U15347 (N_15347,N_15000,N_15083);
xnor U15348 (N_15348,N_15073,N_15012);
xor U15349 (N_15349,N_15079,N_15010);
nand U15350 (N_15350,N_15073,N_15109);
and U15351 (N_15351,N_15029,N_15106);
xor U15352 (N_15352,N_15029,N_15140);
or U15353 (N_15353,N_15058,N_15156);
xor U15354 (N_15354,N_15149,N_15052);
xnor U15355 (N_15355,N_15042,N_15152);
or U15356 (N_15356,N_15119,N_15187);
or U15357 (N_15357,N_15150,N_15053);
nor U15358 (N_15358,N_15079,N_15080);
and U15359 (N_15359,N_15110,N_15190);
and U15360 (N_15360,N_15147,N_15139);
or U15361 (N_15361,N_15193,N_15111);
xnor U15362 (N_15362,N_15149,N_15048);
nand U15363 (N_15363,N_15045,N_15104);
nand U15364 (N_15364,N_15152,N_15178);
xor U15365 (N_15365,N_15143,N_15049);
nor U15366 (N_15366,N_15158,N_15009);
xor U15367 (N_15367,N_15198,N_15066);
and U15368 (N_15368,N_15181,N_15088);
or U15369 (N_15369,N_15016,N_15049);
and U15370 (N_15370,N_15027,N_15178);
nor U15371 (N_15371,N_15060,N_15003);
and U15372 (N_15372,N_15116,N_15002);
or U15373 (N_15373,N_15002,N_15041);
xnor U15374 (N_15374,N_15154,N_15188);
nand U15375 (N_15375,N_15197,N_15149);
xor U15376 (N_15376,N_15136,N_15078);
xor U15377 (N_15377,N_15130,N_15156);
nor U15378 (N_15378,N_15140,N_15154);
nor U15379 (N_15379,N_15004,N_15187);
and U15380 (N_15380,N_15056,N_15165);
nor U15381 (N_15381,N_15040,N_15027);
nand U15382 (N_15382,N_15051,N_15159);
nand U15383 (N_15383,N_15090,N_15028);
xnor U15384 (N_15384,N_15015,N_15122);
nand U15385 (N_15385,N_15082,N_15150);
nand U15386 (N_15386,N_15099,N_15097);
nand U15387 (N_15387,N_15106,N_15057);
nand U15388 (N_15388,N_15172,N_15120);
xor U15389 (N_15389,N_15097,N_15022);
nor U15390 (N_15390,N_15080,N_15094);
xor U15391 (N_15391,N_15146,N_15060);
xor U15392 (N_15392,N_15086,N_15075);
nand U15393 (N_15393,N_15088,N_15028);
xnor U15394 (N_15394,N_15005,N_15179);
nor U15395 (N_15395,N_15140,N_15191);
and U15396 (N_15396,N_15121,N_15195);
nand U15397 (N_15397,N_15156,N_15048);
and U15398 (N_15398,N_15026,N_15082);
xor U15399 (N_15399,N_15055,N_15114);
and U15400 (N_15400,N_15237,N_15298);
nor U15401 (N_15401,N_15349,N_15356);
or U15402 (N_15402,N_15364,N_15346);
xnor U15403 (N_15403,N_15214,N_15244);
or U15404 (N_15404,N_15278,N_15391);
nand U15405 (N_15405,N_15236,N_15361);
xor U15406 (N_15406,N_15305,N_15309);
nand U15407 (N_15407,N_15263,N_15265);
nor U15408 (N_15408,N_15261,N_15310);
xnor U15409 (N_15409,N_15238,N_15251);
and U15410 (N_15410,N_15240,N_15201);
or U15411 (N_15411,N_15387,N_15259);
nor U15412 (N_15412,N_15367,N_15372);
or U15413 (N_15413,N_15258,N_15282);
nand U15414 (N_15414,N_15248,N_15216);
nand U15415 (N_15415,N_15389,N_15245);
nor U15416 (N_15416,N_15229,N_15264);
and U15417 (N_15417,N_15221,N_15250);
nor U15418 (N_15418,N_15392,N_15332);
nor U15419 (N_15419,N_15232,N_15373);
xor U15420 (N_15420,N_15325,N_15218);
nand U15421 (N_15421,N_15351,N_15395);
or U15422 (N_15422,N_15374,N_15225);
or U15423 (N_15423,N_15324,N_15217);
xor U15424 (N_15424,N_15388,N_15357);
or U15425 (N_15425,N_15299,N_15286);
and U15426 (N_15426,N_15350,N_15287);
or U15427 (N_15427,N_15352,N_15386);
nand U15428 (N_15428,N_15215,N_15358);
or U15429 (N_15429,N_15283,N_15380);
or U15430 (N_15430,N_15302,N_15308);
or U15431 (N_15431,N_15219,N_15368);
nor U15432 (N_15432,N_15390,N_15280);
and U15433 (N_15433,N_15329,N_15385);
nand U15434 (N_15434,N_15205,N_15369);
and U15435 (N_15435,N_15353,N_15326);
nand U15436 (N_15436,N_15363,N_15204);
and U15437 (N_15437,N_15262,N_15375);
nor U15438 (N_15438,N_15200,N_15311);
or U15439 (N_15439,N_15397,N_15271);
and U15440 (N_15440,N_15239,N_15365);
and U15441 (N_15441,N_15379,N_15211);
xnor U15442 (N_15442,N_15230,N_15249);
nand U15443 (N_15443,N_15256,N_15378);
nor U15444 (N_15444,N_15371,N_15341);
nor U15445 (N_15445,N_15285,N_15359);
xor U15446 (N_15446,N_15253,N_15235);
and U15447 (N_15447,N_15255,N_15345);
nand U15448 (N_15448,N_15227,N_15366);
nand U15449 (N_15449,N_15399,N_15339);
xnor U15450 (N_15450,N_15394,N_15279);
nor U15451 (N_15451,N_15376,N_15220);
xor U15452 (N_15452,N_15295,N_15344);
and U15453 (N_15453,N_15304,N_15213);
or U15454 (N_15454,N_15223,N_15273);
nor U15455 (N_15455,N_15328,N_15370);
or U15456 (N_15456,N_15336,N_15254);
nand U15457 (N_15457,N_15354,N_15306);
or U15458 (N_15458,N_15355,N_15257);
nand U15459 (N_15459,N_15289,N_15281);
nor U15460 (N_15460,N_15203,N_15334);
and U15461 (N_15461,N_15383,N_15226);
and U15462 (N_15462,N_15342,N_15393);
nor U15463 (N_15463,N_15267,N_15252);
or U15464 (N_15464,N_15323,N_15292);
nand U15465 (N_15465,N_15288,N_15207);
or U15466 (N_15466,N_15347,N_15247);
nor U15467 (N_15467,N_15319,N_15224);
xor U15468 (N_15468,N_15314,N_15290);
and U15469 (N_15469,N_15322,N_15327);
xnor U15470 (N_15470,N_15343,N_15300);
nor U15471 (N_15471,N_15246,N_15315);
xnor U15472 (N_15472,N_15318,N_15231);
or U15473 (N_15473,N_15335,N_15270);
xnor U15474 (N_15474,N_15381,N_15208);
and U15475 (N_15475,N_15277,N_15241);
and U15476 (N_15476,N_15348,N_15398);
xnor U15477 (N_15477,N_15377,N_15321);
or U15478 (N_15478,N_15269,N_15274);
nand U15479 (N_15479,N_15293,N_15338);
nand U15480 (N_15480,N_15396,N_15316);
nor U15481 (N_15481,N_15331,N_15266);
or U15482 (N_15482,N_15210,N_15333);
xor U15483 (N_15483,N_15384,N_15303);
or U15484 (N_15484,N_15212,N_15228);
xor U15485 (N_15485,N_15209,N_15272);
and U15486 (N_15486,N_15260,N_15243);
nand U15487 (N_15487,N_15296,N_15312);
or U15488 (N_15488,N_15330,N_15294);
or U15489 (N_15489,N_15307,N_15242);
nand U15490 (N_15490,N_15340,N_15317);
xnor U15491 (N_15491,N_15233,N_15275);
and U15492 (N_15492,N_15276,N_15222);
nor U15493 (N_15493,N_15268,N_15337);
and U15494 (N_15494,N_15320,N_15202);
nor U15495 (N_15495,N_15234,N_15206);
and U15496 (N_15496,N_15301,N_15382);
nand U15497 (N_15497,N_15284,N_15313);
nand U15498 (N_15498,N_15360,N_15297);
or U15499 (N_15499,N_15291,N_15362);
xor U15500 (N_15500,N_15332,N_15304);
or U15501 (N_15501,N_15365,N_15356);
and U15502 (N_15502,N_15399,N_15353);
xnor U15503 (N_15503,N_15299,N_15354);
nor U15504 (N_15504,N_15391,N_15382);
xor U15505 (N_15505,N_15354,N_15356);
xnor U15506 (N_15506,N_15302,N_15241);
nor U15507 (N_15507,N_15208,N_15363);
xnor U15508 (N_15508,N_15278,N_15223);
or U15509 (N_15509,N_15363,N_15239);
nand U15510 (N_15510,N_15215,N_15338);
xnor U15511 (N_15511,N_15336,N_15313);
xnor U15512 (N_15512,N_15262,N_15216);
or U15513 (N_15513,N_15338,N_15302);
xnor U15514 (N_15514,N_15301,N_15208);
xor U15515 (N_15515,N_15374,N_15213);
or U15516 (N_15516,N_15282,N_15241);
nor U15517 (N_15517,N_15259,N_15378);
nor U15518 (N_15518,N_15239,N_15254);
xor U15519 (N_15519,N_15216,N_15304);
xnor U15520 (N_15520,N_15258,N_15395);
xor U15521 (N_15521,N_15362,N_15220);
nor U15522 (N_15522,N_15230,N_15209);
and U15523 (N_15523,N_15320,N_15358);
nand U15524 (N_15524,N_15370,N_15283);
xor U15525 (N_15525,N_15367,N_15387);
nor U15526 (N_15526,N_15372,N_15296);
nor U15527 (N_15527,N_15369,N_15372);
and U15528 (N_15528,N_15348,N_15288);
xnor U15529 (N_15529,N_15324,N_15360);
nor U15530 (N_15530,N_15263,N_15326);
xor U15531 (N_15531,N_15227,N_15219);
or U15532 (N_15532,N_15375,N_15348);
nand U15533 (N_15533,N_15290,N_15269);
and U15534 (N_15534,N_15362,N_15230);
nor U15535 (N_15535,N_15289,N_15375);
xor U15536 (N_15536,N_15248,N_15319);
nor U15537 (N_15537,N_15298,N_15240);
nand U15538 (N_15538,N_15263,N_15361);
and U15539 (N_15539,N_15303,N_15240);
or U15540 (N_15540,N_15390,N_15356);
xor U15541 (N_15541,N_15330,N_15341);
nand U15542 (N_15542,N_15208,N_15382);
nor U15543 (N_15543,N_15318,N_15223);
nor U15544 (N_15544,N_15359,N_15268);
and U15545 (N_15545,N_15336,N_15368);
nand U15546 (N_15546,N_15307,N_15316);
nor U15547 (N_15547,N_15356,N_15351);
and U15548 (N_15548,N_15344,N_15331);
xor U15549 (N_15549,N_15261,N_15308);
and U15550 (N_15550,N_15223,N_15320);
and U15551 (N_15551,N_15303,N_15243);
xor U15552 (N_15552,N_15330,N_15321);
xnor U15553 (N_15553,N_15273,N_15215);
and U15554 (N_15554,N_15326,N_15378);
xnor U15555 (N_15555,N_15382,N_15342);
xnor U15556 (N_15556,N_15259,N_15398);
xor U15557 (N_15557,N_15391,N_15342);
nand U15558 (N_15558,N_15277,N_15216);
xnor U15559 (N_15559,N_15290,N_15289);
or U15560 (N_15560,N_15335,N_15317);
xnor U15561 (N_15561,N_15329,N_15340);
and U15562 (N_15562,N_15206,N_15348);
nor U15563 (N_15563,N_15237,N_15331);
and U15564 (N_15564,N_15338,N_15311);
xor U15565 (N_15565,N_15341,N_15214);
nor U15566 (N_15566,N_15382,N_15307);
nor U15567 (N_15567,N_15286,N_15261);
and U15568 (N_15568,N_15314,N_15247);
or U15569 (N_15569,N_15348,N_15239);
or U15570 (N_15570,N_15362,N_15387);
and U15571 (N_15571,N_15233,N_15372);
or U15572 (N_15572,N_15399,N_15329);
and U15573 (N_15573,N_15239,N_15385);
nand U15574 (N_15574,N_15345,N_15259);
nor U15575 (N_15575,N_15297,N_15353);
and U15576 (N_15576,N_15205,N_15267);
and U15577 (N_15577,N_15303,N_15312);
and U15578 (N_15578,N_15376,N_15352);
and U15579 (N_15579,N_15383,N_15284);
nor U15580 (N_15580,N_15316,N_15241);
xor U15581 (N_15581,N_15306,N_15237);
xnor U15582 (N_15582,N_15339,N_15233);
and U15583 (N_15583,N_15277,N_15239);
nand U15584 (N_15584,N_15376,N_15388);
or U15585 (N_15585,N_15248,N_15306);
nor U15586 (N_15586,N_15278,N_15212);
and U15587 (N_15587,N_15229,N_15200);
nor U15588 (N_15588,N_15360,N_15372);
and U15589 (N_15589,N_15347,N_15362);
or U15590 (N_15590,N_15286,N_15212);
nor U15591 (N_15591,N_15281,N_15330);
nor U15592 (N_15592,N_15213,N_15292);
nor U15593 (N_15593,N_15322,N_15281);
and U15594 (N_15594,N_15273,N_15237);
or U15595 (N_15595,N_15385,N_15364);
nand U15596 (N_15596,N_15241,N_15219);
or U15597 (N_15597,N_15229,N_15329);
xnor U15598 (N_15598,N_15296,N_15395);
xor U15599 (N_15599,N_15249,N_15200);
nor U15600 (N_15600,N_15544,N_15402);
xor U15601 (N_15601,N_15437,N_15546);
and U15602 (N_15602,N_15579,N_15472);
nor U15603 (N_15603,N_15436,N_15444);
and U15604 (N_15604,N_15547,N_15452);
xor U15605 (N_15605,N_15515,N_15541);
nand U15606 (N_15606,N_15487,N_15599);
or U15607 (N_15607,N_15491,N_15582);
nand U15608 (N_15608,N_15420,N_15403);
xnor U15609 (N_15609,N_15542,N_15584);
nor U15610 (N_15610,N_15555,N_15514);
nand U15611 (N_15611,N_15475,N_15524);
and U15612 (N_15612,N_15496,N_15412);
xnor U15613 (N_15613,N_15500,N_15511);
nand U15614 (N_15614,N_15489,N_15483);
xor U15615 (N_15615,N_15561,N_15520);
xor U15616 (N_15616,N_15509,N_15456);
or U15617 (N_15617,N_15553,N_15481);
xnor U15618 (N_15618,N_15484,N_15554);
nand U15619 (N_15619,N_15537,N_15533);
and U15620 (N_15620,N_15407,N_15536);
nand U15621 (N_15621,N_15516,N_15538);
or U15622 (N_15622,N_15578,N_15519);
and U15623 (N_15623,N_15473,N_15583);
xor U15624 (N_15624,N_15517,N_15461);
nand U15625 (N_15625,N_15462,N_15446);
nor U15626 (N_15626,N_15580,N_15467);
and U15627 (N_15627,N_15508,N_15485);
xor U15628 (N_15628,N_15430,N_15526);
nor U15629 (N_15629,N_15423,N_15528);
or U15630 (N_15630,N_15577,N_15466);
nor U15631 (N_15631,N_15597,N_15505);
nand U15632 (N_15632,N_15545,N_15556);
nand U15633 (N_15633,N_15565,N_15525);
nor U15634 (N_15634,N_15534,N_15426);
nand U15635 (N_15635,N_15558,N_15595);
xnor U15636 (N_15636,N_15571,N_15523);
or U15637 (N_15637,N_15532,N_15576);
nor U15638 (N_15638,N_15465,N_15486);
xnor U15639 (N_15639,N_15596,N_15531);
xnor U15640 (N_15640,N_15506,N_15552);
or U15641 (N_15641,N_15594,N_15476);
nand U15642 (N_15642,N_15419,N_15581);
nand U15643 (N_15643,N_15570,N_15454);
and U15644 (N_15644,N_15405,N_15474);
or U15645 (N_15645,N_15432,N_15557);
nor U15646 (N_15646,N_15439,N_15458);
and U15647 (N_15647,N_15513,N_15471);
or U15648 (N_15648,N_15424,N_15414);
nor U15649 (N_15649,N_15498,N_15453);
or U15650 (N_15650,N_15499,N_15512);
and U15651 (N_15651,N_15566,N_15548);
xnor U15652 (N_15652,N_15497,N_15549);
xor U15653 (N_15653,N_15575,N_15421);
and U15654 (N_15654,N_15477,N_15522);
nand U15655 (N_15655,N_15428,N_15543);
xor U15656 (N_15656,N_15411,N_15404);
nand U15657 (N_15657,N_15455,N_15463);
nand U15658 (N_15658,N_15460,N_15587);
and U15659 (N_15659,N_15588,N_15480);
and U15660 (N_15660,N_15502,N_15589);
nor U15661 (N_15661,N_15429,N_15593);
and U15662 (N_15662,N_15468,N_15442);
or U15663 (N_15663,N_15422,N_15586);
or U15664 (N_15664,N_15493,N_15431);
and U15665 (N_15665,N_15598,N_15401);
nor U15666 (N_15666,N_15521,N_15567);
and U15667 (N_15667,N_15469,N_15441);
nand U15668 (N_15668,N_15518,N_15409);
xnor U15669 (N_15669,N_15572,N_15559);
xor U15670 (N_15670,N_15573,N_15591);
or U15671 (N_15671,N_15427,N_15490);
or U15672 (N_15672,N_15408,N_15551);
nor U15673 (N_15673,N_15563,N_15447);
nand U15674 (N_15674,N_15417,N_15457);
xnor U15675 (N_15675,N_15451,N_15435);
nor U15676 (N_15676,N_15574,N_15479);
or U15677 (N_15677,N_15406,N_15448);
and U15678 (N_15678,N_15585,N_15440);
xor U15679 (N_15679,N_15564,N_15501);
xor U15680 (N_15680,N_15535,N_15507);
or U15681 (N_15681,N_15449,N_15400);
xor U15682 (N_15682,N_15540,N_15562);
and U15683 (N_15683,N_15443,N_15495);
and U15684 (N_15684,N_15529,N_15445);
xor U15685 (N_15685,N_15492,N_15438);
xnor U15686 (N_15686,N_15425,N_15504);
xor U15687 (N_15687,N_15478,N_15592);
or U15688 (N_15688,N_15415,N_15434);
nand U15689 (N_15689,N_15539,N_15470);
or U15690 (N_15690,N_15416,N_15568);
and U15691 (N_15691,N_15527,N_15413);
nand U15692 (N_15692,N_15503,N_15494);
nor U15693 (N_15693,N_15569,N_15459);
and U15694 (N_15694,N_15418,N_15433);
xor U15695 (N_15695,N_15464,N_15550);
xor U15696 (N_15696,N_15482,N_15590);
xnor U15697 (N_15697,N_15488,N_15530);
and U15698 (N_15698,N_15560,N_15450);
or U15699 (N_15699,N_15410,N_15510);
or U15700 (N_15700,N_15476,N_15467);
or U15701 (N_15701,N_15460,N_15444);
or U15702 (N_15702,N_15468,N_15591);
xor U15703 (N_15703,N_15449,N_15508);
or U15704 (N_15704,N_15446,N_15528);
nand U15705 (N_15705,N_15413,N_15528);
xnor U15706 (N_15706,N_15585,N_15400);
nor U15707 (N_15707,N_15428,N_15461);
xnor U15708 (N_15708,N_15524,N_15472);
nor U15709 (N_15709,N_15596,N_15425);
and U15710 (N_15710,N_15503,N_15569);
nor U15711 (N_15711,N_15569,N_15556);
nand U15712 (N_15712,N_15473,N_15421);
nand U15713 (N_15713,N_15521,N_15409);
xnor U15714 (N_15714,N_15496,N_15515);
or U15715 (N_15715,N_15451,N_15439);
nand U15716 (N_15716,N_15542,N_15458);
and U15717 (N_15717,N_15519,N_15411);
xnor U15718 (N_15718,N_15526,N_15598);
or U15719 (N_15719,N_15449,N_15574);
nor U15720 (N_15720,N_15508,N_15597);
and U15721 (N_15721,N_15422,N_15562);
xor U15722 (N_15722,N_15544,N_15424);
nand U15723 (N_15723,N_15489,N_15420);
and U15724 (N_15724,N_15548,N_15520);
and U15725 (N_15725,N_15433,N_15527);
nand U15726 (N_15726,N_15441,N_15553);
nor U15727 (N_15727,N_15556,N_15593);
nor U15728 (N_15728,N_15401,N_15542);
nor U15729 (N_15729,N_15556,N_15495);
nand U15730 (N_15730,N_15439,N_15588);
xnor U15731 (N_15731,N_15482,N_15436);
xnor U15732 (N_15732,N_15455,N_15534);
xnor U15733 (N_15733,N_15549,N_15424);
and U15734 (N_15734,N_15544,N_15514);
nand U15735 (N_15735,N_15548,N_15561);
or U15736 (N_15736,N_15418,N_15531);
xnor U15737 (N_15737,N_15481,N_15449);
or U15738 (N_15738,N_15469,N_15405);
or U15739 (N_15739,N_15551,N_15462);
or U15740 (N_15740,N_15472,N_15453);
nand U15741 (N_15741,N_15435,N_15489);
xnor U15742 (N_15742,N_15515,N_15557);
xor U15743 (N_15743,N_15590,N_15440);
and U15744 (N_15744,N_15466,N_15453);
and U15745 (N_15745,N_15460,N_15451);
nand U15746 (N_15746,N_15406,N_15510);
nand U15747 (N_15747,N_15500,N_15460);
nand U15748 (N_15748,N_15471,N_15579);
or U15749 (N_15749,N_15580,N_15529);
or U15750 (N_15750,N_15406,N_15435);
or U15751 (N_15751,N_15434,N_15457);
nand U15752 (N_15752,N_15483,N_15401);
nand U15753 (N_15753,N_15421,N_15401);
xor U15754 (N_15754,N_15495,N_15510);
nand U15755 (N_15755,N_15537,N_15414);
or U15756 (N_15756,N_15454,N_15484);
and U15757 (N_15757,N_15544,N_15435);
nor U15758 (N_15758,N_15431,N_15426);
nor U15759 (N_15759,N_15451,N_15419);
nand U15760 (N_15760,N_15545,N_15561);
or U15761 (N_15761,N_15538,N_15459);
nand U15762 (N_15762,N_15505,N_15439);
xor U15763 (N_15763,N_15534,N_15429);
and U15764 (N_15764,N_15562,N_15414);
xnor U15765 (N_15765,N_15522,N_15463);
nor U15766 (N_15766,N_15430,N_15500);
nor U15767 (N_15767,N_15546,N_15453);
xor U15768 (N_15768,N_15500,N_15419);
nand U15769 (N_15769,N_15568,N_15511);
nor U15770 (N_15770,N_15482,N_15501);
nor U15771 (N_15771,N_15498,N_15454);
nor U15772 (N_15772,N_15501,N_15494);
and U15773 (N_15773,N_15550,N_15554);
and U15774 (N_15774,N_15411,N_15435);
and U15775 (N_15775,N_15566,N_15499);
and U15776 (N_15776,N_15502,N_15577);
and U15777 (N_15777,N_15461,N_15434);
or U15778 (N_15778,N_15474,N_15580);
xnor U15779 (N_15779,N_15505,N_15499);
nand U15780 (N_15780,N_15507,N_15448);
nand U15781 (N_15781,N_15577,N_15500);
xnor U15782 (N_15782,N_15590,N_15422);
nor U15783 (N_15783,N_15431,N_15515);
or U15784 (N_15784,N_15527,N_15465);
nand U15785 (N_15785,N_15534,N_15503);
nand U15786 (N_15786,N_15505,N_15434);
nand U15787 (N_15787,N_15479,N_15587);
or U15788 (N_15788,N_15447,N_15424);
or U15789 (N_15789,N_15533,N_15405);
and U15790 (N_15790,N_15583,N_15467);
or U15791 (N_15791,N_15433,N_15490);
xor U15792 (N_15792,N_15441,N_15410);
nand U15793 (N_15793,N_15513,N_15481);
nand U15794 (N_15794,N_15567,N_15434);
nor U15795 (N_15795,N_15580,N_15451);
nand U15796 (N_15796,N_15413,N_15457);
nor U15797 (N_15797,N_15438,N_15476);
or U15798 (N_15798,N_15505,N_15501);
and U15799 (N_15799,N_15506,N_15560);
or U15800 (N_15800,N_15639,N_15739);
and U15801 (N_15801,N_15767,N_15768);
xor U15802 (N_15802,N_15717,N_15763);
or U15803 (N_15803,N_15750,N_15760);
nand U15804 (N_15804,N_15791,N_15728);
nand U15805 (N_15805,N_15651,N_15631);
xnor U15806 (N_15806,N_15633,N_15795);
or U15807 (N_15807,N_15744,N_15604);
and U15808 (N_15808,N_15723,N_15673);
nor U15809 (N_15809,N_15688,N_15764);
xnor U15810 (N_15810,N_15692,N_15612);
nand U15811 (N_15811,N_15709,N_15799);
or U15812 (N_15812,N_15691,N_15731);
and U15813 (N_15813,N_15742,N_15664);
nor U15814 (N_15814,N_15652,N_15658);
nor U15815 (N_15815,N_15655,N_15787);
nor U15816 (N_15816,N_15783,N_15666);
and U15817 (N_15817,N_15670,N_15644);
nand U15818 (N_15818,N_15766,N_15672);
nor U15819 (N_15819,N_15732,N_15625);
nor U15820 (N_15820,N_15699,N_15701);
nor U15821 (N_15821,N_15719,N_15754);
or U15822 (N_15822,N_15635,N_15659);
or U15823 (N_15823,N_15778,N_15720);
or U15824 (N_15824,N_15648,N_15789);
or U15825 (N_15825,N_15645,N_15794);
and U15826 (N_15826,N_15657,N_15640);
or U15827 (N_15827,N_15756,N_15653);
and U15828 (N_15828,N_15674,N_15753);
nor U15829 (N_15829,N_15704,N_15602);
and U15830 (N_15830,N_15637,N_15777);
nand U15831 (N_15831,N_15682,N_15618);
nor U15832 (N_15832,N_15622,N_15698);
xor U15833 (N_15833,N_15727,N_15780);
xor U15834 (N_15834,N_15729,N_15738);
and U15835 (N_15835,N_15662,N_15733);
nor U15836 (N_15836,N_15661,N_15788);
and U15837 (N_15837,N_15685,N_15758);
nand U15838 (N_15838,N_15675,N_15703);
nor U15839 (N_15839,N_15748,N_15647);
nor U15840 (N_15840,N_15663,N_15686);
xnor U15841 (N_15841,N_15734,N_15743);
nand U15842 (N_15842,N_15684,N_15683);
nor U15843 (N_15843,N_15718,N_15649);
or U15844 (N_15844,N_15642,N_15679);
xor U15845 (N_15845,N_15715,N_15724);
xnor U15846 (N_15846,N_15707,N_15779);
xnor U15847 (N_15847,N_15740,N_15790);
and U15848 (N_15848,N_15722,N_15601);
nand U15849 (N_15849,N_15693,N_15792);
nand U15850 (N_15850,N_15609,N_15700);
nor U15851 (N_15851,N_15669,N_15615);
or U15852 (N_15852,N_15606,N_15726);
xor U15853 (N_15853,N_15759,N_15628);
or U15854 (N_15854,N_15770,N_15678);
and U15855 (N_15855,N_15775,N_15741);
and U15856 (N_15856,N_15690,N_15751);
and U15857 (N_15857,N_15749,N_15681);
xnor U15858 (N_15858,N_15676,N_15735);
and U15859 (N_15859,N_15621,N_15725);
or U15860 (N_15860,N_15614,N_15773);
nand U15861 (N_15861,N_15708,N_15706);
nand U15862 (N_15862,N_15797,N_15747);
nand U15863 (N_15863,N_15736,N_15757);
nand U15864 (N_15864,N_15607,N_15755);
nand U15865 (N_15865,N_15638,N_15746);
xnor U15866 (N_15866,N_15680,N_15721);
xnor U15867 (N_15867,N_15603,N_15786);
nor U15868 (N_15868,N_15626,N_15782);
nand U15869 (N_15869,N_15713,N_15714);
and U15870 (N_15870,N_15711,N_15776);
and U15871 (N_15871,N_15712,N_15689);
and U15872 (N_15872,N_15696,N_15694);
nor U15873 (N_15873,N_15667,N_15774);
nand U15874 (N_15874,N_15646,N_15769);
or U15875 (N_15875,N_15613,N_15771);
nand U15876 (N_15876,N_15695,N_15761);
nor U15877 (N_15877,N_15697,N_15793);
nand U15878 (N_15878,N_15796,N_15641);
nand U15879 (N_15879,N_15634,N_15710);
xnor U15880 (N_15880,N_15608,N_15730);
and U15881 (N_15881,N_15781,N_15762);
or U15882 (N_15882,N_15702,N_15716);
and U15883 (N_15883,N_15752,N_15671);
nor U15884 (N_15884,N_15616,N_15643);
nor U15885 (N_15885,N_15632,N_15660);
and U15886 (N_15886,N_15665,N_15784);
xor U15887 (N_15887,N_15745,N_15668);
nor U15888 (N_15888,N_15629,N_15630);
and U15889 (N_15889,N_15623,N_15785);
or U15890 (N_15890,N_15765,N_15677);
or U15891 (N_15891,N_15636,N_15619);
nand U15892 (N_15892,N_15656,N_15737);
nand U15893 (N_15893,N_15687,N_15600);
xnor U15894 (N_15894,N_15610,N_15705);
nand U15895 (N_15895,N_15654,N_15798);
or U15896 (N_15896,N_15772,N_15611);
nand U15897 (N_15897,N_15650,N_15627);
nand U15898 (N_15898,N_15624,N_15605);
nor U15899 (N_15899,N_15617,N_15620);
nor U15900 (N_15900,N_15676,N_15661);
or U15901 (N_15901,N_15611,N_15677);
nor U15902 (N_15902,N_15770,N_15764);
xnor U15903 (N_15903,N_15692,N_15667);
and U15904 (N_15904,N_15749,N_15797);
xor U15905 (N_15905,N_15702,N_15620);
and U15906 (N_15906,N_15641,N_15628);
or U15907 (N_15907,N_15722,N_15665);
xor U15908 (N_15908,N_15651,N_15664);
xor U15909 (N_15909,N_15715,N_15716);
and U15910 (N_15910,N_15630,N_15722);
nor U15911 (N_15911,N_15759,N_15713);
and U15912 (N_15912,N_15687,N_15708);
nand U15913 (N_15913,N_15646,N_15650);
xor U15914 (N_15914,N_15713,N_15772);
and U15915 (N_15915,N_15793,N_15630);
xnor U15916 (N_15916,N_15667,N_15714);
nand U15917 (N_15917,N_15751,N_15734);
and U15918 (N_15918,N_15722,N_15677);
and U15919 (N_15919,N_15672,N_15704);
nor U15920 (N_15920,N_15681,N_15697);
xor U15921 (N_15921,N_15788,N_15678);
and U15922 (N_15922,N_15750,N_15659);
or U15923 (N_15923,N_15723,N_15753);
or U15924 (N_15924,N_15623,N_15684);
or U15925 (N_15925,N_15761,N_15778);
and U15926 (N_15926,N_15719,N_15626);
and U15927 (N_15927,N_15622,N_15673);
nor U15928 (N_15928,N_15757,N_15784);
nor U15929 (N_15929,N_15616,N_15717);
and U15930 (N_15930,N_15655,N_15738);
or U15931 (N_15931,N_15654,N_15631);
xnor U15932 (N_15932,N_15734,N_15785);
nor U15933 (N_15933,N_15680,N_15699);
xor U15934 (N_15934,N_15680,N_15708);
and U15935 (N_15935,N_15668,N_15632);
or U15936 (N_15936,N_15717,N_15686);
or U15937 (N_15937,N_15716,N_15649);
and U15938 (N_15938,N_15695,N_15661);
xor U15939 (N_15939,N_15721,N_15689);
nand U15940 (N_15940,N_15666,N_15744);
nor U15941 (N_15941,N_15619,N_15698);
nand U15942 (N_15942,N_15770,N_15701);
nor U15943 (N_15943,N_15681,N_15675);
nand U15944 (N_15944,N_15633,N_15654);
xnor U15945 (N_15945,N_15634,N_15617);
and U15946 (N_15946,N_15609,N_15707);
xor U15947 (N_15947,N_15613,N_15697);
nand U15948 (N_15948,N_15721,N_15765);
and U15949 (N_15949,N_15616,N_15662);
and U15950 (N_15950,N_15722,N_15776);
and U15951 (N_15951,N_15763,N_15729);
xnor U15952 (N_15952,N_15608,N_15655);
or U15953 (N_15953,N_15713,N_15703);
nand U15954 (N_15954,N_15761,N_15628);
xnor U15955 (N_15955,N_15720,N_15728);
nand U15956 (N_15956,N_15602,N_15712);
xor U15957 (N_15957,N_15615,N_15794);
nand U15958 (N_15958,N_15724,N_15733);
xor U15959 (N_15959,N_15783,N_15721);
nor U15960 (N_15960,N_15678,N_15639);
xnor U15961 (N_15961,N_15729,N_15690);
xnor U15962 (N_15962,N_15672,N_15647);
and U15963 (N_15963,N_15613,N_15657);
xor U15964 (N_15964,N_15626,N_15634);
or U15965 (N_15965,N_15650,N_15700);
xnor U15966 (N_15966,N_15694,N_15691);
nor U15967 (N_15967,N_15623,N_15783);
nand U15968 (N_15968,N_15620,N_15731);
xor U15969 (N_15969,N_15715,N_15727);
xnor U15970 (N_15970,N_15747,N_15722);
nand U15971 (N_15971,N_15644,N_15723);
nand U15972 (N_15972,N_15708,N_15779);
or U15973 (N_15973,N_15742,N_15774);
xnor U15974 (N_15974,N_15786,N_15660);
and U15975 (N_15975,N_15666,N_15645);
and U15976 (N_15976,N_15662,N_15702);
nand U15977 (N_15977,N_15756,N_15775);
or U15978 (N_15978,N_15616,N_15712);
nor U15979 (N_15979,N_15686,N_15715);
xnor U15980 (N_15980,N_15616,N_15644);
xnor U15981 (N_15981,N_15715,N_15748);
or U15982 (N_15982,N_15753,N_15687);
xor U15983 (N_15983,N_15782,N_15602);
or U15984 (N_15984,N_15609,N_15606);
or U15985 (N_15985,N_15624,N_15626);
nand U15986 (N_15986,N_15689,N_15704);
and U15987 (N_15987,N_15711,N_15601);
xor U15988 (N_15988,N_15623,N_15602);
nor U15989 (N_15989,N_15772,N_15793);
or U15990 (N_15990,N_15658,N_15684);
nand U15991 (N_15991,N_15634,N_15719);
nor U15992 (N_15992,N_15787,N_15603);
nor U15993 (N_15993,N_15778,N_15725);
nor U15994 (N_15994,N_15689,N_15629);
and U15995 (N_15995,N_15695,N_15728);
nor U15996 (N_15996,N_15606,N_15699);
and U15997 (N_15997,N_15758,N_15734);
nor U15998 (N_15998,N_15662,N_15620);
nand U15999 (N_15999,N_15778,N_15785);
xor U16000 (N_16000,N_15877,N_15982);
nand U16001 (N_16001,N_15914,N_15889);
nor U16002 (N_16002,N_15987,N_15801);
and U16003 (N_16003,N_15851,N_15836);
xor U16004 (N_16004,N_15913,N_15902);
xnor U16005 (N_16005,N_15918,N_15832);
nand U16006 (N_16006,N_15938,N_15948);
nand U16007 (N_16007,N_15890,N_15994);
or U16008 (N_16008,N_15971,N_15924);
or U16009 (N_16009,N_15995,N_15999);
nor U16010 (N_16010,N_15858,N_15867);
or U16011 (N_16011,N_15865,N_15800);
nor U16012 (N_16012,N_15937,N_15952);
and U16013 (N_16013,N_15803,N_15906);
nor U16014 (N_16014,N_15912,N_15864);
nand U16015 (N_16015,N_15961,N_15950);
nor U16016 (N_16016,N_15888,N_15857);
nand U16017 (N_16017,N_15828,N_15977);
or U16018 (N_16018,N_15830,N_15817);
nand U16019 (N_16019,N_15827,N_15835);
or U16020 (N_16020,N_15855,N_15869);
nand U16021 (N_16021,N_15942,N_15845);
nor U16022 (N_16022,N_15842,N_15873);
xor U16023 (N_16023,N_15993,N_15837);
and U16024 (N_16024,N_15926,N_15921);
and U16025 (N_16025,N_15911,N_15949);
nand U16026 (N_16026,N_15820,N_15976);
and U16027 (N_16027,N_15932,N_15881);
nand U16028 (N_16028,N_15829,N_15958);
nor U16029 (N_16029,N_15834,N_15962);
or U16030 (N_16030,N_15894,N_15808);
nor U16031 (N_16031,N_15963,N_15807);
nand U16032 (N_16032,N_15939,N_15998);
or U16033 (N_16033,N_15856,N_15981);
xnor U16034 (N_16034,N_15893,N_15821);
nor U16035 (N_16035,N_15900,N_15879);
nand U16036 (N_16036,N_15805,N_15874);
and U16037 (N_16037,N_15959,N_15984);
xnor U16038 (N_16038,N_15986,N_15996);
nor U16039 (N_16039,N_15839,N_15969);
nand U16040 (N_16040,N_15974,N_15885);
xor U16041 (N_16041,N_15819,N_15980);
xor U16042 (N_16042,N_15871,N_15811);
and U16043 (N_16043,N_15810,N_15957);
and U16044 (N_16044,N_15866,N_15823);
xnor U16045 (N_16045,N_15850,N_15843);
nor U16046 (N_16046,N_15813,N_15804);
nor U16047 (N_16047,N_15951,N_15920);
or U16048 (N_16048,N_15841,N_15972);
xnor U16049 (N_16049,N_15901,N_15973);
nor U16050 (N_16050,N_15929,N_15822);
xnor U16051 (N_16051,N_15824,N_15956);
xnor U16052 (N_16052,N_15891,N_15991);
or U16053 (N_16053,N_15966,N_15935);
nor U16054 (N_16054,N_15988,N_15933);
xnor U16055 (N_16055,N_15979,N_15849);
and U16056 (N_16056,N_15954,N_15947);
and U16057 (N_16057,N_15847,N_15903);
and U16058 (N_16058,N_15990,N_15915);
nor U16059 (N_16059,N_15964,N_15909);
xnor U16060 (N_16060,N_15953,N_15919);
nor U16061 (N_16061,N_15928,N_15838);
nor U16062 (N_16062,N_15814,N_15989);
nand U16063 (N_16063,N_15848,N_15936);
or U16064 (N_16064,N_15944,N_15965);
nor U16065 (N_16065,N_15960,N_15863);
nand U16066 (N_16066,N_15897,N_15923);
nor U16067 (N_16067,N_15852,N_15895);
or U16068 (N_16068,N_15861,N_15868);
and U16069 (N_16069,N_15802,N_15859);
nand U16070 (N_16070,N_15908,N_15955);
nor U16071 (N_16071,N_15883,N_15886);
nand U16072 (N_16072,N_15904,N_15940);
nor U16073 (N_16073,N_15840,N_15978);
xor U16074 (N_16074,N_15816,N_15870);
and U16075 (N_16075,N_15898,N_15882);
nand U16076 (N_16076,N_15872,N_15910);
xor U16077 (N_16077,N_15818,N_15968);
xnor U16078 (N_16078,N_15876,N_15905);
or U16079 (N_16079,N_15916,N_15809);
or U16080 (N_16080,N_15997,N_15930);
or U16081 (N_16081,N_15860,N_15907);
or U16082 (N_16082,N_15878,N_15985);
xor U16083 (N_16083,N_15922,N_15862);
xnor U16084 (N_16084,N_15846,N_15880);
or U16085 (N_16085,N_15853,N_15887);
nand U16086 (N_16086,N_15967,N_15927);
xor U16087 (N_16087,N_15812,N_15892);
xor U16088 (N_16088,N_15831,N_15970);
or U16089 (N_16089,N_15833,N_15983);
and U16090 (N_16090,N_15975,N_15946);
nand U16091 (N_16091,N_15884,N_15931);
xor U16092 (N_16092,N_15943,N_15806);
nor U16093 (N_16093,N_15826,N_15844);
or U16094 (N_16094,N_15917,N_15945);
xor U16095 (N_16095,N_15825,N_15899);
nand U16096 (N_16096,N_15941,N_15854);
or U16097 (N_16097,N_15896,N_15875);
nor U16098 (N_16098,N_15934,N_15815);
nand U16099 (N_16099,N_15925,N_15992);
or U16100 (N_16100,N_15824,N_15865);
or U16101 (N_16101,N_15969,N_15869);
nor U16102 (N_16102,N_15948,N_15983);
or U16103 (N_16103,N_15882,N_15978);
or U16104 (N_16104,N_15800,N_15924);
nand U16105 (N_16105,N_15950,N_15849);
nand U16106 (N_16106,N_15979,N_15952);
nand U16107 (N_16107,N_15896,N_15971);
and U16108 (N_16108,N_15858,N_15856);
nor U16109 (N_16109,N_15838,N_15842);
xor U16110 (N_16110,N_15813,N_15955);
xnor U16111 (N_16111,N_15841,N_15953);
or U16112 (N_16112,N_15931,N_15806);
xnor U16113 (N_16113,N_15818,N_15980);
nand U16114 (N_16114,N_15945,N_15813);
and U16115 (N_16115,N_15888,N_15896);
and U16116 (N_16116,N_15977,N_15967);
xor U16117 (N_16117,N_15968,N_15854);
and U16118 (N_16118,N_15817,N_15819);
xnor U16119 (N_16119,N_15938,N_15846);
xor U16120 (N_16120,N_15822,N_15933);
or U16121 (N_16121,N_15893,N_15883);
and U16122 (N_16122,N_15952,N_15848);
nor U16123 (N_16123,N_15859,N_15882);
or U16124 (N_16124,N_15902,N_15897);
nand U16125 (N_16125,N_15906,N_15919);
nor U16126 (N_16126,N_15840,N_15818);
xnor U16127 (N_16127,N_15909,N_15993);
or U16128 (N_16128,N_15840,N_15882);
xnor U16129 (N_16129,N_15844,N_15934);
nor U16130 (N_16130,N_15824,N_15931);
xor U16131 (N_16131,N_15876,N_15868);
nand U16132 (N_16132,N_15801,N_15955);
or U16133 (N_16133,N_15998,N_15820);
xor U16134 (N_16134,N_15950,N_15940);
or U16135 (N_16135,N_15938,N_15919);
xnor U16136 (N_16136,N_15865,N_15995);
xnor U16137 (N_16137,N_15977,N_15837);
and U16138 (N_16138,N_15824,N_15897);
or U16139 (N_16139,N_15865,N_15807);
or U16140 (N_16140,N_15844,N_15946);
nand U16141 (N_16141,N_15987,N_15976);
and U16142 (N_16142,N_15847,N_15838);
and U16143 (N_16143,N_15918,N_15928);
or U16144 (N_16144,N_15929,N_15987);
xnor U16145 (N_16145,N_15981,N_15901);
nor U16146 (N_16146,N_15920,N_15908);
nor U16147 (N_16147,N_15815,N_15883);
nand U16148 (N_16148,N_15961,N_15816);
nor U16149 (N_16149,N_15858,N_15851);
nand U16150 (N_16150,N_15922,N_15934);
nor U16151 (N_16151,N_15972,N_15963);
and U16152 (N_16152,N_15919,N_15926);
xnor U16153 (N_16153,N_15945,N_15891);
nand U16154 (N_16154,N_15934,N_15881);
nor U16155 (N_16155,N_15950,N_15966);
xnor U16156 (N_16156,N_15932,N_15941);
nand U16157 (N_16157,N_15945,N_15988);
and U16158 (N_16158,N_15988,N_15991);
and U16159 (N_16159,N_15839,N_15909);
or U16160 (N_16160,N_15923,N_15813);
and U16161 (N_16161,N_15925,N_15924);
or U16162 (N_16162,N_15843,N_15989);
or U16163 (N_16163,N_15959,N_15825);
and U16164 (N_16164,N_15892,N_15871);
nor U16165 (N_16165,N_15984,N_15979);
or U16166 (N_16166,N_15867,N_15946);
and U16167 (N_16167,N_15927,N_15900);
and U16168 (N_16168,N_15851,N_15856);
nand U16169 (N_16169,N_15950,N_15960);
and U16170 (N_16170,N_15857,N_15865);
and U16171 (N_16171,N_15877,N_15821);
xnor U16172 (N_16172,N_15910,N_15882);
nand U16173 (N_16173,N_15860,N_15969);
and U16174 (N_16174,N_15900,N_15968);
nand U16175 (N_16175,N_15893,N_15873);
xnor U16176 (N_16176,N_15819,N_15826);
or U16177 (N_16177,N_15865,N_15933);
and U16178 (N_16178,N_15804,N_15829);
xor U16179 (N_16179,N_15823,N_15950);
nand U16180 (N_16180,N_15852,N_15822);
xnor U16181 (N_16181,N_15845,N_15963);
xor U16182 (N_16182,N_15873,N_15966);
nand U16183 (N_16183,N_15882,N_15948);
and U16184 (N_16184,N_15813,N_15805);
or U16185 (N_16185,N_15821,N_15822);
xor U16186 (N_16186,N_15973,N_15904);
nand U16187 (N_16187,N_15892,N_15948);
nor U16188 (N_16188,N_15980,N_15846);
nand U16189 (N_16189,N_15918,N_15989);
nor U16190 (N_16190,N_15826,N_15818);
or U16191 (N_16191,N_15903,N_15865);
or U16192 (N_16192,N_15939,N_15814);
xor U16193 (N_16193,N_15830,N_15931);
and U16194 (N_16194,N_15894,N_15996);
nand U16195 (N_16195,N_15844,N_15984);
or U16196 (N_16196,N_15876,N_15975);
or U16197 (N_16197,N_15811,N_15820);
nand U16198 (N_16198,N_15873,N_15852);
xnor U16199 (N_16199,N_15985,N_15980);
xnor U16200 (N_16200,N_16146,N_16090);
or U16201 (N_16201,N_16152,N_16032);
nor U16202 (N_16202,N_16075,N_16154);
or U16203 (N_16203,N_16134,N_16182);
nor U16204 (N_16204,N_16170,N_16022);
nor U16205 (N_16205,N_16017,N_16161);
xor U16206 (N_16206,N_16093,N_16116);
and U16207 (N_16207,N_16054,N_16163);
nor U16208 (N_16208,N_16003,N_16120);
xnor U16209 (N_16209,N_16119,N_16064);
nor U16210 (N_16210,N_16009,N_16164);
xnor U16211 (N_16211,N_16097,N_16034);
nand U16212 (N_16212,N_16061,N_16013);
and U16213 (N_16213,N_16121,N_16028);
nand U16214 (N_16214,N_16102,N_16157);
and U16215 (N_16215,N_16142,N_16143);
or U16216 (N_16216,N_16124,N_16077);
and U16217 (N_16217,N_16048,N_16010);
or U16218 (N_16218,N_16132,N_16070);
or U16219 (N_16219,N_16079,N_16059);
xnor U16220 (N_16220,N_16108,N_16029);
nor U16221 (N_16221,N_16158,N_16055);
nand U16222 (N_16222,N_16083,N_16072);
nor U16223 (N_16223,N_16160,N_16178);
and U16224 (N_16224,N_16080,N_16033);
or U16225 (N_16225,N_16172,N_16051);
xnor U16226 (N_16226,N_16062,N_16197);
xnor U16227 (N_16227,N_16196,N_16094);
and U16228 (N_16228,N_16128,N_16037);
nand U16229 (N_16229,N_16049,N_16151);
xor U16230 (N_16230,N_16141,N_16006);
xnor U16231 (N_16231,N_16130,N_16195);
xor U16232 (N_16232,N_16100,N_16180);
nor U16233 (N_16233,N_16082,N_16018);
or U16234 (N_16234,N_16042,N_16139);
nor U16235 (N_16235,N_16066,N_16174);
and U16236 (N_16236,N_16117,N_16167);
and U16237 (N_16237,N_16085,N_16004);
nand U16238 (N_16238,N_16112,N_16067);
nor U16239 (N_16239,N_16052,N_16069);
nor U16240 (N_16240,N_16068,N_16145);
and U16241 (N_16241,N_16138,N_16110);
nand U16242 (N_16242,N_16000,N_16104);
or U16243 (N_16243,N_16084,N_16187);
nand U16244 (N_16244,N_16137,N_16191);
xor U16245 (N_16245,N_16183,N_16113);
xnor U16246 (N_16246,N_16162,N_16140);
and U16247 (N_16247,N_16019,N_16041);
and U16248 (N_16248,N_16099,N_16007);
and U16249 (N_16249,N_16098,N_16103);
nor U16250 (N_16250,N_16192,N_16005);
or U16251 (N_16251,N_16115,N_16078);
nor U16252 (N_16252,N_16176,N_16168);
and U16253 (N_16253,N_16107,N_16184);
or U16254 (N_16254,N_16065,N_16091);
nand U16255 (N_16255,N_16111,N_16159);
nand U16256 (N_16256,N_16012,N_16088);
nor U16257 (N_16257,N_16147,N_16060);
or U16258 (N_16258,N_16076,N_16073);
and U16259 (N_16259,N_16135,N_16092);
or U16260 (N_16260,N_16096,N_16122);
xnor U16261 (N_16261,N_16058,N_16189);
nand U16262 (N_16262,N_16074,N_16153);
and U16263 (N_16263,N_16109,N_16125);
and U16264 (N_16264,N_16044,N_16181);
and U16265 (N_16265,N_16021,N_16169);
xnor U16266 (N_16266,N_16001,N_16035);
nand U16267 (N_16267,N_16188,N_16002);
nand U16268 (N_16268,N_16015,N_16045);
nand U16269 (N_16269,N_16105,N_16086);
nand U16270 (N_16270,N_16038,N_16056);
xor U16271 (N_16271,N_16148,N_16123);
and U16272 (N_16272,N_16173,N_16129);
nand U16273 (N_16273,N_16150,N_16190);
nor U16274 (N_16274,N_16185,N_16040);
or U16275 (N_16275,N_16026,N_16016);
nand U16276 (N_16276,N_16063,N_16114);
xnor U16277 (N_16277,N_16199,N_16030);
nor U16278 (N_16278,N_16081,N_16050);
xor U16279 (N_16279,N_16011,N_16101);
nand U16280 (N_16280,N_16027,N_16171);
or U16281 (N_16281,N_16179,N_16046);
xor U16282 (N_16282,N_16057,N_16039);
nor U16283 (N_16283,N_16127,N_16071);
nand U16284 (N_16284,N_16024,N_16095);
nor U16285 (N_16285,N_16025,N_16131);
xor U16286 (N_16286,N_16043,N_16031);
nand U16287 (N_16287,N_16126,N_16144);
or U16288 (N_16288,N_16008,N_16194);
nand U16289 (N_16289,N_16186,N_16014);
and U16290 (N_16290,N_16193,N_16177);
xnor U16291 (N_16291,N_16020,N_16149);
and U16292 (N_16292,N_16053,N_16136);
nand U16293 (N_16293,N_16047,N_16089);
nor U16294 (N_16294,N_16198,N_16118);
and U16295 (N_16295,N_16156,N_16023);
xor U16296 (N_16296,N_16036,N_16175);
xor U16297 (N_16297,N_16133,N_16165);
or U16298 (N_16298,N_16106,N_16166);
nor U16299 (N_16299,N_16155,N_16087);
nor U16300 (N_16300,N_16191,N_16032);
and U16301 (N_16301,N_16050,N_16129);
or U16302 (N_16302,N_16061,N_16156);
nor U16303 (N_16303,N_16029,N_16047);
xnor U16304 (N_16304,N_16041,N_16170);
xor U16305 (N_16305,N_16037,N_16164);
nor U16306 (N_16306,N_16155,N_16073);
or U16307 (N_16307,N_16039,N_16164);
nor U16308 (N_16308,N_16062,N_16149);
nor U16309 (N_16309,N_16134,N_16170);
nor U16310 (N_16310,N_16114,N_16057);
and U16311 (N_16311,N_16025,N_16141);
or U16312 (N_16312,N_16197,N_16032);
nor U16313 (N_16313,N_16178,N_16112);
xnor U16314 (N_16314,N_16118,N_16037);
nor U16315 (N_16315,N_16170,N_16070);
or U16316 (N_16316,N_16191,N_16119);
xor U16317 (N_16317,N_16073,N_16008);
nor U16318 (N_16318,N_16198,N_16101);
xnor U16319 (N_16319,N_16006,N_16099);
and U16320 (N_16320,N_16039,N_16051);
and U16321 (N_16321,N_16139,N_16055);
and U16322 (N_16322,N_16146,N_16194);
nand U16323 (N_16323,N_16167,N_16042);
nor U16324 (N_16324,N_16116,N_16163);
xnor U16325 (N_16325,N_16055,N_16110);
nor U16326 (N_16326,N_16054,N_16057);
nor U16327 (N_16327,N_16098,N_16014);
nand U16328 (N_16328,N_16143,N_16081);
and U16329 (N_16329,N_16011,N_16163);
nor U16330 (N_16330,N_16181,N_16007);
nand U16331 (N_16331,N_16126,N_16163);
and U16332 (N_16332,N_16005,N_16000);
or U16333 (N_16333,N_16186,N_16194);
nand U16334 (N_16334,N_16011,N_16060);
and U16335 (N_16335,N_16175,N_16062);
or U16336 (N_16336,N_16006,N_16179);
and U16337 (N_16337,N_16049,N_16134);
xnor U16338 (N_16338,N_16101,N_16017);
nand U16339 (N_16339,N_16010,N_16197);
and U16340 (N_16340,N_16002,N_16052);
and U16341 (N_16341,N_16141,N_16149);
or U16342 (N_16342,N_16104,N_16018);
or U16343 (N_16343,N_16009,N_16168);
nor U16344 (N_16344,N_16091,N_16014);
or U16345 (N_16345,N_16020,N_16156);
xor U16346 (N_16346,N_16030,N_16042);
or U16347 (N_16347,N_16096,N_16109);
xnor U16348 (N_16348,N_16133,N_16047);
nand U16349 (N_16349,N_16134,N_16043);
nand U16350 (N_16350,N_16146,N_16059);
nor U16351 (N_16351,N_16188,N_16071);
and U16352 (N_16352,N_16027,N_16041);
or U16353 (N_16353,N_16061,N_16087);
and U16354 (N_16354,N_16055,N_16097);
or U16355 (N_16355,N_16055,N_16135);
and U16356 (N_16356,N_16073,N_16080);
nor U16357 (N_16357,N_16185,N_16049);
or U16358 (N_16358,N_16145,N_16092);
nor U16359 (N_16359,N_16069,N_16105);
nand U16360 (N_16360,N_16119,N_16170);
xnor U16361 (N_16361,N_16123,N_16035);
or U16362 (N_16362,N_16133,N_16003);
and U16363 (N_16363,N_16038,N_16178);
or U16364 (N_16364,N_16035,N_16167);
nor U16365 (N_16365,N_16056,N_16103);
and U16366 (N_16366,N_16113,N_16068);
and U16367 (N_16367,N_16098,N_16006);
and U16368 (N_16368,N_16129,N_16077);
and U16369 (N_16369,N_16139,N_16041);
nand U16370 (N_16370,N_16184,N_16139);
nand U16371 (N_16371,N_16064,N_16167);
or U16372 (N_16372,N_16107,N_16040);
nor U16373 (N_16373,N_16091,N_16180);
nand U16374 (N_16374,N_16072,N_16002);
nand U16375 (N_16375,N_16078,N_16113);
and U16376 (N_16376,N_16165,N_16147);
xnor U16377 (N_16377,N_16020,N_16127);
and U16378 (N_16378,N_16177,N_16130);
or U16379 (N_16379,N_16125,N_16061);
and U16380 (N_16380,N_16072,N_16065);
and U16381 (N_16381,N_16065,N_16023);
nand U16382 (N_16382,N_16044,N_16041);
or U16383 (N_16383,N_16133,N_16127);
or U16384 (N_16384,N_16141,N_16074);
or U16385 (N_16385,N_16017,N_16091);
or U16386 (N_16386,N_16042,N_16102);
or U16387 (N_16387,N_16028,N_16179);
nor U16388 (N_16388,N_16125,N_16013);
nor U16389 (N_16389,N_16054,N_16102);
nand U16390 (N_16390,N_16063,N_16181);
nor U16391 (N_16391,N_16089,N_16174);
nand U16392 (N_16392,N_16002,N_16010);
xor U16393 (N_16393,N_16082,N_16130);
xor U16394 (N_16394,N_16079,N_16045);
and U16395 (N_16395,N_16106,N_16003);
or U16396 (N_16396,N_16127,N_16079);
and U16397 (N_16397,N_16004,N_16132);
and U16398 (N_16398,N_16052,N_16059);
and U16399 (N_16399,N_16095,N_16155);
and U16400 (N_16400,N_16356,N_16239);
xnor U16401 (N_16401,N_16231,N_16253);
nand U16402 (N_16402,N_16343,N_16213);
nor U16403 (N_16403,N_16328,N_16291);
nor U16404 (N_16404,N_16273,N_16352);
nand U16405 (N_16405,N_16349,N_16351);
or U16406 (N_16406,N_16218,N_16260);
nor U16407 (N_16407,N_16300,N_16340);
nand U16408 (N_16408,N_16226,N_16211);
nor U16409 (N_16409,N_16290,N_16261);
nand U16410 (N_16410,N_16238,N_16311);
and U16411 (N_16411,N_16358,N_16284);
nor U16412 (N_16412,N_16237,N_16360);
nor U16413 (N_16413,N_16350,N_16301);
nand U16414 (N_16414,N_16299,N_16269);
xnor U16415 (N_16415,N_16287,N_16381);
or U16416 (N_16416,N_16205,N_16251);
and U16417 (N_16417,N_16235,N_16230);
xnor U16418 (N_16418,N_16310,N_16252);
or U16419 (N_16419,N_16225,N_16374);
nor U16420 (N_16420,N_16370,N_16362);
and U16421 (N_16421,N_16314,N_16215);
or U16422 (N_16422,N_16276,N_16308);
nand U16423 (N_16423,N_16289,N_16397);
nand U16424 (N_16424,N_16375,N_16278);
xor U16425 (N_16425,N_16272,N_16206);
xnor U16426 (N_16426,N_16361,N_16382);
nand U16427 (N_16427,N_16214,N_16322);
nand U16428 (N_16428,N_16378,N_16388);
and U16429 (N_16429,N_16280,N_16236);
or U16430 (N_16430,N_16336,N_16248);
and U16431 (N_16431,N_16221,N_16293);
or U16432 (N_16432,N_16354,N_16200);
and U16433 (N_16433,N_16243,N_16249);
nor U16434 (N_16434,N_16304,N_16346);
and U16435 (N_16435,N_16219,N_16371);
nor U16436 (N_16436,N_16222,N_16247);
or U16437 (N_16437,N_16302,N_16357);
or U16438 (N_16438,N_16359,N_16233);
or U16439 (N_16439,N_16394,N_16318);
xor U16440 (N_16440,N_16285,N_16331);
or U16441 (N_16441,N_16320,N_16342);
and U16442 (N_16442,N_16334,N_16244);
nor U16443 (N_16443,N_16212,N_16333);
nand U16444 (N_16444,N_16365,N_16232);
and U16445 (N_16445,N_16377,N_16203);
xor U16446 (N_16446,N_16355,N_16202);
nor U16447 (N_16447,N_16270,N_16345);
nand U16448 (N_16448,N_16325,N_16316);
or U16449 (N_16449,N_16368,N_16242);
and U16450 (N_16450,N_16204,N_16386);
xor U16451 (N_16451,N_16383,N_16353);
xnor U16452 (N_16452,N_16389,N_16312);
xnor U16453 (N_16453,N_16209,N_16305);
or U16454 (N_16454,N_16294,N_16387);
xnor U16455 (N_16455,N_16330,N_16283);
nor U16456 (N_16456,N_16262,N_16347);
xnor U16457 (N_16457,N_16366,N_16391);
and U16458 (N_16458,N_16399,N_16201);
nand U16459 (N_16459,N_16227,N_16220);
or U16460 (N_16460,N_16392,N_16250);
xnor U16461 (N_16461,N_16246,N_16210);
nor U16462 (N_16462,N_16324,N_16315);
nand U16463 (N_16463,N_16376,N_16326);
or U16464 (N_16464,N_16297,N_16337);
or U16465 (N_16465,N_16275,N_16256);
xor U16466 (N_16466,N_16373,N_16228);
or U16467 (N_16467,N_16254,N_16379);
xor U16468 (N_16468,N_16264,N_16319);
and U16469 (N_16469,N_16332,N_16295);
nor U16470 (N_16470,N_16385,N_16288);
and U16471 (N_16471,N_16234,N_16323);
and U16472 (N_16472,N_16281,N_16309);
or U16473 (N_16473,N_16384,N_16207);
or U16474 (N_16474,N_16263,N_16241);
nor U16475 (N_16475,N_16363,N_16372);
or U16476 (N_16476,N_16279,N_16268);
nor U16477 (N_16477,N_16208,N_16321);
nand U16478 (N_16478,N_16395,N_16245);
and U16479 (N_16479,N_16258,N_16292);
xnor U16480 (N_16480,N_16306,N_16229);
and U16481 (N_16481,N_16303,N_16348);
or U16482 (N_16482,N_16296,N_16367);
nor U16483 (N_16483,N_16277,N_16307);
or U16484 (N_16484,N_16398,N_16266);
and U16485 (N_16485,N_16265,N_16390);
nand U16486 (N_16486,N_16335,N_16271);
nand U16487 (N_16487,N_16298,N_16338);
nand U16488 (N_16488,N_16217,N_16286);
and U16489 (N_16489,N_16259,N_16257);
or U16490 (N_16490,N_16224,N_16317);
nor U16491 (N_16491,N_16282,N_16364);
or U16492 (N_16492,N_16341,N_16329);
nand U16493 (N_16493,N_16369,N_16380);
and U16494 (N_16494,N_16339,N_16274);
nor U16495 (N_16495,N_16313,N_16393);
nand U16496 (N_16496,N_16216,N_16267);
nor U16497 (N_16497,N_16396,N_16255);
or U16498 (N_16498,N_16240,N_16327);
or U16499 (N_16499,N_16344,N_16223);
nand U16500 (N_16500,N_16295,N_16369);
nand U16501 (N_16501,N_16289,N_16258);
nor U16502 (N_16502,N_16380,N_16255);
nand U16503 (N_16503,N_16378,N_16272);
nand U16504 (N_16504,N_16334,N_16372);
and U16505 (N_16505,N_16259,N_16390);
nand U16506 (N_16506,N_16335,N_16213);
nand U16507 (N_16507,N_16378,N_16245);
and U16508 (N_16508,N_16243,N_16311);
nand U16509 (N_16509,N_16383,N_16251);
nand U16510 (N_16510,N_16381,N_16234);
nand U16511 (N_16511,N_16390,N_16377);
and U16512 (N_16512,N_16242,N_16371);
nand U16513 (N_16513,N_16260,N_16303);
xor U16514 (N_16514,N_16346,N_16284);
and U16515 (N_16515,N_16386,N_16226);
or U16516 (N_16516,N_16339,N_16368);
or U16517 (N_16517,N_16334,N_16257);
and U16518 (N_16518,N_16340,N_16262);
or U16519 (N_16519,N_16310,N_16257);
nand U16520 (N_16520,N_16301,N_16352);
and U16521 (N_16521,N_16212,N_16224);
or U16522 (N_16522,N_16207,N_16310);
or U16523 (N_16523,N_16378,N_16319);
nor U16524 (N_16524,N_16204,N_16357);
and U16525 (N_16525,N_16211,N_16258);
and U16526 (N_16526,N_16267,N_16305);
nand U16527 (N_16527,N_16295,N_16354);
nand U16528 (N_16528,N_16256,N_16327);
and U16529 (N_16529,N_16301,N_16330);
or U16530 (N_16530,N_16262,N_16302);
nor U16531 (N_16531,N_16343,N_16270);
and U16532 (N_16532,N_16219,N_16354);
nand U16533 (N_16533,N_16394,N_16230);
nand U16534 (N_16534,N_16262,N_16291);
nor U16535 (N_16535,N_16284,N_16291);
nand U16536 (N_16536,N_16392,N_16297);
and U16537 (N_16537,N_16326,N_16361);
or U16538 (N_16538,N_16310,N_16201);
or U16539 (N_16539,N_16327,N_16241);
nand U16540 (N_16540,N_16318,N_16376);
or U16541 (N_16541,N_16279,N_16264);
xor U16542 (N_16542,N_16305,N_16284);
xor U16543 (N_16543,N_16386,N_16367);
and U16544 (N_16544,N_16311,N_16301);
nand U16545 (N_16545,N_16349,N_16214);
or U16546 (N_16546,N_16256,N_16235);
nand U16547 (N_16547,N_16211,N_16374);
and U16548 (N_16548,N_16260,N_16254);
nor U16549 (N_16549,N_16290,N_16213);
or U16550 (N_16550,N_16281,N_16362);
or U16551 (N_16551,N_16247,N_16232);
xnor U16552 (N_16552,N_16226,N_16313);
nand U16553 (N_16553,N_16300,N_16346);
and U16554 (N_16554,N_16227,N_16284);
nand U16555 (N_16555,N_16313,N_16334);
xnor U16556 (N_16556,N_16377,N_16354);
nor U16557 (N_16557,N_16289,N_16228);
or U16558 (N_16558,N_16356,N_16374);
nor U16559 (N_16559,N_16290,N_16279);
or U16560 (N_16560,N_16376,N_16372);
and U16561 (N_16561,N_16385,N_16218);
xnor U16562 (N_16562,N_16249,N_16363);
nor U16563 (N_16563,N_16337,N_16293);
nand U16564 (N_16564,N_16390,N_16262);
nor U16565 (N_16565,N_16288,N_16373);
and U16566 (N_16566,N_16357,N_16318);
xnor U16567 (N_16567,N_16210,N_16346);
xnor U16568 (N_16568,N_16382,N_16356);
and U16569 (N_16569,N_16208,N_16260);
xnor U16570 (N_16570,N_16223,N_16245);
nor U16571 (N_16571,N_16363,N_16254);
and U16572 (N_16572,N_16385,N_16233);
nor U16573 (N_16573,N_16299,N_16245);
nand U16574 (N_16574,N_16363,N_16293);
nand U16575 (N_16575,N_16224,N_16259);
or U16576 (N_16576,N_16368,N_16371);
nor U16577 (N_16577,N_16221,N_16364);
or U16578 (N_16578,N_16317,N_16250);
or U16579 (N_16579,N_16335,N_16302);
nand U16580 (N_16580,N_16264,N_16252);
xor U16581 (N_16581,N_16360,N_16394);
xnor U16582 (N_16582,N_16341,N_16272);
nor U16583 (N_16583,N_16311,N_16383);
or U16584 (N_16584,N_16252,N_16295);
nor U16585 (N_16585,N_16305,N_16344);
nor U16586 (N_16586,N_16329,N_16380);
nor U16587 (N_16587,N_16210,N_16388);
xnor U16588 (N_16588,N_16299,N_16313);
nand U16589 (N_16589,N_16360,N_16263);
xor U16590 (N_16590,N_16289,N_16246);
xor U16591 (N_16591,N_16332,N_16316);
or U16592 (N_16592,N_16201,N_16337);
nor U16593 (N_16593,N_16273,N_16292);
or U16594 (N_16594,N_16237,N_16280);
and U16595 (N_16595,N_16221,N_16273);
nor U16596 (N_16596,N_16291,N_16314);
or U16597 (N_16597,N_16362,N_16229);
xor U16598 (N_16598,N_16338,N_16228);
or U16599 (N_16599,N_16214,N_16396);
and U16600 (N_16600,N_16478,N_16577);
or U16601 (N_16601,N_16513,N_16526);
nor U16602 (N_16602,N_16580,N_16542);
xor U16603 (N_16603,N_16483,N_16406);
xnor U16604 (N_16604,N_16466,N_16461);
nand U16605 (N_16605,N_16424,N_16597);
xor U16606 (N_16606,N_16418,N_16594);
nand U16607 (N_16607,N_16498,N_16431);
nand U16608 (N_16608,N_16447,N_16491);
nor U16609 (N_16609,N_16423,N_16419);
or U16610 (N_16610,N_16598,N_16433);
or U16611 (N_16611,N_16490,N_16479);
and U16612 (N_16612,N_16581,N_16541);
or U16613 (N_16613,N_16485,N_16409);
nand U16614 (N_16614,N_16400,N_16477);
or U16615 (N_16615,N_16476,N_16494);
nor U16616 (N_16616,N_16480,N_16517);
or U16617 (N_16617,N_16556,N_16426);
xnor U16618 (N_16618,N_16511,N_16422);
and U16619 (N_16619,N_16475,N_16536);
xor U16620 (N_16620,N_16495,N_16559);
nand U16621 (N_16621,N_16481,N_16507);
nand U16622 (N_16622,N_16572,N_16545);
xor U16623 (N_16623,N_16544,N_16555);
and U16624 (N_16624,N_16503,N_16413);
or U16625 (N_16625,N_16401,N_16548);
nor U16626 (N_16626,N_16502,N_16560);
nand U16627 (N_16627,N_16529,N_16489);
xor U16628 (N_16628,N_16435,N_16448);
and U16629 (N_16629,N_16404,N_16589);
nor U16630 (N_16630,N_16434,N_16512);
xnor U16631 (N_16631,N_16411,N_16557);
nor U16632 (N_16632,N_16488,N_16452);
or U16633 (N_16633,N_16430,N_16415);
xnor U16634 (N_16634,N_16579,N_16445);
nor U16635 (N_16635,N_16510,N_16595);
xnor U16636 (N_16636,N_16403,N_16407);
or U16637 (N_16637,N_16438,N_16468);
xnor U16638 (N_16638,N_16463,N_16543);
xor U16639 (N_16639,N_16591,N_16514);
nand U16640 (N_16640,N_16496,N_16547);
nor U16641 (N_16641,N_16564,N_16428);
or U16642 (N_16642,N_16539,N_16429);
and U16643 (N_16643,N_16522,N_16528);
or U16644 (N_16644,N_16569,N_16470);
nand U16645 (N_16645,N_16501,N_16492);
or U16646 (N_16646,N_16432,N_16455);
or U16647 (N_16647,N_16558,N_16596);
nor U16648 (N_16648,N_16469,N_16504);
xor U16649 (N_16649,N_16568,N_16530);
nand U16650 (N_16650,N_16578,N_16527);
nor U16651 (N_16651,N_16437,N_16486);
nor U16652 (N_16652,N_16487,N_16570);
and U16653 (N_16653,N_16484,N_16416);
nand U16654 (N_16654,N_16472,N_16464);
nand U16655 (N_16655,N_16450,N_16521);
nand U16656 (N_16656,N_16549,N_16592);
nand U16657 (N_16657,N_16574,N_16458);
xor U16658 (N_16658,N_16590,N_16533);
nor U16659 (N_16659,N_16537,N_16583);
xnor U16660 (N_16660,N_16509,N_16540);
or U16661 (N_16661,N_16499,N_16414);
nand U16662 (N_16662,N_16523,N_16566);
nand U16663 (N_16663,N_16421,N_16473);
or U16664 (N_16664,N_16420,N_16563);
nor U16665 (N_16665,N_16553,N_16567);
and U16666 (N_16666,N_16515,N_16439);
and U16667 (N_16667,N_16457,N_16471);
xnor U16668 (N_16668,N_16554,N_16436);
or U16669 (N_16669,N_16459,N_16442);
and U16670 (N_16670,N_16525,N_16465);
and U16671 (N_16671,N_16546,N_16482);
and U16672 (N_16672,N_16449,N_16518);
xor U16673 (N_16673,N_16582,N_16467);
nor U16674 (N_16674,N_16535,N_16451);
and U16675 (N_16675,N_16454,N_16599);
and U16676 (N_16676,N_16506,N_16508);
xnor U16677 (N_16677,N_16408,N_16500);
xnor U16678 (N_16678,N_16456,N_16516);
nand U16679 (N_16679,N_16425,N_16441);
and U16680 (N_16680,N_16462,N_16588);
or U16681 (N_16681,N_16524,N_16565);
or U16682 (N_16682,N_16443,N_16575);
xnor U16683 (N_16683,N_16497,N_16531);
nand U16684 (N_16684,N_16440,N_16534);
and U16685 (N_16685,N_16584,N_16446);
or U16686 (N_16686,N_16460,N_16538);
and U16687 (N_16687,N_16562,N_16520);
or U16688 (N_16688,N_16576,N_16505);
and U16689 (N_16689,N_16417,N_16552);
or U16690 (N_16690,N_16561,N_16550);
and U16691 (N_16691,N_16474,N_16586);
and U16692 (N_16692,N_16402,N_16571);
or U16693 (N_16693,N_16532,N_16493);
and U16694 (N_16694,N_16405,N_16585);
nor U16695 (N_16695,N_16412,N_16593);
and U16696 (N_16696,N_16573,N_16427);
nand U16697 (N_16697,N_16551,N_16410);
nor U16698 (N_16698,N_16453,N_16519);
nor U16699 (N_16699,N_16444,N_16587);
xor U16700 (N_16700,N_16521,N_16574);
nor U16701 (N_16701,N_16435,N_16468);
nand U16702 (N_16702,N_16469,N_16421);
or U16703 (N_16703,N_16471,N_16482);
nand U16704 (N_16704,N_16402,N_16446);
nor U16705 (N_16705,N_16421,N_16575);
xnor U16706 (N_16706,N_16431,N_16568);
or U16707 (N_16707,N_16490,N_16417);
or U16708 (N_16708,N_16514,N_16413);
nand U16709 (N_16709,N_16489,N_16457);
nor U16710 (N_16710,N_16413,N_16477);
xor U16711 (N_16711,N_16536,N_16474);
nand U16712 (N_16712,N_16566,N_16414);
nor U16713 (N_16713,N_16541,N_16413);
xnor U16714 (N_16714,N_16478,N_16507);
nor U16715 (N_16715,N_16458,N_16571);
or U16716 (N_16716,N_16535,N_16596);
and U16717 (N_16717,N_16421,N_16437);
and U16718 (N_16718,N_16497,N_16597);
or U16719 (N_16719,N_16580,N_16450);
or U16720 (N_16720,N_16558,N_16465);
and U16721 (N_16721,N_16528,N_16412);
nand U16722 (N_16722,N_16551,N_16566);
nor U16723 (N_16723,N_16458,N_16423);
or U16724 (N_16724,N_16589,N_16474);
nor U16725 (N_16725,N_16435,N_16419);
or U16726 (N_16726,N_16546,N_16583);
nor U16727 (N_16727,N_16512,N_16580);
nand U16728 (N_16728,N_16501,N_16565);
or U16729 (N_16729,N_16430,N_16404);
xnor U16730 (N_16730,N_16575,N_16403);
or U16731 (N_16731,N_16591,N_16547);
or U16732 (N_16732,N_16468,N_16462);
or U16733 (N_16733,N_16421,N_16484);
xor U16734 (N_16734,N_16551,N_16506);
nor U16735 (N_16735,N_16599,N_16490);
xnor U16736 (N_16736,N_16575,N_16504);
nor U16737 (N_16737,N_16451,N_16575);
nor U16738 (N_16738,N_16539,N_16439);
and U16739 (N_16739,N_16410,N_16443);
nor U16740 (N_16740,N_16428,N_16527);
xnor U16741 (N_16741,N_16525,N_16587);
nand U16742 (N_16742,N_16565,N_16580);
and U16743 (N_16743,N_16535,N_16586);
and U16744 (N_16744,N_16424,N_16521);
xor U16745 (N_16745,N_16533,N_16501);
and U16746 (N_16746,N_16574,N_16597);
nand U16747 (N_16747,N_16551,N_16464);
nand U16748 (N_16748,N_16478,N_16504);
xor U16749 (N_16749,N_16448,N_16544);
nor U16750 (N_16750,N_16450,N_16467);
and U16751 (N_16751,N_16583,N_16460);
or U16752 (N_16752,N_16413,N_16488);
nand U16753 (N_16753,N_16430,N_16439);
nor U16754 (N_16754,N_16454,N_16580);
nand U16755 (N_16755,N_16548,N_16547);
nand U16756 (N_16756,N_16584,N_16504);
nor U16757 (N_16757,N_16412,N_16516);
nand U16758 (N_16758,N_16400,N_16480);
nand U16759 (N_16759,N_16597,N_16410);
nor U16760 (N_16760,N_16467,N_16549);
nand U16761 (N_16761,N_16407,N_16415);
and U16762 (N_16762,N_16425,N_16586);
nand U16763 (N_16763,N_16499,N_16513);
nand U16764 (N_16764,N_16581,N_16530);
or U16765 (N_16765,N_16455,N_16470);
xor U16766 (N_16766,N_16581,N_16594);
nor U16767 (N_16767,N_16550,N_16493);
xnor U16768 (N_16768,N_16598,N_16465);
or U16769 (N_16769,N_16526,N_16459);
or U16770 (N_16770,N_16506,N_16464);
xor U16771 (N_16771,N_16439,N_16516);
nand U16772 (N_16772,N_16520,N_16543);
nor U16773 (N_16773,N_16537,N_16491);
xnor U16774 (N_16774,N_16472,N_16585);
nor U16775 (N_16775,N_16596,N_16488);
nand U16776 (N_16776,N_16463,N_16437);
or U16777 (N_16777,N_16591,N_16550);
nand U16778 (N_16778,N_16584,N_16437);
or U16779 (N_16779,N_16436,N_16599);
or U16780 (N_16780,N_16492,N_16430);
nand U16781 (N_16781,N_16573,N_16568);
nor U16782 (N_16782,N_16415,N_16514);
nor U16783 (N_16783,N_16447,N_16558);
xnor U16784 (N_16784,N_16511,N_16448);
or U16785 (N_16785,N_16559,N_16570);
nor U16786 (N_16786,N_16447,N_16427);
xnor U16787 (N_16787,N_16437,N_16408);
xor U16788 (N_16788,N_16526,N_16582);
nor U16789 (N_16789,N_16406,N_16535);
nor U16790 (N_16790,N_16580,N_16413);
xnor U16791 (N_16791,N_16599,N_16595);
nand U16792 (N_16792,N_16484,N_16504);
and U16793 (N_16793,N_16467,N_16589);
xnor U16794 (N_16794,N_16554,N_16423);
nor U16795 (N_16795,N_16463,N_16545);
xnor U16796 (N_16796,N_16481,N_16506);
xor U16797 (N_16797,N_16588,N_16520);
and U16798 (N_16798,N_16599,N_16404);
xnor U16799 (N_16799,N_16453,N_16460);
nor U16800 (N_16800,N_16601,N_16721);
nor U16801 (N_16801,N_16697,N_16618);
and U16802 (N_16802,N_16735,N_16726);
and U16803 (N_16803,N_16645,N_16611);
or U16804 (N_16804,N_16699,N_16649);
and U16805 (N_16805,N_16711,N_16724);
xnor U16806 (N_16806,N_16745,N_16623);
nand U16807 (N_16807,N_16755,N_16604);
and U16808 (N_16808,N_16660,N_16790);
xnor U16809 (N_16809,N_16788,N_16610);
or U16810 (N_16810,N_16748,N_16658);
or U16811 (N_16811,N_16680,N_16736);
nand U16812 (N_16812,N_16603,N_16779);
nand U16813 (N_16813,N_16780,N_16741);
nand U16814 (N_16814,N_16714,N_16716);
nand U16815 (N_16815,N_16657,N_16638);
nor U16816 (N_16816,N_16695,N_16734);
nor U16817 (N_16817,N_16605,N_16616);
nor U16818 (N_16818,N_16754,N_16706);
nand U16819 (N_16819,N_16769,N_16630);
or U16820 (N_16820,N_16725,N_16722);
xnor U16821 (N_16821,N_16772,N_16646);
nand U16822 (N_16822,N_16635,N_16617);
nand U16823 (N_16823,N_16723,N_16758);
nor U16824 (N_16824,N_16654,N_16793);
nand U16825 (N_16825,N_16784,N_16651);
xor U16826 (N_16826,N_16691,N_16621);
or U16827 (N_16827,N_16740,N_16674);
and U16828 (N_16828,N_16707,N_16761);
nand U16829 (N_16829,N_16684,N_16762);
nand U16830 (N_16830,N_16719,N_16781);
and U16831 (N_16831,N_16693,N_16760);
nor U16832 (N_16832,N_16648,N_16631);
nor U16833 (N_16833,N_16694,N_16710);
or U16834 (N_16834,N_16770,N_16666);
or U16835 (N_16835,N_16732,N_16730);
nand U16836 (N_16836,N_16692,N_16668);
or U16837 (N_16837,N_16620,N_16681);
and U16838 (N_16838,N_16763,N_16641);
xor U16839 (N_16839,N_16600,N_16700);
or U16840 (N_16840,N_16633,N_16765);
and U16841 (N_16841,N_16798,N_16747);
xor U16842 (N_16842,N_16773,N_16731);
nor U16843 (N_16843,N_16625,N_16717);
nand U16844 (N_16844,N_16789,N_16642);
or U16845 (N_16845,N_16613,N_16656);
and U16846 (N_16846,N_16652,N_16653);
nor U16847 (N_16847,N_16644,N_16713);
or U16848 (N_16848,N_16753,N_16622);
nor U16849 (N_16849,N_16799,N_16796);
xor U16850 (N_16850,N_16709,N_16786);
nor U16851 (N_16851,N_16795,N_16671);
or U16852 (N_16852,N_16702,N_16775);
xnor U16853 (N_16853,N_16669,N_16640);
nor U16854 (N_16854,N_16672,N_16759);
xnor U16855 (N_16855,N_16703,N_16643);
or U16856 (N_16856,N_16767,N_16701);
xnor U16857 (N_16857,N_16637,N_16757);
nand U16858 (N_16858,N_16737,N_16619);
nand U16859 (N_16859,N_16670,N_16708);
nand U16860 (N_16860,N_16739,N_16746);
nand U16861 (N_16861,N_16696,N_16688);
nor U16862 (N_16862,N_16698,N_16627);
and U16863 (N_16863,N_16690,N_16744);
or U16864 (N_16864,N_16686,N_16752);
xor U16865 (N_16865,N_16794,N_16776);
or U16866 (N_16866,N_16639,N_16792);
xnor U16867 (N_16867,N_16607,N_16771);
and U16868 (N_16868,N_16787,N_16727);
and U16869 (N_16869,N_16797,N_16715);
or U16870 (N_16870,N_16636,N_16689);
xor U16871 (N_16871,N_16704,N_16738);
or U16872 (N_16872,N_16661,N_16629);
nand U16873 (N_16873,N_16682,N_16705);
nand U16874 (N_16874,N_16777,N_16663);
nand U16875 (N_16875,N_16687,N_16606);
xnor U16876 (N_16876,N_16733,N_16764);
and U16877 (N_16877,N_16609,N_16679);
nand U16878 (N_16878,N_16712,N_16756);
and U16879 (N_16879,N_16659,N_16783);
nand U16880 (N_16880,N_16628,N_16685);
nand U16881 (N_16881,N_16614,N_16634);
nand U16882 (N_16882,N_16675,N_16632);
xnor U16883 (N_16883,N_16673,N_16662);
and U16884 (N_16884,N_16785,N_16650);
nand U16885 (N_16885,N_16626,N_16729);
or U16886 (N_16886,N_16743,N_16615);
xnor U16887 (N_16887,N_16624,N_16749);
or U16888 (N_16888,N_16751,N_16728);
nand U16889 (N_16889,N_16678,N_16647);
xnor U16890 (N_16890,N_16665,N_16664);
nor U16891 (N_16891,N_16677,N_16655);
nand U16892 (N_16892,N_16791,N_16667);
xor U16893 (N_16893,N_16612,N_16602);
nand U16894 (N_16894,N_16718,N_16774);
xor U16895 (N_16895,N_16782,N_16768);
and U16896 (N_16896,N_16742,N_16720);
nor U16897 (N_16897,N_16608,N_16766);
xnor U16898 (N_16898,N_16750,N_16683);
or U16899 (N_16899,N_16676,N_16778);
nand U16900 (N_16900,N_16779,N_16778);
nand U16901 (N_16901,N_16709,N_16703);
nor U16902 (N_16902,N_16755,N_16652);
or U16903 (N_16903,N_16778,N_16647);
xnor U16904 (N_16904,N_16750,N_16660);
and U16905 (N_16905,N_16720,N_16624);
nand U16906 (N_16906,N_16710,N_16622);
and U16907 (N_16907,N_16663,N_16684);
and U16908 (N_16908,N_16677,N_16720);
nor U16909 (N_16909,N_16666,N_16700);
nor U16910 (N_16910,N_16620,N_16747);
nand U16911 (N_16911,N_16618,N_16726);
and U16912 (N_16912,N_16642,N_16748);
nor U16913 (N_16913,N_16778,N_16738);
and U16914 (N_16914,N_16701,N_16675);
or U16915 (N_16915,N_16793,N_16614);
xnor U16916 (N_16916,N_16700,N_16605);
or U16917 (N_16917,N_16732,N_16717);
nor U16918 (N_16918,N_16747,N_16748);
and U16919 (N_16919,N_16778,N_16796);
xnor U16920 (N_16920,N_16709,N_16683);
nor U16921 (N_16921,N_16769,N_16727);
xor U16922 (N_16922,N_16758,N_16673);
nand U16923 (N_16923,N_16671,N_16672);
and U16924 (N_16924,N_16609,N_16628);
nor U16925 (N_16925,N_16685,N_16797);
or U16926 (N_16926,N_16765,N_16731);
and U16927 (N_16927,N_16759,N_16702);
nor U16928 (N_16928,N_16648,N_16653);
and U16929 (N_16929,N_16743,N_16769);
nor U16930 (N_16930,N_16733,N_16620);
and U16931 (N_16931,N_16623,N_16715);
xor U16932 (N_16932,N_16646,N_16660);
xnor U16933 (N_16933,N_16697,N_16703);
xor U16934 (N_16934,N_16757,N_16656);
or U16935 (N_16935,N_16735,N_16798);
and U16936 (N_16936,N_16731,N_16716);
and U16937 (N_16937,N_16684,N_16727);
nor U16938 (N_16938,N_16635,N_16601);
nand U16939 (N_16939,N_16798,N_16746);
nand U16940 (N_16940,N_16728,N_16623);
or U16941 (N_16941,N_16661,N_16612);
or U16942 (N_16942,N_16726,N_16622);
and U16943 (N_16943,N_16764,N_16667);
nand U16944 (N_16944,N_16641,N_16720);
or U16945 (N_16945,N_16671,N_16691);
and U16946 (N_16946,N_16635,N_16704);
and U16947 (N_16947,N_16675,N_16745);
nor U16948 (N_16948,N_16699,N_16601);
and U16949 (N_16949,N_16617,N_16620);
nand U16950 (N_16950,N_16754,N_16625);
nor U16951 (N_16951,N_16779,N_16784);
xor U16952 (N_16952,N_16646,N_16709);
and U16953 (N_16953,N_16631,N_16632);
xor U16954 (N_16954,N_16655,N_16676);
nand U16955 (N_16955,N_16772,N_16628);
and U16956 (N_16956,N_16624,N_16694);
xnor U16957 (N_16957,N_16757,N_16720);
xor U16958 (N_16958,N_16701,N_16743);
nor U16959 (N_16959,N_16744,N_16634);
and U16960 (N_16960,N_16632,N_16759);
xor U16961 (N_16961,N_16718,N_16658);
or U16962 (N_16962,N_16675,N_16780);
nor U16963 (N_16963,N_16778,N_16737);
nand U16964 (N_16964,N_16716,N_16627);
nand U16965 (N_16965,N_16735,N_16660);
nor U16966 (N_16966,N_16716,N_16774);
nand U16967 (N_16967,N_16705,N_16737);
nand U16968 (N_16968,N_16712,N_16722);
or U16969 (N_16969,N_16647,N_16615);
xnor U16970 (N_16970,N_16672,N_16775);
nor U16971 (N_16971,N_16655,N_16612);
nor U16972 (N_16972,N_16712,N_16627);
nand U16973 (N_16973,N_16676,N_16670);
or U16974 (N_16974,N_16688,N_16715);
or U16975 (N_16975,N_16637,N_16705);
nor U16976 (N_16976,N_16742,N_16640);
xor U16977 (N_16977,N_16751,N_16635);
nor U16978 (N_16978,N_16722,N_16760);
or U16979 (N_16979,N_16784,N_16786);
nor U16980 (N_16980,N_16728,N_16650);
or U16981 (N_16981,N_16789,N_16719);
and U16982 (N_16982,N_16721,N_16619);
xor U16983 (N_16983,N_16651,N_16703);
nand U16984 (N_16984,N_16643,N_16688);
nor U16985 (N_16985,N_16758,N_16791);
nor U16986 (N_16986,N_16634,N_16605);
xnor U16987 (N_16987,N_16793,N_16679);
nor U16988 (N_16988,N_16740,N_16645);
or U16989 (N_16989,N_16679,N_16610);
nand U16990 (N_16990,N_16642,N_16612);
and U16991 (N_16991,N_16741,N_16616);
or U16992 (N_16992,N_16689,N_16746);
nor U16993 (N_16993,N_16677,N_16650);
nand U16994 (N_16994,N_16647,N_16698);
xnor U16995 (N_16995,N_16675,N_16609);
or U16996 (N_16996,N_16714,N_16664);
xor U16997 (N_16997,N_16729,N_16737);
and U16998 (N_16998,N_16616,N_16658);
nor U16999 (N_16999,N_16703,N_16616);
xor U17000 (N_17000,N_16825,N_16938);
nor U17001 (N_17001,N_16816,N_16937);
nand U17002 (N_17002,N_16855,N_16891);
nand U17003 (N_17003,N_16849,N_16908);
xor U17004 (N_17004,N_16857,N_16967);
or U17005 (N_17005,N_16874,N_16911);
nand U17006 (N_17006,N_16821,N_16966);
and U17007 (N_17007,N_16905,N_16927);
and U17008 (N_17008,N_16899,N_16934);
nand U17009 (N_17009,N_16805,N_16812);
nor U17010 (N_17010,N_16854,N_16929);
or U17011 (N_17011,N_16896,N_16815);
or U17012 (N_17012,N_16830,N_16974);
nor U17013 (N_17013,N_16890,N_16933);
and U17014 (N_17014,N_16986,N_16979);
and U17015 (N_17015,N_16800,N_16892);
nor U17016 (N_17016,N_16922,N_16840);
or U17017 (N_17017,N_16829,N_16838);
and U17018 (N_17018,N_16992,N_16880);
xor U17019 (N_17019,N_16846,N_16950);
and U17020 (N_17020,N_16965,N_16914);
and U17021 (N_17021,N_16820,N_16921);
or U17022 (N_17022,N_16902,N_16942);
nand U17023 (N_17023,N_16810,N_16961);
or U17024 (N_17024,N_16894,N_16962);
nand U17025 (N_17025,N_16822,N_16856);
and U17026 (N_17026,N_16888,N_16877);
or U17027 (N_17027,N_16991,N_16819);
or U17028 (N_17028,N_16923,N_16818);
nand U17029 (N_17029,N_16828,N_16955);
nor U17030 (N_17030,N_16906,N_16808);
and U17031 (N_17031,N_16803,N_16882);
and U17032 (N_17032,N_16952,N_16975);
nand U17033 (N_17033,N_16883,N_16873);
and U17034 (N_17034,N_16907,N_16946);
xor U17035 (N_17035,N_16866,N_16999);
or U17036 (N_17036,N_16884,N_16935);
xor U17037 (N_17037,N_16813,N_16931);
or U17038 (N_17038,N_16862,N_16972);
xor U17039 (N_17039,N_16842,N_16903);
nor U17040 (N_17040,N_16878,N_16977);
or U17041 (N_17041,N_16912,N_16981);
and U17042 (N_17042,N_16928,N_16951);
xnor U17043 (N_17043,N_16924,N_16898);
nor U17044 (N_17044,N_16918,N_16801);
and U17045 (N_17045,N_16904,N_16851);
xor U17046 (N_17046,N_16845,N_16833);
xnor U17047 (N_17047,N_16947,N_16958);
xnor U17048 (N_17048,N_16989,N_16945);
xor U17049 (N_17049,N_16811,N_16985);
xor U17050 (N_17050,N_16853,N_16968);
or U17051 (N_17051,N_16936,N_16917);
nor U17052 (N_17052,N_16893,N_16996);
xor U17053 (N_17053,N_16876,N_16848);
nor U17054 (N_17054,N_16881,N_16836);
nor U17055 (N_17055,N_16847,N_16839);
and U17056 (N_17056,N_16832,N_16831);
and U17057 (N_17057,N_16994,N_16943);
and U17058 (N_17058,N_16982,N_16983);
nor U17059 (N_17059,N_16807,N_16915);
or U17060 (N_17060,N_16949,N_16806);
and U17061 (N_17061,N_16867,N_16824);
xor U17062 (N_17062,N_16944,N_16932);
or U17063 (N_17063,N_16858,N_16823);
or U17064 (N_17064,N_16930,N_16963);
or U17065 (N_17065,N_16871,N_16919);
xor U17066 (N_17066,N_16987,N_16885);
nand U17067 (N_17067,N_16901,N_16997);
nand U17068 (N_17068,N_16814,N_16802);
and U17069 (N_17069,N_16872,N_16971);
and U17070 (N_17070,N_16865,N_16850);
nand U17071 (N_17071,N_16889,N_16954);
and U17072 (N_17072,N_16868,N_16969);
or U17073 (N_17073,N_16844,N_16956);
xnor U17074 (N_17074,N_16817,N_16940);
nand U17075 (N_17075,N_16995,N_16948);
or U17076 (N_17076,N_16861,N_16870);
nor U17077 (N_17077,N_16988,N_16864);
nand U17078 (N_17078,N_16869,N_16837);
or U17079 (N_17079,N_16964,N_16976);
nor U17080 (N_17080,N_16852,N_16916);
nand U17081 (N_17081,N_16993,N_16875);
xnor U17082 (N_17082,N_16897,N_16860);
and U17083 (N_17083,N_16957,N_16895);
nand U17084 (N_17084,N_16804,N_16960);
or U17085 (N_17085,N_16990,N_16998);
or U17086 (N_17086,N_16886,N_16859);
and U17087 (N_17087,N_16926,N_16909);
xor U17088 (N_17088,N_16863,N_16843);
nor U17089 (N_17089,N_16959,N_16939);
nor U17090 (N_17090,N_16910,N_16970);
or U17091 (N_17091,N_16973,N_16834);
nor U17092 (N_17092,N_16920,N_16925);
nand U17093 (N_17093,N_16980,N_16984);
and U17094 (N_17094,N_16913,N_16809);
nand U17095 (N_17095,N_16827,N_16900);
nand U17096 (N_17096,N_16953,N_16835);
nand U17097 (N_17097,N_16879,N_16841);
and U17098 (N_17098,N_16941,N_16978);
xnor U17099 (N_17099,N_16887,N_16826);
and U17100 (N_17100,N_16971,N_16837);
xnor U17101 (N_17101,N_16970,N_16824);
xnor U17102 (N_17102,N_16944,N_16868);
or U17103 (N_17103,N_16823,N_16908);
or U17104 (N_17104,N_16947,N_16830);
nor U17105 (N_17105,N_16809,N_16990);
nand U17106 (N_17106,N_16956,N_16837);
xnor U17107 (N_17107,N_16987,N_16810);
or U17108 (N_17108,N_16856,N_16848);
or U17109 (N_17109,N_16941,N_16896);
nand U17110 (N_17110,N_16837,N_16975);
nor U17111 (N_17111,N_16804,N_16997);
or U17112 (N_17112,N_16957,N_16879);
xnor U17113 (N_17113,N_16855,N_16953);
xor U17114 (N_17114,N_16902,N_16997);
or U17115 (N_17115,N_16948,N_16964);
and U17116 (N_17116,N_16987,N_16979);
xor U17117 (N_17117,N_16912,N_16911);
xor U17118 (N_17118,N_16903,N_16885);
nand U17119 (N_17119,N_16954,N_16890);
nand U17120 (N_17120,N_16883,N_16906);
nor U17121 (N_17121,N_16877,N_16946);
nor U17122 (N_17122,N_16829,N_16936);
nor U17123 (N_17123,N_16810,N_16923);
xor U17124 (N_17124,N_16902,N_16929);
xnor U17125 (N_17125,N_16887,N_16811);
nor U17126 (N_17126,N_16961,N_16935);
and U17127 (N_17127,N_16853,N_16987);
nor U17128 (N_17128,N_16884,N_16843);
and U17129 (N_17129,N_16873,N_16849);
or U17130 (N_17130,N_16925,N_16915);
nand U17131 (N_17131,N_16860,N_16842);
or U17132 (N_17132,N_16821,N_16977);
and U17133 (N_17133,N_16842,N_16947);
nand U17134 (N_17134,N_16849,N_16927);
xnor U17135 (N_17135,N_16893,N_16960);
nand U17136 (N_17136,N_16802,N_16870);
nand U17137 (N_17137,N_16880,N_16819);
nand U17138 (N_17138,N_16894,N_16801);
nand U17139 (N_17139,N_16825,N_16915);
nand U17140 (N_17140,N_16860,N_16969);
and U17141 (N_17141,N_16830,N_16850);
xnor U17142 (N_17142,N_16972,N_16831);
xor U17143 (N_17143,N_16897,N_16911);
nand U17144 (N_17144,N_16876,N_16924);
and U17145 (N_17145,N_16837,N_16808);
nand U17146 (N_17146,N_16803,N_16835);
or U17147 (N_17147,N_16835,N_16831);
nor U17148 (N_17148,N_16880,N_16812);
xor U17149 (N_17149,N_16993,N_16915);
nand U17150 (N_17150,N_16941,N_16851);
nand U17151 (N_17151,N_16893,N_16856);
nor U17152 (N_17152,N_16980,N_16896);
nor U17153 (N_17153,N_16998,N_16879);
nor U17154 (N_17154,N_16842,N_16898);
or U17155 (N_17155,N_16974,N_16872);
nand U17156 (N_17156,N_16994,N_16909);
nand U17157 (N_17157,N_16981,N_16927);
nand U17158 (N_17158,N_16939,N_16804);
and U17159 (N_17159,N_16824,N_16877);
and U17160 (N_17160,N_16979,N_16981);
nand U17161 (N_17161,N_16855,N_16839);
nor U17162 (N_17162,N_16977,N_16967);
or U17163 (N_17163,N_16959,N_16980);
xnor U17164 (N_17164,N_16914,N_16879);
or U17165 (N_17165,N_16992,N_16903);
nor U17166 (N_17166,N_16868,N_16804);
nor U17167 (N_17167,N_16918,N_16886);
and U17168 (N_17168,N_16866,N_16801);
xor U17169 (N_17169,N_16852,N_16893);
nor U17170 (N_17170,N_16881,N_16929);
and U17171 (N_17171,N_16970,N_16832);
xnor U17172 (N_17172,N_16904,N_16804);
xor U17173 (N_17173,N_16883,N_16991);
nand U17174 (N_17174,N_16811,N_16938);
nor U17175 (N_17175,N_16860,N_16818);
nand U17176 (N_17176,N_16966,N_16911);
and U17177 (N_17177,N_16977,N_16997);
or U17178 (N_17178,N_16876,N_16861);
xor U17179 (N_17179,N_16849,N_16983);
nand U17180 (N_17180,N_16863,N_16935);
nor U17181 (N_17181,N_16978,N_16874);
nor U17182 (N_17182,N_16965,N_16850);
xnor U17183 (N_17183,N_16916,N_16970);
or U17184 (N_17184,N_16945,N_16805);
nand U17185 (N_17185,N_16822,N_16868);
xnor U17186 (N_17186,N_16986,N_16870);
or U17187 (N_17187,N_16900,N_16925);
and U17188 (N_17188,N_16958,N_16860);
and U17189 (N_17189,N_16978,N_16994);
nor U17190 (N_17190,N_16924,N_16930);
nor U17191 (N_17191,N_16840,N_16868);
nand U17192 (N_17192,N_16885,N_16965);
and U17193 (N_17193,N_16938,N_16943);
and U17194 (N_17194,N_16846,N_16971);
or U17195 (N_17195,N_16960,N_16983);
nor U17196 (N_17196,N_16978,N_16923);
nand U17197 (N_17197,N_16927,N_16989);
xnor U17198 (N_17198,N_16871,N_16867);
nor U17199 (N_17199,N_16996,N_16888);
and U17200 (N_17200,N_17097,N_17083);
and U17201 (N_17201,N_17183,N_17085);
nor U17202 (N_17202,N_17038,N_17118);
nand U17203 (N_17203,N_17071,N_17190);
xnor U17204 (N_17204,N_17060,N_17141);
nor U17205 (N_17205,N_17195,N_17105);
and U17206 (N_17206,N_17077,N_17111);
and U17207 (N_17207,N_17027,N_17155);
or U17208 (N_17208,N_17128,N_17002);
nor U17209 (N_17209,N_17015,N_17169);
and U17210 (N_17210,N_17011,N_17024);
or U17211 (N_17211,N_17177,N_17051);
nand U17212 (N_17212,N_17171,N_17162);
and U17213 (N_17213,N_17055,N_17004);
xnor U17214 (N_17214,N_17025,N_17125);
and U17215 (N_17215,N_17008,N_17166);
xor U17216 (N_17216,N_17021,N_17139);
nor U17217 (N_17217,N_17126,N_17186);
and U17218 (N_17218,N_17044,N_17032);
nand U17219 (N_17219,N_17046,N_17014);
nor U17220 (N_17220,N_17092,N_17040);
and U17221 (N_17221,N_17135,N_17039);
nor U17222 (N_17222,N_17086,N_17007);
xnor U17223 (N_17223,N_17180,N_17100);
nand U17224 (N_17224,N_17065,N_17176);
and U17225 (N_17225,N_17020,N_17189);
or U17226 (N_17226,N_17061,N_17160);
xor U17227 (N_17227,N_17163,N_17017);
and U17228 (N_17228,N_17078,N_17107);
xnor U17229 (N_17229,N_17019,N_17110);
and U17230 (N_17230,N_17016,N_17072);
nor U17231 (N_17231,N_17116,N_17048);
nand U17232 (N_17232,N_17001,N_17074);
nand U17233 (N_17233,N_17143,N_17013);
nor U17234 (N_17234,N_17138,N_17104);
nor U17235 (N_17235,N_17146,N_17120);
nand U17236 (N_17236,N_17037,N_17050);
or U17237 (N_17237,N_17082,N_17114);
and U17238 (N_17238,N_17194,N_17029);
nand U17239 (N_17239,N_17130,N_17041);
or U17240 (N_17240,N_17018,N_17145);
xor U17241 (N_17241,N_17154,N_17150);
and U17242 (N_17242,N_17098,N_17099);
nor U17243 (N_17243,N_17070,N_17106);
nor U17244 (N_17244,N_17022,N_17095);
nand U17245 (N_17245,N_17075,N_17142);
or U17246 (N_17246,N_17043,N_17185);
or U17247 (N_17247,N_17000,N_17134);
or U17248 (N_17248,N_17173,N_17090);
xor U17249 (N_17249,N_17076,N_17133);
or U17250 (N_17250,N_17129,N_17174);
and U17251 (N_17251,N_17047,N_17058);
or U17252 (N_17252,N_17165,N_17198);
nand U17253 (N_17253,N_17164,N_17093);
nand U17254 (N_17254,N_17034,N_17012);
nand U17255 (N_17255,N_17124,N_17188);
or U17256 (N_17256,N_17152,N_17157);
nor U17257 (N_17257,N_17147,N_17035);
nand U17258 (N_17258,N_17172,N_17144);
and U17259 (N_17259,N_17158,N_17094);
nand U17260 (N_17260,N_17108,N_17052);
xor U17261 (N_17261,N_17028,N_17187);
or U17262 (N_17262,N_17087,N_17088);
xor U17263 (N_17263,N_17056,N_17117);
and U17264 (N_17264,N_17010,N_17026);
xnor U17265 (N_17265,N_17042,N_17062);
xor U17266 (N_17266,N_17057,N_17192);
and U17267 (N_17267,N_17064,N_17089);
nand U17268 (N_17268,N_17045,N_17112);
and U17269 (N_17269,N_17113,N_17175);
nand U17270 (N_17270,N_17156,N_17122);
nor U17271 (N_17271,N_17080,N_17030);
nand U17272 (N_17272,N_17084,N_17131);
nor U17273 (N_17273,N_17184,N_17197);
nor U17274 (N_17274,N_17109,N_17023);
or U17275 (N_17275,N_17033,N_17127);
or U17276 (N_17276,N_17182,N_17005);
nand U17277 (N_17277,N_17079,N_17053);
xor U17278 (N_17278,N_17123,N_17073);
and U17279 (N_17279,N_17067,N_17069);
nand U17280 (N_17280,N_17006,N_17179);
xnor U17281 (N_17281,N_17181,N_17049);
or U17282 (N_17282,N_17091,N_17149);
and U17283 (N_17283,N_17140,N_17119);
or U17284 (N_17284,N_17066,N_17031);
or U17285 (N_17285,N_17151,N_17191);
xnor U17286 (N_17286,N_17196,N_17103);
nand U17287 (N_17287,N_17081,N_17009);
xor U17288 (N_17288,N_17054,N_17170);
nand U17289 (N_17289,N_17132,N_17096);
nand U17290 (N_17290,N_17153,N_17068);
xnor U17291 (N_17291,N_17063,N_17003);
or U17292 (N_17292,N_17102,N_17059);
nor U17293 (N_17293,N_17168,N_17036);
nand U17294 (N_17294,N_17193,N_17199);
xor U17295 (N_17295,N_17161,N_17178);
nand U17296 (N_17296,N_17148,N_17101);
and U17297 (N_17297,N_17121,N_17136);
xnor U17298 (N_17298,N_17137,N_17115);
xor U17299 (N_17299,N_17167,N_17159);
or U17300 (N_17300,N_17181,N_17139);
xnor U17301 (N_17301,N_17008,N_17194);
xor U17302 (N_17302,N_17101,N_17078);
xnor U17303 (N_17303,N_17071,N_17053);
or U17304 (N_17304,N_17173,N_17085);
and U17305 (N_17305,N_17167,N_17031);
nand U17306 (N_17306,N_17086,N_17021);
nor U17307 (N_17307,N_17115,N_17037);
and U17308 (N_17308,N_17170,N_17094);
nor U17309 (N_17309,N_17033,N_17125);
nor U17310 (N_17310,N_17030,N_17152);
nand U17311 (N_17311,N_17074,N_17033);
nand U17312 (N_17312,N_17054,N_17103);
or U17313 (N_17313,N_17162,N_17040);
and U17314 (N_17314,N_17106,N_17099);
xnor U17315 (N_17315,N_17180,N_17145);
xnor U17316 (N_17316,N_17017,N_17074);
and U17317 (N_17317,N_17103,N_17101);
or U17318 (N_17318,N_17055,N_17029);
or U17319 (N_17319,N_17122,N_17155);
nor U17320 (N_17320,N_17043,N_17183);
nand U17321 (N_17321,N_17173,N_17166);
or U17322 (N_17322,N_17117,N_17152);
xor U17323 (N_17323,N_17177,N_17118);
nand U17324 (N_17324,N_17017,N_17161);
or U17325 (N_17325,N_17036,N_17166);
or U17326 (N_17326,N_17004,N_17024);
nor U17327 (N_17327,N_17051,N_17159);
nand U17328 (N_17328,N_17185,N_17021);
nor U17329 (N_17329,N_17088,N_17072);
or U17330 (N_17330,N_17076,N_17196);
or U17331 (N_17331,N_17136,N_17047);
nor U17332 (N_17332,N_17112,N_17109);
or U17333 (N_17333,N_17017,N_17160);
nor U17334 (N_17334,N_17130,N_17155);
nor U17335 (N_17335,N_17016,N_17105);
nand U17336 (N_17336,N_17164,N_17009);
or U17337 (N_17337,N_17193,N_17087);
and U17338 (N_17338,N_17169,N_17064);
or U17339 (N_17339,N_17159,N_17095);
nand U17340 (N_17340,N_17192,N_17138);
nor U17341 (N_17341,N_17102,N_17069);
and U17342 (N_17342,N_17037,N_17125);
nor U17343 (N_17343,N_17070,N_17014);
xnor U17344 (N_17344,N_17187,N_17133);
and U17345 (N_17345,N_17163,N_17121);
xnor U17346 (N_17346,N_17184,N_17001);
nand U17347 (N_17347,N_17166,N_17137);
nor U17348 (N_17348,N_17097,N_17099);
nand U17349 (N_17349,N_17172,N_17005);
nor U17350 (N_17350,N_17188,N_17045);
nand U17351 (N_17351,N_17173,N_17004);
and U17352 (N_17352,N_17044,N_17132);
and U17353 (N_17353,N_17102,N_17144);
nand U17354 (N_17354,N_17045,N_17174);
or U17355 (N_17355,N_17069,N_17197);
or U17356 (N_17356,N_17144,N_17087);
nand U17357 (N_17357,N_17014,N_17052);
nor U17358 (N_17358,N_17166,N_17189);
and U17359 (N_17359,N_17192,N_17030);
and U17360 (N_17360,N_17080,N_17088);
nand U17361 (N_17361,N_17040,N_17157);
and U17362 (N_17362,N_17196,N_17024);
nand U17363 (N_17363,N_17181,N_17141);
nor U17364 (N_17364,N_17119,N_17088);
or U17365 (N_17365,N_17188,N_17028);
nand U17366 (N_17366,N_17049,N_17008);
nor U17367 (N_17367,N_17093,N_17135);
nor U17368 (N_17368,N_17063,N_17108);
nand U17369 (N_17369,N_17075,N_17121);
nand U17370 (N_17370,N_17011,N_17010);
xor U17371 (N_17371,N_17119,N_17040);
nor U17372 (N_17372,N_17169,N_17179);
and U17373 (N_17373,N_17176,N_17089);
and U17374 (N_17374,N_17062,N_17110);
or U17375 (N_17375,N_17026,N_17188);
xnor U17376 (N_17376,N_17091,N_17020);
and U17377 (N_17377,N_17086,N_17062);
nor U17378 (N_17378,N_17068,N_17120);
or U17379 (N_17379,N_17143,N_17081);
xor U17380 (N_17380,N_17120,N_17174);
or U17381 (N_17381,N_17036,N_17148);
or U17382 (N_17382,N_17122,N_17191);
or U17383 (N_17383,N_17168,N_17064);
and U17384 (N_17384,N_17119,N_17037);
and U17385 (N_17385,N_17181,N_17175);
and U17386 (N_17386,N_17189,N_17083);
or U17387 (N_17387,N_17122,N_17060);
nand U17388 (N_17388,N_17151,N_17133);
or U17389 (N_17389,N_17164,N_17010);
nor U17390 (N_17390,N_17051,N_17015);
or U17391 (N_17391,N_17094,N_17073);
xor U17392 (N_17392,N_17097,N_17070);
and U17393 (N_17393,N_17055,N_17094);
or U17394 (N_17394,N_17155,N_17127);
and U17395 (N_17395,N_17098,N_17002);
nand U17396 (N_17396,N_17055,N_17123);
or U17397 (N_17397,N_17023,N_17029);
xnor U17398 (N_17398,N_17165,N_17120);
nor U17399 (N_17399,N_17080,N_17172);
or U17400 (N_17400,N_17224,N_17315);
or U17401 (N_17401,N_17310,N_17324);
nor U17402 (N_17402,N_17223,N_17399);
and U17403 (N_17403,N_17263,N_17365);
nor U17404 (N_17404,N_17387,N_17316);
or U17405 (N_17405,N_17379,N_17208);
and U17406 (N_17406,N_17318,N_17375);
nand U17407 (N_17407,N_17236,N_17358);
nand U17408 (N_17408,N_17241,N_17359);
nand U17409 (N_17409,N_17320,N_17322);
and U17410 (N_17410,N_17232,N_17257);
and U17411 (N_17411,N_17344,N_17352);
nand U17412 (N_17412,N_17314,N_17383);
and U17413 (N_17413,N_17242,N_17341);
or U17414 (N_17414,N_17202,N_17378);
or U17415 (N_17415,N_17371,N_17244);
xnor U17416 (N_17416,N_17229,N_17249);
nor U17417 (N_17417,N_17211,N_17312);
xor U17418 (N_17418,N_17277,N_17321);
xnor U17419 (N_17419,N_17271,N_17207);
xor U17420 (N_17420,N_17311,N_17364);
nand U17421 (N_17421,N_17329,N_17396);
or U17422 (N_17422,N_17343,N_17363);
xnor U17423 (N_17423,N_17328,N_17268);
and U17424 (N_17424,N_17309,N_17217);
nor U17425 (N_17425,N_17265,N_17273);
or U17426 (N_17426,N_17376,N_17385);
nor U17427 (N_17427,N_17368,N_17284);
nor U17428 (N_17428,N_17285,N_17326);
xor U17429 (N_17429,N_17302,N_17286);
or U17430 (N_17430,N_17356,N_17215);
xor U17431 (N_17431,N_17209,N_17259);
or U17432 (N_17432,N_17340,N_17353);
and U17433 (N_17433,N_17360,N_17228);
or U17434 (N_17434,N_17346,N_17261);
nand U17435 (N_17435,N_17234,N_17355);
nor U17436 (N_17436,N_17349,N_17380);
xnor U17437 (N_17437,N_17214,N_17243);
and U17438 (N_17438,N_17227,N_17240);
nand U17439 (N_17439,N_17237,N_17304);
xor U17440 (N_17440,N_17275,N_17332);
xor U17441 (N_17441,N_17342,N_17393);
xnor U17442 (N_17442,N_17381,N_17281);
xor U17443 (N_17443,N_17330,N_17398);
nor U17444 (N_17444,N_17231,N_17390);
nand U17445 (N_17445,N_17287,N_17372);
and U17446 (N_17446,N_17303,N_17213);
xor U17447 (N_17447,N_17384,N_17382);
nor U17448 (N_17448,N_17335,N_17313);
nand U17449 (N_17449,N_17388,N_17391);
nand U17450 (N_17450,N_17252,N_17394);
xor U17451 (N_17451,N_17256,N_17200);
and U17452 (N_17452,N_17230,N_17250);
nor U17453 (N_17453,N_17210,N_17377);
and U17454 (N_17454,N_17395,N_17280);
nand U17455 (N_17455,N_17347,N_17266);
and U17456 (N_17456,N_17206,N_17222);
nor U17457 (N_17457,N_17337,N_17269);
or U17458 (N_17458,N_17219,N_17264);
xor U17459 (N_17459,N_17345,N_17258);
nor U17460 (N_17460,N_17246,N_17203);
nor U17461 (N_17461,N_17283,N_17274);
xor U17462 (N_17462,N_17308,N_17218);
nand U17463 (N_17463,N_17221,N_17291);
nand U17464 (N_17464,N_17255,N_17338);
nand U17465 (N_17465,N_17279,N_17317);
nor U17466 (N_17466,N_17362,N_17216);
or U17467 (N_17467,N_17392,N_17386);
xor U17468 (N_17468,N_17293,N_17267);
or U17469 (N_17469,N_17323,N_17270);
or U17470 (N_17470,N_17366,N_17361);
or U17471 (N_17471,N_17233,N_17373);
nor U17472 (N_17472,N_17333,N_17288);
xnor U17473 (N_17473,N_17369,N_17289);
xnor U17474 (N_17474,N_17367,N_17297);
and U17475 (N_17475,N_17290,N_17204);
nor U17476 (N_17476,N_17294,N_17370);
nor U17477 (N_17477,N_17300,N_17350);
nor U17478 (N_17478,N_17374,N_17331);
xnor U17479 (N_17479,N_17319,N_17220);
or U17480 (N_17480,N_17299,N_17292);
or U17481 (N_17481,N_17296,N_17254);
xor U17482 (N_17482,N_17282,N_17339);
and U17483 (N_17483,N_17327,N_17253);
or U17484 (N_17484,N_17239,N_17251);
nand U17485 (N_17485,N_17397,N_17247);
and U17486 (N_17486,N_17212,N_17278);
nand U17487 (N_17487,N_17248,N_17276);
nor U17488 (N_17488,N_17305,N_17298);
xor U17489 (N_17489,N_17357,N_17225);
and U17490 (N_17490,N_17226,N_17235);
or U17491 (N_17491,N_17301,N_17295);
xor U17492 (N_17492,N_17389,N_17272);
nor U17493 (N_17493,N_17201,N_17325);
or U17494 (N_17494,N_17262,N_17306);
or U17495 (N_17495,N_17351,N_17336);
nand U17496 (N_17496,N_17348,N_17205);
xnor U17497 (N_17497,N_17307,N_17354);
and U17498 (N_17498,N_17238,N_17245);
or U17499 (N_17499,N_17260,N_17334);
or U17500 (N_17500,N_17308,N_17273);
nand U17501 (N_17501,N_17232,N_17315);
nand U17502 (N_17502,N_17259,N_17289);
and U17503 (N_17503,N_17379,N_17256);
nor U17504 (N_17504,N_17382,N_17383);
nand U17505 (N_17505,N_17390,N_17225);
xnor U17506 (N_17506,N_17239,N_17390);
and U17507 (N_17507,N_17252,N_17332);
xnor U17508 (N_17508,N_17317,N_17344);
xnor U17509 (N_17509,N_17352,N_17201);
or U17510 (N_17510,N_17301,N_17369);
xor U17511 (N_17511,N_17374,N_17335);
xor U17512 (N_17512,N_17340,N_17244);
and U17513 (N_17513,N_17300,N_17270);
or U17514 (N_17514,N_17387,N_17376);
xor U17515 (N_17515,N_17256,N_17381);
xor U17516 (N_17516,N_17393,N_17240);
nand U17517 (N_17517,N_17243,N_17292);
and U17518 (N_17518,N_17221,N_17266);
xnor U17519 (N_17519,N_17381,N_17371);
nand U17520 (N_17520,N_17268,N_17394);
or U17521 (N_17521,N_17242,N_17327);
and U17522 (N_17522,N_17213,N_17343);
and U17523 (N_17523,N_17354,N_17394);
and U17524 (N_17524,N_17278,N_17203);
nor U17525 (N_17525,N_17201,N_17307);
or U17526 (N_17526,N_17271,N_17369);
xnor U17527 (N_17527,N_17243,N_17212);
and U17528 (N_17528,N_17336,N_17299);
and U17529 (N_17529,N_17227,N_17320);
and U17530 (N_17530,N_17244,N_17222);
and U17531 (N_17531,N_17355,N_17206);
nand U17532 (N_17532,N_17221,N_17305);
xnor U17533 (N_17533,N_17331,N_17347);
nand U17534 (N_17534,N_17261,N_17288);
or U17535 (N_17535,N_17221,N_17200);
or U17536 (N_17536,N_17398,N_17203);
and U17537 (N_17537,N_17236,N_17315);
or U17538 (N_17538,N_17378,N_17239);
or U17539 (N_17539,N_17253,N_17252);
or U17540 (N_17540,N_17314,N_17207);
xor U17541 (N_17541,N_17292,N_17280);
or U17542 (N_17542,N_17380,N_17220);
or U17543 (N_17543,N_17366,N_17306);
and U17544 (N_17544,N_17260,N_17238);
and U17545 (N_17545,N_17272,N_17305);
xor U17546 (N_17546,N_17390,N_17302);
xnor U17547 (N_17547,N_17354,N_17312);
nor U17548 (N_17548,N_17202,N_17270);
and U17549 (N_17549,N_17363,N_17397);
xnor U17550 (N_17550,N_17399,N_17242);
and U17551 (N_17551,N_17227,N_17230);
and U17552 (N_17552,N_17279,N_17261);
nand U17553 (N_17553,N_17363,N_17278);
nand U17554 (N_17554,N_17350,N_17309);
and U17555 (N_17555,N_17296,N_17391);
nand U17556 (N_17556,N_17343,N_17210);
nor U17557 (N_17557,N_17267,N_17211);
and U17558 (N_17558,N_17342,N_17364);
nor U17559 (N_17559,N_17251,N_17202);
nand U17560 (N_17560,N_17209,N_17339);
and U17561 (N_17561,N_17320,N_17229);
or U17562 (N_17562,N_17343,N_17257);
and U17563 (N_17563,N_17273,N_17223);
or U17564 (N_17564,N_17327,N_17200);
xnor U17565 (N_17565,N_17306,N_17289);
nand U17566 (N_17566,N_17361,N_17248);
nor U17567 (N_17567,N_17392,N_17332);
nor U17568 (N_17568,N_17354,N_17239);
or U17569 (N_17569,N_17350,N_17218);
or U17570 (N_17570,N_17363,N_17314);
xnor U17571 (N_17571,N_17276,N_17326);
nand U17572 (N_17572,N_17321,N_17340);
nor U17573 (N_17573,N_17356,N_17274);
nand U17574 (N_17574,N_17293,N_17300);
nand U17575 (N_17575,N_17243,N_17324);
nor U17576 (N_17576,N_17278,N_17353);
nand U17577 (N_17577,N_17320,N_17230);
nand U17578 (N_17578,N_17266,N_17358);
nand U17579 (N_17579,N_17335,N_17371);
nand U17580 (N_17580,N_17382,N_17202);
nor U17581 (N_17581,N_17260,N_17306);
nor U17582 (N_17582,N_17260,N_17383);
xnor U17583 (N_17583,N_17373,N_17241);
nand U17584 (N_17584,N_17237,N_17232);
nor U17585 (N_17585,N_17264,N_17342);
nor U17586 (N_17586,N_17239,N_17370);
nor U17587 (N_17587,N_17284,N_17330);
nor U17588 (N_17588,N_17353,N_17285);
xnor U17589 (N_17589,N_17284,N_17394);
nand U17590 (N_17590,N_17377,N_17272);
nor U17591 (N_17591,N_17234,N_17301);
nor U17592 (N_17592,N_17212,N_17222);
nand U17593 (N_17593,N_17255,N_17305);
nand U17594 (N_17594,N_17332,N_17316);
nand U17595 (N_17595,N_17289,N_17295);
xnor U17596 (N_17596,N_17382,N_17294);
and U17597 (N_17597,N_17390,N_17327);
nor U17598 (N_17598,N_17292,N_17234);
or U17599 (N_17599,N_17262,N_17285);
xnor U17600 (N_17600,N_17458,N_17444);
and U17601 (N_17601,N_17566,N_17422);
xor U17602 (N_17602,N_17576,N_17426);
nor U17603 (N_17603,N_17596,N_17504);
xnor U17604 (N_17604,N_17474,N_17414);
nand U17605 (N_17605,N_17418,N_17515);
and U17606 (N_17606,N_17436,N_17497);
nor U17607 (N_17607,N_17412,N_17518);
nand U17608 (N_17608,N_17472,N_17417);
xnor U17609 (N_17609,N_17523,N_17572);
nor U17610 (N_17610,N_17450,N_17528);
xnor U17611 (N_17611,N_17470,N_17498);
nand U17612 (N_17612,N_17521,N_17540);
nand U17613 (N_17613,N_17456,N_17562);
and U17614 (N_17614,N_17583,N_17505);
nor U17615 (N_17615,N_17533,N_17551);
nor U17616 (N_17616,N_17425,N_17587);
nor U17617 (N_17617,N_17461,N_17558);
xor U17618 (N_17618,N_17559,N_17409);
and U17619 (N_17619,N_17539,N_17594);
nor U17620 (N_17620,N_17452,N_17432);
nor U17621 (N_17621,N_17486,N_17563);
nand U17622 (N_17622,N_17531,N_17479);
nand U17623 (N_17623,N_17541,N_17451);
nand U17624 (N_17624,N_17403,N_17597);
xnor U17625 (N_17625,N_17545,N_17592);
nor U17626 (N_17626,N_17465,N_17549);
and U17627 (N_17627,N_17443,N_17433);
or U17628 (N_17628,N_17481,N_17462);
xnor U17629 (N_17629,N_17509,N_17554);
nor U17630 (N_17630,N_17520,N_17568);
xnor U17631 (N_17631,N_17441,N_17578);
and U17632 (N_17632,N_17502,N_17543);
xnor U17633 (N_17633,N_17435,N_17593);
xnor U17634 (N_17634,N_17471,N_17535);
nand U17635 (N_17635,N_17544,N_17567);
or U17636 (N_17636,N_17582,N_17574);
nand U17637 (N_17637,N_17428,N_17519);
nor U17638 (N_17638,N_17438,N_17410);
and U17639 (N_17639,N_17423,N_17536);
xnor U17640 (N_17640,N_17506,N_17427);
and U17641 (N_17641,N_17512,N_17415);
or U17642 (N_17642,N_17408,N_17495);
nor U17643 (N_17643,N_17575,N_17556);
nor U17644 (N_17644,N_17499,N_17459);
and U17645 (N_17645,N_17577,N_17526);
nor U17646 (N_17646,N_17527,N_17407);
nor U17647 (N_17647,N_17453,N_17421);
and U17648 (N_17648,N_17530,N_17564);
xnor U17649 (N_17649,N_17501,N_17411);
xnor U17650 (N_17650,N_17581,N_17565);
nor U17651 (N_17651,N_17477,N_17442);
nor U17652 (N_17652,N_17516,N_17431);
xnor U17653 (N_17653,N_17448,N_17478);
xor U17654 (N_17654,N_17511,N_17550);
and U17655 (N_17655,N_17494,N_17579);
or U17656 (N_17656,N_17419,N_17555);
and U17657 (N_17657,N_17510,N_17449);
nand U17658 (N_17658,N_17406,N_17416);
nor U17659 (N_17659,N_17500,N_17525);
or U17660 (N_17660,N_17491,N_17586);
nor U17661 (N_17661,N_17404,N_17430);
xor U17662 (N_17662,N_17580,N_17490);
nor U17663 (N_17663,N_17492,N_17517);
xor U17664 (N_17664,N_17538,N_17553);
and U17665 (N_17665,N_17493,N_17420);
and U17666 (N_17666,N_17552,N_17585);
or U17667 (N_17667,N_17557,N_17473);
xnor U17668 (N_17668,N_17476,N_17571);
or U17669 (N_17669,N_17595,N_17591);
xor U17670 (N_17670,N_17485,N_17460);
nand U17671 (N_17671,N_17503,N_17522);
nor U17672 (N_17672,N_17467,N_17524);
or U17673 (N_17673,N_17508,N_17437);
and U17674 (N_17674,N_17546,N_17599);
nand U17675 (N_17675,N_17475,N_17537);
nor U17676 (N_17676,N_17483,N_17542);
or U17677 (N_17677,N_17487,N_17513);
xor U17678 (N_17678,N_17464,N_17514);
nor U17679 (N_17679,N_17589,N_17561);
xnor U17680 (N_17680,N_17598,N_17480);
nand U17681 (N_17681,N_17424,N_17489);
nand U17682 (N_17682,N_17588,N_17440);
nand U17683 (N_17683,N_17455,N_17496);
xor U17684 (N_17684,N_17413,N_17466);
nand U17685 (N_17685,N_17446,N_17469);
nor U17686 (N_17686,N_17445,N_17548);
and U17687 (N_17687,N_17507,N_17529);
or U17688 (N_17688,N_17447,N_17573);
nor U17689 (N_17689,N_17569,N_17570);
and U17690 (N_17690,N_17434,N_17405);
or U17691 (N_17691,N_17482,N_17560);
or U17692 (N_17692,N_17429,N_17463);
or U17693 (N_17693,N_17534,N_17402);
nor U17694 (N_17694,N_17401,N_17454);
and U17695 (N_17695,N_17439,N_17532);
or U17696 (N_17696,N_17584,N_17400);
nor U17697 (N_17697,N_17590,N_17488);
nor U17698 (N_17698,N_17484,N_17468);
xnor U17699 (N_17699,N_17457,N_17547);
and U17700 (N_17700,N_17504,N_17460);
xor U17701 (N_17701,N_17525,N_17591);
nor U17702 (N_17702,N_17569,N_17574);
xor U17703 (N_17703,N_17530,N_17553);
nor U17704 (N_17704,N_17569,N_17430);
xor U17705 (N_17705,N_17413,N_17449);
nor U17706 (N_17706,N_17500,N_17418);
nand U17707 (N_17707,N_17521,N_17497);
xnor U17708 (N_17708,N_17596,N_17438);
xor U17709 (N_17709,N_17560,N_17404);
and U17710 (N_17710,N_17491,N_17472);
nor U17711 (N_17711,N_17519,N_17598);
xnor U17712 (N_17712,N_17451,N_17453);
nor U17713 (N_17713,N_17495,N_17426);
and U17714 (N_17714,N_17537,N_17438);
and U17715 (N_17715,N_17490,N_17527);
or U17716 (N_17716,N_17573,N_17435);
nand U17717 (N_17717,N_17479,N_17406);
nand U17718 (N_17718,N_17444,N_17497);
nand U17719 (N_17719,N_17560,N_17549);
and U17720 (N_17720,N_17526,N_17460);
and U17721 (N_17721,N_17443,N_17494);
nor U17722 (N_17722,N_17556,N_17566);
xnor U17723 (N_17723,N_17563,N_17458);
xnor U17724 (N_17724,N_17445,N_17466);
nor U17725 (N_17725,N_17553,N_17534);
or U17726 (N_17726,N_17524,N_17584);
nor U17727 (N_17727,N_17461,N_17466);
and U17728 (N_17728,N_17545,N_17494);
nand U17729 (N_17729,N_17491,N_17418);
and U17730 (N_17730,N_17554,N_17499);
or U17731 (N_17731,N_17519,N_17480);
or U17732 (N_17732,N_17454,N_17520);
and U17733 (N_17733,N_17435,N_17595);
and U17734 (N_17734,N_17528,N_17557);
xnor U17735 (N_17735,N_17457,N_17594);
xnor U17736 (N_17736,N_17529,N_17525);
xnor U17737 (N_17737,N_17568,N_17446);
nand U17738 (N_17738,N_17481,N_17596);
or U17739 (N_17739,N_17414,N_17472);
or U17740 (N_17740,N_17582,N_17477);
or U17741 (N_17741,N_17547,N_17454);
xor U17742 (N_17742,N_17525,N_17429);
xor U17743 (N_17743,N_17471,N_17560);
xnor U17744 (N_17744,N_17410,N_17406);
xnor U17745 (N_17745,N_17487,N_17576);
and U17746 (N_17746,N_17401,N_17557);
nor U17747 (N_17747,N_17551,N_17549);
or U17748 (N_17748,N_17491,N_17537);
or U17749 (N_17749,N_17407,N_17523);
nor U17750 (N_17750,N_17552,N_17578);
xnor U17751 (N_17751,N_17411,N_17505);
xor U17752 (N_17752,N_17404,N_17536);
or U17753 (N_17753,N_17566,N_17446);
nand U17754 (N_17754,N_17559,N_17487);
nor U17755 (N_17755,N_17594,N_17468);
nand U17756 (N_17756,N_17408,N_17563);
xnor U17757 (N_17757,N_17523,N_17499);
nor U17758 (N_17758,N_17425,N_17492);
nand U17759 (N_17759,N_17489,N_17404);
nor U17760 (N_17760,N_17543,N_17535);
nand U17761 (N_17761,N_17593,N_17469);
or U17762 (N_17762,N_17592,N_17502);
nand U17763 (N_17763,N_17465,N_17520);
or U17764 (N_17764,N_17584,N_17409);
xor U17765 (N_17765,N_17542,N_17421);
or U17766 (N_17766,N_17469,N_17434);
nor U17767 (N_17767,N_17488,N_17563);
nand U17768 (N_17768,N_17559,N_17400);
or U17769 (N_17769,N_17425,N_17588);
nor U17770 (N_17770,N_17591,N_17404);
xnor U17771 (N_17771,N_17475,N_17472);
and U17772 (N_17772,N_17561,N_17555);
nor U17773 (N_17773,N_17526,N_17523);
xor U17774 (N_17774,N_17400,N_17541);
and U17775 (N_17775,N_17442,N_17571);
or U17776 (N_17776,N_17528,N_17430);
xnor U17777 (N_17777,N_17563,N_17560);
nand U17778 (N_17778,N_17412,N_17568);
nand U17779 (N_17779,N_17430,N_17562);
or U17780 (N_17780,N_17462,N_17400);
xnor U17781 (N_17781,N_17520,N_17593);
nand U17782 (N_17782,N_17501,N_17551);
or U17783 (N_17783,N_17525,N_17542);
xnor U17784 (N_17784,N_17448,N_17460);
xor U17785 (N_17785,N_17515,N_17548);
nor U17786 (N_17786,N_17548,N_17523);
and U17787 (N_17787,N_17471,N_17407);
or U17788 (N_17788,N_17533,N_17412);
nor U17789 (N_17789,N_17589,N_17405);
and U17790 (N_17790,N_17562,N_17460);
and U17791 (N_17791,N_17567,N_17519);
and U17792 (N_17792,N_17443,N_17558);
nor U17793 (N_17793,N_17560,N_17524);
nor U17794 (N_17794,N_17444,N_17528);
nand U17795 (N_17795,N_17434,N_17468);
and U17796 (N_17796,N_17548,N_17493);
or U17797 (N_17797,N_17404,N_17455);
or U17798 (N_17798,N_17578,N_17431);
or U17799 (N_17799,N_17500,N_17434);
or U17800 (N_17800,N_17628,N_17641);
xnor U17801 (N_17801,N_17698,N_17753);
nand U17802 (N_17802,N_17623,N_17774);
nor U17803 (N_17803,N_17749,N_17644);
nor U17804 (N_17804,N_17624,N_17704);
xnor U17805 (N_17805,N_17763,N_17744);
or U17806 (N_17806,N_17755,N_17757);
nor U17807 (N_17807,N_17666,N_17741);
nor U17808 (N_17808,N_17664,N_17785);
or U17809 (N_17809,N_17725,N_17632);
and U17810 (N_17810,N_17689,N_17676);
and U17811 (N_17811,N_17608,N_17680);
xnor U17812 (N_17812,N_17708,N_17733);
xnor U17813 (N_17813,N_17653,N_17728);
xnor U17814 (N_17814,N_17773,N_17779);
xor U17815 (N_17815,N_17767,N_17679);
nand U17816 (N_17816,N_17758,N_17713);
xor U17817 (N_17817,N_17724,N_17719);
nor U17818 (N_17818,N_17604,N_17797);
nor U17819 (N_17819,N_17726,N_17621);
nor U17820 (N_17820,N_17788,N_17605);
nor U17821 (N_17821,N_17646,N_17729);
nor U17822 (N_17822,N_17747,N_17671);
xnor U17823 (N_17823,N_17661,N_17791);
or U17824 (N_17824,N_17775,N_17637);
or U17825 (N_17825,N_17638,N_17688);
nor U17826 (N_17826,N_17634,N_17751);
nor U17827 (N_17827,N_17659,N_17610);
and U17828 (N_17828,N_17746,N_17760);
nor U17829 (N_17829,N_17657,N_17798);
and U17830 (N_17830,N_17616,N_17759);
or U17831 (N_17831,N_17672,N_17703);
nor U17832 (N_17832,N_17612,N_17771);
xor U17833 (N_17833,N_17607,N_17740);
nor U17834 (N_17834,N_17777,N_17684);
or U17835 (N_17835,N_17662,N_17640);
nand U17836 (N_17836,N_17602,N_17742);
nand U17837 (N_17837,N_17783,N_17690);
nand U17838 (N_17838,N_17720,N_17776);
or U17839 (N_17839,N_17761,N_17627);
or U17840 (N_17840,N_17642,N_17796);
nand U17841 (N_17841,N_17609,N_17630);
or U17842 (N_17842,N_17691,N_17770);
and U17843 (N_17843,N_17772,N_17613);
nand U17844 (N_17844,N_17606,N_17693);
xor U17845 (N_17845,N_17752,N_17700);
or U17846 (N_17846,N_17625,N_17786);
nor U17847 (N_17847,N_17658,N_17652);
xor U17848 (N_17848,N_17682,N_17732);
nand U17849 (N_17849,N_17631,N_17762);
nand U17850 (N_17850,N_17731,N_17656);
nor U17851 (N_17851,N_17668,N_17790);
and U17852 (N_17852,N_17789,N_17718);
and U17853 (N_17853,N_17667,N_17643);
nor U17854 (N_17854,N_17629,N_17601);
xor U17855 (N_17855,N_17655,N_17717);
nand U17856 (N_17856,N_17648,N_17633);
or U17857 (N_17857,N_17619,N_17692);
and U17858 (N_17858,N_17696,N_17649);
or U17859 (N_17859,N_17603,N_17705);
and U17860 (N_17860,N_17721,N_17681);
nand U17861 (N_17861,N_17739,N_17711);
and U17862 (N_17862,N_17715,N_17635);
and U17863 (N_17863,N_17716,N_17617);
nand U17864 (N_17864,N_17618,N_17722);
xnor U17865 (N_17865,N_17754,N_17673);
and U17866 (N_17866,N_17709,N_17699);
and U17867 (N_17867,N_17714,N_17768);
nor U17868 (N_17868,N_17615,N_17765);
and U17869 (N_17869,N_17600,N_17686);
or U17870 (N_17870,N_17787,N_17685);
and U17871 (N_17871,N_17782,N_17781);
nand U17872 (N_17872,N_17695,N_17674);
xor U17873 (N_17873,N_17793,N_17614);
xor U17874 (N_17874,N_17636,N_17677);
and U17875 (N_17875,N_17647,N_17769);
or U17876 (N_17876,N_17766,N_17622);
nand U17877 (N_17877,N_17727,N_17683);
xnor U17878 (N_17878,N_17712,N_17654);
nor U17879 (N_17879,N_17660,N_17794);
and U17880 (N_17880,N_17734,N_17702);
or U17881 (N_17881,N_17723,N_17650);
nor U17882 (N_17882,N_17738,N_17639);
xnor U17883 (N_17883,N_17651,N_17665);
and U17884 (N_17884,N_17764,N_17670);
nand U17885 (N_17885,N_17710,N_17745);
and U17886 (N_17886,N_17795,N_17707);
nand U17887 (N_17887,N_17697,N_17780);
and U17888 (N_17888,N_17756,N_17620);
nand U17889 (N_17889,N_17694,N_17730);
and U17890 (N_17890,N_17675,N_17799);
or U17891 (N_17891,N_17701,N_17626);
nand U17892 (N_17892,N_17611,N_17678);
and U17893 (N_17893,N_17743,N_17687);
xnor U17894 (N_17894,N_17706,N_17645);
xnor U17895 (N_17895,N_17748,N_17737);
nor U17896 (N_17896,N_17669,N_17736);
or U17897 (N_17897,N_17792,N_17735);
or U17898 (N_17898,N_17750,N_17778);
nand U17899 (N_17899,N_17784,N_17663);
or U17900 (N_17900,N_17787,N_17637);
nor U17901 (N_17901,N_17604,N_17684);
or U17902 (N_17902,N_17675,N_17645);
nand U17903 (N_17903,N_17688,N_17666);
and U17904 (N_17904,N_17705,N_17607);
and U17905 (N_17905,N_17773,N_17693);
nand U17906 (N_17906,N_17679,N_17609);
xnor U17907 (N_17907,N_17790,N_17773);
xor U17908 (N_17908,N_17733,N_17754);
and U17909 (N_17909,N_17628,N_17602);
xnor U17910 (N_17910,N_17605,N_17682);
nor U17911 (N_17911,N_17626,N_17700);
nand U17912 (N_17912,N_17774,N_17689);
and U17913 (N_17913,N_17742,N_17616);
or U17914 (N_17914,N_17741,N_17661);
xor U17915 (N_17915,N_17697,N_17745);
nand U17916 (N_17916,N_17640,N_17650);
nand U17917 (N_17917,N_17680,N_17637);
nand U17918 (N_17918,N_17702,N_17719);
nor U17919 (N_17919,N_17664,N_17633);
nand U17920 (N_17920,N_17660,N_17738);
or U17921 (N_17921,N_17686,N_17715);
nor U17922 (N_17922,N_17735,N_17673);
xnor U17923 (N_17923,N_17792,N_17734);
or U17924 (N_17924,N_17695,N_17614);
nor U17925 (N_17925,N_17685,N_17608);
or U17926 (N_17926,N_17687,N_17794);
nor U17927 (N_17927,N_17620,N_17785);
xnor U17928 (N_17928,N_17785,N_17795);
nand U17929 (N_17929,N_17790,N_17736);
nor U17930 (N_17930,N_17603,N_17660);
nand U17931 (N_17931,N_17797,N_17638);
and U17932 (N_17932,N_17751,N_17716);
or U17933 (N_17933,N_17714,N_17699);
nor U17934 (N_17934,N_17788,N_17622);
xnor U17935 (N_17935,N_17669,N_17757);
nand U17936 (N_17936,N_17775,N_17672);
xnor U17937 (N_17937,N_17703,N_17645);
nor U17938 (N_17938,N_17642,N_17692);
and U17939 (N_17939,N_17703,N_17759);
nor U17940 (N_17940,N_17775,N_17743);
nand U17941 (N_17941,N_17768,N_17752);
nor U17942 (N_17942,N_17614,N_17752);
or U17943 (N_17943,N_17770,N_17602);
xnor U17944 (N_17944,N_17681,N_17643);
xnor U17945 (N_17945,N_17673,N_17641);
xnor U17946 (N_17946,N_17790,N_17707);
and U17947 (N_17947,N_17777,N_17749);
and U17948 (N_17948,N_17643,N_17749);
or U17949 (N_17949,N_17705,N_17615);
nand U17950 (N_17950,N_17641,N_17751);
and U17951 (N_17951,N_17656,N_17635);
xor U17952 (N_17952,N_17703,N_17610);
xor U17953 (N_17953,N_17796,N_17676);
nand U17954 (N_17954,N_17675,N_17726);
nor U17955 (N_17955,N_17713,N_17728);
nor U17956 (N_17956,N_17667,N_17729);
xor U17957 (N_17957,N_17616,N_17709);
xnor U17958 (N_17958,N_17681,N_17703);
xnor U17959 (N_17959,N_17756,N_17764);
nor U17960 (N_17960,N_17615,N_17633);
nor U17961 (N_17961,N_17676,N_17747);
nand U17962 (N_17962,N_17784,N_17765);
nor U17963 (N_17963,N_17781,N_17695);
nand U17964 (N_17964,N_17719,N_17643);
nor U17965 (N_17965,N_17784,N_17763);
xnor U17966 (N_17966,N_17756,N_17629);
nand U17967 (N_17967,N_17652,N_17769);
nand U17968 (N_17968,N_17759,N_17778);
and U17969 (N_17969,N_17710,N_17753);
or U17970 (N_17970,N_17682,N_17742);
xor U17971 (N_17971,N_17688,N_17634);
nor U17972 (N_17972,N_17725,N_17641);
nand U17973 (N_17973,N_17672,N_17705);
or U17974 (N_17974,N_17614,N_17743);
xnor U17975 (N_17975,N_17714,N_17649);
or U17976 (N_17976,N_17620,N_17791);
xnor U17977 (N_17977,N_17721,N_17600);
nor U17978 (N_17978,N_17764,N_17627);
nor U17979 (N_17979,N_17624,N_17761);
nor U17980 (N_17980,N_17780,N_17793);
nand U17981 (N_17981,N_17673,N_17686);
xnor U17982 (N_17982,N_17744,N_17733);
nor U17983 (N_17983,N_17787,N_17794);
xor U17984 (N_17984,N_17754,N_17693);
or U17985 (N_17985,N_17670,N_17720);
xnor U17986 (N_17986,N_17676,N_17797);
nand U17987 (N_17987,N_17681,N_17679);
nor U17988 (N_17988,N_17762,N_17747);
nand U17989 (N_17989,N_17796,N_17770);
xnor U17990 (N_17990,N_17797,N_17714);
or U17991 (N_17991,N_17745,N_17773);
xor U17992 (N_17992,N_17776,N_17636);
nand U17993 (N_17993,N_17693,N_17645);
and U17994 (N_17994,N_17604,N_17657);
or U17995 (N_17995,N_17788,N_17641);
nand U17996 (N_17996,N_17617,N_17633);
or U17997 (N_17997,N_17686,N_17647);
and U17998 (N_17998,N_17681,N_17670);
nor U17999 (N_17999,N_17702,N_17675);
nor U18000 (N_18000,N_17803,N_17944);
and U18001 (N_18001,N_17905,N_17867);
and U18002 (N_18002,N_17871,N_17940);
nand U18003 (N_18003,N_17822,N_17941);
and U18004 (N_18004,N_17876,N_17921);
or U18005 (N_18005,N_17843,N_17999);
nor U18006 (N_18006,N_17989,N_17851);
or U18007 (N_18007,N_17952,N_17899);
and U18008 (N_18008,N_17815,N_17864);
nand U18009 (N_18009,N_17916,N_17947);
nor U18010 (N_18010,N_17942,N_17833);
nand U18011 (N_18011,N_17959,N_17976);
xnor U18012 (N_18012,N_17927,N_17809);
or U18013 (N_18013,N_17813,N_17967);
and U18014 (N_18014,N_17893,N_17934);
xor U18015 (N_18015,N_17885,N_17990);
nand U18016 (N_18016,N_17883,N_17968);
or U18017 (N_18017,N_17849,N_17842);
nor U18018 (N_18018,N_17845,N_17821);
nor U18019 (N_18019,N_17985,N_17907);
nand U18020 (N_18020,N_17856,N_17965);
nand U18021 (N_18021,N_17861,N_17949);
xor U18022 (N_18022,N_17930,N_17848);
or U18023 (N_18023,N_17903,N_17984);
and U18024 (N_18024,N_17844,N_17975);
or U18025 (N_18025,N_17937,N_17924);
and U18026 (N_18026,N_17808,N_17936);
and U18027 (N_18027,N_17805,N_17862);
nor U18028 (N_18028,N_17932,N_17832);
and U18029 (N_18029,N_17824,N_17951);
or U18030 (N_18030,N_17827,N_17973);
nor U18031 (N_18031,N_17854,N_17945);
and U18032 (N_18032,N_17846,N_17869);
nand U18033 (N_18033,N_17841,N_17820);
or U18034 (N_18034,N_17997,N_17982);
xnor U18035 (N_18035,N_17828,N_17962);
xor U18036 (N_18036,N_17906,N_17810);
nor U18037 (N_18037,N_17915,N_17913);
xnor U18038 (N_18038,N_17884,N_17868);
nor U18039 (N_18039,N_17950,N_17819);
or U18040 (N_18040,N_17817,N_17943);
or U18041 (N_18041,N_17960,N_17935);
or U18042 (N_18042,N_17981,N_17858);
and U18043 (N_18043,N_17995,N_17801);
nand U18044 (N_18044,N_17847,N_17926);
xor U18045 (N_18045,N_17928,N_17835);
xor U18046 (N_18046,N_17855,N_17897);
nand U18047 (N_18047,N_17879,N_17972);
nor U18048 (N_18048,N_17958,N_17812);
nor U18049 (N_18049,N_17840,N_17948);
nand U18050 (N_18050,N_17939,N_17831);
nor U18051 (N_18051,N_17909,N_17904);
or U18052 (N_18052,N_17852,N_17863);
nand U18053 (N_18053,N_17900,N_17920);
or U18054 (N_18054,N_17818,N_17823);
or U18055 (N_18055,N_17929,N_17994);
nor U18056 (N_18056,N_17891,N_17898);
and U18057 (N_18057,N_17811,N_17825);
nand U18058 (N_18058,N_17963,N_17918);
and U18059 (N_18059,N_17983,N_17993);
nand U18060 (N_18060,N_17826,N_17908);
or U18061 (N_18061,N_17873,N_17814);
xor U18062 (N_18062,N_17986,N_17922);
or U18063 (N_18063,N_17956,N_17911);
nand U18064 (N_18064,N_17865,N_17838);
nor U18065 (N_18065,N_17955,N_17880);
nor U18066 (N_18066,N_17896,N_17853);
nor U18067 (N_18067,N_17894,N_17837);
xnor U18068 (N_18068,N_17938,N_17850);
xor U18069 (N_18069,N_17980,N_17912);
nor U18070 (N_18070,N_17882,N_17829);
and U18071 (N_18071,N_17866,N_17839);
xor U18072 (N_18072,N_17860,N_17874);
xor U18073 (N_18073,N_17977,N_17919);
or U18074 (N_18074,N_17917,N_17991);
nor U18075 (N_18075,N_17889,N_17979);
nand U18076 (N_18076,N_17870,N_17888);
nand U18077 (N_18077,N_17887,N_17830);
and U18078 (N_18078,N_17923,N_17816);
and U18079 (N_18079,N_17901,N_17998);
nand U18080 (N_18080,N_17987,N_17881);
nand U18081 (N_18081,N_17800,N_17806);
nor U18082 (N_18082,N_17969,N_17914);
nand U18083 (N_18083,N_17978,N_17953);
nand U18084 (N_18084,N_17890,N_17933);
nor U18085 (N_18085,N_17807,N_17875);
and U18086 (N_18086,N_17872,N_17910);
and U18087 (N_18087,N_17996,N_17886);
nor U18088 (N_18088,N_17971,N_17804);
and U18089 (N_18089,N_17988,N_17961);
xor U18090 (N_18090,N_17992,N_17902);
or U18091 (N_18091,N_17859,N_17964);
or U18092 (N_18092,N_17931,N_17802);
xnor U18093 (N_18093,N_17974,N_17836);
or U18094 (N_18094,N_17877,N_17878);
nor U18095 (N_18095,N_17957,N_17857);
nand U18096 (N_18096,N_17895,N_17954);
nand U18097 (N_18097,N_17946,N_17834);
nor U18098 (N_18098,N_17925,N_17970);
and U18099 (N_18099,N_17966,N_17892);
and U18100 (N_18100,N_17802,N_17989);
and U18101 (N_18101,N_17840,N_17818);
and U18102 (N_18102,N_17841,N_17993);
xnor U18103 (N_18103,N_17895,N_17866);
and U18104 (N_18104,N_17949,N_17931);
and U18105 (N_18105,N_17851,N_17873);
or U18106 (N_18106,N_17823,N_17833);
and U18107 (N_18107,N_17869,N_17832);
xor U18108 (N_18108,N_17812,N_17885);
nor U18109 (N_18109,N_17889,N_17930);
nand U18110 (N_18110,N_17991,N_17859);
and U18111 (N_18111,N_17877,N_17972);
or U18112 (N_18112,N_17821,N_17919);
or U18113 (N_18113,N_17940,N_17802);
xor U18114 (N_18114,N_17867,N_17884);
nand U18115 (N_18115,N_17936,N_17996);
nand U18116 (N_18116,N_17856,N_17911);
xor U18117 (N_18117,N_17917,N_17911);
nor U18118 (N_18118,N_17929,N_17881);
and U18119 (N_18119,N_17831,N_17869);
and U18120 (N_18120,N_17909,N_17959);
nand U18121 (N_18121,N_17886,N_17909);
xnor U18122 (N_18122,N_17974,N_17958);
nor U18123 (N_18123,N_17934,N_17909);
xnor U18124 (N_18124,N_17992,N_17829);
nand U18125 (N_18125,N_17982,N_17972);
xor U18126 (N_18126,N_17920,N_17889);
xor U18127 (N_18127,N_17860,N_17914);
nand U18128 (N_18128,N_17952,N_17815);
xor U18129 (N_18129,N_17945,N_17867);
xnor U18130 (N_18130,N_17891,N_17935);
or U18131 (N_18131,N_17981,N_17936);
xnor U18132 (N_18132,N_17921,N_17849);
nand U18133 (N_18133,N_17800,N_17836);
xnor U18134 (N_18134,N_17811,N_17942);
nand U18135 (N_18135,N_17905,N_17948);
or U18136 (N_18136,N_17805,N_17864);
nand U18137 (N_18137,N_17815,N_17854);
nor U18138 (N_18138,N_17881,N_17955);
nand U18139 (N_18139,N_17869,N_17801);
xor U18140 (N_18140,N_17848,N_17888);
nor U18141 (N_18141,N_17803,N_17965);
xor U18142 (N_18142,N_17903,N_17964);
or U18143 (N_18143,N_17827,N_17828);
and U18144 (N_18144,N_17862,N_17910);
nor U18145 (N_18145,N_17988,N_17845);
xor U18146 (N_18146,N_17948,N_17916);
nand U18147 (N_18147,N_17832,N_17811);
and U18148 (N_18148,N_17925,N_17807);
nor U18149 (N_18149,N_17841,N_17999);
nor U18150 (N_18150,N_17960,N_17992);
or U18151 (N_18151,N_17867,N_17908);
nand U18152 (N_18152,N_17809,N_17890);
xnor U18153 (N_18153,N_17974,N_17921);
and U18154 (N_18154,N_17936,N_17864);
nand U18155 (N_18155,N_17878,N_17855);
or U18156 (N_18156,N_17875,N_17859);
nand U18157 (N_18157,N_17984,N_17809);
or U18158 (N_18158,N_17882,N_17925);
or U18159 (N_18159,N_17835,N_17973);
or U18160 (N_18160,N_17888,N_17892);
nand U18161 (N_18161,N_17913,N_17886);
nor U18162 (N_18162,N_17844,N_17834);
and U18163 (N_18163,N_17882,N_17952);
and U18164 (N_18164,N_17925,N_17873);
xor U18165 (N_18165,N_17978,N_17827);
nor U18166 (N_18166,N_17966,N_17802);
nand U18167 (N_18167,N_17893,N_17961);
nor U18168 (N_18168,N_17895,N_17967);
or U18169 (N_18169,N_17816,N_17864);
nand U18170 (N_18170,N_17917,N_17807);
or U18171 (N_18171,N_17871,N_17895);
and U18172 (N_18172,N_17876,N_17964);
nor U18173 (N_18173,N_17951,N_17950);
nand U18174 (N_18174,N_17934,N_17896);
or U18175 (N_18175,N_17915,N_17946);
nor U18176 (N_18176,N_17822,N_17914);
and U18177 (N_18177,N_17925,N_17900);
nor U18178 (N_18178,N_17855,N_17830);
and U18179 (N_18179,N_17984,N_17804);
xor U18180 (N_18180,N_17909,N_17881);
and U18181 (N_18181,N_17817,N_17951);
nor U18182 (N_18182,N_17838,N_17822);
xor U18183 (N_18183,N_17889,N_17948);
and U18184 (N_18184,N_17838,N_17961);
and U18185 (N_18185,N_17899,N_17847);
and U18186 (N_18186,N_17831,N_17935);
or U18187 (N_18187,N_17879,N_17923);
xnor U18188 (N_18188,N_17945,N_17999);
xnor U18189 (N_18189,N_17867,N_17973);
or U18190 (N_18190,N_17937,N_17944);
xor U18191 (N_18191,N_17862,N_17914);
or U18192 (N_18192,N_17866,N_17855);
or U18193 (N_18193,N_17925,N_17986);
or U18194 (N_18194,N_17811,N_17880);
nand U18195 (N_18195,N_17911,N_17849);
and U18196 (N_18196,N_17935,N_17979);
nor U18197 (N_18197,N_17864,N_17851);
nand U18198 (N_18198,N_17878,N_17984);
and U18199 (N_18199,N_17835,N_17825);
or U18200 (N_18200,N_18038,N_18122);
xor U18201 (N_18201,N_18164,N_18185);
and U18202 (N_18202,N_18022,N_18024);
nand U18203 (N_18203,N_18147,N_18137);
nand U18204 (N_18204,N_18199,N_18105);
xnor U18205 (N_18205,N_18091,N_18103);
xnor U18206 (N_18206,N_18014,N_18173);
nor U18207 (N_18207,N_18075,N_18138);
and U18208 (N_18208,N_18002,N_18062);
and U18209 (N_18209,N_18051,N_18080);
or U18210 (N_18210,N_18041,N_18079);
nand U18211 (N_18211,N_18159,N_18025);
nor U18212 (N_18212,N_18174,N_18039);
nor U18213 (N_18213,N_18026,N_18168);
xor U18214 (N_18214,N_18054,N_18176);
nand U18215 (N_18215,N_18195,N_18121);
and U18216 (N_18216,N_18071,N_18037);
xor U18217 (N_18217,N_18089,N_18090);
or U18218 (N_18218,N_18184,N_18048);
nand U18219 (N_18219,N_18156,N_18096);
nor U18220 (N_18220,N_18042,N_18032);
nor U18221 (N_18221,N_18040,N_18072);
and U18222 (N_18222,N_18169,N_18141);
and U18223 (N_18223,N_18009,N_18015);
nor U18224 (N_18224,N_18125,N_18191);
nand U18225 (N_18225,N_18150,N_18019);
or U18226 (N_18226,N_18036,N_18116);
nand U18227 (N_18227,N_18178,N_18110);
and U18228 (N_18228,N_18115,N_18068);
or U18229 (N_18229,N_18175,N_18078);
or U18230 (N_18230,N_18149,N_18183);
or U18231 (N_18231,N_18067,N_18077);
or U18232 (N_18232,N_18070,N_18127);
and U18233 (N_18233,N_18186,N_18189);
or U18234 (N_18234,N_18158,N_18081);
nor U18235 (N_18235,N_18167,N_18058);
or U18236 (N_18236,N_18061,N_18128);
xor U18237 (N_18237,N_18060,N_18082);
nor U18238 (N_18238,N_18064,N_18146);
and U18239 (N_18239,N_18055,N_18131);
xnor U18240 (N_18240,N_18180,N_18047);
xor U18241 (N_18241,N_18117,N_18028);
or U18242 (N_18242,N_18140,N_18165);
nand U18243 (N_18243,N_18119,N_18170);
nor U18244 (N_18244,N_18013,N_18192);
and U18245 (N_18245,N_18144,N_18020);
xnor U18246 (N_18246,N_18107,N_18108);
nor U18247 (N_18247,N_18023,N_18063);
nor U18248 (N_18248,N_18030,N_18123);
nand U18249 (N_18249,N_18021,N_18102);
and U18250 (N_18250,N_18157,N_18053);
nor U18251 (N_18251,N_18076,N_18097);
xnor U18252 (N_18252,N_18008,N_18088);
nor U18253 (N_18253,N_18069,N_18004);
or U18254 (N_18254,N_18109,N_18018);
and U18255 (N_18255,N_18120,N_18151);
and U18256 (N_18256,N_18101,N_18027);
xnor U18257 (N_18257,N_18113,N_18197);
xnor U18258 (N_18258,N_18046,N_18132);
and U18259 (N_18259,N_18066,N_18136);
or U18260 (N_18260,N_18094,N_18172);
xor U18261 (N_18261,N_18056,N_18142);
or U18262 (N_18262,N_18087,N_18112);
nor U18263 (N_18263,N_18126,N_18104);
nor U18264 (N_18264,N_18007,N_18188);
nand U18265 (N_18265,N_18198,N_18065);
nand U18266 (N_18266,N_18153,N_18003);
xnor U18267 (N_18267,N_18074,N_18000);
and U18268 (N_18268,N_18050,N_18034);
nand U18269 (N_18269,N_18052,N_18099);
nor U18270 (N_18270,N_18044,N_18010);
or U18271 (N_18271,N_18017,N_18155);
nand U18272 (N_18272,N_18093,N_18085);
or U18273 (N_18273,N_18049,N_18016);
xor U18274 (N_18274,N_18152,N_18187);
or U18275 (N_18275,N_18190,N_18181);
nand U18276 (N_18276,N_18130,N_18163);
xor U18277 (N_18277,N_18031,N_18012);
nor U18278 (N_18278,N_18114,N_18148);
or U18279 (N_18279,N_18095,N_18134);
or U18280 (N_18280,N_18005,N_18179);
nand U18281 (N_18281,N_18166,N_18143);
and U18282 (N_18282,N_18106,N_18171);
nand U18283 (N_18283,N_18129,N_18135);
nor U18284 (N_18284,N_18160,N_18111);
and U18285 (N_18285,N_18073,N_18177);
and U18286 (N_18286,N_18182,N_18145);
xnor U18287 (N_18287,N_18162,N_18057);
xnor U18288 (N_18288,N_18100,N_18045);
xnor U18289 (N_18289,N_18011,N_18001);
nand U18290 (N_18290,N_18059,N_18118);
nor U18291 (N_18291,N_18029,N_18043);
nand U18292 (N_18292,N_18193,N_18083);
nand U18293 (N_18293,N_18084,N_18154);
nand U18294 (N_18294,N_18194,N_18092);
and U18295 (N_18295,N_18139,N_18133);
nand U18296 (N_18296,N_18161,N_18124);
nand U18297 (N_18297,N_18098,N_18035);
nor U18298 (N_18298,N_18033,N_18006);
and U18299 (N_18299,N_18086,N_18196);
nand U18300 (N_18300,N_18017,N_18066);
and U18301 (N_18301,N_18081,N_18181);
or U18302 (N_18302,N_18133,N_18098);
xnor U18303 (N_18303,N_18031,N_18063);
or U18304 (N_18304,N_18152,N_18081);
and U18305 (N_18305,N_18123,N_18112);
nor U18306 (N_18306,N_18093,N_18087);
or U18307 (N_18307,N_18018,N_18159);
nor U18308 (N_18308,N_18165,N_18127);
or U18309 (N_18309,N_18136,N_18083);
and U18310 (N_18310,N_18185,N_18091);
nand U18311 (N_18311,N_18043,N_18018);
nor U18312 (N_18312,N_18039,N_18130);
and U18313 (N_18313,N_18044,N_18183);
or U18314 (N_18314,N_18014,N_18162);
nor U18315 (N_18315,N_18186,N_18018);
xnor U18316 (N_18316,N_18146,N_18189);
xor U18317 (N_18317,N_18000,N_18084);
or U18318 (N_18318,N_18080,N_18111);
nand U18319 (N_18319,N_18017,N_18003);
and U18320 (N_18320,N_18183,N_18129);
and U18321 (N_18321,N_18067,N_18006);
and U18322 (N_18322,N_18115,N_18061);
xor U18323 (N_18323,N_18070,N_18155);
and U18324 (N_18324,N_18128,N_18171);
or U18325 (N_18325,N_18148,N_18173);
nand U18326 (N_18326,N_18123,N_18041);
or U18327 (N_18327,N_18029,N_18158);
and U18328 (N_18328,N_18138,N_18192);
nor U18329 (N_18329,N_18011,N_18098);
xnor U18330 (N_18330,N_18144,N_18021);
nand U18331 (N_18331,N_18014,N_18168);
nor U18332 (N_18332,N_18065,N_18003);
or U18333 (N_18333,N_18132,N_18076);
nand U18334 (N_18334,N_18120,N_18159);
and U18335 (N_18335,N_18063,N_18194);
and U18336 (N_18336,N_18050,N_18165);
or U18337 (N_18337,N_18048,N_18062);
and U18338 (N_18338,N_18159,N_18130);
nand U18339 (N_18339,N_18076,N_18051);
nor U18340 (N_18340,N_18083,N_18010);
nand U18341 (N_18341,N_18038,N_18060);
or U18342 (N_18342,N_18043,N_18195);
nor U18343 (N_18343,N_18022,N_18093);
xnor U18344 (N_18344,N_18113,N_18120);
and U18345 (N_18345,N_18102,N_18056);
or U18346 (N_18346,N_18069,N_18073);
or U18347 (N_18347,N_18094,N_18116);
nor U18348 (N_18348,N_18038,N_18089);
and U18349 (N_18349,N_18111,N_18117);
nor U18350 (N_18350,N_18137,N_18003);
or U18351 (N_18351,N_18019,N_18183);
nor U18352 (N_18352,N_18044,N_18148);
nor U18353 (N_18353,N_18163,N_18122);
or U18354 (N_18354,N_18138,N_18078);
nand U18355 (N_18355,N_18156,N_18128);
nand U18356 (N_18356,N_18107,N_18123);
nand U18357 (N_18357,N_18061,N_18185);
and U18358 (N_18358,N_18083,N_18120);
nor U18359 (N_18359,N_18152,N_18111);
nor U18360 (N_18360,N_18149,N_18024);
or U18361 (N_18361,N_18198,N_18067);
xnor U18362 (N_18362,N_18046,N_18018);
or U18363 (N_18363,N_18150,N_18177);
and U18364 (N_18364,N_18062,N_18128);
nand U18365 (N_18365,N_18120,N_18177);
and U18366 (N_18366,N_18025,N_18168);
and U18367 (N_18367,N_18103,N_18036);
xnor U18368 (N_18368,N_18062,N_18131);
and U18369 (N_18369,N_18076,N_18163);
nor U18370 (N_18370,N_18098,N_18162);
nor U18371 (N_18371,N_18143,N_18109);
xor U18372 (N_18372,N_18040,N_18067);
nand U18373 (N_18373,N_18097,N_18130);
nand U18374 (N_18374,N_18186,N_18066);
xnor U18375 (N_18375,N_18071,N_18046);
xor U18376 (N_18376,N_18116,N_18010);
or U18377 (N_18377,N_18196,N_18054);
nand U18378 (N_18378,N_18032,N_18113);
nand U18379 (N_18379,N_18140,N_18038);
nand U18380 (N_18380,N_18074,N_18028);
or U18381 (N_18381,N_18190,N_18094);
or U18382 (N_18382,N_18118,N_18065);
and U18383 (N_18383,N_18198,N_18079);
or U18384 (N_18384,N_18151,N_18196);
nor U18385 (N_18385,N_18111,N_18011);
nor U18386 (N_18386,N_18094,N_18084);
nor U18387 (N_18387,N_18002,N_18149);
nor U18388 (N_18388,N_18116,N_18174);
nand U18389 (N_18389,N_18065,N_18149);
nor U18390 (N_18390,N_18126,N_18178);
and U18391 (N_18391,N_18069,N_18072);
and U18392 (N_18392,N_18165,N_18017);
nand U18393 (N_18393,N_18078,N_18004);
nand U18394 (N_18394,N_18014,N_18021);
nor U18395 (N_18395,N_18193,N_18045);
xnor U18396 (N_18396,N_18005,N_18079);
nand U18397 (N_18397,N_18147,N_18152);
xor U18398 (N_18398,N_18133,N_18166);
nor U18399 (N_18399,N_18175,N_18181);
or U18400 (N_18400,N_18266,N_18391);
or U18401 (N_18401,N_18319,N_18358);
nor U18402 (N_18402,N_18379,N_18392);
nand U18403 (N_18403,N_18251,N_18217);
nand U18404 (N_18404,N_18276,N_18261);
nand U18405 (N_18405,N_18343,N_18375);
xor U18406 (N_18406,N_18219,N_18290);
nand U18407 (N_18407,N_18299,N_18317);
nand U18408 (N_18408,N_18389,N_18291);
and U18409 (N_18409,N_18293,N_18374);
xor U18410 (N_18410,N_18275,N_18258);
xor U18411 (N_18411,N_18320,N_18221);
nand U18412 (N_18412,N_18238,N_18370);
and U18413 (N_18413,N_18222,N_18301);
xor U18414 (N_18414,N_18252,N_18287);
nand U18415 (N_18415,N_18386,N_18223);
or U18416 (N_18416,N_18332,N_18333);
or U18417 (N_18417,N_18382,N_18329);
nor U18418 (N_18418,N_18336,N_18200);
or U18419 (N_18419,N_18220,N_18376);
nand U18420 (N_18420,N_18328,N_18260);
nand U18421 (N_18421,N_18216,N_18247);
xor U18422 (N_18422,N_18345,N_18366);
nand U18423 (N_18423,N_18373,N_18321);
nor U18424 (N_18424,N_18241,N_18267);
nand U18425 (N_18425,N_18385,N_18224);
xor U18426 (N_18426,N_18248,N_18339);
or U18427 (N_18427,N_18265,N_18367);
xor U18428 (N_18428,N_18363,N_18364);
or U18429 (N_18429,N_18352,N_18294);
nor U18430 (N_18430,N_18232,N_18323);
and U18431 (N_18431,N_18314,N_18353);
nand U18432 (N_18432,N_18249,N_18213);
or U18433 (N_18433,N_18331,N_18307);
nor U18434 (N_18434,N_18208,N_18225);
nor U18435 (N_18435,N_18322,N_18342);
xnor U18436 (N_18436,N_18348,N_18257);
xor U18437 (N_18437,N_18334,N_18230);
xor U18438 (N_18438,N_18309,N_18354);
nor U18439 (N_18439,N_18242,N_18355);
nor U18440 (N_18440,N_18399,N_18318);
xnor U18441 (N_18441,N_18264,N_18226);
and U18442 (N_18442,N_18227,N_18256);
xor U18443 (N_18443,N_18218,N_18292);
or U18444 (N_18444,N_18233,N_18351);
nor U18445 (N_18445,N_18302,N_18300);
or U18446 (N_18446,N_18346,N_18327);
xor U18447 (N_18447,N_18390,N_18285);
or U18448 (N_18448,N_18202,N_18395);
nor U18449 (N_18449,N_18335,N_18295);
and U18450 (N_18450,N_18337,N_18361);
and U18451 (N_18451,N_18315,N_18387);
nand U18452 (N_18452,N_18371,N_18338);
or U18453 (N_18453,N_18377,N_18255);
or U18454 (N_18454,N_18280,N_18243);
and U18455 (N_18455,N_18305,N_18235);
nand U18456 (N_18456,N_18344,N_18239);
and U18457 (N_18457,N_18326,N_18269);
nor U18458 (N_18458,N_18360,N_18206);
xnor U18459 (N_18459,N_18278,N_18394);
and U18460 (N_18460,N_18362,N_18204);
xor U18461 (N_18461,N_18283,N_18253);
nand U18462 (N_18462,N_18304,N_18214);
or U18463 (N_18463,N_18396,N_18270);
or U18464 (N_18464,N_18262,N_18254);
or U18465 (N_18465,N_18398,N_18350);
xnor U18466 (N_18466,N_18368,N_18341);
nand U18467 (N_18467,N_18286,N_18306);
or U18468 (N_18468,N_18234,N_18274);
or U18469 (N_18469,N_18245,N_18357);
or U18470 (N_18470,N_18347,N_18201);
or U18471 (N_18471,N_18207,N_18237);
nor U18472 (N_18472,N_18288,N_18380);
xor U18473 (N_18473,N_18240,N_18311);
xor U18474 (N_18474,N_18271,N_18210);
nor U18475 (N_18475,N_18303,N_18281);
nand U18476 (N_18476,N_18313,N_18297);
nor U18477 (N_18477,N_18236,N_18284);
and U18478 (N_18478,N_18349,N_18203);
xor U18479 (N_18479,N_18263,N_18298);
nor U18480 (N_18480,N_18324,N_18209);
xnor U18481 (N_18481,N_18215,N_18383);
or U18482 (N_18482,N_18205,N_18372);
xor U18483 (N_18483,N_18356,N_18250);
xor U18484 (N_18484,N_18296,N_18381);
nor U18485 (N_18485,N_18384,N_18397);
nand U18486 (N_18486,N_18340,N_18212);
and U18487 (N_18487,N_18388,N_18365);
xor U18488 (N_18488,N_18308,N_18244);
and U18489 (N_18489,N_18369,N_18272);
and U18490 (N_18490,N_18359,N_18279);
nor U18491 (N_18491,N_18378,N_18273);
or U18492 (N_18492,N_18312,N_18282);
and U18493 (N_18493,N_18229,N_18330);
xor U18494 (N_18494,N_18211,N_18316);
nand U18495 (N_18495,N_18259,N_18228);
nand U18496 (N_18496,N_18393,N_18246);
nand U18497 (N_18497,N_18289,N_18231);
and U18498 (N_18498,N_18310,N_18268);
and U18499 (N_18499,N_18325,N_18277);
xnor U18500 (N_18500,N_18213,N_18301);
nor U18501 (N_18501,N_18230,N_18327);
or U18502 (N_18502,N_18264,N_18270);
and U18503 (N_18503,N_18335,N_18283);
xor U18504 (N_18504,N_18273,N_18224);
or U18505 (N_18505,N_18233,N_18208);
nor U18506 (N_18506,N_18373,N_18386);
nand U18507 (N_18507,N_18370,N_18378);
nor U18508 (N_18508,N_18323,N_18361);
or U18509 (N_18509,N_18398,N_18230);
or U18510 (N_18510,N_18362,N_18348);
and U18511 (N_18511,N_18391,N_18371);
nor U18512 (N_18512,N_18340,N_18337);
nand U18513 (N_18513,N_18289,N_18271);
nor U18514 (N_18514,N_18296,N_18239);
xnor U18515 (N_18515,N_18284,N_18376);
xnor U18516 (N_18516,N_18209,N_18282);
or U18517 (N_18517,N_18289,N_18379);
xnor U18518 (N_18518,N_18214,N_18288);
nor U18519 (N_18519,N_18235,N_18300);
nand U18520 (N_18520,N_18271,N_18338);
xor U18521 (N_18521,N_18221,N_18392);
or U18522 (N_18522,N_18316,N_18267);
and U18523 (N_18523,N_18329,N_18384);
xor U18524 (N_18524,N_18319,N_18247);
nor U18525 (N_18525,N_18320,N_18379);
and U18526 (N_18526,N_18366,N_18310);
and U18527 (N_18527,N_18322,N_18271);
or U18528 (N_18528,N_18282,N_18361);
nand U18529 (N_18529,N_18214,N_18297);
or U18530 (N_18530,N_18381,N_18370);
nor U18531 (N_18531,N_18304,N_18356);
and U18532 (N_18532,N_18311,N_18294);
or U18533 (N_18533,N_18200,N_18367);
nor U18534 (N_18534,N_18322,N_18282);
nand U18535 (N_18535,N_18382,N_18238);
and U18536 (N_18536,N_18243,N_18344);
nor U18537 (N_18537,N_18260,N_18320);
xnor U18538 (N_18538,N_18225,N_18274);
and U18539 (N_18539,N_18290,N_18301);
xnor U18540 (N_18540,N_18273,N_18207);
nand U18541 (N_18541,N_18326,N_18299);
nand U18542 (N_18542,N_18262,N_18337);
or U18543 (N_18543,N_18207,N_18354);
xnor U18544 (N_18544,N_18386,N_18334);
nand U18545 (N_18545,N_18341,N_18222);
nand U18546 (N_18546,N_18362,N_18200);
or U18547 (N_18547,N_18375,N_18262);
xor U18548 (N_18548,N_18374,N_18259);
nor U18549 (N_18549,N_18342,N_18371);
xnor U18550 (N_18550,N_18318,N_18289);
nor U18551 (N_18551,N_18254,N_18251);
nand U18552 (N_18552,N_18286,N_18239);
or U18553 (N_18553,N_18393,N_18248);
or U18554 (N_18554,N_18343,N_18355);
and U18555 (N_18555,N_18238,N_18390);
nand U18556 (N_18556,N_18398,N_18392);
xnor U18557 (N_18557,N_18361,N_18300);
nand U18558 (N_18558,N_18332,N_18327);
nand U18559 (N_18559,N_18372,N_18355);
nor U18560 (N_18560,N_18357,N_18368);
and U18561 (N_18561,N_18256,N_18371);
and U18562 (N_18562,N_18314,N_18388);
or U18563 (N_18563,N_18276,N_18362);
or U18564 (N_18564,N_18275,N_18263);
xor U18565 (N_18565,N_18269,N_18260);
or U18566 (N_18566,N_18353,N_18279);
and U18567 (N_18567,N_18249,N_18345);
and U18568 (N_18568,N_18204,N_18372);
xor U18569 (N_18569,N_18344,N_18290);
nor U18570 (N_18570,N_18202,N_18236);
nor U18571 (N_18571,N_18312,N_18218);
or U18572 (N_18572,N_18275,N_18230);
and U18573 (N_18573,N_18390,N_18300);
xnor U18574 (N_18574,N_18286,N_18230);
nand U18575 (N_18575,N_18262,N_18347);
xnor U18576 (N_18576,N_18287,N_18332);
nor U18577 (N_18577,N_18323,N_18350);
nand U18578 (N_18578,N_18381,N_18365);
xnor U18579 (N_18579,N_18397,N_18338);
xnor U18580 (N_18580,N_18327,N_18328);
and U18581 (N_18581,N_18254,N_18217);
nand U18582 (N_18582,N_18275,N_18268);
nand U18583 (N_18583,N_18316,N_18206);
and U18584 (N_18584,N_18210,N_18221);
or U18585 (N_18585,N_18311,N_18226);
xnor U18586 (N_18586,N_18338,N_18270);
and U18587 (N_18587,N_18361,N_18370);
xnor U18588 (N_18588,N_18226,N_18301);
or U18589 (N_18589,N_18289,N_18309);
and U18590 (N_18590,N_18227,N_18288);
xor U18591 (N_18591,N_18231,N_18307);
and U18592 (N_18592,N_18262,N_18263);
or U18593 (N_18593,N_18213,N_18246);
xor U18594 (N_18594,N_18371,N_18212);
xnor U18595 (N_18595,N_18334,N_18377);
or U18596 (N_18596,N_18391,N_18211);
xor U18597 (N_18597,N_18346,N_18206);
or U18598 (N_18598,N_18237,N_18321);
or U18599 (N_18599,N_18374,N_18380);
and U18600 (N_18600,N_18402,N_18406);
or U18601 (N_18601,N_18530,N_18596);
nand U18602 (N_18602,N_18451,N_18519);
xnor U18603 (N_18603,N_18560,N_18507);
nand U18604 (N_18604,N_18482,N_18520);
nand U18605 (N_18605,N_18450,N_18593);
xor U18606 (N_18606,N_18567,N_18484);
nor U18607 (N_18607,N_18434,N_18432);
or U18608 (N_18608,N_18488,N_18500);
nand U18609 (N_18609,N_18428,N_18509);
xor U18610 (N_18610,N_18581,N_18589);
or U18611 (N_18611,N_18583,N_18590);
nand U18612 (N_18612,N_18407,N_18442);
or U18613 (N_18613,N_18496,N_18457);
and U18614 (N_18614,N_18459,N_18437);
or U18615 (N_18615,N_18541,N_18480);
and U18616 (N_18616,N_18518,N_18400);
nor U18617 (N_18617,N_18591,N_18413);
nor U18618 (N_18618,N_18479,N_18527);
and U18619 (N_18619,N_18462,N_18508);
nor U18620 (N_18620,N_18478,N_18538);
xor U18621 (N_18621,N_18594,N_18515);
nand U18622 (N_18622,N_18526,N_18552);
nand U18623 (N_18623,N_18448,N_18502);
xnor U18624 (N_18624,N_18572,N_18486);
or U18625 (N_18625,N_18592,N_18566);
or U18626 (N_18626,N_18540,N_18458);
and U18627 (N_18627,N_18423,N_18562);
xnor U18628 (N_18628,N_18410,N_18569);
nor U18629 (N_18629,N_18537,N_18582);
nand U18630 (N_18630,N_18564,N_18554);
or U18631 (N_18631,N_18598,N_18467);
or U18632 (N_18632,N_18441,N_18532);
nand U18633 (N_18633,N_18485,N_18439);
nor U18634 (N_18634,N_18573,N_18524);
nor U18635 (N_18635,N_18546,N_18501);
xor U18636 (N_18636,N_18536,N_18525);
nand U18637 (N_18637,N_18542,N_18469);
nand U18638 (N_18638,N_18489,N_18588);
nand U18639 (N_18639,N_18599,N_18559);
nand U18640 (N_18640,N_18403,N_18516);
or U18641 (N_18641,N_18557,N_18440);
nand U18642 (N_18642,N_18495,N_18553);
or U18643 (N_18643,N_18456,N_18419);
or U18644 (N_18644,N_18503,N_18544);
and U18645 (N_18645,N_18504,N_18473);
nand U18646 (N_18646,N_18512,N_18470);
and U18647 (N_18647,N_18521,N_18492);
xnor U18648 (N_18648,N_18422,N_18491);
and U18649 (N_18649,N_18401,N_18424);
xnor U18650 (N_18650,N_18490,N_18597);
and U18651 (N_18651,N_18531,N_18550);
or U18652 (N_18652,N_18412,N_18445);
and U18653 (N_18653,N_18506,N_18463);
and U18654 (N_18654,N_18585,N_18438);
or U18655 (N_18655,N_18558,N_18514);
or U18656 (N_18656,N_18411,N_18426);
nor U18657 (N_18657,N_18427,N_18425);
xor U18658 (N_18658,N_18409,N_18466);
xnor U18659 (N_18659,N_18494,N_18539);
or U18660 (N_18660,N_18580,N_18414);
or U18661 (N_18661,N_18493,N_18433);
and U18662 (N_18662,N_18449,N_18545);
nand U18663 (N_18663,N_18555,N_18416);
xor U18664 (N_18664,N_18579,N_18574);
nor U18665 (N_18665,N_18447,N_18474);
and U18666 (N_18666,N_18571,N_18584);
nor U18667 (N_18667,N_18517,N_18578);
xor U18668 (N_18668,N_18404,N_18513);
or U18669 (N_18669,N_18418,N_18522);
or U18670 (N_18670,N_18529,N_18563);
nand U18671 (N_18671,N_18471,N_18460);
or U18672 (N_18672,N_18595,N_18561);
nor U18673 (N_18673,N_18498,N_18523);
and U18674 (N_18674,N_18547,N_18505);
or U18675 (N_18675,N_18477,N_18430);
and U18676 (N_18676,N_18528,N_18443);
or U18677 (N_18677,N_18468,N_18435);
nand U18678 (N_18678,N_18577,N_18452);
xnor U18679 (N_18679,N_18454,N_18568);
xnor U18680 (N_18680,N_18587,N_18472);
nor U18681 (N_18681,N_18465,N_18455);
xor U18682 (N_18682,N_18415,N_18551);
and U18683 (N_18683,N_18461,N_18510);
xor U18684 (N_18684,N_18431,N_18549);
and U18685 (N_18685,N_18475,N_18429);
or U18686 (N_18686,N_18481,N_18436);
nor U18687 (N_18687,N_18548,N_18408);
or U18688 (N_18688,N_18417,N_18535);
or U18689 (N_18689,N_18464,N_18534);
xor U18690 (N_18690,N_18487,N_18421);
and U18691 (N_18691,N_18556,N_18444);
nor U18692 (N_18692,N_18586,N_18497);
nor U18693 (N_18693,N_18483,N_18576);
xnor U18694 (N_18694,N_18565,N_18543);
nand U18695 (N_18695,N_18499,N_18575);
or U18696 (N_18696,N_18453,N_18533);
or U18697 (N_18697,N_18476,N_18420);
nand U18698 (N_18698,N_18446,N_18405);
nor U18699 (N_18699,N_18570,N_18511);
or U18700 (N_18700,N_18424,N_18476);
nor U18701 (N_18701,N_18534,N_18411);
xor U18702 (N_18702,N_18539,N_18577);
and U18703 (N_18703,N_18412,N_18494);
nand U18704 (N_18704,N_18576,N_18403);
nor U18705 (N_18705,N_18449,N_18556);
and U18706 (N_18706,N_18557,N_18489);
xor U18707 (N_18707,N_18448,N_18454);
or U18708 (N_18708,N_18555,N_18428);
nand U18709 (N_18709,N_18441,N_18483);
or U18710 (N_18710,N_18477,N_18463);
nor U18711 (N_18711,N_18482,N_18471);
xor U18712 (N_18712,N_18453,N_18520);
nor U18713 (N_18713,N_18474,N_18546);
nor U18714 (N_18714,N_18426,N_18446);
and U18715 (N_18715,N_18598,N_18496);
nor U18716 (N_18716,N_18595,N_18484);
xor U18717 (N_18717,N_18433,N_18422);
nand U18718 (N_18718,N_18429,N_18439);
nand U18719 (N_18719,N_18588,N_18484);
nor U18720 (N_18720,N_18478,N_18585);
nor U18721 (N_18721,N_18524,N_18589);
nand U18722 (N_18722,N_18432,N_18502);
nor U18723 (N_18723,N_18574,N_18588);
or U18724 (N_18724,N_18550,N_18538);
or U18725 (N_18725,N_18412,N_18482);
nand U18726 (N_18726,N_18517,N_18556);
nor U18727 (N_18727,N_18447,N_18400);
nor U18728 (N_18728,N_18524,N_18466);
and U18729 (N_18729,N_18460,N_18414);
and U18730 (N_18730,N_18464,N_18434);
and U18731 (N_18731,N_18425,N_18566);
and U18732 (N_18732,N_18459,N_18519);
or U18733 (N_18733,N_18465,N_18566);
xnor U18734 (N_18734,N_18578,N_18537);
nor U18735 (N_18735,N_18409,N_18595);
nand U18736 (N_18736,N_18512,N_18458);
or U18737 (N_18737,N_18400,N_18583);
nand U18738 (N_18738,N_18449,N_18589);
nor U18739 (N_18739,N_18450,N_18548);
nor U18740 (N_18740,N_18508,N_18513);
and U18741 (N_18741,N_18422,N_18595);
or U18742 (N_18742,N_18420,N_18465);
or U18743 (N_18743,N_18510,N_18483);
nand U18744 (N_18744,N_18514,N_18454);
and U18745 (N_18745,N_18444,N_18466);
nand U18746 (N_18746,N_18546,N_18420);
xnor U18747 (N_18747,N_18588,N_18576);
and U18748 (N_18748,N_18402,N_18429);
nor U18749 (N_18749,N_18424,N_18544);
and U18750 (N_18750,N_18442,N_18517);
xnor U18751 (N_18751,N_18433,N_18567);
or U18752 (N_18752,N_18409,N_18520);
or U18753 (N_18753,N_18426,N_18548);
xnor U18754 (N_18754,N_18413,N_18518);
xnor U18755 (N_18755,N_18438,N_18488);
xor U18756 (N_18756,N_18536,N_18415);
or U18757 (N_18757,N_18462,N_18435);
or U18758 (N_18758,N_18427,N_18534);
or U18759 (N_18759,N_18432,N_18526);
and U18760 (N_18760,N_18579,N_18531);
xnor U18761 (N_18761,N_18559,N_18513);
nor U18762 (N_18762,N_18540,N_18589);
or U18763 (N_18763,N_18474,N_18529);
nor U18764 (N_18764,N_18487,N_18506);
nor U18765 (N_18765,N_18490,N_18450);
or U18766 (N_18766,N_18429,N_18443);
xor U18767 (N_18767,N_18556,N_18599);
nand U18768 (N_18768,N_18546,N_18543);
and U18769 (N_18769,N_18565,N_18402);
nand U18770 (N_18770,N_18424,N_18516);
nand U18771 (N_18771,N_18416,N_18459);
nand U18772 (N_18772,N_18578,N_18429);
nand U18773 (N_18773,N_18420,N_18498);
nor U18774 (N_18774,N_18538,N_18521);
and U18775 (N_18775,N_18467,N_18588);
or U18776 (N_18776,N_18463,N_18415);
and U18777 (N_18777,N_18546,N_18586);
or U18778 (N_18778,N_18545,N_18569);
xor U18779 (N_18779,N_18513,N_18402);
nor U18780 (N_18780,N_18568,N_18511);
or U18781 (N_18781,N_18430,N_18520);
and U18782 (N_18782,N_18536,N_18479);
and U18783 (N_18783,N_18408,N_18470);
nor U18784 (N_18784,N_18443,N_18491);
or U18785 (N_18785,N_18550,N_18509);
nor U18786 (N_18786,N_18506,N_18450);
xor U18787 (N_18787,N_18563,N_18503);
or U18788 (N_18788,N_18422,N_18430);
nor U18789 (N_18789,N_18438,N_18477);
or U18790 (N_18790,N_18437,N_18586);
xor U18791 (N_18791,N_18455,N_18495);
nand U18792 (N_18792,N_18531,N_18547);
or U18793 (N_18793,N_18499,N_18446);
or U18794 (N_18794,N_18591,N_18526);
xnor U18795 (N_18795,N_18414,N_18496);
nor U18796 (N_18796,N_18585,N_18430);
or U18797 (N_18797,N_18592,N_18560);
or U18798 (N_18798,N_18469,N_18586);
or U18799 (N_18799,N_18585,N_18545);
and U18800 (N_18800,N_18734,N_18774);
nand U18801 (N_18801,N_18713,N_18697);
or U18802 (N_18802,N_18642,N_18630);
or U18803 (N_18803,N_18624,N_18752);
nor U18804 (N_18804,N_18665,N_18693);
or U18805 (N_18805,N_18668,N_18673);
or U18806 (N_18806,N_18792,N_18634);
and U18807 (N_18807,N_18678,N_18722);
xor U18808 (N_18808,N_18733,N_18637);
or U18809 (N_18809,N_18711,N_18720);
and U18810 (N_18810,N_18756,N_18655);
or U18811 (N_18811,N_18626,N_18645);
nand U18812 (N_18812,N_18747,N_18779);
nand U18813 (N_18813,N_18657,N_18708);
or U18814 (N_18814,N_18788,N_18772);
nor U18815 (N_18815,N_18739,N_18715);
and U18816 (N_18816,N_18729,N_18675);
and U18817 (N_18817,N_18797,N_18652);
and U18818 (N_18818,N_18666,N_18679);
or U18819 (N_18819,N_18707,N_18746);
nor U18820 (N_18820,N_18701,N_18600);
and U18821 (N_18821,N_18609,N_18621);
nand U18822 (N_18822,N_18758,N_18628);
and U18823 (N_18823,N_18755,N_18685);
nor U18824 (N_18824,N_18799,N_18771);
xor U18825 (N_18825,N_18640,N_18727);
nand U18826 (N_18826,N_18648,N_18778);
or U18827 (N_18827,N_18740,N_18632);
xnor U18828 (N_18828,N_18633,N_18623);
or U18829 (N_18829,N_18604,N_18712);
and U18830 (N_18830,N_18647,N_18669);
or U18831 (N_18831,N_18744,N_18680);
and U18832 (N_18832,N_18661,N_18796);
nor U18833 (N_18833,N_18635,N_18664);
xnor U18834 (N_18834,N_18783,N_18718);
nand U18835 (N_18835,N_18775,N_18653);
or U18836 (N_18836,N_18743,N_18646);
xor U18837 (N_18837,N_18631,N_18749);
and U18838 (N_18838,N_18765,N_18753);
or U18839 (N_18839,N_18764,N_18717);
nand U18840 (N_18840,N_18704,N_18617);
xor U18841 (N_18841,N_18798,N_18601);
nor U18842 (N_18842,N_18686,N_18702);
and U18843 (N_18843,N_18638,N_18650);
and U18844 (N_18844,N_18649,N_18723);
xor U18845 (N_18845,N_18670,N_18683);
or U18846 (N_18846,N_18791,N_18793);
nand U18847 (N_18847,N_18687,N_18781);
xor U18848 (N_18848,N_18760,N_18790);
xor U18849 (N_18849,N_18660,N_18745);
or U18850 (N_18850,N_18692,N_18714);
or U18851 (N_18851,N_18751,N_18784);
and U18852 (N_18852,N_18695,N_18651);
nand U18853 (N_18853,N_18659,N_18754);
xor U18854 (N_18854,N_18605,N_18709);
and U18855 (N_18855,N_18730,N_18741);
nand U18856 (N_18856,N_18768,N_18610);
or U18857 (N_18857,N_18611,N_18690);
nand U18858 (N_18858,N_18629,N_18757);
xnor U18859 (N_18859,N_18644,N_18786);
nand U18860 (N_18860,N_18643,N_18607);
nand U18861 (N_18861,N_18620,N_18710);
or U18862 (N_18862,N_18719,N_18766);
or U18863 (N_18863,N_18736,N_18603);
xnor U18864 (N_18864,N_18795,N_18770);
nand U18865 (N_18865,N_18662,N_18671);
or U18866 (N_18866,N_18639,N_18612);
or U18867 (N_18867,N_18732,N_18663);
xnor U18868 (N_18868,N_18636,N_18674);
or U18869 (N_18869,N_18794,N_18667);
or U18870 (N_18870,N_18682,N_18689);
xor U18871 (N_18871,N_18641,N_18615);
or U18872 (N_18872,N_18619,N_18731);
nand U18873 (N_18873,N_18789,N_18785);
or U18874 (N_18874,N_18725,N_18769);
nor U18875 (N_18875,N_18777,N_18762);
and U18876 (N_18876,N_18787,N_18602);
nor U18877 (N_18877,N_18773,N_18684);
xor U18878 (N_18878,N_18694,N_18658);
or U18879 (N_18879,N_18738,N_18696);
nand U18880 (N_18880,N_18672,N_18737);
and U18881 (N_18881,N_18616,N_18699);
nand U18882 (N_18882,N_18700,N_18681);
or U18883 (N_18883,N_18627,N_18759);
nor U18884 (N_18884,N_18625,N_18618);
or U18885 (N_18885,N_18728,N_18608);
and U18886 (N_18886,N_18748,N_18654);
or U18887 (N_18887,N_18780,N_18703);
nand U18888 (N_18888,N_18750,N_18721);
or U18889 (N_18889,N_18761,N_18691);
nand U18890 (N_18890,N_18614,N_18676);
and U18891 (N_18891,N_18613,N_18724);
and U18892 (N_18892,N_18735,N_18742);
xnor U18893 (N_18893,N_18698,N_18606);
nor U18894 (N_18894,N_18776,N_18677);
or U18895 (N_18895,N_18622,N_18656);
and U18896 (N_18896,N_18782,N_18688);
nand U18897 (N_18897,N_18716,N_18706);
nor U18898 (N_18898,N_18726,N_18763);
and U18899 (N_18899,N_18767,N_18705);
nand U18900 (N_18900,N_18618,N_18707);
nor U18901 (N_18901,N_18719,N_18749);
and U18902 (N_18902,N_18762,N_18601);
nand U18903 (N_18903,N_18712,N_18672);
and U18904 (N_18904,N_18756,N_18737);
nand U18905 (N_18905,N_18656,N_18669);
xnor U18906 (N_18906,N_18610,N_18760);
and U18907 (N_18907,N_18679,N_18658);
or U18908 (N_18908,N_18600,N_18779);
nor U18909 (N_18909,N_18642,N_18733);
nor U18910 (N_18910,N_18763,N_18759);
nor U18911 (N_18911,N_18661,N_18793);
xnor U18912 (N_18912,N_18610,N_18736);
and U18913 (N_18913,N_18775,N_18669);
xor U18914 (N_18914,N_18715,N_18793);
nor U18915 (N_18915,N_18729,N_18670);
xor U18916 (N_18916,N_18623,N_18721);
or U18917 (N_18917,N_18683,N_18769);
or U18918 (N_18918,N_18796,N_18676);
or U18919 (N_18919,N_18657,N_18749);
or U18920 (N_18920,N_18789,N_18794);
nand U18921 (N_18921,N_18679,N_18642);
or U18922 (N_18922,N_18611,N_18646);
xor U18923 (N_18923,N_18681,N_18623);
nor U18924 (N_18924,N_18688,N_18646);
nor U18925 (N_18925,N_18607,N_18677);
or U18926 (N_18926,N_18654,N_18614);
nand U18927 (N_18927,N_18684,N_18668);
and U18928 (N_18928,N_18643,N_18788);
nand U18929 (N_18929,N_18699,N_18778);
nor U18930 (N_18930,N_18605,N_18773);
or U18931 (N_18931,N_18615,N_18611);
and U18932 (N_18932,N_18669,N_18785);
nor U18933 (N_18933,N_18779,N_18751);
xor U18934 (N_18934,N_18765,N_18660);
nand U18935 (N_18935,N_18746,N_18624);
nor U18936 (N_18936,N_18726,N_18720);
nand U18937 (N_18937,N_18701,N_18711);
or U18938 (N_18938,N_18757,N_18780);
and U18939 (N_18939,N_18750,N_18648);
xor U18940 (N_18940,N_18615,N_18650);
xnor U18941 (N_18941,N_18701,N_18649);
xnor U18942 (N_18942,N_18614,N_18716);
or U18943 (N_18943,N_18719,N_18704);
xor U18944 (N_18944,N_18752,N_18745);
nand U18945 (N_18945,N_18706,N_18792);
or U18946 (N_18946,N_18677,N_18635);
or U18947 (N_18947,N_18771,N_18641);
nor U18948 (N_18948,N_18605,N_18750);
or U18949 (N_18949,N_18725,N_18635);
and U18950 (N_18950,N_18783,N_18656);
nor U18951 (N_18951,N_18765,N_18795);
and U18952 (N_18952,N_18770,N_18646);
nand U18953 (N_18953,N_18748,N_18681);
nor U18954 (N_18954,N_18741,N_18634);
or U18955 (N_18955,N_18609,N_18658);
or U18956 (N_18956,N_18653,N_18658);
xor U18957 (N_18957,N_18757,N_18746);
xor U18958 (N_18958,N_18756,N_18754);
nand U18959 (N_18959,N_18670,N_18755);
or U18960 (N_18960,N_18783,N_18622);
xnor U18961 (N_18961,N_18735,N_18672);
nand U18962 (N_18962,N_18660,N_18749);
nand U18963 (N_18963,N_18624,N_18601);
nand U18964 (N_18964,N_18737,N_18639);
xnor U18965 (N_18965,N_18720,N_18695);
and U18966 (N_18966,N_18647,N_18680);
nor U18967 (N_18967,N_18634,N_18756);
nand U18968 (N_18968,N_18656,N_18640);
or U18969 (N_18969,N_18622,N_18721);
and U18970 (N_18970,N_18652,N_18766);
and U18971 (N_18971,N_18679,N_18759);
nand U18972 (N_18972,N_18759,N_18645);
and U18973 (N_18973,N_18696,N_18744);
nor U18974 (N_18974,N_18651,N_18770);
nand U18975 (N_18975,N_18648,N_18708);
and U18976 (N_18976,N_18651,N_18755);
nand U18977 (N_18977,N_18756,N_18666);
xor U18978 (N_18978,N_18771,N_18747);
or U18979 (N_18979,N_18684,N_18731);
and U18980 (N_18980,N_18763,N_18611);
nor U18981 (N_18981,N_18786,N_18698);
or U18982 (N_18982,N_18762,N_18735);
xnor U18983 (N_18983,N_18684,N_18615);
nand U18984 (N_18984,N_18787,N_18750);
nand U18985 (N_18985,N_18613,N_18634);
nor U18986 (N_18986,N_18669,N_18768);
nand U18987 (N_18987,N_18656,N_18627);
and U18988 (N_18988,N_18610,N_18638);
nor U18989 (N_18989,N_18701,N_18778);
xnor U18990 (N_18990,N_18724,N_18767);
nor U18991 (N_18991,N_18620,N_18762);
xor U18992 (N_18992,N_18680,N_18768);
nor U18993 (N_18993,N_18755,N_18744);
xor U18994 (N_18994,N_18659,N_18766);
nor U18995 (N_18995,N_18615,N_18751);
nor U18996 (N_18996,N_18731,N_18715);
xor U18997 (N_18997,N_18643,N_18746);
xor U18998 (N_18998,N_18653,N_18654);
nand U18999 (N_18999,N_18668,N_18642);
xnor U19000 (N_19000,N_18819,N_18830);
and U19001 (N_19001,N_18916,N_18980);
nor U19002 (N_19002,N_18908,N_18890);
or U19003 (N_19003,N_18869,N_18887);
xnor U19004 (N_19004,N_18996,N_18837);
or U19005 (N_19005,N_18901,N_18925);
or U19006 (N_19006,N_18967,N_18806);
or U19007 (N_19007,N_18969,N_18891);
nor U19008 (N_19008,N_18818,N_18952);
nand U19009 (N_19009,N_18979,N_18928);
nand U19010 (N_19010,N_18955,N_18807);
and U19011 (N_19011,N_18965,N_18912);
xnor U19012 (N_19012,N_18956,N_18918);
and U19013 (N_19013,N_18898,N_18878);
or U19014 (N_19014,N_18883,N_18886);
xor U19015 (N_19015,N_18958,N_18899);
xor U19016 (N_19016,N_18922,N_18944);
or U19017 (N_19017,N_18850,N_18801);
or U19018 (N_19018,N_18885,N_18931);
xnor U19019 (N_19019,N_18868,N_18810);
and U19020 (N_19020,N_18847,N_18812);
or U19021 (N_19021,N_18917,N_18843);
or U19022 (N_19022,N_18803,N_18968);
xor U19023 (N_19023,N_18932,N_18842);
and U19024 (N_19024,N_18999,N_18892);
xor U19025 (N_19025,N_18904,N_18911);
xnor U19026 (N_19026,N_18848,N_18824);
or U19027 (N_19027,N_18959,N_18838);
nor U19028 (N_19028,N_18948,N_18961);
or U19029 (N_19029,N_18870,N_18945);
and U19030 (N_19030,N_18894,N_18863);
and U19031 (N_19031,N_18920,N_18858);
nor U19032 (N_19032,N_18998,N_18919);
nand U19033 (N_19033,N_18993,N_18835);
nor U19034 (N_19034,N_18888,N_18960);
or U19035 (N_19035,N_18845,N_18989);
and U19036 (N_19036,N_18805,N_18997);
nor U19037 (N_19037,N_18946,N_18926);
and U19038 (N_19038,N_18851,N_18841);
nor U19039 (N_19039,N_18809,N_18934);
or U19040 (N_19040,N_18814,N_18977);
nand U19041 (N_19041,N_18889,N_18984);
xor U19042 (N_19042,N_18896,N_18836);
xnor U19043 (N_19043,N_18895,N_18982);
nor U19044 (N_19044,N_18852,N_18987);
nand U19045 (N_19045,N_18840,N_18902);
or U19046 (N_19046,N_18938,N_18876);
or U19047 (N_19047,N_18981,N_18880);
xor U19048 (N_19048,N_18861,N_18970);
and U19049 (N_19049,N_18913,N_18909);
or U19050 (N_19050,N_18935,N_18940);
nor U19051 (N_19051,N_18834,N_18991);
nand U19052 (N_19052,N_18839,N_18937);
xor U19053 (N_19053,N_18962,N_18846);
nand U19054 (N_19054,N_18828,N_18963);
nor U19055 (N_19055,N_18906,N_18879);
nor U19056 (N_19056,N_18930,N_18910);
or U19057 (N_19057,N_18923,N_18882);
nand U19058 (N_19058,N_18844,N_18856);
nor U19059 (N_19059,N_18831,N_18833);
or U19060 (N_19060,N_18915,N_18914);
or U19061 (N_19061,N_18973,N_18871);
or U19062 (N_19062,N_18823,N_18900);
xor U19063 (N_19063,N_18864,N_18954);
xor U19064 (N_19064,N_18951,N_18854);
nand U19065 (N_19065,N_18893,N_18804);
or U19066 (N_19066,N_18992,N_18903);
nand U19067 (N_19067,N_18942,N_18988);
or U19068 (N_19068,N_18881,N_18816);
nand U19069 (N_19069,N_18985,N_18995);
xnor U19070 (N_19070,N_18978,N_18802);
nor U19071 (N_19071,N_18897,N_18884);
xor U19072 (N_19072,N_18972,N_18949);
nor U19073 (N_19073,N_18867,N_18953);
and U19074 (N_19074,N_18825,N_18950);
or U19075 (N_19075,N_18933,N_18855);
and U19076 (N_19076,N_18865,N_18832);
and U19077 (N_19077,N_18907,N_18815);
xnor U19078 (N_19078,N_18936,N_18872);
or U19079 (N_19079,N_18939,N_18811);
or U19080 (N_19080,N_18983,N_18826);
xnor U19081 (N_19081,N_18866,N_18873);
or U19082 (N_19082,N_18929,N_18941);
or U19083 (N_19083,N_18943,N_18986);
nor U19084 (N_19084,N_18921,N_18808);
nand U19085 (N_19085,N_18817,N_18964);
nand U19086 (N_19086,N_18966,N_18827);
and U19087 (N_19087,N_18976,N_18821);
and U19088 (N_19088,N_18990,N_18947);
nand U19089 (N_19089,N_18957,N_18875);
or U19090 (N_19090,N_18860,N_18874);
nand U19091 (N_19091,N_18859,N_18813);
nand U19092 (N_19092,N_18971,N_18800);
nand U19093 (N_19093,N_18905,N_18924);
nand U19094 (N_19094,N_18994,N_18857);
and U19095 (N_19095,N_18829,N_18862);
xnor U19096 (N_19096,N_18849,N_18927);
or U19097 (N_19097,N_18975,N_18974);
and U19098 (N_19098,N_18853,N_18877);
or U19099 (N_19099,N_18822,N_18820);
or U19100 (N_19100,N_18871,N_18848);
nor U19101 (N_19101,N_18906,N_18819);
or U19102 (N_19102,N_18827,N_18926);
and U19103 (N_19103,N_18858,N_18902);
xor U19104 (N_19104,N_18936,N_18938);
and U19105 (N_19105,N_18944,N_18925);
xor U19106 (N_19106,N_18836,N_18812);
or U19107 (N_19107,N_18975,N_18892);
nand U19108 (N_19108,N_18827,N_18824);
or U19109 (N_19109,N_18809,N_18955);
xor U19110 (N_19110,N_18909,N_18881);
xnor U19111 (N_19111,N_18859,N_18803);
nor U19112 (N_19112,N_18804,N_18934);
xor U19113 (N_19113,N_18857,N_18828);
and U19114 (N_19114,N_18932,N_18973);
nand U19115 (N_19115,N_18813,N_18860);
nor U19116 (N_19116,N_18881,N_18904);
and U19117 (N_19117,N_18861,N_18800);
or U19118 (N_19118,N_18981,N_18892);
xnor U19119 (N_19119,N_18988,N_18898);
nor U19120 (N_19120,N_18893,N_18845);
xor U19121 (N_19121,N_18860,N_18823);
or U19122 (N_19122,N_18880,N_18891);
nand U19123 (N_19123,N_18807,N_18836);
nor U19124 (N_19124,N_18957,N_18934);
xor U19125 (N_19125,N_18869,N_18888);
and U19126 (N_19126,N_18839,N_18938);
nand U19127 (N_19127,N_18829,N_18842);
nand U19128 (N_19128,N_18852,N_18947);
nor U19129 (N_19129,N_18987,N_18911);
nand U19130 (N_19130,N_18823,N_18947);
xor U19131 (N_19131,N_18901,N_18814);
nor U19132 (N_19132,N_18973,N_18923);
nand U19133 (N_19133,N_18872,N_18944);
and U19134 (N_19134,N_18948,N_18862);
xnor U19135 (N_19135,N_18842,N_18864);
and U19136 (N_19136,N_18929,N_18945);
nand U19137 (N_19137,N_18810,N_18817);
nand U19138 (N_19138,N_18855,N_18931);
or U19139 (N_19139,N_18826,N_18886);
xnor U19140 (N_19140,N_18849,N_18987);
xor U19141 (N_19141,N_18809,N_18841);
and U19142 (N_19142,N_18813,N_18975);
or U19143 (N_19143,N_18996,N_18914);
and U19144 (N_19144,N_18888,N_18824);
or U19145 (N_19145,N_18891,N_18877);
and U19146 (N_19146,N_18869,N_18935);
and U19147 (N_19147,N_18925,N_18898);
xnor U19148 (N_19148,N_18810,N_18887);
nand U19149 (N_19149,N_18859,N_18992);
nor U19150 (N_19150,N_18836,N_18837);
xor U19151 (N_19151,N_18907,N_18983);
xnor U19152 (N_19152,N_18987,N_18910);
xnor U19153 (N_19153,N_18963,N_18931);
and U19154 (N_19154,N_18903,N_18826);
nand U19155 (N_19155,N_18927,N_18988);
nor U19156 (N_19156,N_18829,N_18891);
and U19157 (N_19157,N_18810,N_18853);
nor U19158 (N_19158,N_18961,N_18856);
nor U19159 (N_19159,N_18926,N_18812);
or U19160 (N_19160,N_18903,N_18999);
or U19161 (N_19161,N_18984,N_18909);
xor U19162 (N_19162,N_18809,N_18904);
or U19163 (N_19163,N_18859,N_18989);
or U19164 (N_19164,N_18809,N_18873);
or U19165 (N_19165,N_18859,N_18832);
xnor U19166 (N_19166,N_18897,N_18803);
and U19167 (N_19167,N_18861,N_18879);
or U19168 (N_19168,N_18838,N_18975);
or U19169 (N_19169,N_18881,N_18951);
xnor U19170 (N_19170,N_18805,N_18929);
and U19171 (N_19171,N_18894,N_18989);
nand U19172 (N_19172,N_18899,N_18938);
and U19173 (N_19173,N_18817,N_18851);
nor U19174 (N_19174,N_18867,N_18860);
xnor U19175 (N_19175,N_18916,N_18860);
and U19176 (N_19176,N_18810,N_18818);
and U19177 (N_19177,N_18803,N_18847);
and U19178 (N_19178,N_18869,N_18940);
nor U19179 (N_19179,N_18889,N_18999);
nand U19180 (N_19180,N_18960,N_18944);
xnor U19181 (N_19181,N_18878,N_18960);
nor U19182 (N_19182,N_18845,N_18906);
nand U19183 (N_19183,N_18964,N_18922);
xor U19184 (N_19184,N_18937,N_18992);
nor U19185 (N_19185,N_18982,N_18919);
nor U19186 (N_19186,N_18914,N_18846);
or U19187 (N_19187,N_18833,N_18886);
xor U19188 (N_19188,N_18898,N_18981);
nand U19189 (N_19189,N_18992,N_18971);
and U19190 (N_19190,N_18932,N_18887);
xnor U19191 (N_19191,N_18969,N_18957);
xnor U19192 (N_19192,N_18874,N_18817);
nand U19193 (N_19193,N_18852,N_18917);
and U19194 (N_19194,N_18968,N_18929);
xnor U19195 (N_19195,N_18918,N_18840);
xnor U19196 (N_19196,N_18978,N_18957);
xor U19197 (N_19197,N_18899,N_18879);
and U19198 (N_19198,N_18962,N_18928);
or U19199 (N_19199,N_18831,N_18805);
nor U19200 (N_19200,N_19093,N_19083);
or U19201 (N_19201,N_19072,N_19048);
nor U19202 (N_19202,N_19187,N_19071);
nor U19203 (N_19203,N_19011,N_19056);
and U19204 (N_19204,N_19018,N_19198);
xor U19205 (N_19205,N_19184,N_19128);
or U19206 (N_19206,N_19160,N_19163);
nand U19207 (N_19207,N_19015,N_19010);
xor U19208 (N_19208,N_19165,N_19020);
nor U19209 (N_19209,N_19135,N_19067);
or U19210 (N_19210,N_19059,N_19141);
xor U19211 (N_19211,N_19152,N_19191);
xnor U19212 (N_19212,N_19053,N_19029);
xnor U19213 (N_19213,N_19076,N_19132);
xnor U19214 (N_19214,N_19054,N_19147);
xnor U19215 (N_19215,N_19027,N_19004);
nand U19216 (N_19216,N_19116,N_19096);
and U19217 (N_19217,N_19060,N_19088);
or U19218 (N_19218,N_19109,N_19119);
nand U19219 (N_19219,N_19151,N_19002);
and U19220 (N_19220,N_19153,N_19104);
or U19221 (N_19221,N_19057,N_19008);
or U19222 (N_19222,N_19170,N_19155);
nor U19223 (N_19223,N_19085,N_19084);
xor U19224 (N_19224,N_19122,N_19032);
nor U19225 (N_19225,N_19033,N_19194);
and U19226 (N_19226,N_19102,N_19172);
xor U19227 (N_19227,N_19009,N_19098);
and U19228 (N_19228,N_19031,N_19094);
and U19229 (N_19229,N_19006,N_19035);
xor U19230 (N_19230,N_19181,N_19145);
nor U19231 (N_19231,N_19050,N_19196);
and U19232 (N_19232,N_19171,N_19185);
nor U19233 (N_19233,N_19044,N_19188);
and U19234 (N_19234,N_19139,N_19177);
or U19235 (N_19235,N_19156,N_19021);
and U19236 (N_19236,N_19019,N_19065);
nand U19237 (N_19237,N_19061,N_19136);
nand U19238 (N_19238,N_19095,N_19157);
xnor U19239 (N_19239,N_19123,N_19081);
or U19240 (N_19240,N_19164,N_19034);
nor U19241 (N_19241,N_19012,N_19097);
nand U19242 (N_19242,N_19064,N_19111);
xnor U19243 (N_19243,N_19079,N_19073);
nand U19244 (N_19244,N_19052,N_19186);
and U19245 (N_19245,N_19106,N_19195);
nand U19246 (N_19246,N_19068,N_19014);
and U19247 (N_19247,N_19115,N_19007);
nand U19248 (N_19248,N_19023,N_19070);
or U19249 (N_19249,N_19013,N_19161);
nand U19250 (N_19250,N_19114,N_19105);
nand U19251 (N_19251,N_19089,N_19077);
and U19252 (N_19252,N_19125,N_19166);
xor U19253 (N_19253,N_19086,N_19179);
or U19254 (N_19254,N_19154,N_19197);
and U19255 (N_19255,N_19062,N_19180);
and U19256 (N_19256,N_19133,N_19046);
nor U19257 (N_19257,N_19108,N_19099);
or U19258 (N_19258,N_19169,N_19137);
nor U19259 (N_19259,N_19124,N_19022);
nand U19260 (N_19260,N_19131,N_19051);
and U19261 (N_19261,N_19120,N_19080);
nand U19262 (N_19262,N_19142,N_19028);
and U19263 (N_19263,N_19127,N_19075);
nand U19264 (N_19264,N_19178,N_19149);
xor U19265 (N_19265,N_19082,N_19130);
and U19266 (N_19266,N_19016,N_19192);
and U19267 (N_19267,N_19049,N_19158);
nand U19268 (N_19268,N_19017,N_19189);
nor U19269 (N_19269,N_19183,N_19047);
or U19270 (N_19270,N_19100,N_19107);
or U19271 (N_19271,N_19144,N_19182);
and U19272 (N_19272,N_19066,N_19000);
nor U19273 (N_19273,N_19199,N_19038);
nor U19274 (N_19274,N_19055,N_19110);
nor U19275 (N_19275,N_19041,N_19143);
nor U19276 (N_19276,N_19042,N_19148);
nor U19277 (N_19277,N_19140,N_19167);
nor U19278 (N_19278,N_19001,N_19030);
nand U19279 (N_19279,N_19039,N_19025);
nand U19280 (N_19280,N_19058,N_19087);
nor U19281 (N_19281,N_19069,N_19113);
nor U19282 (N_19282,N_19003,N_19168);
xnor U19283 (N_19283,N_19026,N_19126);
nor U19284 (N_19284,N_19045,N_19121);
xor U19285 (N_19285,N_19090,N_19193);
xor U19286 (N_19286,N_19037,N_19150);
nor U19287 (N_19287,N_19146,N_19176);
nor U19288 (N_19288,N_19138,N_19175);
xor U19289 (N_19289,N_19040,N_19103);
or U19290 (N_19290,N_19112,N_19078);
nand U19291 (N_19291,N_19118,N_19036);
or U19292 (N_19292,N_19162,N_19043);
xor U19293 (N_19293,N_19117,N_19063);
xnor U19294 (N_19294,N_19101,N_19129);
xor U19295 (N_19295,N_19092,N_19174);
and U19296 (N_19296,N_19190,N_19074);
or U19297 (N_19297,N_19005,N_19134);
nor U19298 (N_19298,N_19024,N_19173);
nor U19299 (N_19299,N_19159,N_19091);
or U19300 (N_19300,N_19108,N_19029);
and U19301 (N_19301,N_19043,N_19053);
or U19302 (N_19302,N_19040,N_19159);
xnor U19303 (N_19303,N_19105,N_19144);
nand U19304 (N_19304,N_19137,N_19068);
xnor U19305 (N_19305,N_19142,N_19090);
and U19306 (N_19306,N_19021,N_19091);
or U19307 (N_19307,N_19092,N_19035);
nand U19308 (N_19308,N_19094,N_19168);
nand U19309 (N_19309,N_19052,N_19160);
xnor U19310 (N_19310,N_19092,N_19171);
nor U19311 (N_19311,N_19034,N_19165);
or U19312 (N_19312,N_19148,N_19029);
nor U19313 (N_19313,N_19142,N_19064);
nand U19314 (N_19314,N_19059,N_19126);
nor U19315 (N_19315,N_19084,N_19125);
and U19316 (N_19316,N_19029,N_19076);
xnor U19317 (N_19317,N_19111,N_19182);
nand U19318 (N_19318,N_19052,N_19101);
xor U19319 (N_19319,N_19157,N_19067);
nand U19320 (N_19320,N_19058,N_19130);
nand U19321 (N_19321,N_19169,N_19041);
nand U19322 (N_19322,N_19183,N_19010);
nand U19323 (N_19323,N_19102,N_19007);
and U19324 (N_19324,N_19166,N_19151);
nand U19325 (N_19325,N_19117,N_19195);
or U19326 (N_19326,N_19164,N_19118);
and U19327 (N_19327,N_19106,N_19180);
nand U19328 (N_19328,N_19063,N_19064);
nand U19329 (N_19329,N_19183,N_19106);
and U19330 (N_19330,N_19043,N_19069);
nor U19331 (N_19331,N_19008,N_19132);
nor U19332 (N_19332,N_19078,N_19056);
or U19333 (N_19333,N_19189,N_19176);
and U19334 (N_19334,N_19113,N_19183);
and U19335 (N_19335,N_19156,N_19102);
and U19336 (N_19336,N_19141,N_19170);
or U19337 (N_19337,N_19005,N_19044);
nand U19338 (N_19338,N_19178,N_19080);
nand U19339 (N_19339,N_19035,N_19056);
or U19340 (N_19340,N_19191,N_19179);
xor U19341 (N_19341,N_19106,N_19116);
or U19342 (N_19342,N_19172,N_19079);
xnor U19343 (N_19343,N_19110,N_19117);
xnor U19344 (N_19344,N_19111,N_19128);
nor U19345 (N_19345,N_19124,N_19090);
or U19346 (N_19346,N_19066,N_19025);
nand U19347 (N_19347,N_19178,N_19086);
nand U19348 (N_19348,N_19177,N_19074);
xor U19349 (N_19349,N_19050,N_19081);
nor U19350 (N_19350,N_19093,N_19088);
nand U19351 (N_19351,N_19044,N_19026);
nor U19352 (N_19352,N_19137,N_19184);
nor U19353 (N_19353,N_19066,N_19188);
or U19354 (N_19354,N_19122,N_19027);
or U19355 (N_19355,N_19165,N_19167);
and U19356 (N_19356,N_19117,N_19173);
xor U19357 (N_19357,N_19139,N_19056);
or U19358 (N_19358,N_19107,N_19111);
nand U19359 (N_19359,N_19098,N_19083);
or U19360 (N_19360,N_19053,N_19147);
or U19361 (N_19361,N_19143,N_19178);
and U19362 (N_19362,N_19165,N_19189);
or U19363 (N_19363,N_19142,N_19194);
xor U19364 (N_19364,N_19142,N_19072);
or U19365 (N_19365,N_19025,N_19005);
nor U19366 (N_19366,N_19122,N_19120);
xnor U19367 (N_19367,N_19158,N_19065);
xnor U19368 (N_19368,N_19007,N_19124);
nand U19369 (N_19369,N_19053,N_19097);
or U19370 (N_19370,N_19122,N_19005);
nor U19371 (N_19371,N_19162,N_19158);
nand U19372 (N_19372,N_19087,N_19073);
nor U19373 (N_19373,N_19049,N_19088);
and U19374 (N_19374,N_19051,N_19068);
xor U19375 (N_19375,N_19073,N_19136);
nand U19376 (N_19376,N_19013,N_19045);
and U19377 (N_19377,N_19043,N_19111);
xor U19378 (N_19378,N_19024,N_19068);
xor U19379 (N_19379,N_19072,N_19100);
or U19380 (N_19380,N_19021,N_19192);
or U19381 (N_19381,N_19104,N_19197);
nor U19382 (N_19382,N_19071,N_19121);
nor U19383 (N_19383,N_19018,N_19031);
nand U19384 (N_19384,N_19056,N_19105);
nand U19385 (N_19385,N_19184,N_19096);
xor U19386 (N_19386,N_19081,N_19110);
or U19387 (N_19387,N_19104,N_19128);
nor U19388 (N_19388,N_19122,N_19181);
nand U19389 (N_19389,N_19186,N_19057);
xor U19390 (N_19390,N_19039,N_19127);
xor U19391 (N_19391,N_19020,N_19033);
nor U19392 (N_19392,N_19058,N_19005);
nor U19393 (N_19393,N_19080,N_19009);
and U19394 (N_19394,N_19029,N_19165);
xor U19395 (N_19395,N_19013,N_19145);
and U19396 (N_19396,N_19116,N_19174);
nor U19397 (N_19397,N_19120,N_19102);
xor U19398 (N_19398,N_19097,N_19029);
nor U19399 (N_19399,N_19171,N_19088);
nand U19400 (N_19400,N_19308,N_19394);
and U19401 (N_19401,N_19216,N_19241);
and U19402 (N_19402,N_19288,N_19378);
nor U19403 (N_19403,N_19296,N_19212);
nor U19404 (N_19404,N_19312,N_19332);
xor U19405 (N_19405,N_19363,N_19392);
xnor U19406 (N_19406,N_19367,N_19277);
nor U19407 (N_19407,N_19346,N_19356);
nor U19408 (N_19408,N_19359,N_19274);
and U19409 (N_19409,N_19347,N_19328);
nor U19410 (N_19410,N_19223,N_19334);
nor U19411 (N_19411,N_19300,N_19293);
or U19412 (N_19412,N_19201,N_19380);
xor U19413 (N_19413,N_19360,N_19391);
nand U19414 (N_19414,N_19266,N_19203);
and U19415 (N_19415,N_19270,N_19243);
nor U19416 (N_19416,N_19206,N_19321);
xnor U19417 (N_19417,N_19211,N_19306);
xor U19418 (N_19418,N_19204,N_19291);
nor U19419 (N_19419,N_19205,N_19396);
xnor U19420 (N_19420,N_19244,N_19220);
xor U19421 (N_19421,N_19251,N_19264);
or U19422 (N_19422,N_19272,N_19322);
nand U19423 (N_19423,N_19326,N_19325);
nor U19424 (N_19424,N_19222,N_19342);
nand U19425 (N_19425,N_19304,N_19289);
nor U19426 (N_19426,N_19311,N_19388);
or U19427 (N_19427,N_19215,N_19231);
and U19428 (N_19428,N_19250,N_19239);
xor U19429 (N_19429,N_19252,N_19237);
nor U19430 (N_19430,N_19324,N_19278);
or U19431 (N_19431,N_19372,N_19208);
nand U19432 (N_19432,N_19353,N_19207);
xor U19433 (N_19433,N_19302,N_19265);
and U19434 (N_19434,N_19393,N_19294);
nand U19435 (N_19435,N_19268,N_19390);
and U19436 (N_19436,N_19267,N_19316);
or U19437 (N_19437,N_19383,N_19338);
and U19438 (N_19438,N_19336,N_19357);
or U19439 (N_19439,N_19209,N_19318);
nor U19440 (N_19440,N_19249,N_19301);
nand U19441 (N_19441,N_19361,N_19295);
xor U19442 (N_19442,N_19303,N_19213);
or U19443 (N_19443,N_19314,N_19310);
xnor U19444 (N_19444,N_19350,N_19298);
nand U19445 (N_19445,N_19240,N_19370);
or U19446 (N_19446,N_19276,N_19255);
or U19447 (N_19447,N_19235,N_19340);
xor U19448 (N_19448,N_19242,N_19283);
nand U19449 (N_19449,N_19200,N_19327);
nand U19450 (N_19450,N_19232,N_19349);
or U19451 (N_19451,N_19384,N_19245);
and U19452 (N_19452,N_19290,N_19271);
nand U19453 (N_19453,N_19313,N_19233);
nor U19454 (N_19454,N_19224,N_19269);
and U19455 (N_19455,N_19297,N_19238);
nand U19456 (N_19456,N_19248,N_19309);
xor U19457 (N_19457,N_19284,N_19225);
nand U19458 (N_19458,N_19210,N_19364);
nor U19459 (N_19459,N_19263,N_19320);
or U19460 (N_19460,N_19354,N_19234);
xor U19461 (N_19461,N_19330,N_19374);
and U19462 (N_19462,N_19285,N_19262);
nor U19463 (N_19463,N_19398,N_19339);
and U19464 (N_19464,N_19259,N_19292);
nand U19465 (N_19465,N_19315,N_19228);
nand U19466 (N_19466,N_19280,N_19227);
xor U19467 (N_19467,N_19369,N_19366);
nand U19468 (N_19468,N_19254,N_19246);
nand U19469 (N_19469,N_19395,N_19226);
or U19470 (N_19470,N_19273,N_19399);
or U19471 (N_19471,N_19257,N_19218);
or U19472 (N_19472,N_19258,N_19362);
or U19473 (N_19473,N_19345,N_19329);
nor U19474 (N_19474,N_19341,N_19279);
nor U19475 (N_19475,N_19229,N_19343);
and U19476 (N_19476,N_19261,N_19333);
and U19477 (N_19477,N_19379,N_19371);
and U19478 (N_19478,N_19337,N_19373);
nand U19479 (N_19479,N_19387,N_19375);
or U19480 (N_19480,N_19351,N_19260);
nor U19481 (N_19481,N_19281,N_19317);
nand U19482 (N_19482,N_19368,N_19331);
nor U19483 (N_19483,N_19376,N_19221);
or U19484 (N_19484,N_19335,N_19381);
or U19485 (N_19485,N_19214,N_19389);
xnor U19486 (N_19486,N_19275,N_19253);
xnor U19487 (N_19487,N_19247,N_19202);
or U19488 (N_19488,N_19299,N_19319);
xnor U19489 (N_19489,N_19358,N_19344);
or U19490 (N_19490,N_19385,N_19219);
and U19491 (N_19491,N_19365,N_19382);
xnor U19492 (N_19492,N_19217,N_19355);
xor U19493 (N_19493,N_19236,N_19352);
xor U19494 (N_19494,N_19323,N_19286);
nor U19495 (N_19495,N_19397,N_19307);
nor U19496 (N_19496,N_19377,N_19305);
xor U19497 (N_19497,N_19282,N_19386);
nor U19498 (N_19498,N_19287,N_19348);
nor U19499 (N_19499,N_19230,N_19256);
xnor U19500 (N_19500,N_19287,N_19205);
xor U19501 (N_19501,N_19290,N_19253);
nand U19502 (N_19502,N_19394,N_19320);
xor U19503 (N_19503,N_19229,N_19357);
or U19504 (N_19504,N_19246,N_19280);
or U19505 (N_19505,N_19231,N_19218);
nor U19506 (N_19506,N_19370,N_19347);
nor U19507 (N_19507,N_19347,N_19250);
nor U19508 (N_19508,N_19391,N_19273);
and U19509 (N_19509,N_19298,N_19342);
xnor U19510 (N_19510,N_19258,N_19340);
nand U19511 (N_19511,N_19223,N_19290);
nor U19512 (N_19512,N_19306,N_19287);
or U19513 (N_19513,N_19314,N_19285);
nor U19514 (N_19514,N_19381,N_19283);
xor U19515 (N_19515,N_19322,N_19388);
nand U19516 (N_19516,N_19275,N_19375);
or U19517 (N_19517,N_19283,N_19201);
and U19518 (N_19518,N_19340,N_19283);
xnor U19519 (N_19519,N_19318,N_19294);
xor U19520 (N_19520,N_19331,N_19280);
xor U19521 (N_19521,N_19391,N_19326);
nand U19522 (N_19522,N_19204,N_19201);
or U19523 (N_19523,N_19240,N_19292);
and U19524 (N_19524,N_19240,N_19251);
or U19525 (N_19525,N_19309,N_19315);
or U19526 (N_19526,N_19370,N_19293);
and U19527 (N_19527,N_19206,N_19293);
nor U19528 (N_19528,N_19247,N_19384);
or U19529 (N_19529,N_19282,N_19346);
nor U19530 (N_19530,N_19275,N_19262);
nor U19531 (N_19531,N_19289,N_19221);
or U19532 (N_19532,N_19260,N_19212);
nand U19533 (N_19533,N_19307,N_19296);
and U19534 (N_19534,N_19350,N_19399);
or U19535 (N_19535,N_19350,N_19290);
and U19536 (N_19536,N_19345,N_19287);
nand U19537 (N_19537,N_19374,N_19385);
and U19538 (N_19538,N_19363,N_19280);
nor U19539 (N_19539,N_19335,N_19251);
and U19540 (N_19540,N_19272,N_19252);
and U19541 (N_19541,N_19363,N_19209);
or U19542 (N_19542,N_19299,N_19246);
and U19543 (N_19543,N_19279,N_19272);
nor U19544 (N_19544,N_19222,N_19289);
xnor U19545 (N_19545,N_19384,N_19387);
nor U19546 (N_19546,N_19259,N_19397);
or U19547 (N_19547,N_19261,N_19376);
nor U19548 (N_19548,N_19207,N_19229);
and U19549 (N_19549,N_19375,N_19265);
or U19550 (N_19550,N_19354,N_19320);
or U19551 (N_19551,N_19282,N_19355);
and U19552 (N_19552,N_19212,N_19353);
nand U19553 (N_19553,N_19313,N_19266);
or U19554 (N_19554,N_19213,N_19226);
or U19555 (N_19555,N_19349,N_19399);
nand U19556 (N_19556,N_19302,N_19224);
nand U19557 (N_19557,N_19277,N_19338);
or U19558 (N_19558,N_19240,N_19216);
or U19559 (N_19559,N_19284,N_19326);
or U19560 (N_19560,N_19384,N_19238);
xor U19561 (N_19561,N_19310,N_19317);
xnor U19562 (N_19562,N_19238,N_19203);
xnor U19563 (N_19563,N_19227,N_19304);
xor U19564 (N_19564,N_19334,N_19282);
nand U19565 (N_19565,N_19220,N_19348);
xor U19566 (N_19566,N_19384,N_19286);
and U19567 (N_19567,N_19349,N_19301);
xnor U19568 (N_19568,N_19224,N_19346);
nor U19569 (N_19569,N_19351,N_19342);
or U19570 (N_19570,N_19346,N_19338);
or U19571 (N_19571,N_19275,N_19356);
or U19572 (N_19572,N_19228,N_19345);
and U19573 (N_19573,N_19319,N_19345);
nand U19574 (N_19574,N_19280,N_19301);
nand U19575 (N_19575,N_19336,N_19303);
nor U19576 (N_19576,N_19303,N_19370);
nand U19577 (N_19577,N_19362,N_19399);
or U19578 (N_19578,N_19385,N_19333);
and U19579 (N_19579,N_19384,N_19306);
and U19580 (N_19580,N_19225,N_19393);
nor U19581 (N_19581,N_19288,N_19243);
and U19582 (N_19582,N_19233,N_19223);
xor U19583 (N_19583,N_19246,N_19333);
or U19584 (N_19584,N_19358,N_19361);
xor U19585 (N_19585,N_19278,N_19274);
or U19586 (N_19586,N_19225,N_19347);
nor U19587 (N_19587,N_19219,N_19239);
nor U19588 (N_19588,N_19335,N_19206);
or U19589 (N_19589,N_19310,N_19385);
nor U19590 (N_19590,N_19278,N_19206);
nor U19591 (N_19591,N_19323,N_19320);
nor U19592 (N_19592,N_19280,N_19367);
and U19593 (N_19593,N_19263,N_19264);
xor U19594 (N_19594,N_19216,N_19339);
nor U19595 (N_19595,N_19230,N_19211);
nand U19596 (N_19596,N_19317,N_19367);
xnor U19597 (N_19597,N_19377,N_19226);
or U19598 (N_19598,N_19320,N_19241);
and U19599 (N_19599,N_19281,N_19337);
and U19600 (N_19600,N_19400,N_19516);
nor U19601 (N_19601,N_19427,N_19420);
nor U19602 (N_19602,N_19506,N_19578);
nand U19603 (N_19603,N_19589,N_19539);
and U19604 (N_19604,N_19425,N_19435);
or U19605 (N_19605,N_19575,N_19529);
and U19606 (N_19606,N_19556,N_19402);
xor U19607 (N_19607,N_19544,N_19485);
and U19608 (N_19608,N_19585,N_19500);
or U19609 (N_19609,N_19410,N_19525);
and U19610 (N_19610,N_19462,N_19587);
xnor U19611 (N_19611,N_19492,N_19567);
and U19612 (N_19612,N_19482,N_19576);
or U19613 (N_19613,N_19509,N_19561);
nor U19614 (N_19614,N_19433,N_19554);
nor U19615 (N_19615,N_19411,N_19536);
and U19616 (N_19616,N_19495,N_19439);
nor U19617 (N_19617,N_19428,N_19530);
and U19618 (N_19618,N_19552,N_19545);
nor U19619 (N_19619,N_19571,N_19514);
nor U19620 (N_19620,N_19431,N_19437);
or U19621 (N_19621,N_19465,N_19534);
or U19622 (N_19622,N_19555,N_19548);
nand U19623 (N_19623,N_19592,N_19560);
nand U19624 (N_19624,N_19583,N_19542);
and U19625 (N_19625,N_19598,N_19520);
xnor U19626 (N_19626,N_19455,N_19523);
and U19627 (N_19627,N_19527,N_19562);
and U19628 (N_19628,N_19572,N_19450);
nor U19629 (N_19629,N_19564,N_19498);
or U19630 (N_19630,N_19547,N_19593);
and U19631 (N_19631,N_19553,N_19404);
and U19632 (N_19632,N_19401,N_19438);
nand U19633 (N_19633,N_19582,N_19540);
xnor U19634 (N_19634,N_19409,N_19449);
xnor U19635 (N_19635,N_19533,N_19412);
and U19636 (N_19636,N_19568,N_19436);
nand U19637 (N_19637,N_19416,N_19418);
xnor U19638 (N_19638,N_19446,N_19531);
nor U19639 (N_19639,N_19429,N_19467);
xor U19640 (N_19640,N_19508,N_19426);
and U19641 (N_19641,N_19403,N_19565);
nor U19642 (N_19642,N_19470,N_19595);
xor U19643 (N_19643,N_19430,N_19408);
and U19644 (N_19644,N_19457,N_19489);
xnor U19645 (N_19645,N_19473,N_19591);
and U19646 (N_19646,N_19452,N_19468);
nor U19647 (N_19647,N_19524,N_19596);
xnor U19648 (N_19648,N_19479,N_19549);
or U19649 (N_19649,N_19496,N_19494);
xnor U19650 (N_19650,N_19557,N_19484);
xor U19651 (N_19651,N_19488,N_19537);
xnor U19652 (N_19652,N_19415,N_19459);
xor U19653 (N_19653,N_19421,N_19503);
xor U19654 (N_19654,N_19422,N_19458);
or U19655 (N_19655,N_19580,N_19586);
or U19656 (N_19656,N_19518,N_19451);
nor U19657 (N_19657,N_19543,N_19541);
and U19658 (N_19658,N_19413,N_19521);
nor U19659 (N_19659,N_19469,N_19577);
or U19660 (N_19660,N_19442,N_19487);
nor U19661 (N_19661,N_19460,N_19434);
and U19662 (N_19662,N_19502,N_19478);
or U19663 (N_19663,N_19481,N_19483);
and U19664 (N_19664,N_19476,N_19475);
xor U19665 (N_19665,N_19448,N_19574);
nor U19666 (N_19666,N_19546,N_19456);
nand U19667 (N_19667,N_19463,N_19445);
xor U19668 (N_19668,N_19550,N_19581);
nand U19669 (N_19669,N_19535,N_19424);
and U19670 (N_19670,N_19515,N_19490);
nor U19671 (N_19671,N_19480,N_19477);
nand U19672 (N_19672,N_19441,N_19573);
xnor U19673 (N_19673,N_19566,N_19570);
nand U19674 (N_19674,N_19405,N_19497);
or U19675 (N_19675,N_19522,N_19505);
nor U19676 (N_19676,N_19499,N_19528);
or U19677 (N_19677,N_19590,N_19406);
nor U19678 (N_19678,N_19419,N_19519);
nor U19679 (N_19679,N_19510,N_19417);
or U19680 (N_19680,N_19407,N_19471);
nand U19681 (N_19681,N_19551,N_19563);
or U19682 (N_19682,N_19526,N_19512);
nor U19683 (N_19683,N_19466,N_19558);
and U19684 (N_19684,N_19579,N_19472);
nand U19685 (N_19685,N_19559,N_19493);
or U19686 (N_19686,N_19588,N_19440);
nor U19687 (N_19687,N_19423,N_19491);
nor U19688 (N_19688,N_19532,N_19584);
xor U19689 (N_19689,N_19486,N_19507);
xnor U19690 (N_19690,N_19597,N_19511);
or U19691 (N_19691,N_19461,N_19414);
nand U19692 (N_19692,N_19432,N_19569);
and U19693 (N_19693,N_19501,N_19517);
xor U19694 (N_19694,N_19464,N_19447);
xor U19695 (N_19695,N_19594,N_19444);
nor U19696 (N_19696,N_19513,N_19599);
nor U19697 (N_19697,N_19453,N_19454);
and U19698 (N_19698,N_19474,N_19538);
and U19699 (N_19699,N_19443,N_19504);
nor U19700 (N_19700,N_19462,N_19516);
nand U19701 (N_19701,N_19470,N_19432);
xor U19702 (N_19702,N_19468,N_19422);
or U19703 (N_19703,N_19449,N_19514);
and U19704 (N_19704,N_19439,N_19463);
nor U19705 (N_19705,N_19520,N_19431);
and U19706 (N_19706,N_19429,N_19532);
xor U19707 (N_19707,N_19558,N_19525);
and U19708 (N_19708,N_19545,N_19529);
nand U19709 (N_19709,N_19453,N_19446);
nand U19710 (N_19710,N_19596,N_19572);
and U19711 (N_19711,N_19536,N_19558);
xor U19712 (N_19712,N_19567,N_19441);
nand U19713 (N_19713,N_19439,N_19542);
nor U19714 (N_19714,N_19445,N_19412);
or U19715 (N_19715,N_19445,N_19406);
and U19716 (N_19716,N_19532,N_19560);
and U19717 (N_19717,N_19537,N_19518);
or U19718 (N_19718,N_19566,N_19400);
nand U19719 (N_19719,N_19571,N_19558);
nand U19720 (N_19720,N_19477,N_19568);
nand U19721 (N_19721,N_19566,N_19536);
nand U19722 (N_19722,N_19540,N_19520);
and U19723 (N_19723,N_19453,N_19482);
xnor U19724 (N_19724,N_19481,N_19514);
nor U19725 (N_19725,N_19448,N_19523);
xor U19726 (N_19726,N_19565,N_19449);
xor U19727 (N_19727,N_19553,N_19420);
xor U19728 (N_19728,N_19467,N_19432);
nor U19729 (N_19729,N_19522,N_19485);
or U19730 (N_19730,N_19534,N_19584);
or U19731 (N_19731,N_19496,N_19508);
nand U19732 (N_19732,N_19434,N_19487);
xnor U19733 (N_19733,N_19482,N_19545);
nand U19734 (N_19734,N_19495,N_19564);
nor U19735 (N_19735,N_19512,N_19584);
and U19736 (N_19736,N_19506,N_19495);
nand U19737 (N_19737,N_19579,N_19404);
xnor U19738 (N_19738,N_19512,N_19424);
and U19739 (N_19739,N_19595,N_19570);
or U19740 (N_19740,N_19595,N_19572);
nand U19741 (N_19741,N_19557,N_19457);
nand U19742 (N_19742,N_19589,N_19576);
nor U19743 (N_19743,N_19558,N_19553);
and U19744 (N_19744,N_19478,N_19585);
xor U19745 (N_19745,N_19404,N_19582);
nor U19746 (N_19746,N_19491,N_19414);
xnor U19747 (N_19747,N_19477,N_19440);
nor U19748 (N_19748,N_19503,N_19518);
or U19749 (N_19749,N_19406,N_19565);
nor U19750 (N_19750,N_19545,N_19435);
nand U19751 (N_19751,N_19476,N_19538);
or U19752 (N_19752,N_19508,N_19580);
and U19753 (N_19753,N_19515,N_19482);
nor U19754 (N_19754,N_19401,N_19455);
nand U19755 (N_19755,N_19544,N_19434);
and U19756 (N_19756,N_19598,N_19560);
or U19757 (N_19757,N_19486,N_19473);
nand U19758 (N_19758,N_19539,N_19585);
nand U19759 (N_19759,N_19537,N_19578);
nor U19760 (N_19760,N_19401,N_19539);
nand U19761 (N_19761,N_19498,N_19515);
and U19762 (N_19762,N_19456,N_19434);
nor U19763 (N_19763,N_19530,N_19430);
nor U19764 (N_19764,N_19531,N_19430);
xnor U19765 (N_19765,N_19447,N_19469);
nand U19766 (N_19766,N_19434,N_19492);
xor U19767 (N_19767,N_19532,N_19523);
and U19768 (N_19768,N_19459,N_19427);
or U19769 (N_19769,N_19510,N_19472);
or U19770 (N_19770,N_19558,N_19417);
nand U19771 (N_19771,N_19402,N_19567);
xnor U19772 (N_19772,N_19465,N_19510);
or U19773 (N_19773,N_19500,N_19418);
or U19774 (N_19774,N_19444,N_19513);
nor U19775 (N_19775,N_19439,N_19406);
and U19776 (N_19776,N_19571,N_19464);
nor U19777 (N_19777,N_19503,N_19516);
or U19778 (N_19778,N_19589,N_19471);
nand U19779 (N_19779,N_19582,N_19481);
nor U19780 (N_19780,N_19535,N_19532);
xor U19781 (N_19781,N_19476,N_19415);
nand U19782 (N_19782,N_19576,N_19412);
nand U19783 (N_19783,N_19411,N_19504);
xnor U19784 (N_19784,N_19504,N_19576);
or U19785 (N_19785,N_19482,N_19442);
nand U19786 (N_19786,N_19494,N_19553);
and U19787 (N_19787,N_19562,N_19482);
nor U19788 (N_19788,N_19506,N_19417);
nor U19789 (N_19789,N_19409,N_19580);
nor U19790 (N_19790,N_19563,N_19535);
or U19791 (N_19791,N_19402,N_19520);
and U19792 (N_19792,N_19517,N_19584);
nand U19793 (N_19793,N_19475,N_19513);
nand U19794 (N_19794,N_19547,N_19554);
nor U19795 (N_19795,N_19448,N_19463);
or U19796 (N_19796,N_19537,N_19582);
nor U19797 (N_19797,N_19480,N_19553);
or U19798 (N_19798,N_19412,N_19526);
or U19799 (N_19799,N_19529,N_19509);
or U19800 (N_19800,N_19626,N_19604);
and U19801 (N_19801,N_19692,N_19624);
nand U19802 (N_19802,N_19677,N_19690);
xnor U19803 (N_19803,N_19769,N_19618);
or U19804 (N_19804,N_19651,N_19659);
xnor U19805 (N_19805,N_19641,N_19794);
nand U19806 (N_19806,N_19603,N_19731);
nand U19807 (N_19807,N_19774,N_19797);
xor U19808 (N_19808,N_19613,N_19766);
xnor U19809 (N_19809,N_19668,N_19729);
and U19810 (N_19810,N_19699,N_19790);
nor U19811 (N_19811,N_19634,N_19669);
nor U19812 (N_19812,N_19687,N_19702);
or U19813 (N_19813,N_19619,N_19667);
or U19814 (N_19814,N_19673,N_19671);
or U19815 (N_19815,N_19640,N_19761);
xor U19816 (N_19816,N_19765,N_19780);
xnor U19817 (N_19817,N_19726,N_19647);
or U19818 (N_19818,N_19704,N_19628);
xor U19819 (N_19819,N_19674,N_19743);
and U19820 (N_19820,N_19703,N_19611);
nor U19821 (N_19821,N_19662,N_19723);
and U19822 (N_19822,N_19749,N_19772);
nand U19823 (N_19823,N_19676,N_19771);
or U19824 (N_19824,N_19754,N_19784);
or U19825 (N_19825,N_19632,N_19712);
nand U19826 (N_19826,N_19757,N_19742);
and U19827 (N_19827,N_19645,N_19722);
nor U19828 (N_19828,N_19721,N_19635);
xnor U19829 (N_19829,N_19747,N_19796);
nand U19830 (N_19830,N_19751,N_19753);
or U19831 (N_19831,N_19724,N_19629);
or U19832 (N_19832,N_19636,N_19652);
nor U19833 (N_19833,N_19750,N_19606);
and U19834 (N_19834,N_19657,N_19748);
and U19835 (N_19835,N_19786,N_19709);
or U19836 (N_19836,N_19762,N_19678);
nand U19837 (N_19837,N_19773,N_19646);
and U19838 (N_19838,N_19720,N_19658);
and U19839 (N_19839,N_19727,N_19745);
and U19840 (N_19840,N_19679,N_19685);
nor U19841 (N_19841,N_19715,N_19654);
or U19842 (N_19842,N_19610,N_19737);
nor U19843 (N_19843,N_19785,N_19684);
xor U19844 (N_19844,N_19707,N_19608);
xor U19845 (N_19845,N_19601,N_19648);
or U19846 (N_19846,N_19609,N_19710);
nor U19847 (N_19847,N_19717,N_19755);
nand U19848 (N_19848,N_19602,N_19615);
or U19849 (N_19849,N_19728,N_19756);
or U19850 (N_19850,N_19730,N_19693);
nor U19851 (N_19851,N_19622,N_19621);
or U19852 (N_19852,N_19713,N_19695);
xnor U19853 (N_19853,N_19741,N_19653);
or U19854 (N_19854,N_19660,N_19793);
and U19855 (N_19855,N_19643,N_19655);
nor U19856 (N_19856,N_19799,N_19700);
xor U19857 (N_19857,N_19770,N_19639);
xnor U19858 (N_19858,N_19767,N_19688);
or U19859 (N_19859,N_19694,N_19711);
or U19860 (N_19860,N_19738,N_19663);
nor U19861 (N_19861,N_19752,N_19649);
nand U19862 (N_19862,N_19672,N_19779);
or U19863 (N_19863,N_19735,N_19682);
nor U19864 (N_19864,N_19607,N_19787);
nor U19865 (N_19865,N_19656,N_19791);
and U19866 (N_19866,N_19782,N_19675);
xnor U19867 (N_19867,N_19605,N_19759);
xnor U19868 (N_19868,N_19758,N_19666);
nand U19869 (N_19869,N_19705,N_19792);
nand U19870 (N_19870,N_19620,N_19716);
xnor U19871 (N_19871,N_19616,N_19665);
or U19872 (N_19872,N_19733,N_19701);
nand U19873 (N_19873,N_19744,N_19642);
xor U19874 (N_19874,N_19617,N_19718);
nor U19875 (N_19875,N_19708,N_19625);
or U19876 (N_19876,N_19768,N_19706);
and U19877 (N_19877,N_19795,N_19630);
and U19878 (N_19878,N_19697,N_19740);
nor U19879 (N_19879,N_19736,N_19719);
or U19880 (N_19880,N_19789,N_19627);
and U19881 (N_19881,N_19781,N_19638);
or U19882 (N_19882,N_19764,N_19698);
and U19883 (N_19883,N_19691,N_19614);
and U19884 (N_19884,N_19637,N_19650);
and U19885 (N_19885,N_19777,N_19734);
and U19886 (N_19886,N_19623,N_19633);
nand U19887 (N_19887,N_19798,N_19696);
or U19888 (N_19888,N_19644,N_19681);
and U19889 (N_19889,N_19776,N_19661);
or U19890 (N_19890,N_19680,N_19686);
or U19891 (N_19891,N_19689,N_19670);
xor U19892 (N_19892,N_19725,N_19683);
nand U19893 (N_19893,N_19778,N_19746);
and U19894 (N_19894,N_19612,N_19732);
or U19895 (N_19895,N_19775,N_19783);
and U19896 (N_19896,N_19763,N_19760);
or U19897 (N_19897,N_19631,N_19600);
nor U19898 (N_19898,N_19664,N_19788);
and U19899 (N_19899,N_19714,N_19739);
or U19900 (N_19900,N_19708,N_19759);
or U19901 (N_19901,N_19608,N_19673);
or U19902 (N_19902,N_19715,N_19688);
and U19903 (N_19903,N_19799,N_19748);
and U19904 (N_19904,N_19740,N_19656);
nor U19905 (N_19905,N_19620,N_19724);
nor U19906 (N_19906,N_19708,N_19622);
and U19907 (N_19907,N_19785,N_19675);
nand U19908 (N_19908,N_19799,N_19643);
nand U19909 (N_19909,N_19611,N_19773);
xnor U19910 (N_19910,N_19702,N_19618);
nand U19911 (N_19911,N_19600,N_19787);
or U19912 (N_19912,N_19730,N_19637);
xnor U19913 (N_19913,N_19733,N_19718);
or U19914 (N_19914,N_19740,N_19653);
nor U19915 (N_19915,N_19638,N_19744);
nand U19916 (N_19916,N_19660,N_19636);
xor U19917 (N_19917,N_19679,N_19750);
nand U19918 (N_19918,N_19749,N_19626);
and U19919 (N_19919,N_19671,N_19759);
or U19920 (N_19920,N_19776,N_19754);
nor U19921 (N_19921,N_19680,N_19730);
or U19922 (N_19922,N_19762,N_19673);
nor U19923 (N_19923,N_19792,N_19796);
and U19924 (N_19924,N_19795,N_19690);
and U19925 (N_19925,N_19620,N_19692);
nand U19926 (N_19926,N_19673,N_19642);
and U19927 (N_19927,N_19663,N_19792);
nand U19928 (N_19928,N_19734,N_19743);
nand U19929 (N_19929,N_19707,N_19780);
and U19930 (N_19930,N_19658,N_19786);
xnor U19931 (N_19931,N_19747,N_19676);
or U19932 (N_19932,N_19763,N_19751);
xor U19933 (N_19933,N_19679,N_19717);
and U19934 (N_19934,N_19712,N_19638);
nand U19935 (N_19935,N_19665,N_19667);
or U19936 (N_19936,N_19696,N_19680);
or U19937 (N_19937,N_19678,N_19728);
xor U19938 (N_19938,N_19746,N_19638);
or U19939 (N_19939,N_19767,N_19603);
nand U19940 (N_19940,N_19788,N_19674);
and U19941 (N_19941,N_19740,N_19605);
nor U19942 (N_19942,N_19787,N_19739);
nor U19943 (N_19943,N_19741,N_19680);
or U19944 (N_19944,N_19608,N_19737);
xnor U19945 (N_19945,N_19702,N_19616);
and U19946 (N_19946,N_19725,N_19637);
nor U19947 (N_19947,N_19643,N_19779);
nand U19948 (N_19948,N_19777,N_19749);
nor U19949 (N_19949,N_19609,N_19698);
or U19950 (N_19950,N_19617,N_19702);
or U19951 (N_19951,N_19721,N_19772);
nor U19952 (N_19952,N_19603,N_19699);
xnor U19953 (N_19953,N_19603,N_19601);
and U19954 (N_19954,N_19708,N_19716);
xnor U19955 (N_19955,N_19745,N_19612);
nor U19956 (N_19956,N_19771,N_19668);
xnor U19957 (N_19957,N_19764,N_19731);
or U19958 (N_19958,N_19634,N_19632);
xor U19959 (N_19959,N_19617,N_19716);
nand U19960 (N_19960,N_19654,N_19748);
and U19961 (N_19961,N_19729,N_19791);
nand U19962 (N_19962,N_19739,N_19704);
and U19963 (N_19963,N_19794,N_19796);
or U19964 (N_19964,N_19724,N_19601);
xor U19965 (N_19965,N_19776,N_19642);
or U19966 (N_19966,N_19642,N_19721);
xnor U19967 (N_19967,N_19732,N_19651);
or U19968 (N_19968,N_19612,N_19713);
or U19969 (N_19969,N_19754,N_19655);
xor U19970 (N_19970,N_19740,N_19718);
nor U19971 (N_19971,N_19637,N_19700);
nor U19972 (N_19972,N_19668,N_19749);
and U19973 (N_19973,N_19606,N_19621);
xor U19974 (N_19974,N_19685,N_19648);
nand U19975 (N_19975,N_19782,N_19681);
nand U19976 (N_19976,N_19655,N_19743);
and U19977 (N_19977,N_19707,N_19729);
and U19978 (N_19978,N_19689,N_19770);
or U19979 (N_19979,N_19658,N_19604);
or U19980 (N_19980,N_19622,N_19606);
nor U19981 (N_19981,N_19673,N_19614);
nor U19982 (N_19982,N_19742,N_19612);
and U19983 (N_19983,N_19675,N_19715);
and U19984 (N_19984,N_19696,N_19740);
or U19985 (N_19985,N_19773,N_19632);
or U19986 (N_19986,N_19696,N_19613);
or U19987 (N_19987,N_19789,N_19639);
nor U19988 (N_19988,N_19738,N_19661);
nor U19989 (N_19989,N_19747,N_19732);
nor U19990 (N_19990,N_19695,N_19634);
nor U19991 (N_19991,N_19613,N_19647);
and U19992 (N_19992,N_19770,N_19698);
or U19993 (N_19993,N_19796,N_19726);
or U19994 (N_19994,N_19733,N_19601);
or U19995 (N_19995,N_19609,N_19783);
or U19996 (N_19996,N_19736,N_19700);
nor U19997 (N_19997,N_19722,N_19690);
or U19998 (N_19998,N_19617,N_19690);
xor U19999 (N_19999,N_19622,N_19635);
and U20000 (N_20000,N_19935,N_19906);
nor U20001 (N_20001,N_19857,N_19975);
xor U20002 (N_20002,N_19830,N_19923);
nor U20003 (N_20003,N_19957,N_19868);
or U20004 (N_20004,N_19867,N_19989);
or U20005 (N_20005,N_19805,N_19880);
or U20006 (N_20006,N_19921,N_19933);
xor U20007 (N_20007,N_19803,N_19855);
xnor U20008 (N_20008,N_19992,N_19887);
and U20009 (N_20009,N_19823,N_19854);
or U20010 (N_20010,N_19926,N_19990);
or U20011 (N_20011,N_19902,N_19888);
nor U20012 (N_20012,N_19816,N_19968);
nor U20013 (N_20013,N_19988,N_19985);
nand U20014 (N_20014,N_19813,N_19832);
nand U20015 (N_20015,N_19872,N_19905);
and U20016 (N_20016,N_19877,N_19914);
and U20017 (N_20017,N_19860,N_19939);
and U20018 (N_20018,N_19808,N_19831);
xnor U20019 (N_20019,N_19833,N_19814);
or U20020 (N_20020,N_19847,N_19845);
nand U20021 (N_20021,N_19954,N_19922);
nand U20022 (N_20022,N_19991,N_19849);
nor U20023 (N_20023,N_19865,N_19851);
and U20024 (N_20024,N_19873,N_19956);
xor U20025 (N_20025,N_19882,N_19971);
nand U20026 (N_20026,N_19866,N_19800);
or U20027 (N_20027,N_19947,N_19965);
nand U20028 (N_20028,N_19843,N_19815);
and U20029 (N_20029,N_19915,N_19835);
nor U20030 (N_20030,N_19879,N_19824);
nand U20031 (N_20031,N_19959,N_19986);
nor U20032 (N_20032,N_19981,N_19856);
xor U20033 (N_20033,N_19987,N_19810);
nor U20034 (N_20034,N_19972,N_19948);
xor U20035 (N_20035,N_19838,N_19936);
xor U20036 (N_20036,N_19951,N_19916);
or U20037 (N_20037,N_19966,N_19974);
nand U20038 (N_20038,N_19871,N_19897);
xnor U20039 (N_20039,N_19821,N_19932);
or U20040 (N_20040,N_19837,N_19853);
nand U20041 (N_20041,N_19862,N_19907);
nor U20042 (N_20042,N_19804,N_19979);
xor U20043 (N_20043,N_19836,N_19913);
or U20044 (N_20044,N_19812,N_19998);
nor U20045 (N_20045,N_19931,N_19929);
and U20046 (N_20046,N_19994,N_19938);
or U20047 (N_20047,N_19983,N_19909);
xnor U20048 (N_20048,N_19946,N_19852);
nand U20049 (N_20049,N_19917,N_19941);
nand U20050 (N_20050,N_19863,N_19927);
xnor U20051 (N_20051,N_19900,N_19886);
and U20052 (N_20052,N_19898,N_19961);
and U20053 (N_20053,N_19876,N_19858);
or U20054 (N_20054,N_19892,N_19894);
nor U20055 (N_20055,N_19952,N_19910);
nand U20056 (N_20056,N_19955,N_19924);
nand U20057 (N_20057,N_19825,N_19953);
or U20058 (N_20058,N_19885,N_19993);
nor U20059 (N_20059,N_19976,N_19943);
or U20060 (N_20060,N_19802,N_19844);
xor U20061 (N_20061,N_19817,N_19807);
nor U20062 (N_20062,N_19890,N_19970);
xnor U20063 (N_20063,N_19940,N_19945);
nor U20064 (N_20064,N_19818,N_19973);
and U20065 (N_20065,N_19884,N_19811);
nand U20066 (N_20066,N_19999,N_19828);
nor U20067 (N_20067,N_19958,N_19942);
nand U20068 (N_20068,N_19896,N_19997);
xor U20069 (N_20069,N_19978,N_19895);
and U20070 (N_20070,N_19903,N_19904);
and U20071 (N_20071,N_19870,N_19826);
xor U20072 (N_20072,N_19846,N_19850);
nor U20073 (N_20073,N_19864,N_19801);
nand U20074 (N_20074,N_19820,N_19967);
nand U20075 (N_20075,N_19911,N_19893);
or U20076 (N_20076,N_19963,N_19859);
or U20077 (N_20077,N_19878,N_19996);
or U20078 (N_20078,N_19901,N_19875);
or U20079 (N_20079,N_19984,N_19937);
or U20080 (N_20080,N_19995,N_19918);
xor U20081 (N_20081,N_19930,N_19977);
nand U20082 (N_20082,N_19819,N_19934);
xnor U20083 (N_20083,N_19908,N_19834);
nand U20084 (N_20084,N_19925,N_19881);
xor U20085 (N_20085,N_19822,N_19861);
nor U20086 (N_20086,N_19806,N_19827);
xnor U20087 (N_20087,N_19928,N_19891);
or U20088 (N_20088,N_19809,N_19839);
and U20089 (N_20089,N_19969,N_19848);
and U20090 (N_20090,N_19950,N_19841);
nand U20091 (N_20091,N_19883,N_19912);
or U20092 (N_20092,N_19874,N_19829);
nor U20093 (N_20093,N_19960,N_19962);
xor U20094 (N_20094,N_19964,N_19949);
nor U20095 (N_20095,N_19944,N_19919);
nand U20096 (N_20096,N_19920,N_19889);
and U20097 (N_20097,N_19980,N_19899);
and U20098 (N_20098,N_19869,N_19842);
xor U20099 (N_20099,N_19982,N_19840);
and U20100 (N_20100,N_19883,N_19969);
and U20101 (N_20101,N_19927,N_19942);
or U20102 (N_20102,N_19828,N_19884);
xor U20103 (N_20103,N_19965,N_19807);
nor U20104 (N_20104,N_19998,N_19972);
nand U20105 (N_20105,N_19804,N_19953);
nor U20106 (N_20106,N_19945,N_19818);
or U20107 (N_20107,N_19870,N_19966);
nand U20108 (N_20108,N_19868,N_19810);
xor U20109 (N_20109,N_19848,N_19837);
or U20110 (N_20110,N_19911,N_19851);
or U20111 (N_20111,N_19816,N_19864);
nor U20112 (N_20112,N_19920,N_19814);
nor U20113 (N_20113,N_19826,N_19992);
and U20114 (N_20114,N_19843,N_19907);
or U20115 (N_20115,N_19838,N_19962);
nand U20116 (N_20116,N_19952,N_19827);
and U20117 (N_20117,N_19831,N_19825);
xnor U20118 (N_20118,N_19843,N_19847);
and U20119 (N_20119,N_19954,N_19820);
xor U20120 (N_20120,N_19802,N_19993);
or U20121 (N_20121,N_19886,N_19909);
or U20122 (N_20122,N_19991,N_19857);
and U20123 (N_20123,N_19978,N_19832);
nand U20124 (N_20124,N_19930,N_19931);
and U20125 (N_20125,N_19999,N_19815);
and U20126 (N_20126,N_19837,N_19804);
and U20127 (N_20127,N_19982,N_19943);
or U20128 (N_20128,N_19806,N_19988);
or U20129 (N_20129,N_19834,N_19825);
xnor U20130 (N_20130,N_19980,N_19946);
xor U20131 (N_20131,N_19864,N_19813);
xor U20132 (N_20132,N_19839,N_19873);
nor U20133 (N_20133,N_19961,N_19844);
or U20134 (N_20134,N_19954,N_19805);
xor U20135 (N_20135,N_19922,N_19830);
nand U20136 (N_20136,N_19848,N_19991);
and U20137 (N_20137,N_19812,N_19969);
and U20138 (N_20138,N_19847,N_19892);
nand U20139 (N_20139,N_19931,N_19853);
nand U20140 (N_20140,N_19974,N_19864);
xnor U20141 (N_20141,N_19951,N_19810);
or U20142 (N_20142,N_19979,N_19948);
nor U20143 (N_20143,N_19998,N_19965);
and U20144 (N_20144,N_19833,N_19970);
nor U20145 (N_20145,N_19988,N_19956);
and U20146 (N_20146,N_19831,N_19973);
xor U20147 (N_20147,N_19811,N_19924);
and U20148 (N_20148,N_19805,N_19964);
xor U20149 (N_20149,N_19949,N_19820);
and U20150 (N_20150,N_19866,N_19942);
or U20151 (N_20151,N_19807,N_19835);
nor U20152 (N_20152,N_19962,N_19963);
nor U20153 (N_20153,N_19933,N_19850);
nand U20154 (N_20154,N_19908,N_19810);
and U20155 (N_20155,N_19989,N_19934);
nor U20156 (N_20156,N_19961,N_19871);
nand U20157 (N_20157,N_19955,N_19969);
xnor U20158 (N_20158,N_19852,N_19866);
nand U20159 (N_20159,N_19877,N_19913);
or U20160 (N_20160,N_19885,N_19871);
nor U20161 (N_20161,N_19997,N_19915);
xnor U20162 (N_20162,N_19894,N_19879);
and U20163 (N_20163,N_19876,N_19847);
and U20164 (N_20164,N_19897,N_19842);
nor U20165 (N_20165,N_19942,N_19840);
nand U20166 (N_20166,N_19997,N_19812);
xor U20167 (N_20167,N_19997,N_19830);
xnor U20168 (N_20168,N_19890,N_19860);
or U20169 (N_20169,N_19954,N_19936);
xor U20170 (N_20170,N_19808,N_19839);
nor U20171 (N_20171,N_19994,N_19953);
nor U20172 (N_20172,N_19919,N_19809);
and U20173 (N_20173,N_19800,N_19956);
or U20174 (N_20174,N_19942,N_19929);
nand U20175 (N_20175,N_19956,N_19870);
nor U20176 (N_20176,N_19841,N_19887);
and U20177 (N_20177,N_19839,N_19902);
and U20178 (N_20178,N_19830,N_19880);
or U20179 (N_20179,N_19877,N_19936);
nand U20180 (N_20180,N_19905,N_19843);
xnor U20181 (N_20181,N_19818,N_19908);
and U20182 (N_20182,N_19878,N_19971);
or U20183 (N_20183,N_19909,N_19849);
xnor U20184 (N_20184,N_19818,N_19850);
and U20185 (N_20185,N_19963,N_19951);
nor U20186 (N_20186,N_19902,N_19816);
nand U20187 (N_20187,N_19841,N_19920);
and U20188 (N_20188,N_19904,N_19879);
nor U20189 (N_20189,N_19820,N_19854);
and U20190 (N_20190,N_19884,N_19912);
nor U20191 (N_20191,N_19977,N_19983);
and U20192 (N_20192,N_19897,N_19960);
nand U20193 (N_20193,N_19923,N_19828);
xnor U20194 (N_20194,N_19841,N_19952);
and U20195 (N_20195,N_19931,N_19997);
and U20196 (N_20196,N_19837,N_19974);
nand U20197 (N_20197,N_19860,N_19842);
or U20198 (N_20198,N_19801,N_19963);
nor U20199 (N_20199,N_19917,N_19832);
xnor U20200 (N_20200,N_20138,N_20006);
nand U20201 (N_20201,N_20040,N_20008);
xor U20202 (N_20202,N_20096,N_20124);
nand U20203 (N_20203,N_20133,N_20001);
xnor U20204 (N_20204,N_20086,N_20043);
nor U20205 (N_20205,N_20084,N_20112);
xor U20206 (N_20206,N_20173,N_20019);
xnor U20207 (N_20207,N_20120,N_20016);
or U20208 (N_20208,N_20015,N_20183);
and U20209 (N_20209,N_20064,N_20146);
or U20210 (N_20210,N_20017,N_20193);
xnor U20211 (N_20211,N_20185,N_20115);
or U20212 (N_20212,N_20102,N_20167);
and U20213 (N_20213,N_20057,N_20164);
xor U20214 (N_20214,N_20192,N_20059);
nor U20215 (N_20215,N_20093,N_20003);
and U20216 (N_20216,N_20111,N_20116);
xor U20217 (N_20217,N_20094,N_20041);
nor U20218 (N_20218,N_20092,N_20139);
or U20219 (N_20219,N_20065,N_20149);
nor U20220 (N_20220,N_20104,N_20107);
nand U20221 (N_20221,N_20049,N_20091);
or U20222 (N_20222,N_20020,N_20159);
or U20223 (N_20223,N_20103,N_20044);
xnor U20224 (N_20224,N_20089,N_20136);
xnor U20225 (N_20225,N_20154,N_20007);
xnor U20226 (N_20226,N_20031,N_20171);
nor U20227 (N_20227,N_20068,N_20026);
nor U20228 (N_20228,N_20148,N_20128);
or U20229 (N_20229,N_20069,N_20151);
nand U20230 (N_20230,N_20126,N_20119);
nand U20231 (N_20231,N_20052,N_20085);
nand U20232 (N_20232,N_20090,N_20072);
and U20233 (N_20233,N_20143,N_20176);
nor U20234 (N_20234,N_20197,N_20125);
nand U20235 (N_20235,N_20046,N_20060);
nor U20236 (N_20236,N_20177,N_20123);
nand U20237 (N_20237,N_20131,N_20108);
and U20238 (N_20238,N_20137,N_20056);
nor U20239 (N_20239,N_20121,N_20127);
nand U20240 (N_20240,N_20109,N_20032);
and U20241 (N_20241,N_20035,N_20191);
nand U20242 (N_20242,N_20190,N_20074);
nor U20243 (N_20243,N_20101,N_20142);
nand U20244 (N_20244,N_20058,N_20073);
xor U20245 (N_20245,N_20163,N_20135);
or U20246 (N_20246,N_20028,N_20180);
nand U20247 (N_20247,N_20172,N_20005);
and U20248 (N_20248,N_20000,N_20002);
nor U20249 (N_20249,N_20100,N_20134);
nand U20250 (N_20250,N_20118,N_20048);
and U20251 (N_20251,N_20010,N_20029);
nor U20252 (N_20252,N_20114,N_20013);
and U20253 (N_20253,N_20023,N_20199);
or U20254 (N_20254,N_20014,N_20037);
nor U20255 (N_20255,N_20152,N_20082);
nand U20256 (N_20256,N_20165,N_20174);
nand U20257 (N_20257,N_20027,N_20033);
or U20258 (N_20258,N_20099,N_20066);
and U20259 (N_20259,N_20050,N_20051);
or U20260 (N_20260,N_20181,N_20188);
nor U20261 (N_20261,N_20187,N_20144);
nand U20262 (N_20262,N_20129,N_20067);
xor U20263 (N_20263,N_20036,N_20018);
or U20264 (N_20264,N_20153,N_20157);
and U20265 (N_20265,N_20009,N_20087);
xor U20266 (N_20266,N_20160,N_20076);
nor U20267 (N_20267,N_20184,N_20156);
and U20268 (N_20268,N_20178,N_20169);
and U20269 (N_20269,N_20042,N_20055);
or U20270 (N_20270,N_20130,N_20158);
or U20271 (N_20271,N_20147,N_20083);
xor U20272 (N_20272,N_20150,N_20095);
and U20273 (N_20273,N_20011,N_20182);
and U20274 (N_20274,N_20038,N_20024);
nor U20275 (N_20275,N_20141,N_20106);
or U20276 (N_20276,N_20166,N_20021);
nand U20277 (N_20277,N_20195,N_20053);
xnor U20278 (N_20278,N_20077,N_20168);
and U20279 (N_20279,N_20054,N_20022);
and U20280 (N_20280,N_20097,N_20063);
or U20281 (N_20281,N_20132,N_20079);
xor U20282 (N_20282,N_20161,N_20145);
or U20283 (N_20283,N_20140,N_20105);
or U20284 (N_20284,N_20175,N_20162);
or U20285 (N_20285,N_20088,N_20070);
nand U20286 (N_20286,N_20061,N_20194);
nand U20287 (N_20287,N_20186,N_20189);
nor U20288 (N_20288,N_20117,N_20080);
or U20289 (N_20289,N_20030,N_20062);
nor U20290 (N_20290,N_20110,N_20196);
xor U20291 (N_20291,N_20045,N_20198);
and U20292 (N_20292,N_20179,N_20075);
or U20293 (N_20293,N_20004,N_20071);
xor U20294 (N_20294,N_20025,N_20034);
xnor U20295 (N_20295,N_20098,N_20113);
nor U20296 (N_20296,N_20081,N_20078);
xor U20297 (N_20297,N_20122,N_20047);
or U20298 (N_20298,N_20155,N_20170);
nor U20299 (N_20299,N_20039,N_20012);
xnor U20300 (N_20300,N_20083,N_20079);
or U20301 (N_20301,N_20181,N_20034);
xor U20302 (N_20302,N_20035,N_20143);
xnor U20303 (N_20303,N_20080,N_20111);
or U20304 (N_20304,N_20034,N_20050);
nor U20305 (N_20305,N_20147,N_20148);
or U20306 (N_20306,N_20105,N_20025);
or U20307 (N_20307,N_20002,N_20187);
xor U20308 (N_20308,N_20004,N_20066);
nor U20309 (N_20309,N_20049,N_20166);
and U20310 (N_20310,N_20083,N_20137);
nor U20311 (N_20311,N_20146,N_20109);
and U20312 (N_20312,N_20052,N_20082);
and U20313 (N_20313,N_20137,N_20030);
xnor U20314 (N_20314,N_20047,N_20194);
xnor U20315 (N_20315,N_20055,N_20040);
xor U20316 (N_20316,N_20063,N_20033);
nor U20317 (N_20317,N_20165,N_20079);
or U20318 (N_20318,N_20110,N_20031);
and U20319 (N_20319,N_20140,N_20121);
xnor U20320 (N_20320,N_20149,N_20139);
or U20321 (N_20321,N_20020,N_20069);
xnor U20322 (N_20322,N_20179,N_20116);
or U20323 (N_20323,N_20049,N_20131);
xnor U20324 (N_20324,N_20107,N_20113);
and U20325 (N_20325,N_20051,N_20039);
xor U20326 (N_20326,N_20167,N_20060);
xnor U20327 (N_20327,N_20053,N_20045);
xnor U20328 (N_20328,N_20012,N_20134);
and U20329 (N_20329,N_20097,N_20153);
or U20330 (N_20330,N_20186,N_20195);
nand U20331 (N_20331,N_20038,N_20061);
nor U20332 (N_20332,N_20067,N_20136);
xor U20333 (N_20333,N_20159,N_20082);
xor U20334 (N_20334,N_20114,N_20161);
or U20335 (N_20335,N_20055,N_20152);
nor U20336 (N_20336,N_20147,N_20160);
or U20337 (N_20337,N_20052,N_20124);
xnor U20338 (N_20338,N_20187,N_20193);
nand U20339 (N_20339,N_20043,N_20011);
or U20340 (N_20340,N_20065,N_20026);
xor U20341 (N_20341,N_20149,N_20047);
xor U20342 (N_20342,N_20149,N_20173);
nor U20343 (N_20343,N_20051,N_20066);
and U20344 (N_20344,N_20164,N_20126);
and U20345 (N_20345,N_20104,N_20083);
and U20346 (N_20346,N_20125,N_20185);
and U20347 (N_20347,N_20087,N_20165);
and U20348 (N_20348,N_20069,N_20169);
nand U20349 (N_20349,N_20026,N_20105);
nor U20350 (N_20350,N_20142,N_20028);
or U20351 (N_20351,N_20149,N_20089);
xor U20352 (N_20352,N_20034,N_20021);
xnor U20353 (N_20353,N_20112,N_20024);
or U20354 (N_20354,N_20096,N_20031);
or U20355 (N_20355,N_20193,N_20005);
nand U20356 (N_20356,N_20037,N_20173);
xnor U20357 (N_20357,N_20053,N_20072);
nand U20358 (N_20358,N_20188,N_20197);
and U20359 (N_20359,N_20069,N_20083);
nor U20360 (N_20360,N_20127,N_20178);
nor U20361 (N_20361,N_20182,N_20101);
or U20362 (N_20362,N_20092,N_20077);
nand U20363 (N_20363,N_20111,N_20130);
nand U20364 (N_20364,N_20164,N_20071);
nor U20365 (N_20365,N_20037,N_20131);
and U20366 (N_20366,N_20052,N_20055);
nor U20367 (N_20367,N_20178,N_20161);
nor U20368 (N_20368,N_20111,N_20051);
nand U20369 (N_20369,N_20091,N_20190);
nand U20370 (N_20370,N_20093,N_20005);
or U20371 (N_20371,N_20057,N_20073);
or U20372 (N_20372,N_20076,N_20173);
xor U20373 (N_20373,N_20059,N_20136);
and U20374 (N_20374,N_20000,N_20182);
and U20375 (N_20375,N_20169,N_20152);
nand U20376 (N_20376,N_20097,N_20103);
and U20377 (N_20377,N_20157,N_20166);
nand U20378 (N_20378,N_20146,N_20178);
nor U20379 (N_20379,N_20026,N_20014);
nand U20380 (N_20380,N_20144,N_20082);
or U20381 (N_20381,N_20140,N_20149);
xor U20382 (N_20382,N_20012,N_20148);
nand U20383 (N_20383,N_20083,N_20100);
nand U20384 (N_20384,N_20101,N_20029);
and U20385 (N_20385,N_20022,N_20051);
nand U20386 (N_20386,N_20120,N_20191);
and U20387 (N_20387,N_20163,N_20081);
xor U20388 (N_20388,N_20133,N_20152);
nor U20389 (N_20389,N_20162,N_20081);
nor U20390 (N_20390,N_20188,N_20021);
nand U20391 (N_20391,N_20000,N_20012);
or U20392 (N_20392,N_20170,N_20147);
nor U20393 (N_20393,N_20154,N_20192);
and U20394 (N_20394,N_20145,N_20125);
and U20395 (N_20395,N_20178,N_20198);
nand U20396 (N_20396,N_20006,N_20039);
nand U20397 (N_20397,N_20070,N_20187);
and U20398 (N_20398,N_20069,N_20167);
nand U20399 (N_20399,N_20051,N_20155);
nand U20400 (N_20400,N_20350,N_20245);
xor U20401 (N_20401,N_20237,N_20325);
or U20402 (N_20402,N_20234,N_20338);
or U20403 (N_20403,N_20218,N_20215);
xnor U20404 (N_20404,N_20359,N_20375);
nor U20405 (N_20405,N_20315,N_20392);
nor U20406 (N_20406,N_20390,N_20327);
and U20407 (N_20407,N_20381,N_20227);
and U20408 (N_20408,N_20323,N_20251);
and U20409 (N_20409,N_20382,N_20351);
xor U20410 (N_20410,N_20288,N_20280);
or U20411 (N_20411,N_20249,N_20371);
nor U20412 (N_20412,N_20352,N_20310);
xor U20413 (N_20413,N_20263,N_20387);
xnor U20414 (N_20414,N_20283,N_20341);
xnor U20415 (N_20415,N_20357,N_20274);
nand U20416 (N_20416,N_20331,N_20311);
and U20417 (N_20417,N_20329,N_20383);
nor U20418 (N_20418,N_20272,N_20342);
and U20419 (N_20419,N_20242,N_20368);
nor U20420 (N_20420,N_20236,N_20262);
nand U20421 (N_20421,N_20305,N_20285);
xnor U20422 (N_20422,N_20277,N_20303);
nor U20423 (N_20423,N_20235,N_20396);
nand U20424 (N_20424,N_20210,N_20354);
nor U20425 (N_20425,N_20365,N_20246);
nor U20426 (N_20426,N_20349,N_20393);
nor U20427 (N_20427,N_20363,N_20320);
and U20428 (N_20428,N_20355,N_20314);
nor U20429 (N_20429,N_20282,N_20265);
nand U20430 (N_20430,N_20222,N_20239);
xnor U20431 (N_20431,N_20366,N_20254);
or U20432 (N_20432,N_20250,N_20298);
and U20433 (N_20433,N_20394,N_20209);
or U20434 (N_20434,N_20356,N_20213);
xor U20435 (N_20435,N_20228,N_20370);
xnor U20436 (N_20436,N_20240,N_20291);
and U20437 (N_20437,N_20212,N_20289);
and U20438 (N_20438,N_20377,N_20308);
and U20439 (N_20439,N_20214,N_20221);
nand U20440 (N_20440,N_20337,N_20223);
xor U20441 (N_20441,N_20300,N_20296);
xor U20442 (N_20442,N_20276,N_20247);
nand U20443 (N_20443,N_20326,N_20322);
nand U20444 (N_20444,N_20248,N_20367);
xnor U20445 (N_20445,N_20225,N_20379);
nand U20446 (N_20446,N_20292,N_20302);
xor U20447 (N_20447,N_20253,N_20200);
nor U20448 (N_20448,N_20294,N_20226);
and U20449 (N_20449,N_20333,N_20264);
nand U20450 (N_20450,N_20312,N_20231);
nor U20451 (N_20451,N_20238,N_20330);
nand U20452 (N_20452,N_20309,N_20208);
and U20453 (N_20453,N_20270,N_20278);
nor U20454 (N_20454,N_20268,N_20203);
nor U20455 (N_20455,N_20336,N_20399);
nor U20456 (N_20456,N_20229,N_20324);
nor U20457 (N_20457,N_20230,N_20374);
xor U20458 (N_20458,N_20219,N_20241);
xor U20459 (N_20459,N_20206,N_20362);
nor U20460 (N_20460,N_20207,N_20252);
nor U20461 (N_20461,N_20339,N_20385);
or U20462 (N_20462,N_20319,N_20347);
or U20463 (N_20463,N_20232,N_20313);
nand U20464 (N_20464,N_20275,N_20321);
and U20465 (N_20465,N_20334,N_20266);
or U20466 (N_20466,N_20299,N_20345);
and U20467 (N_20467,N_20243,N_20233);
nand U20468 (N_20468,N_20217,N_20306);
or U20469 (N_20469,N_20343,N_20361);
nand U20470 (N_20470,N_20220,N_20360);
nor U20471 (N_20471,N_20358,N_20279);
nor U20472 (N_20472,N_20335,N_20373);
nand U20473 (N_20473,N_20369,N_20391);
and U20474 (N_20474,N_20293,N_20267);
or U20475 (N_20475,N_20332,N_20281);
or U20476 (N_20476,N_20372,N_20301);
and U20477 (N_20477,N_20348,N_20316);
and U20478 (N_20478,N_20304,N_20258);
xnor U20479 (N_20479,N_20201,N_20297);
and U20480 (N_20480,N_20286,N_20290);
xor U20481 (N_20481,N_20376,N_20216);
nand U20482 (N_20482,N_20397,N_20395);
and U20483 (N_20483,N_20259,N_20388);
nor U20484 (N_20484,N_20287,N_20255);
or U20485 (N_20485,N_20205,N_20204);
xor U20486 (N_20486,N_20340,N_20307);
and U20487 (N_20487,N_20284,N_20364);
xor U20488 (N_20488,N_20224,N_20328);
nor U20489 (N_20489,N_20261,N_20344);
nand U20490 (N_20490,N_20260,N_20398);
nand U20491 (N_20491,N_20244,N_20317);
nor U20492 (N_20492,N_20318,N_20257);
nor U20493 (N_20493,N_20295,N_20389);
xor U20494 (N_20494,N_20380,N_20386);
xnor U20495 (N_20495,N_20269,N_20384);
xor U20496 (N_20496,N_20211,N_20256);
nand U20497 (N_20497,N_20202,N_20353);
nand U20498 (N_20498,N_20346,N_20271);
xor U20499 (N_20499,N_20378,N_20273);
nand U20500 (N_20500,N_20341,N_20203);
nor U20501 (N_20501,N_20394,N_20298);
nand U20502 (N_20502,N_20384,N_20220);
nor U20503 (N_20503,N_20274,N_20292);
and U20504 (N_20504,N_20282,N_20237);
xnor U20505 (N_20505,N_20316,N_20295);
nand U20506 (N_20506,N_20258,N_20364);
nor U20507 (N_20507,N_20233,N_20346);
xor U20508 (N_20508,N_20285,N_20376);
and U20509 (N_20509,N_20341,N_20394);
xnor U20510 (N_20510,N_20375,N_20201);
and U20511 (N_20511,N_20342,N_20261);
and U20512 (N_20512,N_20354,N_20287);
and U20513 (N_20513,N_20304,N_20365);
nand U20514 (N_20514,N_20239,N_20384);
nor U20515 (N_20515,N_20389,N_20239);
nor U20516 (N_20516,N_20308,N_20289);
or U20517 (N_20517,N_20367,N_20290);
and U20518 (N_20518,N_20376,N_20343);
nor U20519 (N_20519,N_20322,N_20389);
nor U20520 (N_20520,N_20276,N_20353);
xnor U20521 (N_20521,N_20277,N_20278);
or U20522 (N_20522,N_20224,N_20388);
and U20523 (N_20523,N_20356,N_20247);
or U20524 (N_20524,N_20342,N_20243);
nor U20525 (N_20525,N_20276,N_20322);
nand U20526 (N_20526,N_20341,N_20236);
xnor U20527 (N_20527,N_20235,N_20228);
nor U20528 (N_20528,N_20339,N_20281);
xor U20529 (N_20529,N_20208,N_20374);
xor U20530 (N_20530,N_20359,N_20219);
nand U20531 (N_20531,N_20356,N_20385);
and U20532 (N_20532,N_20304,N_20299);
or U20533 (N_20533,N_20277,N_20334);
or U20534 (N_20534,N_20380,N_20232);
nand U20535 (N_20535,N_20291,N_20340);
nor U20536 (N_20536,N_20300,N_20262);
and U20537 (N_20537,N_20348,N_20333);
and U20538 (N_20538,N_20331,N_20359);
and U20539 (N_20539,N_20203,N_20361);
nand U20540 (N_20540,N_20263,N_20342);
or U20541 (N_20541,N_20391,N_20243);
and U20542 (N_20542,N_20252,N_20224);
xor U20543 (N_20543,N_20371,N_20328);
nor U20544 (N_20544,N_20308,N_20205);
nor U20545 (N_20545,N_20393,N_20223);
xor U20546 (N_20546,N_20251,N_20289);
and U20547 (N_20547,N_20359,N_20239);
nor U20548 (N_20548,N_20305,N_20364);
and U20549 (N_20549,N_20255,N_20254);
and U20550 (N_20550,N_20256,N_20277);
and U20551 (N_20551,N_20361,N_20229);
xnor U20552 (N_20552,N_20215,N_20344);
xor U20553 (N_20553,N_20373,N_20220);
nor U20554 (N_20554,N_20329,N_20357);
nand U20555 (N_20555,N_20394,N_20262);
nor U20556 (N_20556,N_20372,N_20204);
or U20557 (N_20557,N_20364,N_20224);
or U20558 (N_20558,N_20239,N_20380);
nand U20559 (N_20559,N_20268,N_20333);
nor U20560 (N_20560,N_20253,N_20391);
and U20561 (N_20561,N_20349,N_20398);
xor U20562 (N_20562,N_20240,N_20274);
nand U20563 (N_20563,N_20222,N_20229);
nor U20564 (N_20564,N_20390,N_20358);
and U20565 (N_20565,N_20255,N_20263);
or U20566 (N_20566,N_20230,N_20358);
nor U20567 (N_20567,N_20378,N_20242);
xor U20568 (N_20568,N_20210,N_20204);
or U20569 (N_20569,N_20208,N_20259);
nor U20570 (N_20570,N_20220,N_20280);
and U20571 (N_20571,N_20381,N_20325);
nor U20572 (N_20572,N_20308,N_20201);
nand U20573 (N_20573,N_20333,N_20272);
and U20574 (N_20574,N_20383,N_20315);
nor U20575 (N_20575,N_20319,N_20368);
or U20576 (N_20576,N_20351,N_20336);
or U20577 (N_20577,N_20225,N_20212);
nor U20578 (N_20578,N_20380,N_20238);
nand U20579 (N_20579,N_20284,N_20266);
or U20580 (N_20580,N_20227,N_20246);
nand U20581 (N_20581,N_20252,N_20320);
nand U20582 (N_20582,N_20255,N_20368);
and U20583 (N_20583,N_20306,N_20316);
nor U20584 (N_20584,N_20205,N_20257);
xor U20585 (N_20585,N_20336,N_20369);
or U20586 (N_20586,N_20340,N_20384);
xnor U20587 (N_20587,N_20333,N_20260);
nand U20588 (N_20588,N_20219,N_20334);
and U20589 (N_20589,N_20281,N_20344);
nand U20590 (N_20590,N_20347,N_20269);
xnor U20591 (N_20591,N_20394,N_20272);
xnor U20592 (N_20592,N_20292,N_20214);
and U20593 (N_20593,N_20257,N_20229);
nor U20594 (N_20594,N_20368,N_20313);
and U20595 (N_20595,N_20372,N_20290);
and U20596 (N_20596,N_20397,N_20234);
xnor U20597 (N_20597,N_20207,N_20213);
nor U20598 (N_20598,N_20229,N_20334);
or U20599 (N_20599,N_20239,N_20378);
nand U20600 (N_20600,N_20528,N_20498);
or U20601 (N_20601,N_20589,N_20440);
or U20602 (N_20602,N_20441,N_20514);
xor U20603 (N_20603,N_20468,N_20507);
xnor U20604 (N_20604,N_20411,N_20578);
nor U20605 (N_20605,N_20461,N_20499);
xor U20606 (N_20606,N_20410,N_20420);
nand U20607 (N_20607,N_20495,N_20492);
and U20608 (N_20608,N_20597,N_20558);
nand U20609 (N_20609,N_20529,N_20560);
and U20610 (N_20610,N_20573,N_20401);
xnor U20611 (N_20611,N_20442,N_20467);
or U20612 (N_20612,N_20548,N_20424);
or U20613 (N_20613,N_20419,N_20568);
and U20614 (N_20614,N_20474,N_20480);
and U20615 (N_20615,N_20425,N_20470);
nand U20616 (N_20616,N_20590,N_20544);
or U20617 (N_20617,N_20478,N_20554);
xor U20618 (N_20618,N_20562,N_20516);
nor U20619 (N_20619,N_20428,N_20417);
xor U20620 (N_20620,N_20519,N_20407);
nand U20621 (N_20621,N_20592,N_20489);
nor U20622 (N_20622,N_20587,N_20565);
or U20623 (N_20623,N_20582,N_20460);
nand U20624 (N_20624,N_20457,N_20575);
and U20625 (N_20625,N_20459,N_20473);
and U20626 (N_20626,N_20541,N_20415);
nand U20627 (N_20627,N_20563,N_20430);
and U20628 (N_20628,N_20534,N_20408);
nor U20629 (N_20629,N_20572,N_20483);
xnor U20630 (N_20630,N_20452,N_20577);
nand U20631 (N_20631,N_20433,N_20530);
nand U20632 (N_20632,N_20409,N_20463);
or U20633 (N_20633,N_20435,N_20551);
xor U20634 (N_20634,N_20559,N_20538);
nor U20635 (N_20635,N_20412,N_20508);
nand U20636 (N_20636,N_20593,N_20413);
nand U20637 (N_20637,N_20418,N_20518);
or U20638 (N_20638,N_20421,N_20448);
nor U20639 (N_20639,N_20509,N_20423);
xnor U20640 (N_20640,N_20591,N_20505);
nor U20641 (N_20641,N_20438,N_20451);
nand U20642 (N_20642,N_20579,N_20444);
nand U20643 (N_20643,N_20596,N_20556);
nor U20644 (N_20644,N_20501,N_20434);
nor U20645 (N_20645,N_20581,N_20496);
and U20646 (N_20646,N_20553,N_20404);
xor U20647 (N_20647,N_20570,N_20586);
xnor U20648 (N_20648,N_20585,N_20416);
nor U20649 (N_20649,N_20512,N_20406);
and U20650 (N_20650,N_20475,N_20422);
or U20651 (N_20651,N_20469,N_20595);
and U20652 (N_20652,N_20414,N_20598);
xnor U20653 (N_20653,N_20427,N_20439);
nor U20654 (N_20654,N_20531,N_20547);
xor U20655 (N_20655,N_20569,N_20555);
xor U20656 (N_20656,N_20511,N_20447);
and U20657 (N_20657,N_20462,N_20405);
nor U20658 (N_20658,N_20465,N_20520);
or U20659 (N_20659,N_20454,N_20536);
xor U20660 (N_20660,N_20477,N_20588);
nand U20661 (N_20661,N_20523,N_20481);
nor U20662 (N_20662,N_20456,N_20497);
nand U20663 (N_20663,N_20599,N_20561);
and U20664 (N_20664,N_20571,N_20432);
and U20665 (N_20665,N_20527,N_20491);
and U20666 (N_20666,N_20540,N_20539);
nor U20667 (N_20667,N_20521,N_20580);
or U20668 (N_20668,N_20466,N_20506);
nor U20669 (N_20669,N_20566,N_20594);
or U20670 (N_20670,N_20436,N_20524);
xor U20671 (N_20671,N_20537,N_20450);
nor U20672 (N_20672,N_20453,N_20486);
or U20673 (N_20673,N_20449,N_20535);
and U20674 (N_20674,N_20446,N_20471);
nand U20675 (N_20675,N_20458,N_20485);
or U20676 (N_20676,N_20567,N_20517);
xor U20677 (N_20677,N_20543,N_20484);
and U20678 (N_20678,N_20437,N_20546);
xor U20679 (N_20679,N_20488,N_20455);
nor U20680 (N_20680,N_20503,N_20574);
nor U20681 (N_20681,N_20482,N_20490);
xor U20682 (N_20682,N_20576,N_20443);
nor U20683 (N_20683,N_20525,N_20476);
xor U20684 (N_20684,N_20400,N_20504);
nor U20685 (N_20685,N_20494,N_20500);
xor U20686 (N_20686,N_20552,N_20510);
or U20687 (N_20687,N_20429,N_20584);
or U20688 (N_20688,N_20513,N_20533);
nand U20689 (N_20689,N_20402,N_20487);
nand U20690 (N_20690,N_20522,N_20564);
xnor U20691 (N_20691,N_20557,N_20549);
nand U20692 (N_20692,N_20583,N_20431);
or U20693 (N_20693,N_20532,N_20479);
xor U20694 (N_20694,N_20502,N_20464);
and U20695 (N_20695,N_20545,N_20403);
xor U20696 (N_20696,N_20515,N_20526);
xor U20697 (N_20697,N_20472,N_20445);
nand U20698 (N_20698,N_20542,N_20426);
nor U20699 (N_20699,N_20550,N_20493);
or U20700 (N_20700,N_20564,N_20545);
nand U20701 (N_20701,N_20465,N_20491);
nand U20702 (N_20702,N_20451,N_20453);
nand U20703 (N_20703,N_20580,N_20467);
xor U20704 (N_20704,N_20429,N_20442);
or U20705 (N_20705,N_20445,N_20469);
and U20706 (N_20706,N_20420,N_20530);
nor U20707 (N_20707,N_20410,N_20402);
nor U20708 (N_20708,N_20531,N_20417);
or U20709 (N_20709,N_20542,N_20473);
and U20710 (N_20710,N_20547,N_20439);
and U20711 (N_20711,N_20526,N_20431);
or U20712 (N_20712,N_20418,N_20535);
xnor U20713 (N_20713,N_20490,N_20509);
xnor U20714 (N_20714,N_20426,N_20582);
or U20715 (N_20715,N_20552,N_20537);
and U20716 (N_20716,N_20454,N_20537);
nand U20717 (N_20717,N_20564,N_20455);
and U20718 (N_20718,N_20466,N_20456);
nor U20719 (N_20719,N_20574,N_20411);
nor U20720 (N_20720,N_20404,N_20537);
xnor U20721 (N_20721,N_20481,N_20558);
or U20722 (N_20722,N_20595,N_20581);
nor U20723 (N_20723,N_20486,N_20438);
and U20724 (N_20724,N_20450,N_20598);
and U20725 (N_20725,N_20551,N_20493);
nor U20726 (N_20726,N_20454,N_20482);
or U20727 (N_20727,N_20554,N_20572);
nor U20728 (N_20728,N_20577,N_20439);
and U20729 (N_20729,N_20457,N_20562);
nor U20730 (N_20730,N_20489,N_20449);
nor U20731 (N_20731,N_20405,N_20593);
nor U20732 (N_20732,N_20484,N_20520);
nand U20733 (N_20733,N_20555,N_20451);
xnor U20734 (N_20734,N_20505,N_20436);
xor U20735 (N_20735,N_20518,N_20454);
and U20736 (N_20736,N_20543,N_20551);
nand U20737 (N_20737,N_20501,N_20513);
nand U20738 (N_20738,N_20539,N_20400);
or U20739 (N_20739,N_20569,N_20557);
xnor U20740 (N_20740,N_20435,N_20517);
and U20741 (N_20741,N_20526,N_20424);
or U20742 (N_20742,N_20565,N_20501);
xnor U20743 (N_20743,N_20409,N_20565);
nand U20744 (N_20744,N_20595,N_20478);
xnor U20745 (N_20745,N_20562,N_20509);
nand U20746 (N_20746,N_20471,N_20586);
or U20747 (N_20747,N_20498,N_20538);
or U20748 (N_20748,N_20476,N_20594);
xnor U20749 (N_20749,N_20584,N_20565);
and U20750 (N_20750,N_20516,N_20462);
xor U20751 (N_20751,N_20532,N_20570);
or U20752 (N_20752,N_20496,N_20464);
and U20753 (N_20753,N_20503,N_20445);
and U20754 (N_20754,N_20570,N_20410);
and U20755 (N_20755,N_20485,N_20540);
or U20756 (N_20756,N_20533,N_20545);
nor U20757 (N_20757,N_20475,N_20401);
nor U20758 (N_20758,N_20490,N_20413);
xor U20759 (N_20759,N_20569,N_20405);
xnor U20760 (N_20760,N_20505,N_20473);
or U20761 (N_20761,N_20565,N_20458);
nand U20762 (N_20762,N_20432,N_20492);
xor U20763 (N_20763,N_20549,N_20463);
nand U20764 (N_20764,N_20521,N_20458);
and U20765 (N_20765,N_20535,N_20444);
xnor U20766 (N_20766,N_20544,N_20534);
xor U20767 (N_20767,N_20469,N_20553);
and U20768 (N_20768,N_20408,N_20500);
xor U20769 (N_20769,N_20449,N_20406);
and U20770 (N_20770,N_20533,N_20409);
nor U20771 (N_20771,N_20516,N_20403);
xor U20772 (N_20772,N_20480,N_20500);
xor U20773 (N_20773,N_20412,N_20493);
and U20774 (N_20774,N_20585,N_20578);
or U20775 (N_20775,N_20581,N_20431);
nor U20776 (N_20776,N_20596,N_20511);
nand U20777 (N_20777,N_20465,N_20407);
nor U20778 (N_20778,N_20523,N_20448);
nand U20779 (N_20779,N_20557,N_20548);
xor U20780 (N_20780,N_20432,N_20480);
xnor U20781 (N_20781,N_20465,N_20413);
xnor U20782 (N_20782,N_20594,N_20420);
nand U20783 (N_20783,N_20401,N_20557);
nand U20784 (N_20784,N_20535,N_20553);
nand U20785 (N_20785,N_20425,N_20562);
nor U20786 (N_20786,N_20485,N_20581);
or U20787 (N_20787,N_20401,N_20511);
nand U20788 (N_20788,N_20536,N_20540);
xnor U20789 (N_20789,N_20574,N_20576);
and U20790 (N_20790,N_20487,N_20528);
xor U20791 (N_20791,N_20557,N_20463);
xnor U20792 (N_20792,N_20553,N_20530);
nor U20793 (N_20793,N_20535,N_20457);
xor U20794 (N_20794,N_20417,N_20485);
nor U20795 (N_20795,N_20561,N_20475);
xor U20796 (N_20796,N_20498,N_20419);
nor U20797 (N_20797,N_20500,N_20578);
nand U20798 (N_20798,N_20550,N_20522);
and U20799 (N_20799,N_20557,N_20547);
or U20800 (N_20800,N_20754,N_20657);
xnor U20801 (N_20801,N_20646,N_20666);
and U20802 (N_20802,N_20718,N_20693);
and U20803 (N_20803,N_20634,N_20680);
nand U20804 (N_20804,N_20639,N_20720);
nor U20805 (N_20805,N_20791,N_20661);
nand U20806 (N_20806,N_20644,N_20643);
or U20807 (N_20807,N_20678,N_20640);
nor U20808 (N_20808,N_20618,N_20713);
or U20809 (N_20809,N_20743,N_20746);
or U20810 (N_20810,N_20740,N_20626);
nand U20811 (N_20811,N_20691,N_20773);
nor U20812 (N_20812,N_20765,N_20648);
nand U20813 (N_20813,N_20721,N_20630);
or U20814 (N_20814,N_20797,N_20716);
nor U20815 (N_20815,N_20745,N_20629);
and U20816 (N_20816,N_20785,N_20724);
xnor U20817 (N_20817,N_20605,N_20756);
nor U20818 (N_20818,N_20735,N_20623);
nor U20819 (N_20819,N_20794,N_20604);
and U20820 (N_20820,N_20631,N_20652);
xor U20821 (N_20821,N_20700,N_20706);
or U20822 (N_20822,N_20798,N_20766);
xnor U20823 (N_20823,N_20655,N_20674);
xor U20824 (N_20824,N_20614,N_20650);
xnor U20825 (N_20825,N_20719,N_20664);
xor U20826 (N_20826,N_20679,N_20627);
and U20827 (N_20827,N_20733,N_20772);
xnor U20828 (N_20828,N_20774,N_20695);
or U20829 (N_20829,N_20600,N_20654);
xnor U20830 (N_20830,N_20758,N_20762);
nand U20831 (N_20831,N_20789,N_20698);
nand U20832 (N_20832,N_20676,N_20726);
and U20833 (N_20833,N_20729,N_20686);
or U20834 (N_20834,N_20703,N_20778);
and U20835 (N_20835,N_20753,N_20705);
or U20836 (N_20836,N_20731,N_20741);
and U20837 (N_20837,N_20611,N_20704);
xor U20838 (N_20838,N_20739,N_20633);
nand U20839 (N_20839,N_20671,N_20768);
or U20840 (N_20840,N_20625,N_20659);
xnor U20841 (N_20841,N_20635,N_20622);
xnor U20842 (N_20842,N_20793,N_20669);
nor U20843 (N_20843,N_20653,N_20711);
xor U20844 (N_20844,N_20734,N_20736);
or U20845 (N_20845,N_20744,N_20672);
nand U20846 (N_20846,N_20621,N_20790);
and U20847 (N_20847,N_20781,N_20760);
nand U20848 (N_20848,N_20795,N_20662);
and U20849 (N_20849,N_20777,N_20699);
or U20850 (N_20850,N_20670,N_20761);
nor U20851 (N_20851,N_20682,N_20602);
and U20852 (N_20852,N_20668,N_20701);
xor U20853 (N_20853,N_20750,N_20722);
nand U20854 (N_20854,N_20663,N_20742);
nor U20855 (N_20855,N_20628,N_20632);
xnor U20856 (N_20856,N_20641,N_20619);
and U20857 (N_20857,N_20707,N_20799);
nor U20858 (N_20858,N_20769,N_20787);
nor U20859 (N_20859,N_20732,N_20606);
nor U20860 (N_20860,N_20609,N_20776);
nand U20861 (N_20861,N_20752,N_20624);
nand U20862 (N_20862,N_20688,N_20642);
xnor U20863 (N_20863,N_20685,N_20748);
and U20864 (N_20864,N_20690,N_20755);
nor U20865 (N_20865,N_20771,N_20749);
nor U20866 (N_20866,N_20647,N_20782);
nor U20867 (N_20867,N_20660,N_20651);
or U20868 (N_20868,N_20649,N_20764);
nand U20869 (N_20869,N_20747,N_20613);
nor U20870 (N_20870,N_20687,N_20788);
or U20871 (N_20871,N_20786,N_20675);
xnor U20872 (N_20872,N_20612,N_20796);
nor U20873 (N_20873,N_20616,N_20710);
xor U20874 (N_20874,N_20709,N_20702);
xor U20875 (N_20875,N_20775,N_20607);
nand U20876 (N_20876,N_20677,N_20637);
nand U20877 (N_20877,N_20615,N_20694);
or U20878 (N_20878,N_20738,N_20683);
nor U20879 (N_20879,N_20725,N_20783);
nor U20880 (N_20880,N_20608,N_20770);
and U20881 (N_20881,N_20723,N_20692);
or U20882 (N_20882,N_20645,N_20603);
or U20883 (N_20883,N_20656,N_20712);
or U20884 (N_20884,N_20714,N_20784);
or U20885 (N_20885,N_20715,N_20759);
nor U20886 (N_20886,N_20708,N_20610);
nand U20887 (N_20887,N_20767,N_20751);
and U20888 (N_20888,N_20665,N_20684);
and U20889 (N_20889,N_20617,N_20620);
nand U20890 (N_20890,N_20601,N_20636);
nor U20891 (N_20891,N_20638,N_20681);
nor U20892 (N_20892,N_20730,N_20763);
and U20893 (N_20893,N_20727,N_20779);
or U20894 (N_20894,N_20757,N_20792);
xor U20895 (N_20895,N_20728,N_20689);
nor U20896 (N_20896,N_20697,N_20673);
xnor U20897 (N_20897,N_20737,N_20658);
or U20898 (N_20898,N_20667,N_20717);
nor U20899 (N_20899,N_20780,N_20696);
and U20900 (N_20900,N_20782,N_20794);
and U20901 (N_20901,N_20760,N_20693);
and U20902 (N_20902,N_20712,N_20717);
and U20903 (N_20903,N_20705,N_20709);
and U20904 (N_20904,N_20611,N_20610);
nand U20905 (N_20905,N_20769,N_20763);
nor U20906 (N_20906,N_20762,N_20678);
xnor U20907 (N_20907,N_20705,N_20755);
nor U20908 (N_20908,N_20689,N_20793);
nand U20909 (N_20909,N_20767,N_20785);
or U20910 (N_20910,N_20719,N_20601);
nor U20911 (N_20911,N_20790,N_20639);
nor U20912 (N_20912,N_20746,N_20620);
and U20913 (N_20913,N_20749,N_20785);
xnor U20914 (N_20914,N_20667,N_20741);
or U20915 (N_20915,N_20621,N_20735);
nand U20916 (N_20916,N_20641,N_20784);
nand U20917 (N_20917,N_20674,N_20773);
and U20918 (N_20918,N_20722,N_20738);
nand U20919 (N_20919,N_20616,N_20767);
xor U20920 (N_20920,N_20658,N_20733);
or U20921 (N_20921,N_20797,N_20692);
nand U20922 (N_20922,N_20710,N_20646);
nor U20923 (N_20923,N_20604,N_20757);
xnor U20924 (N_20924,N_20775,N_20730);
or U20925 (N_20925,N_20662,N_20641);
nor U20926 (N_20926,N_20678,N_20634);
or U20927 (N_20927,N_20631,N_20760);
nand U20928 (N_20928,N_20711,N_20683);
nor U20929 (N_20929,N_20660,N_20619);
or U20930 (N_20930,N_20642,N_20628);
nand U20931 (N_20931,N_20762,N_20771);
nor U20932 (N_20932,N_20759,N_20737);
xor U20933 (N_20933,N_20744,N_20740);
and U20934 (N_20934,N_20784,N_20632);
nor U20935 (N_20935,N_20786,N_20631);
and U20936 (N_20936,N_20790,N_20609);
and U20937 (N_20937,N_20778,N_20770);
nand U20938 (N_20938,N_20653,N_20614);
nand U20939 (N_20939,N_20766,N_20635);
or U20940 (N_20940,N_20675,N_20785);
nand U20941 (N_20941,N_20795,N_20774);
nor U20942 (N_20942,N_20792,N_20788);
and U20943 (N_20943,N_20625,N_20728);
nand U20944 (N_20944,N_20696,N_20778);
nor U20945 (N_20945,N_20729,N_20732);
or U20946 (N_20946,N_20654,N_20655);
or U20947 (N_20947,N_20658,N_20667);
and U20948 (N_20948,N_20741,N_20717);
nand U20949 (N_20949,N_20757,N_20784);
xnor U20950 (N_20950,N_20727,N_20622);
nor U20951 (N_20951,N_20737,N_20690);
and U20952 (N_20952,N_20746,N_20635);
or U20953 (N_20953,N_20677,N_20782);
or U20954 (N_20954,N_20667,N_20606);
nand U20955 (N_20955,N_20745,N_20783);
nor U20956 (N_20956,N_20722,N_20786);
or U20957 (N_20957,N_20656,N_20671);
xnor U20958 (N_20958,N_20652,N_20617);
or U20959 (N_20959,N_20695,N_20658);
nand U20960 (N_20960,N_20668,N_20741);
nand U20961 (N_20961,N_20617,N_20787);
or U20962 (N_20962,N_20718,N_20781);
and U20963 (N_20963,N_20626,N_20796);
xnor U20964 (N_20964,N_20644,N_20695);
or U20965 (N_20965,N_20640,N_20605);
nor U20966 (N_20966,N_20669,N_20746);
and U20967 (N_20967,N_20611,N_20757);
xor U20968 (N_20968,N_20783,N_20775);
xor U20969 (N_20969,N_20782,N_20701);
nand U20970 (N_20970,N_20706,N_20645);
nor U20971 (N_20971,N_20790,N_20625);
nor U20972 (N_20972,N_20748,N_20745);
or U20973 (N_20973,N_20644,N_20774);
or U20974 (N_20974,N_20650,N_20686);
or U20975 (N_20975,N_20734,N_20719);
nor U20976 (N_20976,N_20642,N_20614);
xnor U20977 (N_20977,N_20744,N_20634);
xor U20978 (N_20978,N_20733,N_20660);
nand U20979 (N_20979,N_20706,N_20786);
nor U20980 (N_20980,N_20628,N_20671);
or U20981 (N_20981,N_20666,N_20765);
xnor U20982 (N_20982,N_20748,N_20669);
nor U20983 (N_20983,N_20667,N_20648);
nor U20984 (N_20984,N_20668,N_20764);
nand U20985 (N_20985,N_20627,N_20682);
or U20986 (N_20986,N_20712,N_20746);
or U20987 (N_20987,N_20679,N_20707);
or U20988 (N_20988,N_20794,N_20678);
nor U20989 (N_20989,N_20616,N_20696);
xor U20990 (N_20990,N_20637,N_20634);
and U20991 (N_20991,N_20623,N_20723);
nand U20992 (N_20992,N_20687,N_20682);
and U20993 (N_20993,N_20704,N_20728);
xnor U20994 (N_20994,N_20649,N_20718);
or U20995 (N_20995,N_20779,N_20771);
or U20996 (N_20996,N_20636,N_20748);
or U20997 (N_20997,N_20669,N_20777);
nor U20998 (N_20998,N_20786,N_20781);
or U20999 (N_20999,N_20679,N_20737);
xor U21000 (N_21000,N_20849,N_20983);
and U21001 (N_21001,N_20853,N_20908);
or U21002 (N_21002,N_20976,N_20898);
nor U21003 (N_21003,N_20906,N_20991);
or U21004 (N_21004,N_20930,N_20875);
and U21005 (N_21005,N_20862,N_20847);
nor U21006 (N_21006,N_20865,N_20841);
xnor U21007 (N_21007,N_20842,N_20843);
or U21008 (N_21008,N_20901,N_20947);
nand U21009 (N_21009,N_20848,N_20942);
and U21010 (N_21010,N_20850,N_20851);
nor U21011 (N_21011,N_20870,N_20982);
or U21012 (N_21012,N_20860,N_20832);
and U21013 (N_21013,N_20855,N_20888);
and U21014 (N_21014,N_20964,N_20931);
xnor U21015 (N_21015,N_20846,N_20915);
nand U21016 (N_21016,N_20935,N_20872);
xnor U21017 (N_21017,N_20899,N_20918);
xor U21018 (N_21018,N_20834,N_20940);
or U21019 (N_21019,N_20929,N_20943);
or U21020 (N_21020,N_20928,N_20936);
xnor U21021 (N_21021,N_20809,N_20957);
nand U21022 (N_21022,N_20977,N_20953);
nor U21023 (N_21023,N_20934,N_20965);
nand U21024 (N_21024,N_20959,N_20987);
nand U21025 (N_21025,N_20954,N_20919);
nor U21026 (N_21026,N_20980,N_20817);
nor U21027 (N_21027,N_20973,N_20812);
xor U21028 (N_21028,N_20814,N_20894);
and U21029 (N_21029,N_20966,N_20978);
or U21030 (N_21030,N_20926,N_20994);
or U21031 (N_21031,N_20944,N_20968);
nor U21032 (N_21032,N_20884,N_20825);
xor U21033 (N_21033,N_20844,N_20858);
or U21034 (N_21034,N_20808,N_20949);
xor U21035 (N_21035,N_20854,N_20986);
nand U21036 (N_21036,N_20920,N_20877);
nor U21037 (N_21037,N_20995,N_20989);
and U21038 (N_21038,N_20880,N_20904);
nand U21039 (N_21039,N_20826,N_20951);
or U21040 (N_21040,N_20800,N_20829);
nor U21041 (N_21041,N_20891,N_20861);
nand U21042 (N_21042,N_20893,N_20878);
xnor U21043 (N_21043,N_20967,N_20801);
or U21044 (N_21044,N_20903,N_20958);
or U21045 (N_21045,N_20909,N_20837);
and U21046 (N_21046,N_20955,N_20911);
and U21047 (N_21047,N_20938,N_20916);
nand U21048 (N_21048,N_20839,N_20981);
and U21049 (N_21049,N_20913,N_20892);
xor U21050 (N_21050,N_20910,N_20863);
nor U21051 (N_21051,N_20946,N_20927);
or U21052 (N_21052,N_20912,N_20859);
nand U21053 (N_21053,N_20974,N_20886);
nand U21054 (N_21054,N_20962,N_20924);
nor U21055 (N_21055,N_20961,N_20992);
xnor U21056 (N_21056,N_20900,N_20869);
and U21057 (N_21057,N_20804,N_20887);
nand U21058 (N_21058,N_20970,N_20822);
or U21059 (N_21059,N_20811,N_20838);
nor U21060 (N_21060,N_20998,N_20835);
nor U21061 (N_21061,N_20882,N_20895);
and U21062 (N_21062,N_20883,N_20917);
nor U21063 (N_21063,N_20879,N_20856);
nand U21064 (N_21064,N_20914,N_20950);
or U21065 (N_21065,N_20802,N_20840);
and U21066 (N_21066,N_20867,N_20828);
or U21067 (N_21067,N_20821,N_20945);
xnor U21068 (N_21068,N_20923,N_20993);
and U21069 (N_21069,N_20960,N_20939);
or U21070 (N_21070,N_20988,N_20823);
or U21071 (N_21071,N_20999,N_20824);
nand U21072 (N_21072,N_20815,N_20881);
xnor U21073 (N_21073,N_20810,N_20890);
xnor U21074 (N_21074,N_20874,N_20933);
xor U21075 (N_21075,N_20818,N_20922);
and U21076 (N_21076,N_20975,N_20819);
nand U21077 (N_21077,N_20845,N_20857);
xor U21078 (N_21078,N_20984,N_20990);
and U21079 (N_21079,N_20830,N_20925);
and U21080 (N_21080,N_20803,N_20816);
nand U21081 (N_21081,N_20831,N_20852);
and U21082 (N_21082,N_20807,N_20820);
nand U21083 (N_21083,N_20905,N_20827);
nand U21084 (N_21084,N_20805,N_20907);
nor U21085 (N_21085,N_20996,N_20969);
or U21086 (N_21086,N_20921,N_20937);
or U21087 (N_21087,N_20972,N_20889);
xor U21088 (N_21088,N_20932,N_20864);
nor U21089 (N_21089,N_20896,N_20897);
or U21090 (N_21090,N_20806,N_20873);
nor U21091 (N_21091,N_20979,N_20971);
xor U21092 (N_21092,N_20902,N_20866);
nand U21093 (N_21093,N_20836,N_20876);
xor U21094 (N_21094,N_20997,N_20813);
nor U21095 (N_21095,N_20963,N_20952);
or U21096 (N_21096,N_20948,N_20868);
xor U21097 (N_21097,N_20941,N_20956);
or U21098 (N_21098,N_20885,N_20833);
and U21099 (N_21099,N_20871,N_20985);
or U21100 (N_21100,N_20929,N_20947);
or U21101 (N_21101,N_20841,N_20860);
xnor U21102 (N_21102,N_20902,N_20803);
nor U21103 (N_21103,N_20982,N_20871);
nand U21104 (N_21104,N_20950,N_20838);
nor U21105 (N_21105,N_20989,N_20867);
nand U21106 (N_21106,N_20829,N_20857);
and U21107 (N_21107,N_20922,N_20964);
and U21108 (N_21108,N_20903,N_20991);
xnor U21109 (N_21109,N_20852,N_20858);
or U21110 (N_21110,N_20943,N_20939);
xor U21111 (N_21111,N_20846,N_20862);
nor U21112 (N_21112,N_20953,N_20919);
xor U21113 (N_21113,N_20991,N_20899);
or U21114 (N_21114,N_20977,N_20938);
nor U21115 (N_21115,N_20889,N_20862);
nand U21116 (N_21116,N_20999,N_20907);
or U21117 (N_21117,N_20866,N_20841);
or U21118 (N_21118,N_20860,N_20936);
or U21119 (N_21119,N_20815,N_20889);
nor U21120 (N_21120,N_20887,N_20813);
or U21121 (N_21121,N_20902,N_20855);
and U21122 (N_21122,N_20988,N_20999);
and U21123 (N_21123,N_20839,N_20872);
and U21124 (N_21124,N_20954,N_20941);
or U21125 (N_21125,N_20880,N_20921);
nor U21126 (N_21126,N_20962,N_20956);
and U21127 (N_21127,N_20828,N_20909);
nor U21128 (N_21128,N_20861,N_20951);
nand U21129 (N_21129,N_20960,N_20857);
nand U21130 (N_21130,N_20872,N_20824);
and U21131 (N_21131,N_20969,N_20902);
nor U21132 (N_21132,N_20878,N_20956);
xor U21133 (N_21133,N_20837,N_20865);
nor U21134 (N_21134,N_20826,N_20967);
xor U21135 (N_21135,N_20845,N_20839);
nor U21136 (N_21136,N_20892,N_20985);
or U21137 (N_21137,N_20972,N_20949);
and U21138 (N_21138,N_20860,N_20818);
nand U21139 (N_21139,N_20984,N_20825);
nand U21140 (N_21140,N_20818,N_20945);
or U21141 (N_21141,N_20821,N_20885);
or U21142 (N_21142,N_20843,N_20918);
and U21143 (N_21143,N_20948,N_20989);
or U21144 (N_21144,N_20867,N_20878);
xor U21145 (N_21145,N_20866,N_20920);
nor U21146 (N_21146,N_20941,N_20923);
and U21147 (N_21147,N_20998,N_20937);
or U21148 (N_21148,N_20890,N_20844);
or U21149 (N_21149,N_20948,N_20885);
xor U21150 (N_21150,N_20822,N_20805);
nor U21151 (N_21151,N_20939,N_20929);
and U21152 (N_21152,N_20834,N_20968);
xor U21153 (N_21153,N_20821,N_20814);
nand U21154 (N_21154,N_20968,N_20883);
or U21155 (N_21155,N_20923,N_20825);
or U21156 (N_21156,N_20921,N_20801);
nand U21157 (N_21157,N_20976,N_20875);
xor U21158 (N_21158,N_20816,N_20979);
xor U21159 (N_21159,N_20838,N_20921);
nor U21160 (N_21160,N_20800,N_20852);
or U21161 (N_21161,N_20801,N_20927);
nor U21162 (N_21162,N_20803,N_20813);
nand U21163 (N_21163,N_20956,N_20868);
nor U21164 (N_21164,N_20900,N_20847);
or U21165 (N_21165,N_20966,N_20989);
nor U21166 (N_21166,N_20869,N_20905);
xor U21167 (N_21167,N_20956,N_20947);
nand U21168 (N_21168,N_20975,N_20853);
and U21169 (N_21169,N_20953,N_20910);
nand U21170 (N_21170,N_20914,N_20952);
or U21171 (N_21171,N_20825,N_20834);
and U21172 (N_21172,N_20866,N_20835);
xor U21173 (N_21173,N_20960,N_20888);
xnor U21174 (N_21174,N_20823,N_20930);
nand U21175 (N_21175,N_20844,N_20822);
nor U21176 (N_21176,N_20808,N_20934);
nor U21177 (N_21177,N_20913,N_20831);
or U21178 (N_21178,N_20881,N_20840);
nor U21179 (N_21179,N_20979,N_20818);
nor U21180 (N_21180,N_20836,N_20877);
nand U21181 (N_21181,N_20869,N_20974);
or U21182 (N_21182,N_20823,N_20946);
nor U21183 (N_21183,N_20800,N_20834);
nor U21184 (N_21184,N_20931,N_20891);
xnor U21185 (N_21185,N_20878,N_20923);
xor U21186 (N_21186,N_20884,N_20998);
nor U21187 (N_21187,N_20972,N_20998);
nand U21188 (N_21188,N_20957,N_20980);
nor U21189 (N_21189,N_20965,N_20966);
nor U21190 (N_21190,N_20915,N_20887);
and U21191 (N_21191,N_20947,N_20960);
nor U21192 (N_21192,N_20867,N_20836);
and U21193 (N_21193,N_20834,N_20844);
or U21194 (N_21194,N_20802,N_20903);
nand U21195 (N_21195,N_20825,N_20935);
or U21196 (N_21196,N_20865,N_20842);
nand U21197 (N_21197,N_20969,N_20858);
nand U21198 (N_21198,N_20990,N_20851);
nand U21199 (N_21199,N_20947,N_20936);
xor U21200 (N_21200,N_21006,N_21031);
nor U21201 (N_21201,N_21129,N_21010);
and U21202 (N_21202,N_21159,N_21099);
nor U21203 (N_21203,N_21045,N_21098);
nor U21204 (N_21204,N_21147,N_21197);
or U21205 (N_21205,N_21057,N_21151);
nor U21206 (N_21206,N_21005,N_21106);
or U21207 (N_21207,N_21108,N_21164);
or U21208 (N_21208,N_21107,N_21175);
nand U21209 (N_21209,N_21195,N_21160);
nor U21210 (N_21210,N_21067,N_21027);
nand U21211 (N_21211,N_21021,N_21174);
nor U21212 (N_21212,N_21130,N_21192);
nor U21213 (N_21213,N_21181,N_21198);
nand U21214 (N_21214,N_21056,N_21121);
and U21215 (N_21215,N_21112,N_21154);
or U21216 (N_21216,N_21120,N_21061);
or U21217 (N_21217,N_21033,N_21051);
or U21218 (N_21218,N_21125,N_21178);
or U21219 (N_21219,N_21109,N_21059);
xor U21220 (N_21220,N_21104,N_21017);
or U21221 (N_21221,N_21105,N_21141);
nor U21222 (N_21222,N_21144,N_21070);
xor U21223 (N_21223,N_21042,N_21179);
and U21224 (N_21224,N_21124,N_21187);
xor U21225 (N_21225,N_21188,N_21193);
xnor U21226 (N_21226,N_21052,N_21012);
xor U21227 (N_21227,N_21158,N_21172);
nor U21228 (N_21228,N_21035,N_21093);
nand U21229 (N_21229,N_21189,N_21115);
nor U21230 (N_21230,N_21134,N_21149);
and U21231 (N_21231,N_21122,N_21153);
nand U21232 (N_21232,N_21110,N_21022);
or U21233 (N_21233,N_21183,N_21039);
nor U21234 (N_21234,N_21028,N_21139);
or U21235 (N_21235,N_21029,N_21169);
xnor U21236 (N_21236,N_21150,N_21173);
nand U21237 (N_21237,N_21111,N_21080);
or U21238 (N_21238,N_21043,N_21020);
nand U21239 (N_21239,N_21199,N_21090);
xor U21240 (N_21240,N_21085,N_21162);
nor U21241 (N_21241,N_21068,N_21089);
and U21242 (N_21242,N_21170,N_21165);
xor U21243 (N_21243,N_21001,N_21152);
nor U21244 (N_21244,N_21076,N_21184);
xor U21245 (N_21245,N_21077,N_21015);
or U21246 (N_21246,N_21000,N_21131);
and U21247 (N_21247,N_21163,N_21074);
nand U21248 (N_21248,N_21040,N_21008);
nand U21249 (N_21249,N_21185,N_21123);
nor U21250 (N_21250,N_21142,N_21171);
or U21251 (N_21251,N_21023,N_21078);
and U21252 (N_21252,N_21100,N_21018);
nand U21253 (N_21253,N_21087,N_21191);
or U21254 (N_21254,N_21048,N_21086);
nand U21255 (N_21255,N_21146,N_21116);
nand U21256 (N_21256,N_21166,N_21194);
nor U21257 (N_21257,N_21011,N_21156);
or U21258 (N_21258,N_21113,N_21084);
or U21259 (N_21259,N_21063,N_21066);
and U21260 (N_21260,N_21126,N_21128);
nand U21261 (N_21261,N_21135,N_21047);
xor U21262 (N_21262,N_21054,N_21167);
xor U21263 (N_21263,N_21025,N_21155);
and U21264 (N_21264,N_21058,N_21081);
or U21265 (N_21265,N_21182,N_21132);
xnor U21266 (N_21266,N_21038,N_21024);
nor U21267 (N_21267,N_21036,N_21095);
xor U21268 (N_21268,N_21050,N_21065);
xnor U21269 (N_21269,N_21055,N_21136);
or U21270 (N_21270,N_21082,N_21196);
nand U21271 (N_21271,N_21137,N_21034);
xor U21272 (N_21272,N_21114,N_21083);
nor U21273 (N_21273,N_21003,N_21037);
xnor U21274 (N_21274,N_21140,N_21049);
xor U21275 (N_21275,N_21133,N_21026);
xnor U21276 (N_21276,N_21002,N_21186);
nand U21277 (N_21277,N_21072,N_21177);
nor U21278 (N_21278,N_21019,N_21161);
xnor U21279 (N_21279,N_21071,N_21117);
xnor U21280 (N_21280,N_21064,N_21102);
or U21281 (N_21281,N_21079,N_21046);
and U21282 (N_21282,N_21180,N_21053);
nor U21283 (N_21283,N_21096,N_21075);
nor U21284 (N_21284,N_21176,N_21013);
or U21285 (N_21285,N_21118,N_21069);
and U21286 (N_21286,N_21138,N_21007);
xor U21287 (N_21287,N_21143,N_21119);
nor U21288 (N_21288,N_21016,N_21101);
xor U21289 (N_21289,N_21088,N_21148);
xor U21290 (N_21290,N_21168,N_21157);
or U21291 (N_21291,N_21062,N_21094);
or U21292 (N_21292,N_21103,N_21190);
or U21293 (N_21293,N_21097,N_21060);
and U21294 (N_21294,N_21073,N_21030);
or U21295 (N_21295,N_21009,N_21092);
or U21296 (N_21296,N_21145,N_21127);
nand U21297 (N_21297,N_21032,N_21014);
xor U21298 (N_21298,N_21004,N_21044);
nand U21299 (N_21299,N_21091,N_21041);
nor U21300 (N_21300,N_21047,N_21144);
nand U21301 (N_21301,N_21194,N_21100);
and U21302 (N_21302,N_21112,N_21064);
nand U21303 (N_21303,N_21198,N_21096);
and U21304 (N_21304,N_21149,N_21048);
xor U21305 (N_21305,N_21199,N_21087);
or U21306 (N_21306,N_21090,N_21048);
nor U21307 (N_21307,N_21016,N_21116);
and U21308 (N_21308,N_21166,N_21185);
nor U21309 (N_21309,N_21178,N_21045);
xor U21310 (N_21310,N_21044,N_21189);
and U21311 (N_21311,N_21000,N_21017);
xor U21312 (N_21312,N_21072,N_21082);
xnor U21313 (N_21313,N_21158,N_21123);
nand U21314 (N_21314,N_21067,N_21091);
nor U21315 (N_21315,N_21055,N_21183);
xor U21316 (N_21316,N_21188,N_21149);
xnor U21317 (N_21317,N_21095,N_21061);
nor U21318 (N_21318,N_21089,N_21134);
nand U21319 (N_21319,N_21105,N_21010);
xnor U21320 (N_21320,N_21194,N_21097);
nand U21321 (N_21321,N_21074,N_21024);
or U21322 (N_21322,N_21168,N_21004);
or U21323 (N_21323,N_21092,N_21190);
and U21324 (N_21324,N_21197,N_21198);
nand U21325 (N_21325,N_21085,N_21086);
xnor U21326 (N_21326,N_21125,N_21035);
nand U21327 (N_21327,N_21168,N_21138);
xnor U21328 (N_21328,N_21025,N_21129);
nor U21329 (N_21329,N_21134,N_21015);
and U21330 (N_21330,N_21151,N_21181);
and U21331 (N_21331,N_21146,N_21123);
and U21332 (N_21332,N_21111,N_21127);
and U21333 (N_21333,N_21066,N_21093);
or U21334 (N_21334,N_21119,N_21166);
and U21335 (N_21335,N_21127,N_21141);
xnor U21336 (N_21336,N_21180,N_21192);
or U21337 (N_21337,N_21013,N_21038);
nor U21338 (N_21338,N_21016,N_21093);
and U21339 (N_21339,N_21153,N_21090);
xnor U21340 (N_21340,N_21154,N_21095);
xnor U21341 (N_21341,N_21107,N_21016);
xor U21342 (N_21342,N_21094,N_21144);
nor U21343 (N_21343,N_21023,N_21136);
and U21344 (N_21344,N_21029,N_21196);
nand U21345 (N_21345,N_21065,N_21033);
nor U21346 (N_21346,N_21194,N_21018);
and U21347 (N_21347,N_21010,N_21181);
xnor U21348 (N_21348,N_21159,N_21137);
nand U21349 (N_21349,N_21040,N_21189);
nor U21350 (N_21350,N_21144,N_21097);
or U21351 (N_21351,N_21094,N_21183);
and U21352 (N_21352,N_21119,N_21151);
nor U21353 (N_21353,N_21101,N_21136);
nor U21354 (N_21354,N_21092,N_21010);
and U21355 (N_21355,N_21111,N_21099);
nor U21356 (N_21356,N_21096,N_21124);
nor U21357 (N_21357,N_21137,N_21119);
or U21358 (N_21358,N_21159,N_21088);
nor U21359 (N_21359,N_21019,N_21091);
xnor U21360 (N_21360,N_21135,N_21098);
nand U21361 (N_21361,N_21169,N_21138);
nor U21362 (N_21362,N_21101,N_21002);
or U21363 (N_21363,N_21059,N_21173);
nor U21364 (N_21364,N_21165,N_21104);
nor U21365 (N_21365,N_21012,N_21030);
or U21366 (N_21366,N_21037,N_21106);
or U21367 (N_21367,N_21038,N_21041);
or U21368 (N_21368,N_21068,N_21184);
nand U21369 (N_21369,N_21169,N_21089);
nand U21370 (N_21370,N_21148,N_21096);
xor U21371 (N_21371,N_21046,N_21024);
nor U21372 (N_21372,N_21074,N_21160);
nand U21373 (N_21373,N_21041,N_21036);
and U21374 (N_21374,N_21162,N_21031);
xnor U21375 (N_21375,N_21093,N_21101);
or U21376 (N_21376,N_21119,N_21046);
nor U21377 (N_21377,N_21108,N_21183);
and U21378 (N_21378,N_21131,N_21178);
nand U21379 (N_21379,N_21033,N_21138);
or U21380 (N_21380,N_21121,N_21183);
nand U21381 (N_21381,N_21091,N_21011);
nor U21382 (N_21382,N_21160,N_21061);
and U21383 (N_21383,N_21163,N_21076);
nand U21384 (N_21384,N_21124,N_21023);
or U21385 (N_21385,N_21067,N_21062);
nand U21386 (N_21386,N_21042,N_21182);
nand U21387 (N_21387,N_21068,N_21001);
and U21388 (N_21388,N_21189,N_21080);
nor U21389 (N_21389,N_21147,N_21120);
or U21390 (N_21390,N_21096,N_21009);
xor U21391 (N_21391,N_21180,N_21073);
or U21392 (N_21392,N_21006,N_21044);
or U21393 (N_21393,N_21168,N_21009);
nor U21394 (N_21394,N_21173,N_21087);
nor U21395 (N_21395,N_21132,N_21045);
nand U21396 (N_21396,N_21011,N_21056);
or U21397 (N_21397,N_21171,N_21109);
nor U21398 (N_21398,N_21133,N_21199);
xnor U21399 (N_21399,N_21077,N_21183);
xnor U21400 (N_21400,N_21281,N_21232);
and U21401 (N_21401,N_21378,N_21311);
nand U21402 (N_21402,N_21258,N_21295);
xnor U21403 (N_21403,N_21356,N_21204);
or U21404 (N_21404,N_21273,N_21323);
or U21405 (N_21405,N_21301,N_21335);
nor U21406 (N_21406,N_21360,N_21332);
nand U21407 (N_21407,N_21297,N_21251);
nand U21408 (N_21408,N_21381,N_21256);
and U21409 (N_21409,N_21326,N_21220);
nand U21410 (N_21410,N_21364,N_21352);
nand U21411 (N_21411,N_21219,N_21346);
and U21412 (N_21412,N_21261,N_21336);
nand U21413 (N_21413,N_21398,N_21361);
or U21414 (N_21414,N_21298,N_21280);
nand U21415 (N_21415,N_21215,N_21321);
xnor U21416 (N_21416,N_21284,N_21319);
or U21417 (N_21417,N_21268,N_21337);
or U21418 (N_21418,N_21371,N_21314);
nand U21419 (N_21419,N_21317,N_21262);
and U21420 (N_21420,N_21286,N_21302);
nor U21421 (N_21421,N_21228,N_21222);
nand U21422 (N_21422,N_21207,N_21265);
and U21423 (N_21423,N_21342,N_21217);
or U21424 (N_21424,N_21316,N_21376);
or U21425 (N_21425,N_21201,N_21283);
nand U21426 (N_21426,N_21328,N_21329);
xor U21427 (N_21427,N_21287,N_21386);
nor U21428 (N_21428,N_21389,N_21291);
nor U21429 (N_21429,N_21213,N_21293);
nand U21430 (N_21430,N_21210,N_21212);
and U21431 (N_21431,N_21282,N_21277);
xor U21432 (N_21432,N_21245,N_21373);
and U21433 (N_21433,N_21312,N_21351);
and U21434 (N_21434,N_21309,N_21365);
nand U21435 (N_21435,N_21271,N_21338);
nand U21436 (N_21436,N_21266,N_21345);
and U21437 (N_21437,N_21252,N_21230);
and U21438 (N_21438,N_21358,N_21366);
nor U21439 (N_21439,N_21226,N_21390);
xor U21440 (N_21440,N_21237,N_21362);
xor U21441 (N_21441,N_21272,N_21203);
or U21442 (N_21442,N_21348,N_21289);
or U21443 (N_21443,N_21285,N_21322);
nor U21444 (N_21444,N_21385,N_21339);
nand U21445 (N_21445,N_21372,N_21233);
nor U21446 (N_21446,N_21341,N_21227);
and U21447 (N_21447,N_21259,N_21308);
or U21448 (N_21448,N_21238,N_21391);
or U21449 (N_21449,N_21324,N_21347);
xnor U21450 (N_21450,N_21320,N_21369);
nand U21451 (N_21451,N_21264,N_21206);
nand U21452 (N_21452,N_21396,N_21246);
nor U21453 (N_21453,N_21205,N_21236);
nor U21454 (N_21454,N_21257,N_21394);
or U21455 (N_21455,N_21292,N_21343);
and U21456 (N_21456,N_21325,N_21380);
xnor U21457 (N_21457,N_21388,N_21225);
or U21458 (N_21458,N_21235,N_21310);
xnor U21459 (N_21459,N_21242,N_21216);
and U21460 (N_21460,N_21229,N_21375);
nand U21461 (N_21461,N_21334,N_21374);
or U21462 (N_21462,N_21241,N_21353);
nor U21463 (N_21463,N_21303,N_21202);
xnor U21464 (N_21464,N_21255,N_21368);
nor U21465 (N_21465,N_21208,N_21355);
and U21466 (N_21466,N_21244,N_21397);
xor U21467 (N_21467,N_21275,N_21218);
nand U21468 (N_21468,N_21399,N_21248);
or U21469 (N_21469,N_21340,N_21223);
or U21470 (N_21470,N_21363,N_21367);
nand U21471 (N_21471,N_21247,N_21370);
and U21472 (N_21472,N_21263,N_21200);
nand U21473 (N_21473,N_21269,N_21327);
and U21474 (N_21474,N_21253,N_21279);
nand U21475 (N_21475,N_21315,N_21243);
xnor U21476 (N_21476,N_21331,N_21211);
nor U21477 (N_21477,N_21270,N_21209);
or U21478 (N_21478,N_21296,N_21350);
xnor U21479 (N_21479,N_21304,N_21318);
or U21480 (N_21480,N_21393,N_21240);
or U21481 (N_21481,N_21234,N_21214);
nor U21482 (N_21482,N_21224,N_21290);
and U21483 (N_21483,N_21278,N_21383);
xnor U21484 (N_21484,N_21349,N_21387);
and U21485 (N_21485,N_21344,N_21231);
or U21486 (N_21486,N_21239,N_21306);
nand U21487 (N_21487,N_21395,N_21249);
nand U21488 (N_21488,N_21313,N_21305);
and U21489 (N_21489,N_21274,N_21300);
nand U21490 (N_21490,N_21359,N_21254);
nand U21491 (N_21491,N_21276,N_21267);
nor U21492 (N_21492,N_21382,N_21377);
or U21493 (N_21493,N_21299,N_21288);
xnor U21494 (N_21494,N_21384,N_21354);
or U21495 (N_21495,N_21357,N_21221);
xnor U21496 (N_21496,N_21307,N_21330);
nor U21497 (N_21497,N_21250,N_21379);
and U21498 (N_21498,N_21392,N_21294);
and U21499 (N_21499,N_21333,N_21260);
xnor U21500 (N_21500,N_21222,N_21337);
and U21501 (N_21501,N_21382,N_21203);
xnor U21502 (N_21502,N_21218,N_21363);
nand U21503 (N_21503,N_21398,N_21369);
nor U21504 (N_21504,N_21222,N_21343);
and U21505 (N_21505,N_21240,N_21267);
nand U21506 (N_21506,N_21238,N_21255);
or U21507 (N_21507,N_21307,N_21335);
xnor U21508 (N_21508,N_21232,N_21252);
or U21509 (N_21509,N_21263,N_21340);
xor U21510 (N_21510,N_21236,N_21211);
nor U21511 (N_21511,N_21374,N_21311);
nor U21512 (N_21512,N_21284,N_21265);
xor U21513 (N_21513,N_21213,N_21306);
and U21514 (N_21514,N_21228,N_21300);
nand U21515 (N_21515,N_21387,N_21326);
and U21516 (N_21516,N_21386,N_21242);
nor U21517 (N_21517,N_21341,N_21216);
and U21518 (N_21518,N_21200,N_21221);
or U21519 (N_21519,N_21278,N_21230);
xnor U21520 (N_21520,N_21392,N_21201);
xnor U21521 (N_21521,N_21363,N_21386);
nor U21522 (N_21522,N_21309,N_21301);
xnor U21523 (N_21523,N_21350,N_21327);
or U21524 (N_21524,N_21320,N_21247);
nor U21525 (N_21525,N_21222,N_21347);
nor U21526 (N_21526,N_21379,N_21329);
nand U21527 (N_21527,N_21209,N_21367);
or U21528 (N_21528,N_21388,N_21277);
nand U21529 (N_21529,N_21255,N_21251);
nand U21530 (N_21530,N_21348,N_21327);
nor U21531 (N_21531,N_21356,N_21289);
and U21532 (N_21532,N_21386,N_21351);
nor U21533 (N_21533,N_21354,N_21390);
or U21534 (N_21534,N_21315,N_21256);
and U21535 (N_21535,N_21270,N_21207);
xor U21536 (N_21536,N_21316,N_21332);
and U21537 (N_21537,N_21285,N_21361);
or U21538 (N_21538,N_21320,N_21354);
or U21539 (N_21539,N_21392,N_21352);
nand U21540 (N_21540,N_21375,N_21325);
nand U21541 (N_21541,N_21238,N_21226);
nor U21542 (N_21542,N_21353,N_21296);
nor U21543 (N_21543,N_21276,N_21207);
nand U21544 (N_21544,N_21357,N_21353);
and U21545 (N_21545,N_21373,N_21209);
xnor U21546 (N_21546,N_21270,N_21332);
or U21547 (N_21547,N_21224,N_21255);
and U21548 (N_21548,N_21201,N_21339);
xnor U21549 (N_21549,N_21349,N_21350);
and U21550 (N_21550,N_21360,N_21348);
nand U21551 (N_21551,N_21302,N_21279);
nand U21552 (N_21552,N_21250,N_21283);
nand U21553 (N_21553,N_21336,N_21341);
and U21554 (N_21554,N_21224,N_21267);
xor U21555 (N_21555,N_21243,N_21310);
and U21556 (N_21556,N_21257,N_21262);
nand U21557 (N_21557,N_21251,N_21338);
xor U21558 (N_21558,N_21309,N_21335);
nand U21559 (N_21559,N_21256,N_21294);
or U21560 (N_21560,N_21247,N_21261);
or U21561 (N_21561,N_21398,N_21207);
and U21562 (N_21562,N_21231,N_21202);
nor U21563 (N_21563,N_21384,N_21203);
or U21564 (N_21564,N_21341,N_21396);
and U21565 (N_21565,N_21320,N_21204);
nor U21566 (N_21566,N_21289,N_21380);
nand U21567 (N_21567,N_21256,N_21353);
nand U21568 (N_21568,N_21228,N_21245);
xnor U21569 (N_21569,N_21280,N_21330);
or U21570 (N_21570,N_21260,N_21305);
nor U21571 (N_21571,N_21376,N_21209);
xnor U21572 (N_21572,N_21357,N_21276);
and U21573 (N_21573,N_21234,N_21363);
and U21574 (N_21574,N_21245,N_21284);
nand U21575 (N_21575,N_21220,N_21339);
or U21576 (N_21576,N_21272,N_21275);
nor U21577 (N_21577,N_21205,N_21348);
or U21578 (N_21578,N_21251,N_21240);
nor U21579 (N_21579,N_21346,N_21307);
or U21580 (N_21580,N_21234,N_21254);
or U21581 (N_21581,N_21220,N_21234);
and U21582 (N_21582,N_21235,N_21360);
xnor U21583 (N_21583,N_21320,N_21259);
nor U21584 (N_21584,N_21268,N_21202);
nand U21585 (N_21585,N_21201,N_21285);
or U21586 (N_21586,N_21282,N_21328);
or U21587 (N_21587,N_21248,N_21331);
nor U21588 (N_21588,N_21359,N_21356);
or U21589 (N_21589,N_21385,N_21344);
xor U21590 (N_21590,N_21291,N_21219);
and U21591 (N_21591,N_21304,N_21376);
and U21592 (N_21592,N_21231,N_21286);
nor U21593 (N_21593,N_21279,N_21252);
nand U21594 (N_21594,N_21331,N_21263);
or U21595 (N_21595,N_21378,N_21299);
nand U21596 (N_21596,N_21233,N_21281);
nand U21597 (N_21597,N_21204,N_21309);
and U21598 (N_21598,N_21338,N_21355);
xor U21599 (N_21599,N_21364,N_21348);
or U21600 (N_21600,N_21553,N_21495);
or U21601 (N_21601,N_21492,N_21562);
and U21602 (N_21602,N_21501,N_21528);
nor U21603 (N_21603,N_21555,N_21558);
nor U21604 (N_21604,N_21508,N_21448);
xor U21605 (N_21605,N_21420,N_21453);
and U21606 (N_21606,N_21596,N_21529);
or U21607 (N_21607,N_21469,N_21456);
and U21608 (N_21608,N_21527,N_21570);
nand U21609 (N_21609,N_21526,N_21407);
or U21610 (N_21610,N_21512,N_21592);
nor U21611 (N_21611,N_21466,N_21455);
nand U21612 (N_21612,N_21540,N_21462);
nand U21613 (N_21613,N_21416,N_21591);
or U21614 (N_21614,N_21408,N_21468);
nor U21615 (N_21615,N_21490,N_21538);
xnor U21616 (N_21616,N_21424,N_21521);
xnor U21617 (N_21617,N_21594,N_21535);
nand U21618 (N_21618,N_21584,N_21496);
xnor U21619 (N_21619,N_21557,N_21589);
and U21620 (N_21620,N_21545,N_21411);
nand U21621 (N_21621,N_21532,N_21426);
nor U21622 (N_21622,N_21568,N_21465);
nand U21623 (N_21623,N_21428,N_21518);
xnor U21624 (N_21624,N_21597,N_21579);
or U21625 (N_21625,N_21457,N_21461);
or U21626 (N_21626,N_21498,N_21503);
xnor U21627 (N_21627,N_21410,N_21542);
nand U21628 (N_21628,N_21506,N_21452);
or U21629 (N_21629,N_21511,N_21515);
and U21630 (N_21630,N_21406,N_21563);
and U21631 (N_21631,N_21583,N_21487);
nand U21632 (N_21632,N_21401,N_21483);
or U21633 (N_21633,N_21470,N_21547);
or U21634 (N_21634,N_21544,N_21421);
nand U21635 (N_21635,N_21516,N_21444);
and U21636 (N_21636,N_21432,N_21485);
nand U21637 (N_21637,N_21441,N_21463);
or U21638 (N_21638,N_21572,N_21478);
xor U21639 (N_21639,N_21443,N_21510);
xnor U21640 (N_21640,N_21405,N_21476);
and U21641 (N_21641,N_21522,N_21445);
or U21642 (N_21642,N_21433,N_21585);
or U21643 (N_21643,N_21595,N_21413);
nand U21644 (N_21644,N_21414,N_21430);
and U21645 (N_21645,N_21412,N_21451);
nand U21646 (N_21646,N_21530,N_21507);
nand U21647 (N_21647,N_21582,N_21409);
xor U21648 (N_21648,N_21404,N_21574);
and U21649 (N_21649,N_21520,N_21442);
xor U21650 (N_21650,N_21590,N_21473);
and U21651 (N_21651,N_21477,N_21434);
nand U21652 (N_21652,N_21436,N_21580);
xnor U21653 (N_21653,N_21427,N_21559);
xnor U21654 (N_21654,N_21549,N_21536);
xnor U21655 (N_21655,N_21588,N_21598);
or U21656 (N_21656,N_21577,N_21482);
nand U21657 (N_21657,N_21519,N_21446);
and U21658 (N_21658,N_21593,N_21440);
nand U21659 (N_21659,N_21474,N_21419);
or U21660 (N_21660,N_21415,N_21576);
nand U21661 (N_21661,N_21587,N_21537);
nand U21662 (N_21662,N_21479,N_21548);
nor U21663 (N_21663,N_21450,N_21534);
or U21664 (N_21664,N_21586,N_21565);
nand U21665 (N_21665,N_21417,N_21431);
nor U21666 (N_21666,N_21472,N_21567);
nand U21667 (N_21667,N_21569,N_21581);
or U21668 (N_21668,N_21454,N_21514);
nor U21669 (N_21669,N_21403,N_21460);
and U21670 (N_21670,N_21422,N_21546);
nor U21671 (N_21671,N_21423,N_21513);
or U21672 (N_21672,N_21539,N_21400);
or U21673 (N_21673,N_21475,N_21481);
and U21674 (N_21674,N_21480,N_21502);
and U21675 (N_21675,N_21517,N_21599);
or U21676 (N_21676,N_21575,N_21573);
or U21677 (N_21677,N_21551,N_21524);
nand U21678 (N_21678,N_21458,N_21402);
nor U21679 (N_21679,N_21439,N_21484);
xor U21680 (N_21680,N_21491,N_21493);
nor U21681 (N_21681,N_21488,N_21429);
nor U21682 (N_21682,N_21564,N_21571);
or U21683 (N_21683,N_21509,N_21435);
and U21684 (N_21684,N_21525,N_21505);
and U21685 (N_21685,N_21467,N_21471);
nor U21686 (N_21686,N_21556,N_21554);
and U21687 (N_21687,N_21504,N_21464);
nand U21688 (N_21688,N_21578,N_21561);
nor U21689 (N_21689,N_21437,N_21497);
nand U21690 (N_21690,N_21486,N_21438);
or U21691 (N_21691,N_21499,N_21447);
and U21692 (N_21692,N_21459,N_21523);
and U21693 (N_21693,N_21531,N_21489);
and U21694 (N_21694,N_21418,N_21541);
nor U21695 (N_21695,N_21500,N_21543);
xor U21696 (N_21696,N_21550,N_21533);
nor U21697 (N_21697,N_21566,N_21425);
nand U21698 (N_21698,N_21560,N_21552);
xor U21699 (N_21699,N_21449,N_21494);
or U21700 (N_21700,N_21484,N_21579);
nand U21701 (N_21701,N_21476,N_21499);
xor U21702 (N_21702,N_21500,N_21427);
or U21703 (N_21703,N_21533,N_21541);
or U21704 (N_21704,N_21425,N_21579);
nor U21705 (N_21705,N_21536,N_21457);
xnor U21706 (N_21706,N_21502,N_21591);
xor U21707 (N_21707,N_21570,N_21533);
nand U21708 (N_21708,N_21532,N_21480);
and U21709 (N_21709,N_21423,N_21446);
xnor U21710 (N_21710,N_21579,N_21558);
and U21711 (N_21711,N_21585,N_21513);
and U21712 (N_21712,N_21493,N_21425);
xnor U21713 (N_21713,N_21576,N_21476);
or U21714 (N_21714,N_21525,N_21442);
nand U21715 (N_21715,N_21588,N_21433);
nand U21716 (N_21716,N_21476,N_21462);
xor U21717 (N_21717,N_21534,N_21508);
nand U21718 (N_21718,N_21533,N_21574);
nor U21719 (N_21719,N_21411,N_21466);
nand U21720 (N_21720,N_21588,N_21543);
nand U21721 (N_21721,N_21564,N_21411);
and U21722 (N_21722,N_21559,N_21440);
nand U21723 (N_21723,N_21544,N_21522);
nor U21724 (N_21724,N_21434,N_21554);
xnor U21725 (N_21725,N_21475,N_21596);
nor U21726 (N_21726,N_21502,N_21549);
or U21727 (N_21727,N_21594,N_21555);
nand U21728 (N_21728,N_21567,N_21483);
and U21729 (N_21729,N_21512,N_21583);
nor U21730 (N_21730,N_21438,N_21565);
and U21731 (N_21731,N_21444,N_21589);
nand U21732 (N_21732,N_21515,N_21418);
nor U21733 (N_21733,N_21439,N_21438);
and U21734 (N_21734,N_21591,N_21493);
nand U21735 (N_21735,N_21524,N_21422);
xor U21736 (N_21736,N_21473,N_21564);
xnor U21737 (N_21737,N_21504,N_21410);
xnor U21738 (N_21738,N_21489,N_21420);
nand U21739 (N_21739,N_21470,N_21410);
nand U21740 (N_21740,N_21408,N_21441);
nor U21741 (N_21741,N_21478,N_21513);
nand U21742 (N_21742,N_21439,N_21489);
and U21743 (N_21743,N_21487,N_21513);
nand U21744 (N_21744,N_21535,N_21455);
and U21745 (N_21745,N_21420,N_21477);
nor U21746 (N_21746,N_21413,N_21563);
nor U21747 (N_21747,N_21562,N_21450);
and U21748 (N_21748,N_21493,N_21410);
and U21749 (N_21749,N_21508,N_21572);
and U21750 (N_21750,N_21541,N_21526);
and U21751 (N_21751,N_21542,N_21505);
or U21752 (N_21752,N_21499,N_21430);
and U21753 (N_21753,N_21503,N_21476);
or U21754 (N_21754,N_21415,N_21441);
or U21755 (N_21755,N_21547,N_21401);
nand U21756 (N_21756,N_21485,N_21594);
xor U21757 (N_21757,N_21446,N_21454);
nor U21758 (N_21758,N_21585,N_21409);
and U21759 (N_21759,N_21590,N_21549);
and U21760 (N_21760,N_21482,N_21534);
or U21761 (N_21761,N_21535,N_21585);
nor U21762 (N_21762,N_21457,N_21437);
or U21763 (N_21763,N_21428,N_21540);
or U21764 (N_21764,N_21440,N_21580);
nor U21765 (N_21765,N_21514,N_21540);
or U21766 (N_21766,N_21470,N_21464);
or U21767 (N_21767,N_21547,N_21550);
and U21768 (N_21768,N_21504,N_21443);
xor U21769 (N_21769,N_21545,N_21583);
and U21770 (N_21770,N_21422,N_21527);
and U21771 (N_21771,N_21529,N_21533);
nor U21772 (N_21772,N_21428,N_21522);
or U21773 (N_21773,N_21431,N_21452);
xor U21774 (N_21774,N_21511,N_21406);
and U21775 (N_21775,N_21491,N_21485);
nand U21776 (N_21776,N_21498,N_21552);
nand U21777 (N_21777,N_21438,N_21519);
nand U21778 (N_21778,N_21508,N_21539);
nor U21779 (N_21779,N_21491,N_21511);
and U21780 (N_21780,N_21542,N_21465);
or U21781 (N_21781,N_21408,N_21406);
nand U21782 (N_21782,N_21444,N_21553);
and U21783 (N_21783,N_21493,N_21436);
nand U21784 (N_21784,N_21407,N_21415);
nor U21785 (N_21785,N_21521,N_21531);
nand U21786 (N_21786,N_21562,N_21509);
nor U21787 (N_21787,N_21542,N_21463);
nand U21788 (N_21788,N_21503,N_21545);
nor U21789 (N_21789,N_21588,N_21451);
or U21790 (N_21790,N_21449,N_21524);
and U21791 (N_21791,N_21430,N_21508);
and U21792 (N_21792,N_21416,N_21430);
and U21793 (N_21793,N_21420,N_21536);
xnor U21794 (N_21794,N_21570,N_21564);
nor U21795 (N_21795,N_21434,N_21559);
nand U21796 (N_21796,N_21512,N_21509);
or U21797 (N_21797,N_21544,N_21508);
nand U21798 (N_21798,N_21518,N_21539);
xnor U21799 (N_21799,N_21417,N_21577);
nor U21800 (N_21800,N_21603,N_21672);
or U21801 (N_21801,N_21718,N_21751);
xnor U21802 (N_21802,N_21626,N_21758);
and U21803 (N_21803,N_21727,N_21605);
nand U21804 (N_21804,N_21662,N_21713);
and U21805 (N_21805,N_21664,N_21634);
or U21806 (N_21806,N_21686,N_21682);
nor U21807 (N_21807,N_21668,N_21723);
nor U21808 (N_21808,N_21691,N_21705);
nand U21809 (N_21809,N_21671,N_21740);
nor U21810 (N_21810,N_21708,N_21677);
nor U21811 (N_21811,N_21607,N_21726);
nand U21812 (N_21812,N_21648,N_21709);
nand U21813 (N_21813,N_21788,N_21661);
nand U21814 (N_21814,N_21780,N_21742);
or U21815 (N_21815,N_21630,N_21619);
xor U21816 (N_21816,N_21635,N_21666);
xor U21817 (N_21817,N_21745,N_21657);
nand U21818 (N_21818,N_21748,N_21636);
nor U21819 (N_21819,N_21711,N_21743);
xor U21820 (N_21820,N_21791,N_21656);
and U21821 (N_21821,N_21757,N_21645);
nor U21822 (N_21822,N_21675,N_21651);
nand U21823 (N_21823,N_21608,N_21716);
xor U21824 (N_21824,N_21735,N_21699);
and U21825 (N_21825,N_21683,N_21752);
or U21826 (N_21826,N_21773,N_21617);
xor U21827 (N_21827,N_21698,N_21710);
and U21828 (N_21828,N_21674,N_21725);
nand U21829 (N_21829,N_21613,N_21775);
and U21830 (N_21830,N_21642,N_21736);
and U21831 (N_21831,N_21640,N_21777);
and U21832 (N_21832,N_21782,N_21712);
and U21833 (N_21833,N_21625,N_21793);
nor U21834 (N_21834,N_21749,N_21754);
nor U21835 (N_21835,N_21770,N_21797);
and U21836 (N_21836,N_21799,N_21706);
or U21837 (N_21837,N_21679,N_21781);
xnor U21838 (N_21838,N_21728,N_21750);
xor U21839 (N_21839,N_21611,N_21704);
nand U21840 (N_21840,N_21796,N_21787);
and U21841 (N_21841,N_21637,N_21643);
xnor U21842 (N_21842,N_21700,N_21612);
or U21843 (N_21843,N_21618,N_21663);
nand U21844 (N_21844,N_21676,N_21702);
xor U21845 (N_21845,N_21768,N_21692);
xnor U21846 (N_21846,N_21628,N_21707);
and U21847 (N_21847,N_21769,N_21732);
and U21848 (N_21848,N_21766,N_21703);
nand U21849 (N_21849,N_21792,N_21715);
nand U21850 (N_21850,N_21776,N_21685);
and U21851 (N_21851,N_21681,N_21647);
and U21852 (N_21852,N_21695,N_21653);
nor U21853 (N_21853,N_21697,N_21688);
xor U21854 (N_21854,N_21667,N_21623);
nor U21855 (N_21855,N_21655,N_21600);
and U21856 (N_21856,N_21763,N_21690);
and U21857 (N_21857,N_21624,N_21627);
or U21858 (N_21858,N_21650,N_21772);
or U21859 (N_21859,N_21601,N_21784);
and U21860 (N_21860,N_21610,N_21765);
xnor U21861 (N_21861,N_21602,N_21670);
or U21862 (N_21862,N_21795,N_21646);
or U21863 (N_21863,N_21778,N_21761);
xnor U21864 (N_21864,N_21696,N_21660);
and U21865 (N_21865,N_21669,N_21629);
xnor U21866 (N_21866,N_21738,N_21762);
and U21867 (N_21867,N_21730,N_21759);
nor U21868 (N_21868,N_21771,N_21684);
xor U21869 (N_21869,N_21641,N_21638);
nand U21870 (N_21870,N_21734,N_21639);
xor U21871 (N_21871,N_21659,N_21609);
nor U21872 (N_21872,N_21722,N_21694);
nor U21873 (N_21873,N_21654,N_21652);
and U21874 (N_21874,N_21714,N_21614);
or U21875 (N_21875,N_21798,N_21622);
xor U21876 (N_21876,N_21737,N_21658);
xnor U21877 (N_21877,N_21621,N_21632);
xor U21878 (N_21878,N_21721,N_21774);
nor U21879 (N_21879,N_21680,N_21786);
nand U21880 (N_21880,N_21729,N_21606);
and U21881 (N_21881,N_21741,N_21689);
and U21882 (N_21882,N_21756,N_21719);
or U21883 (N_21883,N_21724,N_21767);
or U21884 (N_21884,N_21665,N_21701);
and U21885 (N_21885,N_21755,N_21644);
nor U21886 (N_21886,N_21747,N_21616);
or U21887 (N_21887,N_21794,N_21744);
and U21888 (N_21888,N_21687,N_21790);
xor U21889 (N_21889,N_21649,N_21760);
nand U21890 (N_21890,N_21720,N_21785);
and U21891 (N_21891,N_21604,N_21779);
nor U21892 (N_21892,N_21746,N_21733);
or U21893 (N_21893,N_21717,N_21764);
nor U21894 (N_21894,N_21620,N_21739);
nand U21895 (N_21895,N_21783,N_21753);
nand U21896 (N_21896,N_21673,N_21731);
and U21897 (N_21897,N_21789,N_21693);
xnor U21898 (N_21898,N_21631,N_21633);
or U21899 (N_21899,N_21678,N_21615);
nand U21900 (N_21900,N_21774,N_21706);
and U21901 (N_21901,N_21727,N_21738);
xor U21902 (N_21902,N_21784,N_21631);
nand U21903 (N_21903,N_21686,N_21629);
nor U21904 (N_21904,N_21710,N_21728);
or U21905 (N_21905,N_21646,N_21797);
nor U21906 (N_21906,N_21736,N_21740);
or U21907 (N_21907,N_21794,N_21755);
or U21908 (N_21908,N_21652,N_21767);
nand U21909 (N_21909,N_21665,N_21768);
nand U21910 (N_21910,N_21725,N_21678);
nor U21911 (N_21911,N_21603,N_21794);
nor U21912 (N_21912,N_21654,N_21720);
nand U21913 (N_21913,N_21776,N_21702);
xnor U21914 (N_21914,N_21754,N_21686);
or U21915 (N_21915,N_21675,N_21778);
nand U21916 (N_21916,N_21684,N_21720);
xor U21917 (N_21917,N_21770,N_21615);
xor U21918 (N_21918,N_21661,N_21783);
nor U21919 (N_21919,N_21677,N_21632);
xnor U21920 (N_21920,N_21689,N_21666);
nand U21921 (N_21921,N_21616,N_21723);
xor U21922 (N_21922,N_21695,N_21627);
nor U21923 (N_21923,N_21625,N_21648);
xnor U21924 (N_21924,N_21734,N_21704);
nor U21925 (N_21925,N_21796,N_21752);
nor U21926 (N_21926,N_21697,N_21797);
or U21927 (N_21927,N_21766,N_21784);
nand U21928 (N_21928,N_21732,N_21770);
and U21929 (N_21929,N_21627,N_21705);
xnor U21930 (N_21930,N_21771,N_21707);
nand U21931 (N_21931,N_21635,N_21767);
and U21932 (N_21932,N_21780,N_21608);
xor U21933 (N_21933,N_21625,N_21736);
nand U21934 (N_21934,N_21797,N_21651);
and U21935 (N_21935,N_21603,N_21753);
and U21936 (N_21936,N_21737,N_21740);
or U21937 (N_21937,N_21666,N_21659);
nand U21938 (N_21938,N_21629,N_21695);
or U21939 (N_21939,N_21640,N_21604);
nor U21940 (N_21940,N_21651,N_21647);
and U21941 (N_21941,N_21686,N_21637);
and U21942 (N_21942,N_21664,N_21613);
or U21943 (N_21943,N_21655,N_21742);
nor U21944 (N_21944,N_21707,N_21672);
nand U21945 (N_21945,N_21730,N_21615);
nand U21946 (N_21946,N_21729,N_21708);
xor U21947 (N_21947,N_21740,N_21622);
or U21948 (N_21948,N_21748,N_21727);
xor U21949 (N_21949,N_21618,N_21674);
nor U21950 (N_21950,N_21733,N_21609);
or U21951 (N_21951,N_21773,N_21772);
nor U21952 (N_21952,N_21680,N_21699);
xnor U21953 (N_21953,N_21651,N_21732);
nand U21954 (N_21954,N_21630,N_21617);
nand U21955 (N_21955,N_21743,N_21741);
or U21956 (N_21956,N_21676,N_21778);
nand U21957 (N_21957,N_21796,N_21791);
and U21958 (N_21958,N_21727,N_21639);
xnor U21959 (N_21959,N_21602,N_21632);
xor U21960 (N_21960,N_21645,N_21740);
nor U21961 (N_21961,N_21707,N_21669);
or U21962 (N_21962,N_21647,N_21625);
nor U21963 (N_21963,N_21757,N_21754);
nand U21964 (N_21964,N_21635,N_21705);
nand U21965 (N_21965,N_21755,N_21640);
xnor U21966 (N_21966,N_21682,N_21669);
or U21967 (N_21967,N_21636,N_21784);
or U21968 (N_21968,N_21778,N_21671);
nand U21969 (N_21969,N_21683,N_21611);
nand U21970 (N_21970,N_21611,N_21638);
or U21971 (N_21971,N_21676,N_21639);
xnor U21972 (N_21972,N_21650,N_21664);
or U21973 (N_21973,N_21724,N_21779);
nand U21974 (N_21974,N_21645,N_21678);
xor U21975 (N_21975,N_21734,N_21664);
nor U21976 (N_21976,N_21715,N_21647);
nor U21977 (N_21977,N_21696,N_21765);
or U21978 (N_21978,N_21747,N_21628);
and U21979 (N_21979,N_21626,N_21735);
or U21980 (N_21980,N_21715,N_21782);
xnor U21981 (N_21981,N_21638,N_21717);
and U21982 (N_21982,N_21759,N_21620);
nand U21983 (N_21983,N_21677,N_21643);
or U21984 (N_21984,N_21623,N_21705);
or U21985 (N_21985,N_21790,N_21647);
and U21986 (N_21986,N_21781,N_21653);
nand U21987 (N_21987,N_21764,N_21659);
xor U21988 (N_21988,N_21774,N_21692);
xor U21989 (N_21989,N_21785,N_21624);
nor U21990 (N_21990,N_21723,N_21674);
and U21991 (N_21991,N_21617,N_21632);
nor U21992 (N_21992,N_21676,N_21644);
and U21993 (N_21993,N_21788,N_21789);
xor U21994 (N_21994,N_21627,N_21639);
xor U21995 (N_21995,N_21603,N_21699);
and U21996 (N_21996,N_21694,N_21709);
xor U21997 (N_21997,N_21729,N_21635);
and U21998 (N_21998,N_21714,N_21794);
nand U21999 (N_21999,N_21624,N_21674);
or U22000 (N_22000,N_21933,N_21989);
xor U22001 (N_22001,N_21954,N_21929);
or U22002 (N_22002,N_21909,N_21948);
xor U22003 (N_22003,N_21993,N_21949);
or U22004 (N_22004,N_21934,N_21880);
nand U22005 (N_22005,N_21960,N_21847);
nand U22006 (N_22006,N_21869,N_21808);
nor U22007 (N_22007,N_21829,N_21913);
xor U22008 (N_22008,N_21977,N_21853);
nor U22009 (N_22009,N_21930,N_21824);
or U22010 (N_22010,N_21961,N_21839);
nor U22011 (N_22011,N_21863,N_21932);
nor U22012 (N_22012,N_21816,N_21941);
nor U22013 (N_22013,N_21935,N_21838);
xnor U22014 (N_22014,N_21857,N_21823);
nor U22015 (N_22015,N_21819,N_21895);
or U22016 (N_22016,N_21859,N_21806);
or U22017 (N_22017,N_21979,N_21896);
or U22018 (N_22018,N_21887,N_21910);
and U22019 (N_22019,N_21902,N_21959);
and U22020 (N_22020,N_21963,N_21939);
and U22021 (N_22021,N_21956,N_21992);
nor U22022 (N_22022,N_21912,N_21876);
nand U22023 (N_22023,N_21858,N_21833);
and U22024 (N_22024,N_21968,N_21974);
and U22025 (N_22025,N_21976,N_21879);
xnor U22026 (N_22026,N_21872,N_21882);
nand U22027 (N_22027,N_21918,N_21985);
or U22028 (N_22028,N_21831,N_21850);
xor U22029 (N_22029,N_21969,N_21825);
and U22030 (N_22030,N_21978,N_21984);
and U22031 (N_22031,N_21893,N_21826);
nor U22032 (N_22032,N_21860,N_21990);
nor U22033 (N_22033,N_21862,N_21972);
xnor U22034 (N_22034,N_21973,N_21904);
xnor U22035 (N_22035,N_21938,N_21925);
or U22036 (N_22036,N_21878,N_21921);
nor U22037 (N_22037,N_21950,N_21818);
nor U22038 (N_22038,N_21817,N_21805);
nand U22039 (N_22039,N_21946,N_21994);
and U22040 (N_22040,N_21940,N_21865);
and U22041 (N_22041,N_21966,N_21811);
nand U22042 (N_22042,N_21828,N_21856);
nand U22043 (N_22043,N_21927,N_21982);
xnor U22044 (N_22044,N_21892,N_21911);
nand U22045 (N_22045,N_21945,N_21957);
and U22046 (N_22046,N_21834,N_21964);
nand U22047 (N_22047,N_21849,N_21883);
nor U22048 (N_22048,N_21958,N_21822);
nor U22049 (N_22049,N_21846,N_21801);
nor U22050 (N_22050,N_21890,N_21844);
nor U22051 (N_22051,N_21955,N_21814);
and U22052 (N_22052,N_21965,N_21988);
or U22053 (N_22053,N_21886,N_21802);
nand U22054 (N_22054,N_21908,N_21804);
nor U22055 (N_22055,N_21813,N_21922);
nor U22056 (N_22056,N_21970,N_21914);
nor U22057 (N_22057,N_21810,N_21837);
and U22058 (N_22058,N_21821,N_21916);
nand U22059 (N_22059,N_21943,N_21840);
xnor U22060 (N_22060,N_21815,N_21907);
nand U22061 (N_22061,N_21962,N_21967);
or U22062 (N_22062,N_21953,N_21931);
nor U22063 (N_22063,N_21845,N_21851);
nor U22064 (N_22064,N_21881,N_21900);
and U22065 (N_22065,N_21871,N_21873);
or U22066 (N_22066,N_21868,N_21919);
xor U22067 (N_22067,N_21812,N_21986);
and U22068 (N_22068,N_21920,N_21996);
and U22069 (N_22069,N_21991,N_21981);
nand U22070 (N_22070,N_21889,N_21842);
nand U22071 (N_22071,N_21874,N_21894);
or U22072 (N_22072,N_21923,N_21809);
and U22073 (N_22073,N_21928,N_21897);
nor U22074 (N_22074,N_21999,N_21937);
or U22075 (N_22075,N_21877,N_21942);
or U22076 (N_22076,N_21980,N_21854);
or U22077 (N_22077,N_21848,N_21803);
xor U22078 (N_22078,N_21807,N_21917);
nand U22079 (N_22079,N_21915,N_21898);
or U22080 (N_22080,N_21841,N_21926);
or U22081 (N_22081,N_21952,N_21830);
or U22082 (N_22082,N_21820,N_21906);
nand U22083 (N_22083,N_21870,N_21998);
nand U22084 (N_22084,N_21951,N_21901);
nor U22085 (N_22085,N_21875,N_21947);
xnor U22086 (N_22086,N_21971,N_21866);
nor U22087 (N_22087,N_21975,N_21936);
nand U22088 (N_22088,N_21924,N_21867);
nor U22089 (N_22089,N_21903,N_21995);
nand U22090 (N_22090,N_21861,N_21987);
nand U22091 (N_22091,N_21983,N_21852);
or U22092 (N_22092,N_21800,N_21855);
nor U22093 (N_22093,N_21827,N_21891);
xnor U22094 (N_22094,N_21864,N_21843);
or U22095 (N_22095,N_21836,N_21944);
nand U22096 (N_22096,N_21835,N_21905);
xnor U22097 (N_22097,N_21832,N_21885);
nand U22098 (N_22098,N_21997,N_21888);
nand U22099 (N_22099,N_21899,N_21884);
xnor U22100 (N_22100,N_21884,N_21915);
xnor U22101 (N_22101,N_21967,N_21819);
and U22102 (N_22102,N_21801,N_21952);
xor U22103 (N_22103,N_21943,N_21923);
nor U22104 (N_22104,N_21875,N_21815);
nand U22105 (N_22105,N_21952,N_21959);
xor U22106 (N_22106,N_21876,N_21871);
and U22107 (N_22107,N_21960,N_21887);
and U22108 (N_22108,N_21812,N_21982);
nand U22109 (N_22109,N_21861,N_21971);
xnor U22110 (N_22110,N_21905,N_21809);
xnor U22111 (N_22111,N_21861,N_21929);
or U22112 (N_22112,N_21809,N_21844);
nor U22113 (N_22113,N_21958,N_21909);
nand U22114 (N_22114,N_21809,N_21816);
or U22115 (N_22115,N_21873,N_21963);
nand U22116 (N_22116,N_21871,N_21913);
nor U22117 (N_22117,N_21845,N_21824);
xnor U22118 (N_22118,N_21902,N_21857);
or U22119 (N_22119,N_21804,N_21938);
and U22120 (N_22120,N_21974,N_21914);
and U22121 (N_22121,N_21878,N_21910);
xnor U22122 (N_22122,N_21968,N_21914);
nor U22123 (N_22123,N_21897,N_21902);
and U22124 (N_22124,N_21852,N_21869);
nand U22125 (N_22125,N_21941,N_21801);
nor U22126 (N_22126,N_21803,N_21974);
and U22127 (N_22127,N_21953,N_21824);
and U22128 (N_22128,N_21965,N_21929);
and U22129 (N_22129,N_21974,N_21818);
nor U22130 (N_22130,N_21961,N_21891);
nand U22131 (N_22131,N_21829,N_21986);
nor U22132 (N_22132,N_21852,N_21871);
nand U22133 (N_22133,N_21976,N_21852);
xor U22134 (N_22134,N_21850,N_21859);
nor U22135 (N_22135,N_21863,N_21986);
or U22136 (N_22136,N_21941,N_21966);
nor U22137 (N_22137,N_21887,N_21962);
or U22138 (N_22138,N_21893,N_21891);
nand U22139 (N_22139,N_21955,N_21877);
nor U22140 (N_22140,N_21881,N_21802);
nand U22141 (N_22141,N_21906,N_21861);
nor U22142 (N_22142,N_21834,N_21925);
nand U22143 (N_22143,N_21944,N_21890);
nand U22144 (N_22144,N_21878,N_21816);
and U22145 (N_22145,N_21916,N_21857);
nand U22146 (N_22146,N_21850,N_21851);
or U22147 (N_22147,N_21898,N_21835);
nor U22148 (N_22148,N_21943,N_21946);
nor U22149 (N_22149,N_21845,N_21970);
nand U22150 (N_22150,N_21882,N_21879);
nand U22151 (N_22151,N_21879,N_21818);
or U22152 (N_22152,N_21963,N_21804);
and U22153 (N_22153,N_21923,N_21860);
and U22154 (N_22154,N_21996,N_21887);
xor U22155 (N_22155,N_21954,N_21875);
nor U22156 (N_22156,N_21981,N_21913);
nor U22157 (N_22157,N_21910,N_21835);
xor U22158 (N_22158,N_21868,N_21989);
xor U22159 (N_22159,N_21997,N_21852);
nor U22160 (N_22160,N_21859,N_21967);
and U22161 (N_22161,N_21993,N_21958);
and U22162 (N_22162,N_21998,N_21823);
nor U22163 (N_22163,N_21947,N_21855);
or U22164 (N_22164,N_21984,N_21955);
or U22165 (N_22165,N_21991,N_21830);
nand U22166 (N_22166,N_21942,N_21977);
xnor U22167 (N_22167,N_21960,N_21899);
and U22168 (N_22168,N_21898,N_21964);
and U22169 (N_22169,N_21954,N_21807);
or U22170 (N_22170,N_21925,N_21809);
nor U22171 (N_22171,N_21876,N_21962);
nor U22172 (N_22172,N_21825,N_21874);
xor U22173 (N_22173,N_21841,N_21883);
nand U22174 (N_22174,N_21956,N_21954);
or U22175 (N_22175,N_21819,N_21986);
or U22176 (N_22176,N_21822,N_21842);
or U22177 (N_22177,N_21923,N_21841);
nand U22178 (N_22178,N_21914,N_21865);
xor U22179 (N_22179,N_21892,N_21990);
and U22180 (N_22180,N_21844,N_21992);
nor U22181 (N_22181,N_21964,N_21974);
nand U22182 (N_22182,N_21964,N_21986);
nor U22183 (N_22183,N_21836,N_21989);
xor U22184 (N_22184,N_21824,N_21959);
and U22185 (N_22185,N_21994,N_21814);
and U22186 (N_22186,N_21818,N_21930);
nand U22187 (N_22187,N_21967,N_21996);
or U22188 (N_22188,N_21927,N_21814);
or U22189 (N_22189,N_21853,N_21821);
xnor U22190 (N_22190,N_21972,N_21976);
or U22191 (N_22191,N_21808,N_21929);
nor U22192 (N_22192,N_21893,N_21813);
xnor U22193 (N_22193,N_21964,N_21959);
nand U22194 (N_22194,N_21915,N_21902);
nand U22195 (N_22195,N_21846,N_21961);
and U22196 (N_22196,N_21898,N_21817);
or U22197 (N_22197,N_21878,N_21922);
or U22198 (N_22198,N_21884,N_21988);
nor U22199 (N_22199,N_21850,N_21808);
nor U22200 (N_22200,N_22160,N_22154);
nand U22201 (N_22201,N_22024,N_22135);
xnor U22202 (N_22202,N_22131,N_22048);
nand U22203 (N_22203,N_22157,N_22130);
nor U22204 (N_22204,N_22122,N_22136);
or U22205 (N_22205,N_22041,N_22017);
xor U22206 (N_22206,N_22146,N_22014);
xnor U22207 (N_22207,N_22061,N_22089);
nor U22208 (N_22208,N_22194,N_22110);
nand U22209 (N_22209,N_22035,N_22166);
nor U22210 (N_22210,N_22104,N_22056);
or U22211 (N_22211,N_22071,N_22027);
or U22212 (N_22212,N_22054,N_22178);
or U22213 (N_22213,N_22044,N_22016);
xnor U22214 (N_22214,N_22198,N_22137);
nor U22215 (N_22215,N_22064,N_22097);
nand U22216 (N_22216,N_22013,N_22032);
xnor U22217 (N_22217,N_22195,N_22175);
or U22218 (N_22218,N_22078,N_22021);
xnor U22219 (N_22219,N_22028,N_22163);
or U22220 (N_22220,N_22039,N_22069);
xor U22221 (N_22221,N_22192,N_22004);
nor U22222 (N_22222,N_22076,N_22180);
and U22223 (N_22223,N_22031,N_22019);
or U22224 (N_22224,N_22162,N_22077);
nand U22225 (N_22225,N_22118,N_22108);
xor U22226 (N_22226,N_22156,N_22119);
xnor U22227 (N_22227,N_22124,N_22100);
nor U22228 (N_22228,N_22121,N_22058);
xor U22229 (N_22229,N_22172,N_22082);
nor U22230 (N_22230,N_22188,N_22010);
nand U22231 (N_22231,N_22183,N_22053);
xor U22232 (N_22232,N_22063,N_22057);
xor U22233 (N_22233,N_22143,N_22102);
nand U22234 (N_22234,N_22085,N_22006);
and U22235 (N_22235,N_22185,N_22099);
xor U22236 (N_22236,N_22134,N_22020);
or U22237 (N_22237,N_22083,N_22126);
nand U22238 (N_22238,N_22144,N_22141);
and U22239 (N_22239,N_22115,N_22033);
and U22240 (N_22240,N_22109,N_22092);
or U22241 (N_22241,N_22184,N_22171);
nand U22242 (N_22242,N_22008,N_22059);
and U22243 (N_22243,N_22161,N_22111);
nand U22244 (N_22244,N_22009,N_22081);
xnor U22245 (N_22245,N_22070,N_22176);
nor U22246 (N_22246,N_22158,N_22128);
xnor U22247 (N_22247,N_22036,N_22065);
nor U22248 (N_22248,N_22129,N_22095);
xor U22249 (N_22249,N_22153,N_22011);
xor U22250 (N_22250,N_22155,N_22101);
and U22251 (N_22251,N_22113,N_22073);
xor U22252 (N_22252,N_22152,N_22148);
xnor U22253 (N_22253,N_22132,N_22096);
nand U22254 (N_22254,N_22138,N_22164);
xnor U22255 (N_22255,N_22116,N_22186);
nor U22256 (N_22256,N_22117,N_22051);
xor U22257 (N_22257,N_22120,N_22103);
and U22258 (N_22258,N_22139,N_22079);
nor U22259 (N_22259,N_22149,N_22000);
nor U22260 (N_22260,N_22106,N_22142);
xnor U22261 (N_22261,N_22191,N_22022);
or U22262 (N_22262,N_22127,N_22075);
xor U22263 (N_22263,N_22030,N_22159);
xor U22264 (N_22264,N_22040,N_22168);
or U22265 (N_22265,N_22047,N_22147);
and U22266 (N_22266,N_22133,N_22174);
xor U22267 (N_22267,N_22190,N_22034);
nand U22268 (N_22268,N_22060,N_22001);
nor U22269 (N_22269,N_22052,N_22187);
nand U22270 (N_22270,N_22066,N_22043);
or U22271 (N_22271,N_22112,N_22145);
xnor U22272 (N_22272,N_22196,N_22179);
or U22273 (N_22273,N_22072,N_22046);
xor U22274 (N_22274,N_22197,N_22094);
xnor U22275 (N_22275,N_22090,N_22026);
and U22276 (N_22276,N_22062,N_22087);
nor U22277 (N_22277,N_22193,N_22012);
nand U22278 (N_22278,N_22049,N_22042);
and U22279 (N_22279,N_22105,N_22025);
nor U22280 (N_22280,N_22091,N_22199);
nand U22281 (N_22281,N_22093,N_22086);
and U22282 (N_22282,N_22007,N_22055);
nand U22283 (N_22283,N_22023,N_22181);
or U22284 (N_22284,N_22169,N_22074);
nand U22285 (N_22285,N_22038,N_22125);
or U22286 (N_22286,N_22173,N_22088);
nor U22287 (N_22287,N_22165,N_22015);
or U22288 (N_22288,N_22177,N_22151);
and U22289 (N_22289,N_22114,N_22150);
xor U22290 (N_22290,N_22045,N_22098);
and U22291 (N_22291,N_22189,N_22068);
or U22292 (N_22292,N_22140,N_22080);
or U22293 (N_22293,N_22084,N_22037);
nor U22294 (N_22294,N_22002,N_22123);
or U22295 (N_22295,N_22167,N_22029);
or U22296 (N_22296,N_22170,N_22005);
and U22297 (N_22297,N_22050,N_22182);
and U22298 (N_22298,N_22067,N_22003);
and U22299 (N_22299,N_22107,N_22018);
xor U22300 (N_22300,N_22062,N_22007);
nand U22301 (N_22301,N_22000,N_22134);
nand U22302 (N_22302,N_22049,N_22106);
nand U22303 (N_22303,N_22168,N_22004);
and U22304 (N_22304,N_22175,N_22096);
nand U22305 (N_22305,N_22139,N_22121);
and U22306 (N_22306,N_22073,N_22182);
or U22307 (N_22307,N_22046,N_22036);
nor U22308 (N_22308,N_22138,N_22038);
nand U22309 (N_22309,N_22180,N_22023);
and U22310 (N_22310,N_22090,N_22075);
nor U22311 (N_22311,N_22050,N_22021);
xor U22312 (N_22312,N_22088,N_22142);
nand U22313 (N_22313,N_22172,N_22178);
xor U22314 (N_22314,N_22135,N_22187);
xnor U22315 (N_22315,N_22007,N_22029);
nor U22316 (N_22316,N_22094,N_22129);
xor U22317 (N_22317,N_22105,N_22015);
xor U22318 (N_22318,N_22024,N_22021);
or U22319 (N_22319,N_22003,N_22000);
nand U22320 (N_22320,N_22145,N_22089);
nand U22321 (N_22321,N_22157,N_22018);
nand U22322 (N_22322,N_22017,N_22141);
xnor U22323 (N_22323,N_22127,N_22035);
xor U22324 (N_22324,N_22160,N_22018);
nor U22325 (N_22325,N_22064,N_22109);
and U22326 (N_22326,N_22085,N_22122);
nand U22327 (N_22327,N_22133,N_22166);
or U22328 (N_22328,N_22103,N_22115);
and U22329 (N_22329,N_22187,N_22101);
and U22330 (N_22330,N_22165,N_22197);
and U22331 (N_22331,N_22192,N_22132);
nand U22332 (N_22332,N_22107,N_22158);
nand U22333 (N_22333,N_22102,N_22006);
nand U22334 (N_22334,N_22186,N_22106);
nor U22335 (N_22335,N_22079,N_22135);
and U22336 (N_22336,N_22187,N_22065);
nand U22337 (N_22337,N_22196,N_22040);
xor U22338 (N_22338,N_22007,N_22041);
nand U22339 (N_22339,N_22006,N_22071);
nor U22340 (N_22340,N_22048,N_22030);
nor U22341 (N_22341,N_22102,N_22109);
and U22342 (N_22342,N_22133,N_22171);
nand U22343 (N_22343,N_22041,N_22003);
and U22344 (N_22344,N_22175,N_22113);
and U22345 (N_22345,N_22026,N_22160);
xnor U22346 (N_22346,N_22130,N_22190);
xor U22347 (N_22347,N_22162,N_22006);
and U22348 (N_22348,N_22049,N_22116);
nor U22349 (N_22349,N_22162,N_22107);
or U22350 (N_22350,N_22038,N_22025);
nand U22351 (N_22351,N_22049,N_22069);
and U22352 (N_22352,N_22105,N_22092);
or U22353 (N_22353,N_22046,N_22043);
nor U22354 (N_22354,N_22124,N_22064);
or U22355 (N_22355,N_22056,N_22124);
and U22356 (N_22356,N_22017,N_22171);
or U22357 (N_22357,N_22059,N_22092);
or U22358 (N_22358,N_22034,N_22115);
nand U22359 (N_22359,N_22152,N_22120);
nor U22360 (N_22360,N_22107,N_22015);
nand U22361 (N_22361,N_22169,N_22119);
nand U22362 (N_22362,N_22161,N_22194);
nand U22363 (N_22363,N_22186,N_22005);
nor U22364 (N_22364,N_22179,N_22022);
or U22365 (N_22365,N_22184,N_22028);
or U22366 (N_22366,N_22128,N_22090);
nand U22367 (N_22367,N_22109,N_22088);
xnor U22368 (N_22368,N_22150,N_22151);
nor U22369 (N_22369,N_22102,N_22120);
xor U22370 (N_22370,N_22179,N_22127);
and U22371 (N_22371,N_22010,N_22129);
and U22372 (N_22372,N_22070,N_22181);
or U22373 (N_22373,N_22062,N_22167);
xnor U22374 (N_22374,N_22091,N_22075);
and U22375 (N_22375,N_22160,N_22079);
nand U22376 (N_22376,N_22153,N_22196);
xor U22377 (N_22377,N_22142,N_22013);
xor U22378 (N_22378,N_22058,N_22095);
and U22379 (N_22379,N_22141,N_22180);
nor U22380 (N_22380,N_22115,N_22024);
nor U22381 (N_22381,N_22159,N_22052);
xor U22382 (N_22382,N_22148,N_22010);
or U22383 (N_22383,N_22159,N_22103);
xnor U22384 (N_22384,N_22016,N_22050);
or U22385 (N_22385,N_22143,N_22072);
xnor U22386 (N_22386,N_22164,N_22117);
xnor U22387 (N_22387,N_22030,N_22148);
nor U22388 (N_22388,N_22171,N_22190);
xnor U22389 (N_22389,N_22132,N_22002);
xor U22390 (N_22390,N_22050,N_22179);
xnor U22391 (N_22391,N_22198,N_22122);
xnor U22392 (N_22392,N_22068,N_22197);
or U22393 (N_22393,N_22058,N_22129);
xor U22394 (N_22394,N_22058,N_22041);
nor U22395 (N_22395,N_22086,N_22175);
and U22396 (N_22396,N_22131,N_22139);
and U22397 (N_22397,N_22072,N_22092);
or U22398 (N_22398,N_22069,N_22009);
nor U22399 (N_22399,N_22165,N_22037);
nor U22400 (N_22400,N_22213,N_22337);
or U22401 (N_22401,N_22313,N_22260);
nor U22402 (N_22402,N_22206,N_22203);
nor U22403 (N_22403,N_22365,N_22385);
and U22404 (N_22404,N_22323,N_22208);
and U22405 (N_22405,N_22397,N_22379);
xor U22406 (N_22406,N_22223,N_22282);
nor U22407 (N_22407,N_22295,N_22225);
xnor U22408 (N_22408,N_22265,N_22211);
and U22409 (N_22409,N_22392,N_22274);
or U22410 (N_22410,N_22219,N_22239);
nor U22411 (N_22411,N_22288,N_22372);
nand U22412 (N_22412,N_22373,N_22244);
nor U22413 (N_22413,N_22259,N_22364);
nor U22414 (N_22414,N_22387,N_22331);
xor U22415 (N_22415,N_22328,N_22354);
and U22416 (N_22416,N_22312,N_22353);
and U22417 (N_22417,N_22386,N_22215);
and U22418 (N_22418,N_22240,N_22252);
and U22419 (N_22419,N_22201,N_22230);
or U22420 (N_22420,N_22281,N_22324);
or U22421 (N_22421,N_22358,N_22227);
nand U22422 (N_22422,N_22224,N_22394);
nand U22423 (N_22423,N_22381,N_22375);
nand U22424 (N_22424,N_22367,N_22299);
and U22425 (N_22425,N_22391,N_22303);
or U22426 (N_22426,N_22356,N_22396);
and U22427 (N_22427,N_22298,N_22280);
nor U22428 (N_22428,N_22256,N_22200);
nor U22429 (N_22429,N_22261,N_22236);
or U22430 (N_22430,N_22220,N_22359);
nor U22431 (N_22431,N_22348,N_22376);
nor U22432 (N_22432,N_22246,N_22306);
and U22433 (N_22433,N_22279,N_22322);
and U22434 (N_22434,N_22234,N_22368);
or U22435 (N_22435,N_22316,N_22320);
nor U22436 (N_22436,N_22339,N_22380);
and U22437 (N_22437,N_22302,N_22271);
or U22438 (N_22438,N_22383,N_22305);
and U22439 (N_22439,N_22267,N_22273);
or U22440 (N_22440,N_22245,N_22300);
nor U22441 (N_22441,N_22366,N_22222);
nor U22442 (N_22442,N_22350,N_22333);
nor U22443 (N_22443,N_22238,N_22241);
and U22444 (N_22444,N_22228,N_22395);
nor U22445 (N_22445,N_22370,N_22361);
xor U22446 (N_22446,N_22317,N_22226);
or U22447 (N_22447,N_22388,N_22291);
nor U22448 (N_22448,N_22263,N_22344);
xor U22449 (N_22449,N_22360,N_22377);
nor U22450 (N_22450,N_22268,N_22275);
nor U22451 (N_22451,N_22218,N_22216);
xor U22452 (N_22452,N_22314,N_22209);
nor U22453 (N_22453,N_22286,N_22311);
nor U22454 (N_22454,N_22293,N_22307);
xor U22455 (N_22455,N_22251,N_22340);
or U22456 (N_22456,N_22231,N_22232);
nand U22457 (N_22457,N_22390,N_22341);
or U22458 (N_22458,N_22315,N_22276);
or U22459 (N_22459,N_22378,N_22389);
nand U22460 (N_22460,N_22229,N_22371);
xor U22461 (N_22461,N_22352,N_22253);
nand U22462 (N_22462,N_22217,N_22334);
xnor U22463 (N_22463,N_22285,N_22235);
xor U22464 (N_22464,N_22205,N_22290);
nand U22465 (N_22465,N_22297,N_22248);
xor U22466 (N_22466,N_22258,N_22342);
and U22467 (N_22467,N_22250,N_22257);
nand U22468 (N_22468,N_22301,N_22351);
or U22469 (N_22469,N_22272,N_22262);
and U22470 (N_22470,N_22332,N_22343);
and U22471 (N_22471,N_22212,N_22336);
or U22472 (N_22472,N_22349,N_22346);
or U22473 (N_22473,N_22269,N_22308);
nand U22474 (N_22474,N_22327,N_22330);
nor U22475 (N_22475,N_22210,N_22335);
or U22476 (N_22476,N_22319,N_22318);
nand U22477 (N_22477,N_22363,N_22321);
xnor U22478 (N_22478,N_22214,N_22393);
nand U22479 (N_22479,N_22362,N_22338);
and U22480 (N_22480,N_22233,N_22398);
nor U22481 (N_22481,N_22255,N_22289);
and U22482 (N_22482,N_22202,N_22384);
nand U22483 (N_22483,N_22292,N_22329);
or U22484 (N_22484,N_22355,N_22247);
nor U22485 (N_22485,N_22357,N_22249);
and U22486 (N_22486,N_22345,N_22264);
and U22487 (N_22487,N_22294,N_22237);
and U22488 (N_22488,N_22242,N_22254);
or U22489 (N_22489,N_22304,N_22326);
nor U22490 (N_22490,N_22399,N_22310);
xor U22491 (N_22491,N_22221,N_22325);
xnor U22492 (N_22492,N_22309,N_22243);
or U22493 (N_22493,N_22369,N_22283);
and U22494 (N_22494,N_22270,N_22374);
nand U22495 (N_22495,N_22287,N_22296);
nor U22496 (N_22496,N_22204,N_22207);
nand U22497 (N_22497,N_22277,N_22266);
or U22498 (N_22498,N_22347,N_22284);
or U22499 (N_22499,N_22382,N_22278);
nand U22500 (N_22500,N_22231,N_22271);
nand U22501 (N_22501,N_22336,N_22273);
nor U22502 (N_22502,N_22334,N_22312);
and U22503 (N_22503,N_22308,N_22368);
nand U22504 (N_22504,N_22358,N_22284);
and U22505 (N_22505,N_22307,N_22383);
or U22506 (N_22506,N_22310,N_22217);
xor U22507 (N_22507,N_22348,N_22216);
or U22508 (N_22508,N_22230,N_22381);
nor U22509 (N_22509,N_22360,N_22346);
nand U22510 (N_22510,N_22374,N_22323);
and U22511 (N_22511,N_22246,N_22335);
xnor U22512 (N_22512,N_22354,N_22393);
nor U22513 (N_22513,N_22276,N_22362);
xnor U22514 (N_22514,N_22251,N_22365);
nand U22515 (N_22515,N_22292,N_22226);
nand U22516 (N_22516,N_22386,N_22342);
nor U22517 (N_22517,N_22206,N_22271);
nor U22518 (N_22518,N_22219,N_22328);
and U22519 (N_22519,N_22240,N_22339);
or U22520 (N_22520,N_22220,N_22327);
xor U22521 (N_22521,N_22384,N_22322);
nor U22522 (N_22522,N_22237,N_22367);
and U22523 (N_22523,N_22218,N_22313);
or U22524 (N_22524,N_22376,N_22323);
xnor U22525 (N_22525,N_22251,N_22381);
xor U22526 (N_22526,N_22391,N_22252);
and U22527 (N_22527,N_22243,N_22298);
xnor U22528 (N_22528,N_22373,N_22222);
and U22529 (N_22529,N_22296,N_22273);
or U22530 (N_22530,N_22398,N_22211);
nand U22531 (N_22531,N_22319,N_22276);
nand U22532 (N_22532,N_22277,N_22216);
nor U22533 (N_22533,N_22348,N_22365);
nand U22534 (N_22534,N_22330,N_22339);
and U22535 (N_22535,N_22296,N_22239);
and U22536 (N_22536,N_22359,N_22391);
xor U22537 (N_22537,N_22366,N_22392);
nand U22538 (N_22538,N_22222,N_22295);
or U22539 (N_22539,N_22211,N_22332);
xor U22540 (N_22540,N_22317,N_22248);
and U22541 (N_22541,N_22358,N_22300);
xnor U22542 (N_22542,N_22244,N_22224);
or U22543 (N_22543,N_22262,N_22296);
xnor U22544 (N_22544,N_22227,N_22383);
xnor U22545 (N_22545,N_22360,N_22216);
nor U22546 (N_22546,N_22223,N_22212);
and U22547 (N_22547,N_22290,N_22303);
and U22548 (N_22548,N_22341,N_22337);
or U22549 (N_22549,N_22243,N_22344);
xnor U22550 (N_22550,N_22360,N_22251);
nor U22551 (N_22551,N_22252,N_22207);
nand U22552 (N_22552,N_22309,N_22379);
nor U22553 (N_22553,N_22228,N_22270);
and U22554 (N_22554,N_22301,N_22362);
xnor U22555 (N_22555,N_22280,N_22278);
nor U22556 (N_22556,N_22357,N_22380);
nand U22557 (N_22557,N_22366,N_22273);
nand U22558 (N_22558,N_22331,N_22266);
and U22559 (N_22559,N_22293,N_22378);
nand U22560 (N_22560,N_22372,N_22237);
nor U22561 (N_22561,N_22278,N_22235);
nor U22562 (N_22562,N_22271,N_22383);
and U22563 (N_22563,N_22273,N_22297);
nand U22564 (N_22564,N_22316,N_22311);
nand U22565 (N_22565,N_22215,N_22345);
or U22566 (N_22566,N_22271,N_22310);
and U22567 (N_22567,N_22246,N_22370);
nor U22568 (N_22568,N_22373,N_22381);
xnor U22569 (N_22569,N_22263,N_22369);
nand U22570 (N_22570,N_22247,N_22269);
xnor U22571 (N_22571,N_22335,N_22234);
xor U22572 (N_22572,N_22241,N_22225);
xor U22573 (N_22573,N_22244,N_22305);
and U22574 (N_22574,N_22359,N_22356);
nand U22575 (N_22575,N_22369,N_22392);
xor U22576 (N_22576,N_22362,N_22313);
nand U22577 (N_22577,N_22232,N_22385);
or U22578 (N_22578,N_22381,N_22252);
xor U22579 (N_22579,N_22264,N_22216);
xnor U22580 (N_22580,N_22353,N_22261);
nor U22581 (N_22581,N_22296,N_22222);
nor U22582 (N_22582,N_22282,N_22201);
nor U22583 (N_22583,N_22303,N_22200);
xnor U22584 (N_22584,N_22263,N_22350);
and U22585 (N_22585,N_22353,N_22255);
and U22586 (N_22586,N_22274,N_22331);
nand U22587 (N_22587,N_22364,N_22354);
nand U22588 (N_22588,N_22357,N_22397);
nor U22589 (N_22589,N_22352,N_22368);
or U22590 (N_22590,N_22328,N_22341);
xor U22591 (N_22591,N_22267,N_22380);
xor U22592 (N_22592,N_22247,N_22287);
xor U22593 (N_22593,N_22275,N_22353);
nand U22594 (N_22594,N_22368,N_22290);
and U22595 (N_22595,N_22304,N_22293);
and U22596 (N_22596,N_22260,N_22390);
nand U22597 (N_22597,N_22211,N_22201);
xor U22598 (N_22598,N_22364,N_22303);
nand U22599 (N_22599,N_22320,N_22329);
xor U22600 (N_22600,N_22535,N_22500);
nand U22601 (N_22601,N_22417,N_22420);
and U22602 (N_22602,N_22528,N_22568);
xor U22603 (N_22603,N_22590,N_22541);
nor U22604 (N_22604,N_22427,N_22518);
or U22605 (N_22605,N_22573,N_22591);
or U22606 (N_22606,N_22524,N_22433);
xnor U22607 (N_22607,N_22428,N_22487);
nand U22608 (N_22608,N_22585,N_22468);
nand U22609 (N_22609,N_22421,N_22509);
nor U22610 (N_22610,N_22526,N_22593);
nor U22611 (N_22611,N_22478,N_22501);
and U22612 (N_22612,N_22533,N_22586);
xnor U22613 (N_22613,N_22592,N_22547);
nand U22614 (N_22614,N_22440,N_22446);
or U22615 (N_22615,N_22424,N_22456);
and U22616 (N_22616,N_22581,N_22466);
nand U22617 (N_22617,N_22572,N_22411);
and U22618 (N_22618,N_22452,N_22574);
nor U22619 (N_22619,N_22447,N_22489);
xor U22620 (N_22620,N_22510,N_22415);
xnor U22621 (N_22621,N_22596,N_22543);
xnor U22622 (N_22622,N_22537,N_22464);
or U22623 (N_22623,N_22463,N_22579);
nand U22624 (N_22624,N_22474,N_22408);
and U22625 (N_22625,N_22546,N_22529);
xnor U22626 (N_22626,N_22584,N_22549);
nand U22627 (N_22627,N_22550,N_22462);
nor U22628 (N_22628,N_22483,N_22407);
nor U22629 (N_22629,N_22517,N_22409);
nor U22630 (N_22630,N_22443,N_22511);
and U22631 (N_22631,N_22454,N_22571);
xnor U22632 (N_22632,N_22522,N_22414);
xnor U22633 (N_22633,N_22540,N_22458);
xnor U22634 (N_22634,N_22558,N_22472);
nor U22635 (N_22635,N_22423,N_22429);
xor U22636 (N_22636,N_22406,N_22453);
and U22637 (N_22637,N_22513,N_22444);
and U22638 (N_22638,N_22476,N_22597);
nand U22639 (N_22639,N_22555,N_22514);
nor U22640 (N_22640,N_22402,N_22479);
and U22641 (N_22641,N_22507,N_22403);
nand U22642 (N_22642,N_22439,N_22565);
or U22643 (N_22643,N_22499,N_22577);
and U22644 (N_22644,N_22416,N_22508);
nor U22645 (N_22645,N_22425,N_22467);
nor U22646 (N_22646,N_22552,N_22490);
and U22647 (N_22647,N_22544,N_22588);
or U22648 (N_22648,N_22548,N_22488);
nor U22649 (N_22649,N_22480,N_22580);
nand U22650 (N_22650,N_22523,N_22494);
nand U22651 (N_22651,N_22595,N_22422);
nor U22652 (N_22652,N_22412,N_22450);
nor U22653 (N_22653,N_22438,N_22471);
nand U22654 (N_22654,N_22562,N_22598);
and U22655 (N_22655,N_22459,N_22451);
and U22656 (N_22656,N_22559,N_22542);
xnor U22657 (N_22657,N_22564,N_22503);
nor U22658 (N_22658,N_22569,N_22538);
nand U22659 (N_22659,N_22437,N_22566);
and U22660 (N_22660,N_22525,N_22469);
and U22661 (N_22661,N_22418,N_22589);
and U22662 (N_22662,N_22401,N_22492);
nor U22663 (N_22663,N_22504,N_22436);
nor U22664 (N_22664,N_22410,N_22495);
xnor U22665 (N_22665,N_22587,N_22570);
xnor U22666 (N_22666,N_22404,N_22455);
or U22667 (N_22667,N_22491,N_22519);
and U22668 (N_22668,N_22553,N_22515);
and U22669 (N_22669,N_22431,N_22485);
xor U22670 (N_22670,N_22400,N_22545);
nand U22671 (N_22671,N_22460,N_22556);
nor U22672 (N_22672,N_22505,N_22516);
xnor U22673 (N_22673,N_22563,N_22521);
xnor U22674 (N_22674,N_22484,N_22434);
xnor U22675 (N_22675,N_22486,N_22497);
nand U22676 (N_22676,N_22578,N_22473);
nand U22677 (N_22677,N_22477,N_22405);
or U22678 (N_22678,N_22534,N_22594);
and U22679 (N_22679,N_22442,N_22430);
or U22680 (N_22680,N_22582,N_22496);
and U22681 (N_22681,N_22512,N_22560);
nand U22682 (N_22682,N_22465,N_22493);
nor U22683 (N_22683,N_22441,N_22498);
nand U22684 (N_22684,N_22536,N_22482);
or U22685 (N_22685,N_22575,N_22432);
or U22686 (N_22686,N_22448,N_22413);
nor U22687 (N_22687,N_22445,N_22475);
and U22688 (N_22688,N_22426,N_22502);
xor U22689 (N_22689,N_22551,N_22530);
xnor U22690 (N_22690,N_22449,N_22557);
nor U22691 (N_22691,N_22539,N_22561);
nand U22692 (N_22692,N_22554,N_22419);
and U22693 (N_22693,N_22567,N_22470);
nand U22694 (N_22694,N_22532,N_22457);
xnor U22695 (N_22695,N_22520,N_22481);
nand U22696 (N_22696,N_22583,N_22527);
xor U22697 (N_22697,N_22461,N_22599);
or U22698 (N_22698,N_22531,N_22576);
and U22699 (N_22699,N_22506,N_22435);
and U22700 (N_22700,N_22535,N_22499);
nand U22701 (N_22701,N_22531,N_22442);
or U22702 (N_22702,N_22503,N_22436);
or U22703 (N_22703,N_22496,N_22491);
nand U22704 (N_22704,N_22511,N_22485);
nand U22705 (N_22705,N_22592,N_22425);
and U22706 (N_22706,N_22550,N_22534);
nand U22707 (N_22707,N_22543,N_22434);
and U22708 (N_22708,N_22515,N_22482);
nand U22709 (N_22709,N_22496,N_22517);
nor U22710 (N_22710,N_22515,N_22578);
xor U22711 (N_22711,N_22464,N_22449);
and U22712 (N_22712,N_22540,N_22497);
and U22713 (N_22713,N_22467,N_22536);
nand U22714 (N_22714,N_22593,N_22569);
or U22715 (N_22715,N_22590,N_22475);
xnor U22716 (N_22716,N_22531,N_22504);
or U22717 (N_22717,N_22479,N_22412);
nand U22718 (N_22718,N_22474,N_22438);
and U22719 (N_22719,N_22469,N_22567);
nand U22720 (N_22720,N_22456,N_22525);
nand U22721 (N_22721,N_22566,N_22587);
or U22722 (N_22722,N_22541,N_22492);
or U22723 (N_22723,N_22574,N_22556);
nor U22724 (N_22724,N_22437,N_22480);
and U22725 (N_22725,N_22451,N_22502);
or U22726 (N_22726,N_22409,N_22479);
nor U22727 (N_22727,N_22493,N_22495);
xor U22728 (N_22728,N_22437,N_22462);
nand U22729 (N_22729,N_22549,N_22534);
nand U22730 (N_22730,N_22413,N_22477);
and U22731 (N_22731,N_22587,N_22544);
or U22732 (N_22732,N_22495,N_22476);
nor U22733 (N_22733,N_22591,N_22547);
nor U22734 (N_22734,N_22470,N_22435);
nor U22735 (N_22735,N_22590,N_22529);
nor U22736 (N_22736,N_22445,N_22581);
nand U22737 (N_22737,N_22569,N_22521);
and U22738 (N_22738,N_22402,N_22593);
nand U22739 (N_22739,N_22577,N_22568);
xor U22740 (N_22740,N_22516,N_22445);
xor U22741 (N_22741,N_22427,N_22420);
and U22742 (N_22742,N_22596,N_22573);
nor U22743 (N_22743,N_22497,N_22474);
nor U22744 (N_22744,N_22457,N_22535);
or U22745 (N_22745,N_22595,N_22588);
nor U22746 (N_22746,N_22434,N_22513);
or U22747 (N_22747,N_22438,N_22560);
or U22748 (N_22748,N_22568,N_22417);
nor U22749 (N_22749,N_22455,N_22416);
or U22750 (N_22750,N_22469,N_22585);
nor U22751 (N_22751,N_22582,N_22414);
xor U22752 (N_22752,N_22511,N_22522);
or U22753 (N_22753,N_22428,N_22486);
or U22754 (N_22754,N_22441,N_22406);
xor U22755 (N_22755,N_22596,N_22408);
or U22756 (N_22756,N_22570,N_22445);
or U22757 (N_22757,N_22568,N_22593);
xor U22758 (N_22758,N_22513,N_22573);
nand U22759 (N_22759,N_22583,N_22599);
nor U22760 (N_22760,N_22497,N_22484);
or U22761 (N_22761,N_22533,N_22410);
or U22762 (N_22762,N_22422,N_22464);
nor U22763 (N_22763,N_22421,N_22427);
xor U22764 (N_22764,N_22429,N_22514);
xor U22765 (N_22765,N_22474,N_22435);
nand U22766 (N_22766,N_22513,N_22479);
nand U22767 (N_22767,N_22561,N_22424);
nor U22768 (N_22768,N_22512,N_22454);
xnor U22769 (N_22769,N_22586,N_22513);
and U22770 (N_22770,N_22493,N_22445);
and U22771 (N_22771,N_22599,N_22571);
and U22772 (N_22772,N_22594,N_22529);
nor U22773 (N_22773,N_22538,N_22556);
nor U22774 (N_22774,N_22456,N_22433);
xor U22775 (N_22775,N_22495,N_22479);
xnor U22776 (N_22776,N_22407,N_22525);
nor U22777 (N_22777,N_22453,N_22512);
xnor U22778 (N_22778,N_22465,N_22450);
nand U22779 (N_22779,N_22493,N_22563);
nor U22780 (N_22780,N_22596,N_22410);
xor U22781 (N_22781,N_22572,N_22494);
nor U22782 (N_22782,N_22505,N_22490);
or U22783 (N_22783,N_22422,N_22548);
xnor U22784 (N_22784,N_22521,N_22430);
or U22785 (N_22785,N_22508,N_22528);
nor U22786 (N_22786,N_22539,N_22589);
xor U22787 (N_22787,N_22452,N_22510);
nor U22788 (N_22788,N_22438,N_22445);
nor U22789 (N_22789,N_22439,N_22487);
and U22790 (N_22790,N_22543,N_22401);
or U22791 (N_22791,N_22468,N_22445);
nand U22792 (N_22792,N_22548,N_22426);
nor U22793 (N_22793,N_22411,N_22578);
nand U22794 (N_22794,N_22455,N_22441);
xnor U22795 (N_22795,N_22578,N_22532);
or U22796 (N_22796,N_22552,N_22454);
and U22797 (N_22797,N_22496,N_22487);
xor U22798 (N_22798,N_22551,N_22474);
and U22799 (N_22799,N_22585,N_22418);
nor U22800 (N_22800,N_22731,N_22666);
nand U22801 (N_22801,N_22707,N_22695);
or U22802 (N_22802,N_22694,N_22661);
xnor U22803 (N_22803,N_22676,N_22613);
nand U22804 (N_22804,N_22644,N_22652);
and U22805 (N_22805,N_22693,N_22785);
and U22806 (N_22806,N_22793,N_22630);
or U22807 (N_22807,N_22679,N_22773);
or U22808 (N_22808,N_22664,N_22637);
nand U22809 (N_22809,N_22635,N_22761);
nand U22810 (N_22810,N_22677,N_22674);
xnor U22811 (N_22811,N_22739,N_22702);
nand U22812 (N_22812,N_22600,N_22659);
nand U22813 (N_22813,N_22604,N_22714);
xor U22814 (N_22814,N_22766,N_22689);
and U22815 (N_22815,N_22625,N_22696);
nand U22816 (N_22816,N_22764,N_22788);
and U22817 (N_22817,N_22723,N_22657);
xnor U22818 (N_22818,N_22701,N_22781);
or U22819 (N_22819,N_22726,N_22720);
or U22820 (N_22820,N_22783,N_22605);
nor U22821 (N_22821,N_22636,N_22607);
and U22822 (N_22822,N_22698,N_22759);
and U22823 (N_22823,N_22757,N_22665);
or U22824 (N_22824,N_22648,N_22735);
nand U22825 (N_22825,N_22794,N_22745);
or U22826 (N_22826,N_22670,N_22712);
xor U22827 (N_22827,N_22634,N_22631);
or U22828 (N_22828,N_22621,N_22615);
and U22829 (N_22829,N_22704,N_22620);
nor U22830 (N_22830,N_22639,N_22612);
nand U22831 (N_22831,N_22705,N_22609);
or U22832 (N_22832,N_22624,N_22688);
nor U22833 (N_22833,N_22775,N_22683);
nand U22834 (N_22834,N_22730,N_22716);
nand U22835 (N_22835,N_22606,N_22741);
nand U22836 (N_22836,N_22654,N_22711);
nand U22837 (N_22837,N_22641,N_22709);
or U22838 (N_22838,N_22697,N_22672);
or U22839 (N_22839,N_22771,N_22673);
nand U22840 (N_22840,N_22601,N_22755);
or U22841 (N_22841,N_22776,N_22645);
or U22842 (N_22842,N_22718,N_22765);
xnor U22843 (N_22843,N_22682,N_22721);
nand U22844 (N_22844,N_22728,N_22749);
nand U22845 (N_22845,N_22792,N_22725);
nand U22846 (N_22846,N_22758,N_22640);
xnor U22847 (N_22847,N_22713,N_22727);
nor U22848 (N_22848,N_22797,N_22602);
nor U22849 (N_22849,N_22633,N_22743);
or U22850 (N_22850,N_22622,N_22710);
xnor U22851 (N_22851,N_22616,N_22778);
or U22852 (N_22852,N_22772,N_22603);
nand U22853 (N_22853,N_22746,N_22732);
nand U22854 (N_22854,N_22717,N_22729);
or U22855 (N_22855,N_22791,N_22687);
or U22856 (N_22856,N_22638,N_22774);
nand U22857 (N_22857,N_22678,N_22692);
nor U22858 (N_22858,N_22686,N_22690);
nand U22859 (N_22859,N_22628,N_22706);
and U22860 (N_22860,N_22782,N_22650);
and U22861 (N_22861,N_22614,N_22660);
nand U22862 (N_22862,N_22653,N_22769);
xnor U22863 (N_22863,N_22667,N_22799);
and U22864 (N_22864,N_22787,N_22617);
nor U22865 (N_22865,N_22647,N_22608);
xnor U22866 (N_22866,N_22681,N_22629);
or U22867 (N_22867,N_22722,N_22632);
or U22868 (N_22868,N_22733,N_22747);
nand U22869 (N_22869,N_22763,N_22724);
xnor U22870 (N_22870,N_22779,N_22751);
xor U22871 (N_22871,N_22626,N_22753);
or U22872 (N_22872,N_22784,N_22643);
or U22873 (N_22873,N_22684,N_22740);
and U22874 (N_22874,N_22744,N_22699);
or U22875 (N_22875,N_22658,N_22685);
xor U22876 (N_22876,N_22703,N_22708);
and U22877 (N_22877,N_22646,N_22796);
nand U22878 (N_22878,N_22790,N_22770);
xnor U22879 (N_22879,N_22669,N_22752);
xnor U22880 (N_22880,N_22627,N_22671);
nor U22881 (N_22881,N_22675,N_22777);
nand U22882 (N_22882,N_22619,N_22668);
xnor U22883 (N_22883,N_22789,N_22662);
and U22884 (N_22884,N_22737,N_22715);
nor U22885 (N_22885,N_22786,N_22610);
nor U22886 (N_22886,N_22623,N_22719);
nand U22887 (N_22887,N_22767,N_22642);
nand U22888 (N_22888,N_22780,N_22768);
nor U22889 (N_22889,N_22734,N_22655);
xnor U22890 (N_22890,N_22680,N_22649);
xor U22891 (N_22891,N_22762,N_22663);
or U22892 (N_22892,N_22700,N_22795);
nand U22893 (N_22893,N_22618,N_22760);
xor U22894 (N_22894,N_22691,N_22651);
xnor U22895 (N_22895,N_22798,N_22742);
nor U22896 (N_22896,N_22611,N_22738);
or U22897 (N_22897,N_22756,N_22750);
or U22898 (N_22898,N_22754,N_22736);
or U22899 (N_22899,N_22748,N_22656);
or U22900 (N_22900,N_22623,N_22695);
xor U22901 (N_22901,N_22757,N_22773);
or U22902 (N_22902,N_22731,N_22699);
and U22903 (N_22903,N_22650,N_22682);
nor U22904 (N_22904,N_22671,N_22799);
nor U22905 (N_22905,N_22624,N_22676);
or U22906 (N_22906,N_22650,N_22790);
nor U22907 (N_22907,N_22764,N_22770);
and U22908 (N_22908,N_22683,N_22685);
xor U22909 (N_22909,N_22769,N_22689);
nand U22910 (N_22910,N_22792,N_22774);
xor U22911 (N_22911,N_22762,N_22688);
or U22912 (N_22912,N_22653,N_22614);
xor U22913 (N_22913,N_22606,N_22665);
and U22914 (N_22914,N_22672,N_22794);
or U22915 (N_22915,N_22644,N_22666);
xnor U22916 (N_22916,N_22643,N_22754);
and U22917 (N_22917,N_22676,N_22622);
xnor U22918 (N_22918,N_22725,N_22668);
nor U22919 (N_22919,N_22783,N_22686);
or U22920 (N_22920,N_22706,N_22616);
nor U22921 (N_22921,N_22736,N_22621);
xor U22922 (N_22922,N_22687,N_22643);
and U22923 (N_22923,N_22730,N_22667);
nor U22924 (N_22924,N_22655,N_22616);
xor U22925 (N_22925,N_22746,N_22716);
nor U22926 (N_22926,N_22671,N_22782);
nor U22927 (N_22927,N_22612,N_22781);
xnor U22928 (N_22928,N_22791,N_22788);
or U22929 (N_22929,N_22676,N_22712);
nor U22930 (N_22930,N_22618,N_22735);
and U22931 (N_22931,N_22635,N_22751);
and U22932 (N_22932,N_22714,N_22603);
or U22933 (N_22933,N_22710,N_22611);
or U22934 (N_22934,N_22722,N_22651);
or U22935 (N_22935,N_22747,N_22765);
and U22936 (N_22936,N_22663,N_22646);
nor U22937 (N_22937,N_22620,N_22651);
or U22938 (N_22938,N_22649,N_22667);
or U22939 (N_22939,N_22783,N_22746);
and U22940 (N_22940,N_22681,N_22791);
and U22941 (N_22941,N_22622,N_22707);
or U22942 (N_22942,N_22700,N_22762);
xnor U22943 (N_22943,N_22674,N_22622);
nor U22944 (N_22944,N_22793,N_22765);
nand U22945 (N_22945,N_22757,N_22723);
nor U22946 (N_22946,N_22722,N_22760);
or U22947 (N_22947,N_22776,N_22770);
nand U22948 (N_22948,N_22696,N_22661);
xor U22949 (N_22949,N_22619,N_22787);
xor U22950 (N_22950,N_22700,N_22613);
nor U22951 (N_22951,N_22739,N_22647);
xor U22952 (N_22952,N_22696,N_22776);
xor U22953 (N_22953,N_22670,N_22619);
or U22954 (N_22954,N_22668,N_22735);
xnor U22955 (N_22955,N_22653,N_22731);
nor U22956 (N_22956,N_22766,N_22704);
nand U22957 (N_22957,N_22712,N_22612);
or U22958 (N_22958,N_22773,N_22739);
and U22959 (N_22959,N_22660,N_22635);
or U22960 (N_22960,N_22698,N_22717);
xor U22961 (N_22961,N_22744,N_22724);
nor U22962 (N_22962,N_22663,N_22603);
or U22963 (N_22963,N_22663,N_22771);
nand U22964 (N_22964,N_22799,N_22744);
nand U22965 (N_22965,N_22675,N_22669);
nor U22966 (N_22966,N_22744,N_22694);
or U22967 (N_22967,N_22638,N_22745);
nor U22968 (N_22968,N_22639,N_22690);
xnor U22969 (N_22969,N_22726,N_22601);
xor U22970 (N_22970,N_22645,N_22671);
xnor U22971 (N_22971,N_22636,N_22606);
nor U22972 (N_22972,N_22787,N_22688);
xnor U22973 (N_22973,N_22730,N_22605);
or U22974 (N_22974,N_22624,N_22605);
and U22975 (N_22975,N_22774,N_22713);
or U22976 (N_22976,N_22608,N_22610);
or U22977 (N_22977,N_22720,N_22636);
or U22978 (N_22978,N_22617,N_22611);
or U22979 (N_22979,N_22711,N_22616);
and U22980 (N_22980,N_22701,N_22648);
xor U22981 (N_22981,N_22734,N_22750);
xnor U22982 (N_22982,N_22664,N_22749);
nor U22983 (N_22983,N_22627,N_22729);
and U22984 (N_22984,N_22744,N_22738);
nand U22985 (N_22985,N_22703,N_22735);
and U22986 (N_22986,N_22776,N_22740);
nor U22987 (N_22987,N_22727,N_22629);
xor U22988 (N_22988,N_22677,N_22622);
xnor U22989 (N_22989,N_22761,N_22799);
nand U22990 (N_22990,N_22652,N_22766);
or U22991 (N_22991,N_22679,N_22685);
and U22992 (N_22992,N_22797,N_22768);
or U22993 (N_22993,N_22766,N_22682);
nand U22994 (N_22994,N_22638,N_22601);
or U22995 (N_22995,N_22648,N_22723);
and U22996 (N_22996,N_22698,N_22608);
nor U22997 (N_22997,N_22783,N_22778);
xor U22998 (N_22998,N_22760,N_22690);
nor U22999 (N_22999,N_22734,N_22633);
and U23000 (N_23000,N_22922,N_22878);
nand U23001 (N_23001,N_22903,N_22951);
or U23002 (N_23002,N_22916,N_22861);
nand U23003 (N_23003,N_22843,N_22906);
and U23004 (N_23004,N_22968,N_22883);
or U23005 (N_23005,N_22858,N_22945);
nor U23006 (N_23006,N_22831,N_22868);
nor U23007 (N_23007,N_22851,N_22876);
xor U23008 (N_23008,N_22840,N_22897);
xor U23009 (N_23009,N_22869,N_22873);
xnor U23010 (N_23010,N_22854,N_22904);
nor U23011 (N_23011,N_22894,N_22834);
and U23012 (N_23012,N_22957,N_22862);
and U23013 (N_23013,N_22847,N_22935);
and U23014 (N_23014,N_22824,N_22817);
nor U23015 (N_23015,N_22888,N_22837);
or U23016 (N_23016,N_22812,N_22933);
nor U23017 (N_23017,N_22956,N_22838);
or U23018 (N_23018,N_22971,N_22908);
and U23019 (N_23019,N_22842,N_22885);
and U23020 (N_23020,N_22990,N_22928);
nand U23021 (N_23021,N_22926,N_22895);
xor U23022 (N_23022,N_22949,N_22932);
xnor U23023 (N_23023,N_22818,N_22921);
nor U23024 (N_23024,N_22811,N_22911);
or U23025 (N_23025,N_22986,N_22820);
and U23026 (N_23026,N_22823,N_22961);
nand U23027 (N_23027,N_22970,N_22808);
xnor U23028 (N_23028,N_22844,N_22856);
and U23029 (N_23029,N_22942,N_22985);
and U23030 (N_23030,N_22946,N_22972);
nor U23031 (N_23031,N_22827,N_22890);
or U23032 (N_23032,N_22919,N_22828);
and U23033 (N_23033,N_22874,N_22999);
nor U23034 (N_23034,N_22802,N_22830);
or U23035 (N_23035,N_22886,N_22845);
or U23036 (N_23036,N_22816,N_22966);
nand U23037 (N_23037,N_22965,N_22998);
xnor U23038 (N_23038,N_22829,N_22804);
nand U23039 (N_23039,N_22898,N_22944);
nor U23040 (N_23040,N_22953,N_22914);
xnor U23041 (N_23041,N_22870,N_22963);
or U23042 (N_23042,N_22969,N_22880);
nor U23043 (N_23043,N_22836,N_22989);
xor U23044 (N_23044,N_22887,N_22825);
and U23045 (N_23045,N_22846,N_22979);
or U23046 (N_23046,N_22915,N_22934);
nand U23047 (N_23047,N_22841,N_22967);
nor U23048 (N_23048,N_22864,N_22987);
nor U23049 (N_23049,N_22991,N_22884);
nand U23050 (N_23050,N_22859,N_22850);
nand U23051 (N_23051,N_22832,N_22980);
nor U23052 (N_23052,N_22924,N_22923);
or U23053 (N_23053,N_22994,N_22964);
nand U23054 (N_23054,N_22978,N_22867);
xor U23055 (N_23055,N_22900,N_22974);
nand U23056 (N_23056,N_22940,N_22973);
xor U23057 (N_23057,N_22930,N_22819);
nand U23058 (N_23058,N_22893,N_22860);
or U23059 (N_23059,N_22981,N_22917);
nor U23060 (N_23060,N_22805,N_22835);
xor U23061 (N_23061,N_22954,N_22849);
or U23062 (N_23062,N_22905,N_22902);
and U23063 (N_23063,N_22803,N_22892);
nor U23064 (N_23064,N_22976,N_22992);
and U23065 (N_23065,N_22800,N_22826);
nor U23066 (N_23066,N_22814,N_22807);
nor U23067 (N_23067,N_22853,N_22806);
nand U23068 (N_23068,N_22815,N_22996);
nand U23069 (N_23069,N_22863,N_22855);
nor U23070 (N_23070,N_22848,N_22983);
nand U23071 (N_23071,N_22913,N_22857);
and U23072 (N_23072,N_22889,N_22901);
nor U23073 (N_23073,N_22907,N_22960);
xor U23074 (N_23074,N_22984,N_22821);
nor U23075 (N_23075,N_22950,N_22877);
or U23076 (N_23076,N_22822,N_22918);
or U23077 (N_23077,N_22959,N_22801);
nand U23078 (N_23078,N_22982,N_22955);
xor U23079 (N_23079,N_22937,N_22912);
and U23080 (N_23080,N_22852,N_22993);
nand U23081 (N_23081,N_22941,N_22962);
nor U23082 (N_23082,N_22997,N_22975);
xor U23083 (N_23083,N_22939,N_22810);
xor U23084 (N_23084,N_22943,N_22875);
nand U23085 (N_23085,N_22833,N_22925);
nand U23086 (N_23086,N_22910,N_22977);
nand U23087 (N_23087,N_22995,N_22881);
or U23088 (N_23088,N_22866,N_22865);
or U23089 (N_23089,N_22871,N_22891);
or U23090 (N_23090,N_22938,N_22879);
or U23091 (N_23091,N_22813,N_22929);
xnor U23092 (N_23092,N_22931,N_22988);
nor U23093 (N_23093,N_22899,N_22882);
xnor U23094 (N_23094,N_22936,N_22952);
nand U23095 (N_23095,N_22839,N_22920);
nand U23096 (N_23096,N_22809,N_22958);
and U23097 (N_23097,N_22947,N_22896);
nor U23098 (N_23098,N_22872,N_22927);
or U23099 (N_23099,N_22948,N_22909);
or U23100 (N_23100,N_22930,N_22862);
nor U23101 (N_23101,N_22978,N_22880);
nand U23102 (N_23102,N_22900,N_22822);
and U23103 (N_23103,N_22985,N_22821);
nand U23104 (N_23104,N_22956,N_22964);
nand U23105 (N_23105,N_22923,N_22893);
or U23106 (N_23106,N_22836,N_22946);
or U23107 (N_23107,N_22875,N_22820);
nand U23108 (N_23108,N_22871,N_22942);
nor U23109 (N_23109,N_22943,N_22862);
or U23110 (N_23110,N_22847,N_22891);
or U23111 (N_23111,N_22802,N_22883);
or U23112 (N_23112,N_22862,N_22949);
nor U23113 (N_23113,N_22931,N_22994);
and U23114 (N_23114,N_22852,N_22934);
nand U23115 (N_23115,N_22879,N_22980);
nor U23116 (N_23116,N_22972,N_22917);
nor U23117 (N_23117,N_22952,N_22977);
nor U23118 (N_23118,N_22937,N_22860);
nand U23119 (N_23119,N_22813,N_22811);
nand U23120 (N_23120,N_22800,N_22824);
and U23121 (N_23121,N_22923,N_22950);
nand U23122 (N_23122,N_22809,N_22887);
nor U23123 (N_23123,N_22993,N_22801);
nor U23124 (N_23124,N_22978,N_22930);
nor U23125 (N_23125,N_22993,N_22967);
xor U23126 (N_23126,N_22949,N_22885);
xnor U23127 (N_23127,N_22997,N_22892);
nor U23128 (N_23128,N_22893,N_22925);
or U23129 (N_23129,N_22928,N_22915);
xor U23130 (N_23130,N_22947,N_22836);
nor U23131 (N_23131,N_22952,N_22931);
xnor U23132 (N_23132,N_22968,N_22963);
and U23133 (N_23133,N_22950,N_22894);
or U23134 (N_23134,N_22844,N_22880);
xor U23135 (N_23135,N_22982,N_22851);
nand U23136 (N_23136,N_22929,N_22828);
nand U23137 (N_23137,N_22847,N_22802);
and U23138 (N_23138,N_22819,N_22811);
nor U23139 (N_23139,N_22864,N_22806);
xnor U23140 (N_23140,N_22891,N_22962);
or U23141 (N_23141,N_22934,N_22820);
and U23142 (N_23142,N_22973,N_22853);
or U23143 (N_23143,N_22936,N_22972);
xnor U23144 (N_23144,N_22941,N_22925);
and U23145 (N_23145,N_22822,N_22930);
or U23146 (N_23146,N_22941,N_22875);
nor U23147 (N_23147,N_22936,N_22941);
nand U23148 (N_23148,N_22870,N_22950);
and U23149 (N_23149,N_22834,N_22949);
or U23150 (N_23150,N_22902,N_22848);
or U23151 (N_23151,N_22836,N_22810);
or U23152 (N_23152,N_22818,N_22904);
xor U23153 (N_23153,N_22847,N_22998);
nor U23154 (N_23154,N_22855,N_22824);
or U23155 (N_23155,N_22826,N_22991);
and U23156 (N_23156,N_22983,N_22880);
or U23157 (N_23157,N_22905,N_22953);
nand U23158 (N_23158,N_22928,N_22955);
nor U23159 (N_23159,N_22925,N_22892);
nand U23160 (N_23160,N_22882,N_22987);
xnor U23161 (N_23161,N_22969,N_22803);
xor U23162 (N_23162,N_22936,N_22915);
and U23163 (N_23163,N_22821,N_22891);
xnor U23164 (N_23164,N_22812,N_22822);
or U23165 (N_23165,N_22914,N_22969);
and U23166 (N_23166,N_22988,N_22896);
nor U23167 (N_23167,N_22865,N_22902);
nor U23168 (N_23168,N_22822,N_22992);
xor U23169 (N_23169,N_22946,N_22986);
nor U23170 (N_23170,N_22937,N_22925);
nor U23171 (N_23171,N_22834,N_22820);
or U23172 (N_23172,N_22894,N_22911);
xnor U23173 (N_23173,N_22813,N_22949);
xnor U23174 (N_23174,N_22880,N_22836);
xor U23175 (N_23175,N_22861,N_22993);
xnor U23176 (N_23176,N_22804,N_22916);
or U23177 (N_23177,N_22870,N_22936);
nor U23178 (N_23178,N_22824,N_22869);
and U23179 (N_23179,N_22869,N_22863);
nor U23180 (N_23180,N_22981,N_22857);
nor U23181 (N_23181,N_22898,N_22810);
or U23182 (N_23182,N_22949,N_22973);
nand U23183 (N_23183,N_22871,N_22973);
and U23184 (N_23184,N_22842,N_22890);
nand U23185 (N_23185,N_22944,N_22849);
or U23186 (N_23186,N_22841,N_22961);
and U23187 (N_23187,N_22987,N_22920);
nand U23188 (N_23188,N_22949,N_22894);
or U23189 (N_23189,N_22933,N_22929);
and U23190 (N_23190,N_22995,N_22867);
nand U23191 (N_23191,N_22801,N_22846);
nand U23192 (N_23192,N_22871,N_22850);
nand U23193 (N_23193,N_22858,N_22873);
and U23194 (N_23194,N_22948,N_22838);
and U23195 (N_23195,N_22936,N_22812);
nand U23196 (N_23196,N_22938,N_22968);
or U23197 (N_23197,N_22842,N_22902);
xor U23198 (N_23198,N_22944,N_22821);
or U23199 (N_23199,N_22957,N_22994);
nor U23200 (N_23200,N_23159,N_23162);
nand U23201 (N_23201,N_23099,N_23060);
and U23202 (N_23202,N_23116,N_23119);
nor U23203 (N_23203,N_23141,N_23085);
nand U23204 (N_23204,N_23192,N_23071);
nor U23205 (N_23205,N_23164,N_23024);
nor U23206 (N_23206,N_23032,N_23165);
nand U23207 (N_23207,N_23109,N_23007);
xnor U23208 (N_23208,N_23076,N_23149);
and U23209 (N_23209,N_23057,N_23104);
nor U23210 (N_23210,N_23087,N_23114);
or U23211 (N_23211,N_23118,N_23144);
nor U23212 (N_23212,N_23124,N_23137);
or U23213 (N_23213,N_23107,N_23133);
nor U23214 (N_23214,N_23061,N_23058);
or U23215 (N_23215,N_23113,N_23028);
nand U23216 (N_23216,N_23129,N_23139);
and U23217 (N_23217,N_23054,N_23105);
nand U23218 (N_23218,N_23095,N_23112);
and U23219 (N_23219,N_23140,N_23166);
xnor U23220 (N_23220,N_23169,N_23163);
nand U23221 (N_23221,N_23182,N_23186);
or U23222 (N_23222,N_23016,N_23046);
xor U23223 (N_23223,N_23147,N_23062);
and U23224 (N_23224,N_23027,N_23185);
xnor U23225 (N_23225,N_23089,N_23083);
and U23226 (N_23226,N_23088,N_23020);
nand U23227 (N_23227,N_23100,N_23151);
or U23228 (N_23228,N_23050,N_23036);
or U23229 (N_23229,N_23106,N_23053);
or U23230 (N_23230,N_23191,N_23037);
nand U23231 (N_23231,N_23115,N_23157);
nand U23232 (N_23232,N_23011,N_23065);
xor U23233 (N_23233,N_23148,N_23193);
xor U23234 (N_23234,N_23091,N_23030);
and U23235 (N_23235,N_23097,N_23103);
or U23236 (N_23236,N_23029,N_23072);
and U23237 (N_23237,N_23015,N_23023);
and U23238 (N_23238,N_23063,N_23171);
xor U23239 (N_23239,N_23123,N_23013);
nand U23240 (N_23240,N_23194,N_23008);
nor U23241 (N_23241,N_23174,N_23045);
and U23242 (N_23242,N_23128,N_23012);
xnor U23243 (N_23243,N_23134,N_23146);
and U23244 (N_23244,N_23073,N_23075);
nor U23245 (N_23245,N_23096,N_23183);
or U23246 (N_23246,N_23077,N_23035);
and U23247 (N_23247,N_23055,N_23040);
nor U23248 (N_23248,N_23160,N_23066);
or U23249 (N_23249,N_23181,N_23189);
nor U23250 (N_23250,N_23130,N_23158);
xor U23251 (N_23251,N_23131,N_23017);
and U23252 (N_23252,N_23051,N_23120);
or U23253 (N_23253,N_23003,N_23168);
or U23254 (N_23254,N_23167,N_23180);
or U23255 (N_23255,N_23086,N_23000);
nor U23256 (N_23256,N_23173,N_23143);
and U23257 (N_23257,N_23154,N_23177);
nor U23258 (N_23258,N_23047,N_23111);
nor U23259 (N_23259,N_23197,N_23175);
nor U23260 (N_23260,N_23138,N_23110);
or U23261 (N_23261,N_23127,N_23042);
nor U23262 (N_23262,N_23067,N_23125);
or U23263 (N_23263,N_23102,N_23018);
and U23264 (N_23264,N_23108,N_23092);
xnor U23265 (N_23265,N_23025,N_23005);
nor U23266 (N_23266,N_23082,N_23049);
nor U23267 (N_23267,N_23198,N_23084);
and U23268 (N_23268,N_23121,N_23033);
nand U23269 (N_23269,N_23039,N_23135);
or U23270 (N_23270,N_23142,N_23009);
or U23271 (N_23271,N_23064,N_23031);
xnor U23272 (N_23272,N_23021,N_23122);
xnor U23273 (N_23273,N_23172,N_23152);
nand U23274 (N_23274,N_23044,N_23019);
or U23275 (N_23275,N_23070,N_23014);
nor U23276 (N_23276,N_23170,N_23093);
or U23277 (N_23277,N_23199,N_23145);
nor U23278 (N_23278,N_23034,N_23136);
nor U23279 (N_23279,N_23190,N_23074);
nand U23280 (N_23280,N_23187,N_23078);
nand U23281 (N_23281,N_23069,N_23038);
and U23282 (N_23282,N_23188,N_23068);
nor U23283 (N_23283,N_23001,N_23079);
xnor U23284 (N_23284,N_23090,N_23196);
or U23285 (N_23285,N_23081,N_23150);
or U23286 (N_23286,N_23094,N_23126);
nor U23287 (N_23287,N_23002,N_23153);
nor U23288 (N_23288,N_23117,N_23052);
nor U23289 (N_23289,N_23006,N_23179);
and U23290 (N_23290,N_23184,N_23080);
nand U23291 (N_23291,N_23176,N_23195);
nor U23292 (N_23292,N_23098,N_23156);
and U23293 (N_23293,N_23048,N_23026);
xor U23294 (N_23294,N_23041,N_23004);
nor U23295 (N_23295,N_23101,N_23022);
xor U23296 (N_23296,N_23056,N_23043);
xnor U23297 (N_23297,N_23178,N_23155);
or U23298 (N_23298,N_23010,N_23059);
nand U23299 (N_23299,N_23132,N_23161);
or U23300 (N_23300,N_23056,N_23030);
nor U23301 (N_23301,N_23180,N_23176);
or U23302 (N_23302,N_23129,N_23183);
and U23303 (N_23303,N_23176,N_23062);
or U23304 (N_23304,N_23156,N_23147);
xor U23305 (N_23305,N_23095,N_23008);
and U23306 (N_23306,N_23038,N_23145);
nor U23307 (N_23307,N_23117,N_23109);
nor U23308 (N_23308,N_23185,N_23022);
and U23309 (N_23309,N_23032,N_23077);
and U23310 (N_23310,N_23160,N_23025);
nor U23311 (N_23311,N_23109,N_23091);
and U23312 (N_23312,N_23081,N_23034);
nor U23313 (N_23313,N_23043,N_23131);
xor U23314 (N_23314,N_23144,N_23122);
and U23315 (N_23315,N_23150,N_23043);
xnor U23316 (N_23316,N_23009,N_23014);
nor U23317 (N_23317,N_23054,N_23126);
xor U23318 (N_23318,N_23086,N_23056);
nand U23319 (N_23319,N_23008,N_23093);
xor U23320 (N_23320,N_23076,N_23162);
nor U23321 (N_23321,N_23152,N_23138);
and U23322 (N_23322,N_23178,N_23139);
and U23323 (N_23323,N_23033,N_23040);
nand U23324 (N_23324,N_23181,N_23138);
nor U23325 (N_23325,N_23060,N_23096);
or U23326 (N_23326,N_23022,N_23105);
nor U23327 (N_23327,N_23034,N_23005);
and U23328 (N_23328,N_23192,N_23135);
and U23329 (N_23329,N_23157,N_23006);
xnor U23330 (N_23330,N_23111,N_23133);
xor U23331 (N_23331,N_23199,N_23189);
nand U23332 (N_23332,N_23082,N_23053);
and U23333 (N_23333,N_23001,N_23182);
nand U23334 (N_23334,N_23076,N_23034);
nand U23335 (N_23335,N_23074,N_23118);
nor U23336 (N_23336,N_23190,N_23126);
xnor U23337 (N_23337,N_23167,N_23022);
xor U23338 (N_23338,N_23168,N_23153);
nand U23339 (N_23339,N_23117,N_23196);
and U23340 (N_23340,N_23068,N_23084);
and U23341 (N_23341,N_23096,N_23070);
nand U23342 (N_23342,N_23049,N_23062);
xnor U23343 (N_23343,N_23004,N_23044);
and U23344 (N_23344,N_23068,N_23118);
nand U23345 (N_23345,N_23170,N_23148);
nand U23346 (N_23346,N_23148,N_23027);
xor U23347 (N_23347,N_23048,N_23057);
or U23348 (N_23348,N_23041,N_23073);
xor U23349 (N_23349,N_23071,N_23122);
and U23350 (N_23350,N_23102,N_23024);
and U23351 (N_23351,N_23067,N_23135);
and U23352 (N_23352,N_23158,N_23045);
nand U23353 (N_23353,N_23066,N_23030);
and U23354 (N_23354,N_23050,N_23154);
nor U23355 (N_23355,N_23143,N_23013);
or U23356 (N_23356,N_23178,N_23101);
xor U23357 (N_23357,N_23145,N_23036);
or U23358 (N_23358,N_23033,N_23151);
or U23359 (N_23359,N_23072,N_23031);
or U23360 (N_23360,N_23102,N_23038);
nor U23361 (N_23361,N_23058,N_23076);
nor U23362 (N_23362,N_23056,N_23174);
xor U23363 (N_23363,N_23041,N_23103);
nand U23364 (N_23364,N_23138,N_23014);
or U23365 (N_23365,N_23102,N_23161);
or U23366 (N_23366,N_23138,N_23047);
and U23367 (N_23367,N_23186,N_23084);
nand U23368 (N_23368,N_23070,N_23079);
or U23369 (N_23369,N_23015,N_23109);
nand U23370 (N_23370,N_23071,N_23041);
and U23371 (N_23371,N_23068,N_23018);
nand U23372 (N_23372,N_23180,N_23066);
and U23373 (N_23373,N_23043,N_23177);
nor U23374 (N_23374,N_23112,N_23010);
or U23375 (N_23375,N_23176,N_23015);
nor U23376 (N_23376,N_23123,N_23141);
nand U23377 (N_23377,N_23078,N_23114);
nor U23378 (N_23378,N_23120,N_23044);
xnor U23379 (N_23379,N_23191,N_23087);
nor U23380 (N_23380,N_23180,N_23033);
xnor U23381 (N_23381,N_23121,N_23129);
xnor U23382 (N_23382,N_23039,N_23099);
or U23383 (N_23383,N_23184,N_23116);
nand U23384 (N_23384,N_23161,N_23159);
and U23385 (N_23385,N_23011,N_23004);
and U23386 (N_23386,N_23162,N_23160);
or U23387 (N_23387,N_23011,N_23057);
nor U23388 (N_23388,N_23042,N_23059);
nor U23389 (N_23389,N_23098,N_23090);
and U23390 (N_23390,N_23039,N_23013);
nor U23391 (N_23391,N_23057,N_23114);
or U23392 (N_23392,N_23143,N_23040);
and U23393 (N_23393,N_23144,N_23002);
nand U23394 (N_23394,N_23090,N_23150);
xnor U23395 (N_23395,N_23029,N_23107);
nand U23396 (N_23396,N_23020,N_23070);
or U23397 (N_23397,N_23185,N_23189);
and U23398 (N_23398,N_23139,N_23155);
xnor U23399 (N_23399,N_23010,N_23113);
nand U23400 (N_23400,N_23392,N_23324);
nand U23401 (N_23401,N_23266,N_23245);
xor U23402 (N_23402,N_23312,N_23293);
or U23403 (N_23403,N_23378,N_23387);
xnor U23404 (N_23404,N_23320,N_23232);
xnor U23405 (N_23405,N_23230,N_23244);
nand U23406 (N_23406,N_23253,N_23247);
xnor U23407 (N_23407,N_23398,N_23295);
and U23408 (N_23408,N_23305,N_23338);
and U23409 (N_23409,N_23233,N_23348);
and U23410 (N_23410,N_23228,N_23306);
and U23411 (N_23411,N_23269,N_23379);
and U23412 (N_23412,N_23214,N_23393);
xor U23413 (N_23413,N_23291,N_23208);
xor U23414 (N_23414,N_23209,N_23224);
nand U23415 (N_23415,N_23268,N_23328);
nor U23416 (N_23416,N_23376,N_23234);
and U23417 (N_23417,N_23263,N_23221);
or U23418 (N_23418,N_23301,N_23210);
nand U23419 (N_23419,N_23369,N_23389);
and U23420 (N_23420,N_23396,N_23300);
nor U23421 (N_23421,N_23342,N_23215);
nand U23422 (N_23422,N_23202,N_23226);
or U23423 (N_23423,N_23397,N_23371);
xor U23424 (N_23424,N_23279,N_23203);
or U23425 (N_23425,N_23211,N_23345);
or U23426 (N_23426,N_23283,N_23204);
nand U23427 (N_23427,N_23256,N_23351);
and U23428 (N_23428,N_23257,N_23331);
and U23429 (N_23429,N_23260,N_23304);
nor U23430 (N_23430,N_23242,N_23274);
nor U23431 (N_23431,N_23217,N_23358);
nor U23432 (N_23432,N_23282,N_23354);
nor U23433 (N_23433,N_23308,N_23325);
or U23434 (N_23434,N_23319,N_23243);
nor U23435 (N_23435,N_23276,N_23307);
or U23436 (N_23436,N_23288,N_23265);
nor U23437 (N_23437,N_23363,N_23316);
or U23438 (N_23438,N_23380,N_23314);
xor U23439 (N_23439,N_23362,N_23258);
nand U23440 (N_23440,N_23322,N_23366);
nand U23441 (N_23441,N_23240,N_23361);
and U23442 (N_23442,N_23241,N_23278);
nand U23443 (N_23443,N_23273,N_23235);
or U23444 (N_23444,N_23332,N_23231);
xor U23445 (N_23445,N_23277,N_23333);
or U23446 (N_23446,N_23252,N_23310);
xnor U23447 (N_23447,N_23355,N_23374);
or U23448 (N_23448,N_23286,N_23311);
and U23449 (N_23449,N_23329,N_23299);
and U23450 (N_23450,N_23343,N_23254);
nand U23451 (N_23451,N_23272,N_23297);
nand U23452 (N_23452,N_23349,N_23261);
or U23453 (N_23453,N_23386,N_23302);
nand U23454 (N_23454,N_23384,N_23394);
nand U23455 (N_23455,N_23359,N_23372);
or U23456 (N_23456,N_23216,N_23227);
nand U23457 (N_23457,N_23340,N_23367);
xor U23458 (N_23458,N_23284,N_23344);
xor U23459 (N_23459,N_23287,N_23236);
or U23460 (N_23460,N_23303,N_23341);
nand U23461 (N_23461,N_23205,N_23270);
nand U23462 (N_23462,N_23326,N_23220);
xor U23463 (N_23463,N_23225,N_23330);
xnor U23464 (N_23464,N_23296,N_23370);
nand U23465 (N_23465,N_23289,N_23334);
xnor U23466 (N_23466,N_23201,N_23381);
xnor U23467 (N_23467,N_23388,N_23347);
nor U23468 (N_23468,N_23360,N_23375);
xor U23469 (N_23469,N_23391,N_23364);
or U23470 (N_23470,N_23327,N_23281);
nor U23471 (N_23471,N_23238,N_23353);
xor U23472 (N_23472,N_23346,N_23222);
nor U23473 (N_23473,N_23382,N_23350);
nor U23474 (N_23474,N_23294,N_23280);
nand U23475 (N_23475,N_23352,N_23219);
nor U23476 (N_23476,N_23356,N_23390);
or U23477 (N_23477,N_23317,N_23218);
or U23478 (N_23478,N_23239,N_23250);
nor U23479 (N_23479,N_23290,N_23323);
nand U23480 (N_23480,N_23251,N_23259);
nand U23481 (N_23481,N_23377,N_23249);
nor U23482 (N_23482,N_23212,N_23385);
xor U23483 (N_23483,N_23335,N_23336);
nor U23484 (N_23484,N_23267,N_23207);
nand U23485 (N_23485,N_23365,N_23339);
and U23486 (N_23486,N_23368,N_23262);
nor U23487 (N_23487,N_23275,N_23399);
and U23488 (N_23488,N_23298,N_23285);
nor U23489 (N_23489,N_23264,N_23313);
and U23490 (N_23490,N_23206,N_23292);
xnor U23491 (N_23491,N_23223,N_23321);
xor U23492 (N_23492,N_23337,N_23357);
or U23493 (N_23493,N_23200,N_23318);
or U23494 (N_23494,N_23383,N_23271);
xor U23495 (N_23495,N_23248,N_23255);
and U23496 (N_23496,N_23395,N_23213);
and U23497 (N_23497,N_23229,N_23315);
nor U23498 (N_23498,N_23309,N_23373);
xor U23499 (N_23499,N_23246,N_23237);
xor U23500 (N_23500,N_23301,N_23328);
xor U23501 (N_23501,N_23306,N_23385);
or U23502 (N_23502,N_23360,N_23332);
or U23503 (N_23503,N_23335,N_23219);
or U23504 (N_23504,N_23250,N_23335);
and U23505 (N_23505,N_23395,N_23320);
and U23506 (N_23506,N_23387,N_23381);
or U23507 (N_23507,N_23240,N_23367);
or U23508 (N_23508,N_23329,N_23231);
and U23509 (N_23509,N_23363,N_23274);
nand U23510 (N_23510,N_23355,N_23251);
nand U23511 (N_23511,N_23233,N_23360);
and U23512 (N_23512,N_23254,N_23315);
and U23513 (N_23513,N_23313,N_23293);
nor U23514 (N_23514,N_23240,N_23315);
nor U23515 (N_23515,N_23265,N_23230);
and U23516 (N_23516,N_23279,N_23359);
or U23517 (N_23517,N_23238,N_23339);
and U23518 (N_23518,N_23374,N_23219);
and U23519 (N_23519,N_23317,N_23375);
nor U23520 (N_23520,N_23359,N_23274);
xnor U23521 (N_23521,N_23323,N_23310);
nor U23522 (N_23522,N_23221,N_23273);
nor U23523 (N_23523,N_23214,N_23326);
nand U23524 (N_23524,N_23357,N_23222);
and U23525 (N_23525,N_23221,N_23286);
nand U23526 (N_23526,N_23294,N_23278);
nand U23527 (N_23527,N_23367,N_23238);
and U23528 (N_23528,N_23244,N_23294);
nor U23529 (N_23529,N_23364,N_23378);
nand U23530 (N_23530,N_23207,N_23373);
or U23531 (N_23531,N_23260,N_23315);
nor U23532 (N_23532,N_23323,N_23376);
or U23533 (N_23533,N_23223,N_23349);
nor U23534 (N_23534,N_23396,N_23320);
xnor U23535 (N_23535,N_23267,N_23273);
nor U23536 (N_23536,N_23287,N_23274);
and U23537 (N_23537,N_23324,N_23306);
and U23538 (N_23538,N_23326,N_23370);
nor U23539 (N_23539,N_23323,N_23210);
nand U23540 (N_23540,N_23376,N_23213);
nand U23541 (N_23541,N_23374,N_23232);
nor U23542 (N_23542,N_23369,N_23336);
or U23543 (N_23543,N_23364,N_23300);
xor U23544 (N_23544,N_23270,N_23279);
xor U23545 (N_23545,N_23205,N_23220);
xor U23546 (N_23546,N_23364,N_23287);
or U23547 (N_23547,N_23222,N_23368);
xor U23548 (N_23548,N_23236,N_23322);
and U23549 (N_23549,N_23355,N_23295);
and U23550 (N_23550,N_23219,N_23310);
nor U23551 (N_23551,N_23222,N_23260);
nor U23552 (N_23552,N_23339,N_23289);
nor U23553 (N_23553,N_23266,N_23344);
xnor U23554 (N_23554,N_23369,N_23257);
nand U23555 (N_23555,N_23389,N_23338);
or U23556 (N_23556,N_23241,N_23284);
or U23557 (N_23557,N_23256,N_23337);
or U23558 (N_23558,N_23368,N_23315);
xnor U23559 (N_23559,N_23384,N_23269);
xnor U23560 (N_23560,N_23352,N_23269);
or U23561 (N_23561,N_23293,N_23365);
or U23562 (N_23562,N_23241,N_23343);
xnor U23563 (N_23563,N_23217,N_23352);
nor U23564 (N_23564,N_23353,N_23347);
xor U23565 (N_23565,N_23215,N_23236);
and U23566 (N_23566,N_23203,N_23211);
or U23567 (N_23567,N_23300,N_23272);
or U23568 (N_23568,N_23259,N_23213);
and U23569 (N_23569,N_23306,N_23323);
xnor U23570 (N_23570,N_23393,N_23368);
or U23571 (N_23571,N_23231,N_23398);
or U23572 (N_23572,N_23298,N_23357);
and U23573 (N_23573,N_23374,N_23302);
nand U23574 (N_23574,N_23392,N_23270);
nor U23575 (N_23575,N_23375,N_23382);
nand U23576 (N_23576,N_23201,N_23383);
xor U23577 (N_23577,N_23265,N_23271);
nand U23578 (N_23578,N_23213,N_23277);
or U23579 (N_23579,N_23399,N_23243);
xor U23580 (N_23580,N_23391,N_23256);
xnor U23581 (N_23581,N_23363,N_23383);
xnor U23582 (N_23582,N_23363,N_23336);
nor U23583 (N_23583,N_23282,N_23205);
nand U23584 (N_23584,N_23275,N_23363);
or U23585 (N_23585,N_23290,N_23236);
and U23586 (N_23586,N_23396,N_23282);
or U23587 (N_23587,N_23213,N_23297);
or U23588 (N_23588,N_23363,N_23217);
and U23589 (N_23589,N_23308,N_23218);
or U23590 (N_23590,N_23323,N_23361);
nor U23591 (N_23591,N_23227,N_23385);
and U23592 (N_23592,N_23380,N_23384);
nand U23593 (N_23593,N_23303,N_23236);
and U23594 (N_23594,N_23393,N_23384);
xnor U23595 (N_23595,N_23368,N_23273);
or U23596 (N_23596,N_23346,N_23319);
nand U23597 (N_23597,N_23210,N_23366);
nand U23598 (N_23598,N_23209,N_23202);
nor U23599 (N_23599,N_23317,N_23269);
or U23600 (N_23600,N_23559,N_23414);
xnor U23601 (N_23601,N_23532,N_23522);
or U23602 (N_23602,N_23549,N_23484);
or U23603 (N_23603,N_23579,N_23431);
nand U23604 (N_23604,N_23539,N_23439);
nand U23605 (N_23605,N_23401,N_23483);
or U23606 (N_23606,N_23402,N_23450);
nand U23607 (N_23607,N_23419,N_23470);
nand U23608 (N_23608,N_23500,N_23516);
and U23609 (N_23609,N_23437,N_23517);
nor U23610 (N_23610,N_23475,N_23507);
and U23611 (N_23611,N_23413,N_23472);
xnor U23612 (N_23612,N_23540,N_23432);
nand U23613 (N_23613,N_23546,N_23508);
nor U23614 (N_23614,N_23423,N_23447);
and U23615 (N_23615,N_23511,N_23596);
or U23616 (N_23616,N_23462,N_23573);
xor U23617 (N_23617,N_23427,N_23459);
nand U23618 (N_23618,N_23551,N_23561);
nor U23619 (N_23619,N_23407,N_23587);
nand U23620 (N_23620,N_23405,N_23542);
or U23621 (N_23621,N_23461,N_23456);
or U23622 (N_23622,N_23533,N_23486);
nand U23623 (N_23623,N_23481,N_23592);
and U23624 (N_23624,N_23543,N_23482);
nor U23625 (N_23625,N_23526,N_23473);
nand U23626 (N_23626,N_23564,N_23452);
nand U23627 (N_23627,N_23502,N_23535);
nor U23628 (N_23628,N_23442,N_23444);
or U23629 (N_23629,N_23440,N_23411);
xor U23630 (N_23630,N_23460,N_23446);
or U23631 (N_23631,N_23585,N_23420);
and U23632 (N_23632,N_23488,N_23465);
xor U23633 (N_23633,N_23479,N_23586);
nand U23634 (N_23634,N_23572,N_23489);
xnor U23635 (N_23635,N_23513,N_23448);
nor U23636 (N_23636,N_23578,N_23429);
or U23637 (N_23637,N_23471,N_23415);
and U23638 (N_23638,N_23593,N_23518);
or U23639 (N_23639,N_23436,N_23555);
nor U23640 (N_23640,N_23428,N_23597);
nand U23641 (N_23641,N_23476,N_23443);
xnor U23642 (N_23642,N_23544,N_23469);
nor U23643 (N_23643,N_23480,N_23589);
nor U23644 (N_23644,N_23523,N_23410);
nor U23645 (N_23645,N_23501,N_23531);
and U23646 (N_23646,N_23556,N_23527);
nor U23647 (N_23647,N_23591,N_23455);
nor U23648 (N_23648,N_23541,N_23421);
or U23649 (N_23649,N_23406,N_23468);
nand U23650 (N_23650,N_23441,N_23566);
and U23651 (N_23651,N_23494,N_23477);
and U23652 (N_23652,N_23560,N_23525);
and U23653 (N_23653,N_23520,N_23451);
nor U23654 (N_23654,N_23409,N_23514);
nand U23655 (N_23655,N_23598,N_23403);
xor U23656 (N_23656,N_23503,N_23550);
xor U23657 (N_23657,N_23487,N_23464);
and U23658 (N_23658,N_23595,N_23568);
nand U23659 (N_23659,N_23498,N_23445);
nand U23660 (N_23660,N_23493,N_23426);
or U23661 (N_23661,N_23485,N_23492);
or U23662 (N_23662,N_23569,N_23529);
nor U23663 (N_23663,N_23580,N_23496);
nor U23664 (N_23664,N_23534,N_23495);
nor U23665 (N_23665,N_23562,N_23416);
or U23666 (N_23666,N_23537,N_23557);
and U23667 (N_23667,N_23575,N_23599);
xnor U23668 (N_23668,N_23418,N_23491);
xnor U23669 (N_23669,N_23454,N_23425);
xnor U23670 (N_23670,N_23417,N_23530);
and U23671 (N_23671,N_23565,N_23582);
nor U23672 (N_23672,N_23504,N_23548);
nand U23673 (N_23673,N_23553,N_23430);
and U23674 (N_23674,N_23515,N_23490);
nor U23675 (N_23675,N_23571,N_23524);
nor U23676 (N_23676,N_23510,N_23554);
or U23677 (N_23677,N_23588,N_23519);
or U23678 (N_23678,N_23552,N_23458);
nor U23679 (N_23679,N_23577,N_23467);
or U23680 (N_23680,N_23558,N_23422);
nand U23681 (N_23681,N_23435,N_23453);
xor U23682 (N_23682,N_23576,N_23434);
or U23683 (N_23683,N_23412,N_23438);
and U23684 (N_23684,N_23474,N_23466);
nand U23685 (N_23685,N_23424,N_23570);
nor U23686 (N_23686,N_23528,N_23583);
or U23687 (N_23687,N_23400,N_23433);
or U23688 (N_23688,N_23478,N_23538);
and U23689 (N_23689,N_23512,N_23499);
or U23690 (N_23690,N_23521,N_23536);
xnor U23691 (N_23691,N_23567,N_23590);
nand U23692 (N_23692,N_23545,N_23497);
nand U23693 (N_23693,N_23404,N_23574);
or U23694 (N_23694,N_23463,N_23457);
nor U23695 (N_23695,N_23449,N_23506);
and U23696 (N_23696,N_23581,N_23505);
nor U23697 (N_23697,N_23509,N_23584);
nor U23698 (N_23698,N_23408,N_23547);
nand U23699 (N_23699,N_23594,N_23563);
nand U23700 (N_23700,N_23569,N_23455);
nor U23701 (N_23701,N_23466,N_23465);
and U23702 (N_23702,N_23404,N_23535);
nor U23703 (N_23703,N_23484,N_23423);
nor U23704 (N_23704,N_23586,N_23407);
nand U23705 (N_23705,N_23587,N_23538);
nand U23706 (N_23706,N_23408,N_23598);
nor U23707 (N_23707,N_23572,N_23549);
or U23708 (N_23708,N_23482,N_23417);
nand U23709 (N_23709,N_23465,N_23580);
nor U23710 (N_23710,N_23485,N_23458);
nor U23711 (N_23711,N_23416,N_23488);
and U23712 (N_23712,N_23504,N_23418);
and U23713 (N_23713,N_23520,N_23423);
nand U23714 (N_23714,N_23514,N_23459);
nor U23715 (N_23715,N_23569,N_23471);
nand U23716 (N_23716,N_23571,N_23429);
nor U23717 (N_23717,N_23420,N_23453);
and U23718 (N_23718,N_23536,N_23553);
nand U23719 (N_23719,N_23500,N_23546);
nand U23720 (N_23720,N_23463,N_23554);
and U23721 (N_23721,N_23564,N_23474);
and U23722 (N_23722,N_23457,N_23476);
xor U23723 (N_23723,N_23529,N_23583);
and U23724 (N_23724,N_23446,N_23470);
or U23725 (N_23725,N_23424,N_23461);
and U23726 (N_23726,N_23467,N_23576);
or U23727 (N_23727,N_23461,N_23413);
xor U23728 (N_23728,N_23588,N_23443);
nand U23729 (N_23729,N_23590,N_23446);
nand U23730 (N_23730,N_23462,N_23443);
or U23731 (N_23731,N_23474,N_23443);
nand U23732 (N_23732,N_23523,N_23420);
nor U23733 (N_23733,N_23453,N_23510);
or U23734 (N_23734,N_23486,N_23447);
and U23735 (N_23735,N_23563,N_23404);
xor U23736 (N_23736,N_23419,N_23566);
xnor U23737 (N_23737,N_23456,N_23594);
or U23738 (N_23738,N_23576,N_23523);
xnor U23739 (N_23739,N_23589,N_23481);
nor U23740 (N_23740,N_23454,N_23576);
nor U23741 (N_23741,N_23432,N_23442);
and U23742 (N_23742,N_23523,N_23547);
nand U23743 (N_23743,N_23420,N_23520);
nor U23744 (N_23744,N_23494,N_23424);
nand U23745 (N_23745,N_23536,N_23448);
nand U23746 (N_23746,N_23431,N_23520);
and U23747 (N_23747,N_23475,N_23561);
xor U23748 (N_23748,N_23427,N_23565);
xnor U23749 (N_23749,N_23582,N_23405);
nand U23750 (N_23750,N_23464,N_23591);
and U23751 (N_23751,N_23517,N_23459);
xnor U23752 (N_23752,N_23503,N_23568);
nand U23753 (N_23753,N_23454,N_23509);
nand U23754 (N_23754,N_23559,N_23587);
nand U23755 (N_23755,N_23469,N_23507);
or U23756 (N_23756,N_23475,N_23551);
xnor U23757 (N_23757,N_23412,N_23437);
xor U23758 (N_23758,N_23480,N_23424);
xor U23759 (N_23759,N_23519,N_23438);
nand U23760 (N_23760,N_23598,N_23584);
xor U23761 (N_23761,N_23447,N_23402);
or U23762 (N_23762,N_23417,N_23514);
nand U23763 (N_23763,N_23463,N_23464);
nand U23764 (N_23764,N_23570,N_23430);
or U23765 (N_23765,N_23556,N_23432);
xnor U23766 (N_23766,N_23498,N_23403);
nor U23767 (N_23767,N_23429,N_23531);
and U23768 (N_23768,N_23447,N_23445);
nor U23769 (N_23769,N_23509,N_23423);
or U23770 (N_23770,N_23562,N_23502);
and U23771 (N_23771,N_23526,N_23524);
nand U23772 (N_23772,N_23539,N_23401);
nand U23773 (N_23773,N_23592,N_23407);
and U23774 (N_23774,N_23595,N_23460);
nand U23775 (N_23775,N_23568,N_23417);
nand U23776 (N_23776,N_23400,N_23516);
xor U23777 (N_23777,N_23589,N_23568);
nand U23778 (N_23778,N_23475,N_23586);
and U23779 (N_23779,N_23406,N_23554);
and U23780 (N_23780,N_23440,N_23537);
xnor U23781 (N_23781,N_23562,N_23471);
or U23782 (N_23782,N_23543,N_23411);
nand U23783 (N_23783,N_23590,N_23571);
nand U23784 (N_23784,N_23561,N_23443);
and U23785 (N_23785,N_23420,N_23437);
nor U23786 (N_23786,N_23400,N_23427);
xor U23787 (N_23787,N_23417,N_23488);
and U23788 (N_23788,N_23592,N_23408);
and U23789 (N_23789,N_23404,N_23576);
xor U23790 (N_23790,N_23470,N_23589);
and U23791 (N_23791,N_23439,N_23447);
nand U23792 (N_23792,N_23496,N_23503);
nand U23793 (N_23793,N_23401,N_23443);
or U23794 (N_23794,N_23537,N_23589);
nor U23795 (N_23795,N_23484,N_23461);
xor U23796 (N_23796,N_23505,N_23573);
xnor U23797 (N_23797,N_23462,N_23542);
xor U23798 (N_23798,N_23427,N_23515);
xor U23799 (N_23799,N_23544,N_23561);
nand U23800 (N_23800,N_23693,N_23645);
nand U23801 (N_23801,N_23759,N_23756);
xor U23802 (N_23802,N_23714,N_23644);
xor U23803 (N_23803,N_23605,N_23637);
nand U23804 (N_23804,N_23619,N_23667);
and U23805 (N_23805,N_23792,N_23701);
nor U23806 (N_23806,N_23652,N_23633);
or U23807 (N_23807,N_23776,N_23696);
nor U23808 (N_23808,N_23683,N_23799);
nand U23809 (N_23809,N_23695,N_23775);
nand U23810 (N_23810,N_23718,N_23682);
or U23811 (N_23811,N_23630,N_23697);
nor U23812 (N_23812,N_23657,N_23716);
nor U23813 (N_23813,N_23684,N_23741);
and U23814 (N_23814,N_23774,N_23734);
and U23815 (N_23815,N_23761,N_23733);
nor U23816 (N_23816,N_23770,N_23677);
nor U23817 (N_23817,N_23664,N_23738);
nor U23818 (N_23818,N_23732,N_23692);
nand U23819 (N_23819,N_23791,N_23671);
and U23820 (N_23820,N_23726,N_23700);
nand U23821 (N_23821,N_23609,N_23778);
xor U23822 (N_23822,N_23647,N_23681);
xor U23823 (N_23823,N_23705,N_23604);
nor U23824 (N_23824,N_23602,N_23629);
and U23825 (N_23825,N_23612,N_23639);
nand U23826 (N_23826,N_23690,N_23663);
or U23827 (N_23827,N_23781,N_23653);
and U23828 (N_23828,N_23796,N_23650);
xor U23829 (N_23829,N_23707,N_23751);
or U23830 (N_23830,N_23721,N_23728);
nor U23831 (N_23831,N_23782,N_23676);
and U23832 (N_23832,N_23606,N_23669);
and U23833 (N_23833,N_23698,N_23632);
xnor U23834 (N_23834,N_23764,N_23725);
nor U23835 (N_23835,N_23720,N_23771);
nand U23836 (N_23836,N_23739,N_23643);
xnor U23837 (N_23837,N_23731,N_23797);
and U23838 (N_23838,N_23788,N_23742);
and U23839 (N_23839,N_23628,N_23710);
nand U23840 (N_23840,N_23793,N_23687);
or U23841 (N_23841,N_23747,N_23786);
nor U23842 (N_23842,N_23621,N_23755);
nand U23843 (N_23843,N_23625,N_23635);
and U23844 (N_23844,N_23724,N_23757);
nand U23845 (N_23845,N_23668,N_23631);
xor U23846 (N_23846,N_23743,N_23679);
and U23847 (N_23847,N_23624,N_23712);
or U23848 (N_23848,N_23740,N_23749);
xnor U23849 (N_23849,N_23766,N_23616);
nor U23850 (N_23850,N_23750,N_23779);
xnor U23851 (N_23851,N_23758,N_23654);
xnor U23852 (N_23852,N_23620,N_23672);
or U23853 (N_23853,N_23660,N_23662);
or U23854 (N_23854,N_23691,N_23623);
nor U23855 (N_23855,N_23675,N_23610);
or U23856 (N_23856,N_23754,N_23685);
nor U23857 (N_23857,N_23736,N_23706);
xor U23858 (N_23858,N_23789,N_23636);
nor U23859 (N_23859,N_23790,N_23702);
nand U23860 (N_23860,N_23600,N_23648);
and U23861 (N_23861,N_23634,N_23794);
xnor U23862 (N_23862,N_23787,N_23638);
nor U23863 (N_23863,N_23753,N_23780);
nand U23864 (N_23864,N_23666,N_23646);
nand U23865 (N_23865,N_23613,N_23703);
nor U23866 (N_23866,N_23708,N_23608);
xor U23867 (N_23867,N_23615,N_23649);
xor U23868 (N_23868,N_23689,N_23735);
nand U23869 (N_23869,N_23772,N_23680);
nand U23870 (N_23870,N_23711,N_23723);
or U23871 (N_23871,N_23762,N_23763);
nor U23872 (N_23872,N_23611,N_23730);
nor U23873 (N_23873,N_23719,N_23670);
and U23874 (N_23874,N_23785,N_23642);
and U23875 (N_23875,N_23704,N_23744);
and U23876 (N_23876,N_23607,N_23627);
nor U23877 (N_23877,N_23688,N_23614);
and U23878 (N_23878,N_23665,N_23699);
nor U23879 (N_23879,N_23765,N_23717);
or U23880 (N_23880,N_23769,N_23641);
and U23881 (N_23881,N_23694,N_23783);
xor U23882 (N_23882,N_23722,N_23746);
xnor U23883 (N_23883,N_23777,N_23678);
nor U23884 (N_23884,N_23727,N_23674);
and U23885 (N_23885,N_23661,N_23798);
xor U23886 (N_23886,N_23640,N_23773);
nand U23887 (N_23887,N_23686,N_23655);
or U23888 (N_23888,N_23673,N_23745);
nand U23889 (N_23889,N_23748,N_23626);
or U23890 (N_23890,N_23601,N_23656);
nor U23891 (N_23891,N_23752,N_23729);
xnor U23892 (N_23892,N_23618,N_23617);
nand U23893 (N_23893,N_23760,N_23709);
xor U23894 (N_23894,N_23713,N_23767);
xor U23895 (N_23895,N_23603,N_23715);
or U23896 (N_23896,N_23651,N_23737);
and U23897 (N_23897,N_23622,N_23784);
nor U23898 (N_23898,N_23658,N_23768);
nor U23899 (N_23899,N_23795,N_23659);
or U23900 (N_23900,N_23601,N_23668);
and U23901 (N_23901,N_23707,N_23651);
nor U23902 (N_23902,N_23743,N_23654);
or U23903 (N_23903,N_23678,N_23702);
and U23904 (N_23904,N_23611,N_23757);
and U23905 (N_23905,N_23615,N_23735);
or U23906 (N_23906,N_23612,N_23775);
and U23907 (N_23907,N_23699,N_23766);
or U23908 (N_23908,N_23757,N_23713);
nor U23909 (N_23909,N_23741,N_23690);
xor U23910 (N_23910,N_23704,N_23734);
xor U23911 (N_23911,N_23619,N_23757);
nor U23912 (N_23912,N_23633,N_23644);
and U23913 (N_23913,N_23636,N_23650);
nor U23914 (N_23914,N_23750,N_23798);
nand U23915 (N_23915,N_23630,N_23646);
nor U23916 (N_23916,N_23747,N_23692);
nand U23917 (N_23917,N_23737,N_23750);
or U23918 (N_23918,N_23611,N_23617);
xor U23919 (N_23919,N_23781,N_23674);
and U23920 (N_23920,N_23678,N_23641);
or U23921 (N_23921,N_23796,N_23695);
nand U23922 (N_23922,N_23707,N_23671);
nor U23923 (N_23923,N_23725,N_23706);
nand U23924 (N_23924,N_23725,N_23709);
or U23925 (N_23925,N_23759,N_23645);
or U23926 (N_23926,N_23799,N_23749);
and U23927 (N_23927,N_23713,N_23739);
nand U23928 (N_23928,N_23723,N_23661);
nor U23929 (N_23929,N_23760,N_23781);
and U23930 (N_23930,N_23756,N_23795);
xor U23931 (N_23931,N_23757,N_23651);
and U23932 (N_23932,N_23622,N_23697);
and U23933 (N_23933,N_23668,N_23798);
xnor U23934 (N_23934,N_23701,N_23780);
and U23935 (N_23935,N_23639,N_23627);
and U23936 (N_23936,N_23658,N_23709);
or U23937 (N_23937,N_23634,N_23686);
and U23938 (N_23938,N_23658,N_23607);
or U23939 (N_23939,N_23630,N_23722);
nor U23940 (N_23940,N_23743,N_23676);
and U23941 (N_23941,N_23712,N_23670);
nor U23942 (N_23942,N_23790,N_23703);
nor U23943 (N_23943,N_23698,N_23783);
nor U23944 (N_23944,N_23617,N_23791);
or U23945 (N_23945,N_23620,N_23777);
and U23946 (N_23946,N_23686,N_23632);
or U23947 (N_23947,N_23756,N_23708);
nand U23948 (N_23948,N_23685,N_23759);
nor U23949 (N_23949,N_23692,N_23643);
and U23950 (N_23950,N_23705,N_23606);
and U23951 (N_23951,N_23631,N_23764);
or U23952 (N_23952,N_23747,N_23795);
xnor U23953 (N_23953,N_23792,N_23735);
nor U23954 (N_23954,N_23626,N_23773);
nor U23955 (N_23955,N_23682,N_23701);
xnor U23956 (N_23956,N_23672,N_23638);
xor U23957 (N_23957,N_23685,N_23786);
or U23958 (N_23958,N_23752,N_23770);
nor U23959 (N_23959,N_23768,N_23661);
xor U23960 (N_23960,N_23731,N_23759);
and U23961 (N_23961,N_23708,N_23795);
xnor U23962 (N_23962,N_23727,N_23773);
nand U23963 (N_23963,N_23620,N_23692);
nand U23964 (N_23964,N_23655,N_23737);
or U23965 (N_23965,N_23741,N_23735);
and U23966 (N_23966,N_23625,N_23613);
xnor U23967 (N_23967,N_23716,N_23603);
or U23968 (N_23968,N_23654,N_23716);
nand U23969 (N_23969,N_23773,N_23694);
nand U23970 (N_23970,N_23642,N_23621);
and U23971 (N_23971,N_23640,N_23724);
nor U23972 (N_23972,N_23738,N_23730);
nor U23973 (N_23973,N_23678,N_23782);
nor U23974 (N_23974,N_23765,N_23747);
nand U23975 (N_23975,N_23798,N_23629);
or U23976 (N_23976,N_23770,N_23783);
nand U23977 (N_23977,N_23737,N_23707);
xnor U23978 (N_23978,N_23651,N_23614);
nand U23979 (N_23979,N_23737,N_23652);
nor U23980 (N_23980,N_23775,N_23649);
and U23981 (N_23981,N_23775,N_23779);
nand U23982 (N_23982,N_23613,N_23778);
xor U23983 (N_23983,N_23680,N_23760);
nand U23984 (N_23984,N_23672,N_23732);
xnor U23985 (N_23985,N_23646,N_23726);
nor U23986 (N_23986,N_23757,N_23754);
or U23987 (N_23987,N_23617,N_23646);
and U23988 (N_23988,N_23631,N_23698);
and U23989 (N_23989,N_23699,N_23797);
nor U23990 (N_23990,N_23610,N_23783);
xor U23991 (N_23991,N_23663,N_23627);
nor U23992 (N_23992,N_23649,N_23798);
xnor U23993 (N_23993,N_23722,N_23775);
xor U23994 (N_23994,N_23773,N_23608);
nor U23995 (N_23995,N_23654,N_23715);
nand U23996 (N_23996,N_23665,N_23773);
nand U23997 (N_23997,N_23715,N_23698);
xnor U23998 (N_23998,N_23773,N_23742);
nand U23999 (N_23999,N_23766,N_23774);
xor U24000 (N_24000,N_23894,N_23832);
nand U24001 (N_24001,N_23955,N_23882);
or U24002 (N_24002,N_23885,N_23961);
nor U24003 (N_24003,N_23845,N_23982);
and U24004 (N_24004,N_23820,N_23991);
nor U24005 (N_24005,N_23985,N_23976);
xnor U24006 (N_24006,N_23898,N_23887);
or U24007 (N_24007,N_23997,N_23859);
xor U24008 (N_24008,N_23804,N_23877);
nand U24009 (N_24009,N_23974,N_23865);
xor U24010 (N_24010,N_23841,N_23917);
and U24011 (N_24011,N_23920,N_23844);
and U24012 (N_24012,N_23937,N_23881);
xor U24013 (N_24013,N_23999,N_23809);
nand U24014 (N_24014,N_23984,N_23812);
nand U24015 (N_24015,N_23831,N_23970);
or U24016 (N_24016,N_23880,N_23862);
xor U24017 (N_24017,N_23957,N_23945);
and U24018 (N_24018,N_23822,N_23901);
xnor U24019 (N_24019,N_23939,N_23929);
nor U24020 (N_24020,N_23825,N_23936);
and U24021 (N_24021,N_23883,N_23817);
xor U24022 (N_24022,N_23871,N_23872);
and U24023 (N_24023,N_23989,N_23931);
nor U24024 (N_24024,N_23923,N_23904);
xnor U24025 (N_24025,N_23839,N_23916);
nand U24026 (N_24026,N_23824,N_23861);
xnor U24027 (N_24027,N_23846,N_23981);
and U24028 (N_24028,N_23857,N_23966);
or U24029 (N_24029,N_23884,N_23821);
nand U24030 (N_24030,N_23949,N_23912);
or U24031 (N_24031,N_23956,N_23930);
xnor U24032 (N_24032,N_23876,N_23826);
xor U24033 (N_24033,N_23899,N_23962);
and U24034 (N_24034,N_23996,N_23992);
and U24035 (N_24035,N_23867,N_23906);
nand U24036 (N_24036,N_23915,N_23874);
and U24037 (N_24037,N_23828,N_23807);
nor U24038 (N_24038,N_23958,N_23918);
xnor U24039 (N_24039,N_23907,N_23837);
xor U24040 (N_24040,N_23902,N_23995);
nand U24041 (N_24041,N_23944,N_23941);
nand U24042 (N_24042,N_23870,N_23935);
nand U24043 (N_24043,N_23965,N_23842);
nand U24044 (N_24044,N_23924,N_23803);
xor U24045 (N_24045,N_23927,N_23895);
nor U24046 (N_24046,N_23951,N_23878);
nor U24047 (N_24047,N_23819,N_23897);
or U24048 (N_24048,N_23848,N_23813);
and U24049 (N_24049,N_23834,N_23814);
xnor U24050 (N_24050,N_23973,N_23856);
or U24051 (N_24051,N_23980,N_23942);
or U24052 (N_24052,N_23922,N_23811);
and U24053 (N_24053,N_23806,N_23964);
and U24054 (N_24054,N_23875,N_23911);
and U24055 (N_24055,N_23863,N_23928);
or U24056 (N_24056,N_23827,N_23851);
xnor U24057 (N_24057,N_23890,N_23823);
or U24058 (N_24058,N_23879,N_23829);
nand U24059 (N_24059,N_23919,N_23843);
xor U24060 (N_24060,N_23903,N_23840);
and U24061 (N_24061,N_23900,N_23810);
or U24062 (N_24062,N_23971,N_23866);
nor U24063 (N_24063,N_23816,N_23946);
and U24064 (N_24064,N_23943,N_23979);
and U24065 (N_24065,N_23913,N_23987);
and U24066 (N_24066,N_23994,N_23926);
or U24067 (N_24067,N_23977,N_23892);
and U24068 (N_24068,N_23852,N_23934);
and U24069 (N_24069,N_23808,N_23853);
and U24070 (N_24070,N_23800,N_23932);
xor U24071 (N_24071,N_23909,N_23815);
nor U24072 (N_24072,N_23908,N_23886);
or U24073 (N_24073,N_23802,N_23869);
xnor U24074 (N_24074,N_23873,N_23805);
nor U24075 (N_24075,N_23959,N_23954);
and U24076 (N_24076,N_23978,N_23910);
or U24077 (N_24077,N_23975,N_23891);
nor U24078 (N_24078,N_23967,N_23938);
or U24079 (N_24079,N_23864,N_23963);
nand U24080 (N_24080,N_23940,N_23925);
or U24081 (N_24081,N_23921,N_23858);
nor U24082 (N_24082,N_23854,N_23836);
nand U24083 (N_24083,N_23993,N_23801);
xnor U24084 (N_24084,N_23868,N_23893);
nor U24085 (N_24085,N_23969,N_23947);
xnor U24086 (N_24086,N_23860,N_23960);
nor U24087 (N_24087,N_23933,N_23968);
or U24088 (N_24088,N_23914,N_23850);
and U24089 (N_24089,N_23953,N_23986);
nand U24090 (N_24090,N_23998,N_23948);
nor U24091 (N_24091,N_23833,N_23905);
nand U24092 (N_24092,N_23830,N_23888);
and U24093 (N_24093,N_23889,N_23983);
and U24094 (N_24094,N_23847,N_23838);
and U24095 (N_24095,N_23952,N_23818);
and U24096 (N_24096,N_23849,N_23950);
nor U24097 (N_24097,N_23990,N_23988);
and U24098 (N_24098,N_23855,N_23835);
or U24099 (N_24099,N_23896,N_23972);
and U24100 (N_24100,N_23945,N_23846);
nand U24101 (N_24101,N_23815,N_23903);
nor U24102 (N_24102,N_23892,N_23851);
nor U24103 (N_24103,N_23915,N_23826);
or U24104 (N_24104,N_23875,N_23820);
nor U24105 (N_24105,N_23855,N_23873);
nor U24106 (N_24106,N_23981,N_23875);
and U24107 (N_24107,N_23909,N_23830);
and U24108 (N_24108,N_23879,N_23838);
or U24109 (N_24109,N_23843,N_23831);
and U24110 (N_24110,N_23810,N_23827);
and U24111 (N_24111,N_23902,N_23964);
nor U24112 (N_24112,N_23885,N_23908);
nand U24113 (N_24113,N_23947,N_23927);
or U24114 (N_24114,N_23984,N_23946);
and U24115 (N_24115,N_23965,N_23922);
nand U24116 (N_24116,N_23853,N_23955);
and U24117 (N_24117,N_23933,N_23874);
xor U24118 (N_24118,N_23901,N_23965);
xor U24119 (N_24119,N_23944,N_23845);
or U24120 (N_24120,N_23934,N_23859);
nor U24121 (N_24121,N_23809,N_23955);
and U24122 (N_24122,N_23987,N_23915);
and U24123 (N_24123,N_23883,N_23939);
and U24124 (N_24124,N_23930,N_23877);
and U24125 (N_24125,N_23910,N_23951);
nand U24126 (N_24126,N_23992,N_23925);
and U24127 (N_24127,N_23927,N_23808);
or U24128 (N_24128,N_23883,N_23816);
or U24129 (N_24129,N_23917,N_23845);
or U24130 (N_24130,N_23819,N_23814);
and U24131 (N_24131,N_23845,N_23834);
nand U24132 (N_24132,N_23993,N_23940);
and U24133 (N_24133,N_23865,N_23916);
nor U24134 (N_24134,N_23943,N_23870);
and U24135 (N_24135,N_23987,N_23956);
or U24136 (N_24136,N_23997,N_23856);
nor U24137 (N_24137,N_23959,N_23911);
nand U24138 (N_24138,N_23870,N_23881);
and U24139 (N_24139,N_23865,N_23815);
xor U24140 (N_24140,N_23998,N_23843);
xnor U24141 (N_24141,N_23809,N_23935);
xor U24142 (N_24142,N_23876,N_23938);
nand U24143 (N_24143,N_23825,N_23998);
and U24144 (N_24144,N_23987,N_23802);
or U24145 (N_24145,N_23867,N_23896);
nor U24146 (N_24146,N_23850,N_23973);
nor U24147 (N_24147,N_23882,N_23988);
nand U24148 (N_24148,N_23905,N_23958);
nor U24149 (N_24149,N_23855,N_23977);
nand U24150 (N_24150,N_23916,N_23875);
and U24151 (N_24151,N_23916,N_23802);
or U24152 (N_24152,N_23802,N_23853);
nand U24153 (N_24153,N_23913,N_23962);
nor U24154 (N_24154,N_23899,N_23906);
nor U24155 (N_24155,N_23924,N_23936);
xor U24156 (N_24156,N_23951,N_23999);
nand U24157 (N_24157,N_23868,N_23933);
and U24158 (N_24158,N_23986,N_23811);
nand U24159 (N_24159,N_23858,N_23965);
and U24160 (N_24160,N_23998,N_23837);
xnor U24161 (N_24161,N_23955,N_23999);
xor U24162 (N_24162,N_23906,N_23893);
and U24163 (N_24163,N_23930,N_23938);
or U24164 (N_24164,N_23984,N_23942);
xnor U24165 (N_24165,N_23815,N_23986);
and U24166 (N_24166,N_23938,N_23986);
nor U24167 (N_24167,N_23824,N_23943);
or U24168 (N_24168,N_23911,N_23843);
nor U24169 (N_24169,N_23990,N_23874);
or U24170 (N_24170,N_23899,N_23870);
nand U24171 (N_24171,N_23925,N_23820);
nor U24172 (N_24172,N_23918,N_23959);
nand U24173 (N_24173,N_23887,N_23940);
and U24174 (N_24174,N_23880,N_23889);
and U24175 (N_24175,N_23941,N_23853);
nor U24176 (N_24176,N_23857,N_23846);
xor U24177 (N_24177,N_23968,N_23934);
nor U24178 (N_24178,N_23874,N_23896);
and U24179 (N_24179,N_23989,N_23837);
and U24180 (N_24180,N_23812,N_23871);
and U24181 (N_24181,N_23886,N_23990);
xor U24182 (N_24182,N_23921,N_23891);
and U24183 (N_24183,N_23811,N_23951);
nand U24184 (N_24184,N_23917,N_23964);
xnor U24185 (N_24185,N_23919,N_23901);
nand U24186 (N_24186,N_23888,N_23994);
or U24187 (N_24187,N_23911,N_23949);
xor U24188 (N_24188,N_23892,N_23919);
and U24189 (N_24189,N_23953,N_23837);
nand U24190 (N_24190,N_23906,N_23915);
or U24191 (N_24191,N_23969,N_23811);
and U24192 (N_24192,N_23806,N_23867);
or U24193 (N_24193,N_23907,N_23906);
nor U24194 (N_24194,N_23950,N_23834);
nor U24195 (N_24195,N_23816,N_23851);
or U24196 (N_24196,N_23842,N_23820);
nand U24197 (N_24197,N_23816,N_23807);
or U24198 (N_24198,N_23936,N_23899);
or U24199 (N_24199,N_23950,N_23862);
or U24200 (N_24200,N_24148,N_24074);
nand U24201 (N_24201,N_24184,N_24071);
xor U24202 (N_24202,N_24199,N_24058);
nand U24203 (N_24203,N_24124,N_24185);
nand U24204 (N_24204,N_24103,N_24030);
nor U24205 (N_24205,N_24079,N_24091);
xnor U24206 (N_24206,N_24178,N_24152);
and U24207 (N_24207,N_24115,N_24020);
nor U24208 (N_24208,N_24006,N_24097);
xor U24209 (N_24209,N_24029,N_24171);
nor U24210 (N_24210,N_24126,N_24149);
nor U24211 (N_24211,N_24141,N_24121);
and U24212 (N_24212,N_24038,N_24198);
xor U24213 (N_24213,N_24009,N_24052);
and U24214 (N_24214,N_24092,N_24179);
xor U24215 (N_24215,N_24143,N_24080);
nand U24216 (N_24216,N_24047,N_24162);
nand U24217 (N_24217,N_24085,N_24005);
and U24218 (N_24218,N_24193,N_24145);
nand U24219 (N_24219,N_24134,N_24054);
nor U24220 (N_24220,N_24131,N_24151);
and U24221 (N_24221,N_24161,N_24012);
nand U24222 (N_24222,N_24046,N_24122);
and U24223 (N_24223,N_24107,N_24083);
xnor U24224 (N_24224,N_24077,N_24111);
xnor U24225 (N_24225,N_24064,N_24167);
or U24226 (N_24226,N_24105,N_24144);
nor U24227 (N_24227,N_24041,N_24166);
or U24228 (N_24228,N_24036,N_24073);
xnor U24229 (N_24229,N_24173,N_24156);
xor U24230 (N_24230,N_24067,N_24118);
nor U24231 (N_24231,N_24004,N_24048);
and U24232 (N_24232,N_24088,N_24060);
nor U24233 (N_24233,N_24086,N_24158);
and U24234 (N_24234,N_24076,N_24026);
nor U24235 (N_24235,N_24159,N_24096);
and U24236 (N_24236,N_24062,N_24120);
nand U24237 (N_24237,N_24190,N_24057);
nor U24238 (N_24238,N_24010,N_24129);
xnor U24239 (N_24239,N_24195,N_24128);
nor U24240 (N_24240,N_24139,N_24017);
and U24241 (N_24241,N_24133,N_24110);
or U24242 (N_24242,N_24093,N_24053);
nand U24243 (N_24243,N_24163,N_24114);
xor U24244 (N_24244,N_24150,N_24176);
nor U24245 (N_24245,N_24015,N_24069);
or U24246 (N_24246,N_24087,N_24055);
xor U24247 (N_24247,N_24197,N_24075);
xnor U24248 (N_24248,N_24169,N_24008);
and U24249 (N_24249,N_24138,N_24065);
xnor U24250 (N_24250,N_24136,N_24040);
and U24251 (N_24251,N_24089,N_24090);
xor U24252 (N_24252,N_24094,N_24021);
xnor U24253 (N_24253,N_24051,N_24172);
xnor U24254 (N_24254,N_24045,N_24153);
xor U24255 (N_24255,N_24066,N_24186);
or U24256 (N_24256,N_24028,N_24157);
and U24257 (N_24257,N_24192,N_24130);
xnor U24258 (N_24258,N_24098,N_24101);
and U24259 (N_24259,N_24180,N_24019);
or U24260 (N_24260,N_24194,N_24160);
nand U24261 (N_24261,N_24049,N_24137);
xnor U24262 (N_24262,N_24147,N_24146);
nor U24263 (N_24263,N_24104,N_24177);
nor U24264 (N_24264,N_24032,N_24025);
nand U24265 (N_24265,N_24007,N_24174);
nand U24266 (N_24266,N_24196,N_24082);
xnor U24267 (N_24267,N_24001,N_24003);
nand U24268 (N_24268,N_24044,N_24095);
and U24269 (N_24269,N_24135,N_24154);
nand U24270 (N_24270,N_24039,N_24070);
xnor U24271 (N_24271,N_24119,N_24013);
nand U24272 (N_24272,N_24031,N_24022);
nand U24273 (N_24273,N_24181,N_24109);
and U24274 (N_24274,N_24018,N_24187);
xor U24275 (N_24275,N_24059,N_24165);
nor U24276 (N_24276,N_24188,N_24011);
or U24277 (N_24277,N_24127,N_24034);
or U24278 (N_24278,N_24099,N_24170);
nand U24279 (N_24279,N_24072,N_24033);
and U24280 (N_24280,N_24164,N_24182);
xor U24281 (N_24281,N_24132,N_24168);
and U24282 (N_24282,N_24081,N_24042);
nand U24283 (N_24283,N_24043,N_24056);
or U24284 (N_24284,N_24027,N_24189);
or U24285 (N_24285,N_24191,N_24023);
or U24286 (N_24286,N_24050,N_24142);
xnor U24287 (N_24287,N_24016,N_24108);
or U24288 (N_24288,N_24100,N_24102);
nand U24289 (N_24289,N_24037,N_24116);
nor U24290 (N_24290,N_24024,N_24183);
nand U24291 (N_24291,N_24002,N_24113);
or U24292 (N_24292,N_24084,N_24117);
nor U24293 (N_24293,N_24112,N_24035);
nor U24294 (N_24294,N_24068,N_24061);
and U24295 (N_24295,N_24140,N_24078);
xor U24296 (N_24296,N_24175,N_24106);
nand U24297 (N_24297,N_24123,N_24155);
nor U24298 (N_24298,N_24125,N_24000);
nand U24299 (N_24299,N_24014,N_24063);
and U24300 (N_24300,N_24167,N_24191);
or U24301 (N_24301,N_24094,N_24068);
or U24302 (N_24302,N_24163,N_24144);
nand U24303 (N_24303,N_24058,N_24175);
nand U24304 (N_24304,N_24098,N_24154);
nand U24305 (N_24305,N_24170,N_24075);
and U24306 (N_24306,N_24018,N_24095);
nand U24307 (N_24307,N_24106,N_24069);
nand U24308 (N_24308,N_24079,N_24098);
and U24309 (N_24309,N_24136,N_24015);
xor U24310 (N_24310,N_24086,N_24149);
nand U24311 (N_24311,N_24133,N_24121);
and U24312 (N_24312,N_24196,N_24152);
xor U24313 (N_24313,N_24066,N_24073);
or U24314 (N_24314,N_24165,N_24162);
nand U24315 (N_24315,N_24121,N_24006);
or U24316 (N_24316,N_24188,N_24008);
xnor U24317 (N_24317,N_24196,N_24074);
xnor U24318 (N_24318,N_24012,N_24060);
nand U24319 (N_24319,N_24101,N_24096);
nand U24320 (N_24320,N_24036,N_24059);
nor U24321 (N_24321,N_24124,N_24187);
or U24322 (N_24322,N_24168,N_24082);
nor U24323 (N_24323,N_24046,N_24038);
and U24324 (N_24324,N_24116,N_24013);
nand U24325 (N_24325,N_24088,N_24068);
nor U24326 (N_24326,N_24025,N_24179);
nor U24327 (N_24327,N_24118,N_24010);
or U24328 (N_24328,N_24197,N_24157);
or U24329 (N_24329,N_24065,N_24140);
nor U24330 (N_24330,N_24035,N_24069);
xnor U24331 (N_24331,N_24192,N_24121);
and U24332 (N_24332,N_24008,N_24190);
nor U24333 (N_24333,N_24171,N_24024);
nor U24334 (N_24334,N_24127,N_24003);
xnor U24335 (N_24335,N_24094,N_24162);
and U24336 (N_24336,N_24068,N_24076);
xor U24337 (N_24337,N_24026,N_24048);
and U24338 (N_24338,N_24028,N_24022);
nor U24339 (N_24339,N_24184,N_24199);
and U24340 (N_24340,N_24133,N_24032);
and U24341 (N_24341,N_24193,N_24028);
nand U24342 (N_24342,N_24057,N_24169);
nand U24343 (N_24343,N_24188,N_24121);
and U24344 (N_24344,N_24125,N_24004);
nand U24345 (N_24345,N_24050,N_24118);
nor U24346 (N_24346,N_24014,N_24062);
nand U24347 (N_24347,N_24110,N_24042);
nor U24348 (N_24348,N_24098,N_24135);
nor U24349 (N_24349,N_24036,N_24038);
nand U24350 (N_24350,N_24018,N_24087);
nor U24351 (N_24351,N_24080,N_24191);
nor U24352 (N_24352,N_24008,N_24195);
nor U24353 (N_24353,N_24088,N_24188);
or U24354 (N_24354,N_24110,N_24030);
nor U24355 (N_24355,N_24187,N_24010);
and U24356 (N_24356,N_24084,N_24092);
nand U24357 (N_24357,N_24061,N_24041);
xor U24358 (N_24358,N_24056,N_24136);
nor U24359 (N_24359,N_24167,N_24072);
or U24360 (N_24360,N_24078,N_24061);
and U24361 (N_24361,N_24031,N_24179);
or U24362 (N_24362,N_24170,N_24118);
nand U24363 (N_24363,N_24161,N_24159);
nand U24364 (N_24364,N_24071,N_24165);
nor U24365 (N_24365,N_24166,N_24026);
and U24366 (N_24366,N_24038,N_24193);
and U24367 (N_24367,N_24178,N_24119);
nor U24368 (N_24368,N_24028,N_24084);
xnor U24369 (N_24369,N_24042,N_24102);
xor U24370 (N_24370,N_24016,N_24182);
xor U24371 (N_24371,N_24124,N_24056);
or U24372 (N_24372,N_24028,N_24038);
xor U24373 (N_24373,N_24029,N_24095);
or U24374 (N_24374,N_24139,N_24197);
and U24375 (N_24375,N_24164,N_24170);
nor U24376 (N_24376,N_24107,N_24066);
and U24377 (N_24377,N_24012,N_24108);
or U24378 (N_24378,N_24168,N_24034);
and U24379 (N_24379,N_24002,N_24107);
nand U24380 (N_24380,N_24010,N_24197);
or U24381 (N_24381,N_24084,N_24189);
xor U24382 (N_24382,N_24073,N_24158);
and U24383 (N_24383,N_24111,N_24104);
nand U24384 (N_24384,N_24059,N_24169);
xnor U24385 (N_24385,N_24197,N_24022);
nand U24386 (N_24386,N_24122,N_24080);
or U24387 (N_24387,N_24044,N_24174);
nand U24388 (N_24388,N_24021,N_24182);
nand U24389 (N_24389,N_24075,N_24083);
or U24390 (N_24390,N_24089,N_24113);
xor U24391 (N_24391,N_24104,N_24165);
and U24392 (N_24392,N_24050,N_24150);
or U24393 (N_24393,N_24155,N_24076);
or U24394 (N_24394,N_24073,N_24132);
nand U24395 (N_24395,N_24160,N_24095);
nor U24396 (N_24396,N_24105,N_24023);
xnor U24397 (N_24397,N_24174,N_24160);
nand U24398 (N_24398,N_24148,N_24177);
or U24399 (N_24399,N_24177,N_24163);
nor U24400 (N_24400,N_24291,N_24377);
nor U24401 (N_24401,N_24307,N_24369);
and U24402 (N_24402,N_24223,N_24208);
or U24403 (N_24403,N_24359,N_24367);
xor U24404 (N_24404,N_24381,N_24248);
or U24405 (N_24405,N_24247,N_24279);
xnor U24406 (N_24406,N_24396,N_24224);
xnor U24407 (N_24407,N_24316,N_24204);
or U24408 (N_24408,N_24234,N_24380);
xnor U24409 (N_24409,N_24350,N_24249);
nand U24410 (N_24410,N_24206,N_24363);
xor U24411 (N_24411,N_24244,N_24256);
nand U24412 (N_24412,N_24375,N_24276);
nor U24413 (N_24413,N_24322,N_24216);
xor U24414 (N_24414,N_24211,N_24225);
and U24415 (N_24415,N_24356,N_24203);
nand U24416 (N_24416,N_24376,N_24399);
or U24417 (N_24417,N_24320,N_24352);
and U24418 (N_24418,N_24347,N_24295);
and U24419 (N_24419,N_24288,N_24318);
or U24420 (N_24420,N_24338,N_24258);
and U24421 (N_24421,N_24240,N_24342);
xor U24422 (N_24422,N_24314,N_24372);
nor U24423 (N_24423,N_24236,N_24230);
and U24424 (N_24424,N_24280,N_24393);
nand U24425 (N_24425,N_24286,N_24302);
nand U24426 (N_24426,N_24210,N_24214);
and U24427 (N_24427,N_24219,N_24293);
nor U24428 (N_24428,N_24228,N_24389);
nand U24429 (N_24429,N_24289,N_24353);
or U24430 (N_24430,N_24227,N_24262);
xnor U24431 (N_24431,N_24284,N_24315);
xnor U24432 (N_24432,N_24296,N_24213);
nor U24433 (N_24433,N_24305,N_24266);
xor U24434 (N_24434,N_24365,N_24332);
or U24435 (N_24435,N_24283,N_24311);
and U24436 (N_24436,N_24253,N_24222);
nor U24437 (N_24437,N_24226,N_24310);
nor U24438 (N_24438,N_24220,N_24218);
xor U24439 (N_24439,N_24264,N_24301);
nand U24440 (N_24440,N_24290,N_24265);
xor U24441 (N_24441,N_24202,N_24207);
nor U24442 (N_24442,N_24382,N_24200);
nand U24443 (N_24443,N_24340,N_24394);
or U24444 (N_24444,N_24309,N_24341);
nor U24445 (N_24445,N_24368,N_24278);
or U24446 (N_24446,N_24242,N_24261);
and U24447 (N_24447,N_24237,N_24298);
or U24448 (N_24448,N_24395,N_24312);
or U24449 (N_24449,N_24324,N_24308);
nand U24450 (N_24450,N_24345,N_24260);
and U24451 (N_24451,N_24327,N_24362);
nor U24452 (N_24452,N_24360,N_24233);
or U24453 (N_24453,N_24201,N_24205);
or U24454 (N_24454,N_24370,N_24217);
nand U24455 (N_24455,N_24373,N_24209);
and U24456 (N_24456,N_24357,N_24245);
nand U24457 (N_24457,N_24398,N_24255);
or U24458 (N_24458,N_24331,N_24270);
nand U24459 (N_24459,N_24231,N_24325);
nor U24460 (N_24460,N_24383,N_24297);
nor U24461 (N_24461,N_24386,N_24323);
xor U24462 (N_24462,N_24326,N_24273);
or U24463 (N_24463,N_24337,N_24303);
xor U24464 (N_24464,N_24321,N_24238);
or U24465 (N_24465,N_24246,N_24251);
or U24466 (N_24466,N_24285,N_24387);
and U24467 (N_24467,N_24287,N_24319);
or U24468 (N_24468,N_24384,N_24268);
nor U24469 (N_24469,N_24364,N_24335);
xnor U24470 (N_24470,N_24271,N_24277);
nor U24471 (N_24471,N_24348,N_24259);
or U24472 (N_24472,N_24306,N_24392);
and U24473 (N_24473,N_24275,N_24339);
nor U24474 (N_24474,N_24304,N_24294);
xnor U24475 (N_24475,N_24215,N_24232);
xor U24476 (N_24476,N_24274,N_24317);
or U24477 (N_24477,N_24328,N_24333);
nor U24478 (N_24478,N_24391,N_24330);
nand U24479 (N_24479,N_24221,N_24351);
nand U24480 (N_24480,N_24241,N_24346);
and U24481 (N_24481,N_24354,N_24272);
nor U24482 (N_24482,N_24371,N_24374);
or U24483 (N_24483,N_24300,N_24267);
or U24484 (N_24484,N_24358,N_24361);
nand U24485 (N_24485,N_24390,N_24269);
nor U24486 (N_24486,N_24349,N_24379);
and U24487 (N_24487,N_24329,N_24281);
nand U24488 (N_24488,N_24263,N_24334);
or U24489 (N_24489,N_24344,N_24313);
or U24490 (N_24490,N_24252,N_24250);
xnor U24491 (N_24491,N_24229,N_24235);
nor U24492 (N_24492,N_24336,N_24282);
nor U24493 (N_24493,N_24257,N_24299);
nand U24494 (N_24494,N_24243,N_24385);
nor U24495 (N_24495,N_24378,N_24397);
xor U24496 (N_24496,N_24388,N_24355);
nand U24497 (N_24497,N_24343,N_24239);
nor U24498 (N_24498,N_24212,N_24292);
xor U24499 (N_24499,N_24254,N_24366);
nand U24500 (N_24500,N_24200,N_24240);
and U24501 (N_24501,N_24323,N_24353);
or U24502 (N_24502,N_24388,N_24360);
nand U24503 (N_24503,N_24328,N_24342);
nor U24504 (N_24504,N_24378,N_24239);
xor U24505 (N_24505,N_24363,N_24307);
or U24506 (N_24506,N_24259,N_24307);
and U24507 (N_24507,N_24294,N_24379);
and U24508 (N_24508,N_24330,N_24284);
nand U24509 (N_24509,N_24377,N_24280);
nor U24510 (N_24510,N_24348,N_24274);
xnor U24511 (N_24511,N_24226,N_24286);
nor U24512 (N_24512,N_24289,N_24340);
nor U24513 (N_24513,N_24285,N_24239);
and U24514 (N_24514,N_24392,N_24260);
and U24515 (N_24515,N_24372,N_24223);
xnor U24516 (N_24516,N_24359,N_24290);
nor U24517 (N_24517,N_24387,N_24210);
or U24518 (N_24518,N_24367,N_24277);
nor U24519 (N_24519,N_24346,N_24255);
nor U24520 (N_24520,N_24292,N_24237);
xor U24521 (N_24521,N_24207,N_24367);
nor U24522 (N_24522,N_24382,N_24247);
nor U24523 (N_24523,N_24242,N_24202);
nor U24524 (N_24524,N_24276,N_24202);
nor U24525 (N_24525,N_24306,N_24343);
and U24526 (N_24526,N_24220,N_24307);
nor U24527 (N_24527,N_24335,N_24260);
nor U24528 (N_24528,N_24264,N_24220);
nor U24529 (N_24529,N_24272,N_24323);
xnor U24530 (N_24530,N_24372,N_24370);
nand U24531 (N_24531,N_24293,N_24350);
and U24532 (N_24532,N_24308,N_24330);
nand U24533 (N_24533,N_24236,N_24398);
nand U24534 (N_24534,N_24376,N_24323);
nor U24535 (N_24535,N_24205,N_24335);
and U24536 (N_24536,N_24369,N_24231);
or U24537 (N_24537,N_24324,N_24227);
and U24538 (N_24538,N_24272,N_24315);
or U24539 (N_24539,N_24239,N_24383);
and U24540 (N_24540,N_24270,N_24396);
nand U24541 (N_24541,N_24359,N_24376);
and U24542 (N_24542,N_24252,N_24212);
nand U24543 (N_24543,N_24221,N_24288);
nand U24544 (N_24544,N_24217,N_24277);
or U24545 (N_24545,N_24386,N_24362);
nor U24546 (N_24546,N_24297,N_24349);
nand U24547 (N_24547,N_24243,N_24391);
xor U24548 (N_24548,N_24256,N_24229);
xor U24549 (N_24549,N_24338,N_24275);
xnor U24550 (N_24550,N_24255,N_24224);
or U24551 (N_24551,N_24324,N_24240);
nor U24552 (N_24552,N_24359,N_24337);
xor U24553 (N_24553,N_24376,N_24237);
and U24554 (N_24554,N_24262,N_24360);
nand U24555 (N_24555,N_24334,N_24392);
or U24556 (N_24556,N_24202,N_24375);
and U24557 (N_24557,N_24202,N_24362);
or U24558 (N_24558,N_24390,N_24291);
nor U24559 (N_24559,N_24326,N_24348);
nand U24560 (N_24560,N_24220,N_24217);
nand U24561 (N_24561,N_24288,N_24242);
xnor U24562 (N_24562,N_24302,N_24377);
nor U24563 (N_24563,N_24330,N_24286);
nor U24564 (N_24564,N_24267,N_24372);
xnor U24565 (N_24565,N_24351,N_24225);
nand U24566 (N_24566,N_24267,N_24385);
xnor U24567 (N_24567,N_24343,N_24300);
xor U24568 (N_24568,N_24367,N_24221);
xnor U24569 (N_24569,N_24258,N_24250);
and U24570 (N_24570,N_24349,N_24248);
xor U24571 (N_24571,N_24221,N_24233);
and U24572 (N_24572,N_24349,N_24383);
nand U24573 (N_24573,N_24395,N_24360);
or U24574 (N_24574,N_24251,N_24306);
and U24575 (N_24575,N_24360,N_24240);
and U24576 (N_24576,N_24277,N_24254);
xor U24577 (N_24577,N_24393,N_24378);
xnor U24578 (N_24578,N_24234,N_24212);
nand U24579 (N_24579,N_24289,N_24306);
nor U24580 (N_24580,N_24372,N_24384);
nor U24581 (N_24581,N_24308,N_24254);
and U24582 (N_24582,N_24384,N_24203);
or U24583 (N_24583,N_24343,N_24241);
and U24584 (N_24584,N_24229,N_24387);
nor U24585 (N_24585,N_24363,N_24297);
nor U24586 (N_24586,N_24391,N_24228);
and U24587 (N_24587,N_24346,N_24327);
nor U24588 (N_24588,N_24398,N_24335);
or U24589 (N_24589,N_24387,N_24259);
nor U24590 (N_24590,N_24386,N_24200);
nor U24591 (N_24591,N_24274,N_24214);
xor U24592 (N_24592,N_24343,N_24324);
nor U24593 (N_24593,N_24303,N_24275);
nand U24594 (N_24594,N_24385,N_24313);
or U24595 (N_24595,N_24398,N_24362);
xnor U24596 (N_24596,N_24218,N_24379);
xnor U24597 (N_24597,N_24274,N_24258);
or U24598 (N_24598,N_24246,N_24210);
nand U24599 (N_24599,N_24219,N_24317);
and U24600 (N_24600,N_24598,N_24528);
xnor U24601 (N_24601,N_24449,N_24413);
nand U24602 (N_24602,N_24555,N_24507);
xnor U24603 (N_24603,N_24578,N_24589);
and U24604 (N_24604,N_24572,N_24597);
and U24605 (N_24605,N_24490,N_24510);
nand U24606 (N_24606,N_24501,N_24423);
nor U24607 (N_24607,N_24525,N_24472);
or U24608 (N_24608,N_24406,N_24473);
xnor U24609 (N_24609,N_24411,N_24431);
nand U24610 (N_24610,N_24557,N_24479);
and U24611 (N_24611,N_24586,N_24531);
nand U24612 (N_24612,N_24454,N_24434);
and U24613 (N_24613,N_24551,N_24493);
nor U24614 (N_24614,N_24455,N_24486);
nand U24615 (N_24615,N_24542,N_24566);
xnor U24616 (N_24616,N_24569,N_24556);
or U24617 (N_24617,N_24446,N_24595);
xor U24618 (N_24618,N_24456,N_24488);
nor U24619 (N_24619,N_24429,N_24538);
xor U24620 (N_24620,N_24422,N_24487);
and U24621 (N_24621,N_24530,N_24483);
nand U24622 (N_24622,N_24546,N_24513);
xnor U24623 (N_24623,N_24432,N_24596);
nor U24624 (N_24624,N_24509,N_24448);
nor U24625 (N_24625,N_24420,N_24405);
or U24626 (N_24626,N_24447,N_24465);
xnor U24627 (N_24627,N_24553,N_24492);
or U24628 (N_24628,N_24599,N_24476);
or U24629 (N_24629,N_24444,N_24451);
or U24630 (N_24630,N_24505,N_24503);
and U24631 (N_24631,N_24539,N_24498);
nor U24632 (N_24632,N_24435,N_24443);
or U24633 (N_24633,N_24532,N_24552);
and U24634 (N_24634,N_24562,N_24494);
nand U24635 (N_24635,N_24561,N_24577);
and U24636 (N_24636,N_24523,N_24550);
nor U24637 (N_24637,N_24401,N_24594);
or U24638 (N_24638,N_24426,N_24407);
and U24639 (N_24639,N_24558,N_24529);
nand U24640 (N_24640,N_24414,N_24504);
or U24641 (N_24641,N_24592,N_24588);
nor U24642 (N_24642,N_24459,N_24575);
nor U24643 (N_24643,N_24527,N_24425);
nand U24644 (N_24644,N_24461,N_24526);
or U24645 (N_24645,N_24506,N_24502);
nor U24646 (N_24646,N_24587,N_24478);
nor U24647 (N_24647,N_24433,N_24421);
xor U24648 (N_24648,N_24418,N_24417);
nor U24649 (N_24649,N_24593,N_24519);
or U24650 (N_24650,N_24464,N_24474);
and U24651 (N_24651,N_24565,N_24524);
nor U24652 (N_24652,N_24591,N_24583);
or U24653 (N_24653,N_24496,N_24437);
nor U24654 (N_24654,N_24475,N_24497);
and U24655 (N_24655,N_24515,N_24452);
and U24656 (N_24656,N_24585,N_24581);
nand U24657 (N_24657,N_24511,N_24580);
xnor U24658 (N_24658,N_24590,N_24516);
nor U24659 (N_24659,N_24564,N_24537);
or U24660 (N_24660,N_24574,N_24442);
nor U24661 (N_24661,N_24579,N_24549);
nand U24662 (N_24662,N_24554,N_24402);
and U24663 (N_24663,N_24543,N_24441);
and U24664 (N_24664,N_24477,N_24436);
and U24665 (N_24665,N_24427,N_24471);
nand U24666 (N_24666,N_24570,N_24584);
and U24667 (N_24667,N_24484,N_24518);
nand U24668 (N_24668,N_24535,N_24440);
nand U24669 (N_24669,N_24428,N_24544);
nand U24670 (N_24670,N_24495,N_24568);
xnor U24671 (N_24671,N_24457,N_24485);
nor U24672 (N_24672,N_24521,N_24412);
xnor U24673 (N_24673,N_24450,N_24439);
nand U24674 (N_24674,N_24512,N_24548);
and U24675 (N_24675,N_24508,N_24491);
nand U24676 (N_24676,N_24469,N_24467);
nor U24677 (N_24677,N_24480,N_24482);
xor U24678 (N_24678,N_24403,N_24522);
nand U24679 (N_24679,N_24567,N_24463);
nor U24680 (N_24680,N_24453,N_24563);
nor U24681 (N_24681,N_24560,N_24534);
and U24682 (N_24682,N_24460,N_24533);
and U24683 (N_24683,N_24462,N_24416);
xnor U24684 (N_24684,N_24445,N_24545);
or U24685 (N_24685,N_24514,N_24415);
and U24686 (N_24686,N_24400,N_24408);
and U24687 (N_24687,N_24547,N_24536);
xor U24688 (N_24688,N_24540,N_24430);
nor U24689 (N_24689,N_24424,N_24520);
nor U24690 (N_24690,N_24582,N_24409);
and U24691 (N_24691,N_24559,N_24466);
and U24692 (N_24692,N_24458,N_24404);
xor U24693 (N_24693,N_24517,N_24438);
xnor U24694 (N_24694,N_24489,N_24500);
xnor U24695 (N_24695,N_24541,N_24410);
and U24696 (N_24696,N_24468,N_24470);
and U24697 (N_24697,N_24481,N_24419);
nand U24698 (N_24698,N_24571,N_24576);
xor U24699 (N_24699,N_24573,N_24499);
nand U24700 (N_24700,N_24485,N_24439);
or U24701 (N_24701,N_24430,N_24574);
and U24702 (N_24702,N_24516,N_24428);
or U24703 (N_24703,N_24405,N_24486);
nor U24704 (N_24704,N_24524,N_24567);
and U24705 (N_24705,N_24524,N_24549);
nor U24706 (N_24706,N_24417,N_24580);
or U24707 (N_24707,N_24412,N_24515);
xor U24708 (N_24708,N_24475,N_24588);
xor U24709 (N_24709,N_24500,N_24583);
or U24710 (N_24710,N_24444,N_24465);
and U24711 (N_24711,N_24402,N_24507);
nor U24712 (N_24712,N_24458,N_24453);
nand U24713 (N_24713,N_24435,N_24573);
xor U24714 (N_24714,N_24598,N_24538);
nand U24715 (N_24715,N_24515,N_24496);
xor U24716 (N_24716,N_24547,N_24535);
and U24717 (N_24717,N_24551,N_24496);
nand U24718 (N_24718,N_24450,N_24477);
nand U24719 (N_24719,N_24484,N_24559);
and U24720 (N_24720,N_24580,N_24431);
and U24721 (N_24721,N_24426,N_24578);
nand U24722 (N_24722,N_24448,N_24444);
xnor U24723 (N_24723,N_24426,N_24561);
or U24724 (N_24724,N_24587,N_24484);
or U24725 (N_24725,N_24498,N_24514);
nand U24726 (N_24726,N_24568,N_24594);
nor U24727 (N_24727,N_24538,N_24583);
nor U24728 (N_24728,N_24522,N_24441);
and U24729 (N_24729,N_24427,N_24474);
nand U24730 (N_24730,N_24448,N_24402);
nand U24731 (N_24731,N_24432,N_24508);
nor U24732 (N_24732,N_24498,N_24535);
nand U24733 (N_24733,N_24422,N_24545);
nor U24734 (N_24734,N_24529,N_24439);
and U24735 (N_24735,N_24596,N_24479);
and U24736 (N_24736,N_24487,N_24452);
nand U24737 (N_24737,N_24469,N_24479);
nand U24738 (N_24738,N_24429,N_24431);
and U24739 (N_24739,N_24450,N_24559);
nor U24740 (N_24740,N_24432,N_24446);
xor U24741 (N_24741,N_24454,N_24470);
or U24742 (N_24742,N_24430,N_24425);
and U24743 (N_24743,N_24420,N_24438);
and U24744 (N_24744,N_24515,N_24443);
and U24745 (N_24745,N_24538,N_24430);
and U24746 (N_24746,N_24594,N_24428);
nor U24747 (N_24747,N_24422,N_24515);
and U24748 (N_24748,N_24582,N_24450);
nor U24749 (N_24749,N_24510,N_24488);
or U24750 (N_24750,N_24528,N_24433);
xor U24751 (N_24751,N_24536,N_24432);
nand U24752 (N_24752,N_24485,N_24484);
or U24753 (N_24753,N_24454,N_24548);
or U24754 (N_24754,N_24467,N_24576);
or U24755 (N_24755,N_24452,N_24419);
nand U24756 (N_24756,N_24453,N_24528);
or U24757 (N_24757,N_24541,N_24427);
nand U24758 (N_24758,N_24458,N_24468);
nor U24759 (N_24759,N_24592,N_24422);
nor U24760 (N_24760,N_24494,N_24450);
xnor U24761 (N_24761,N_24593,N_24424);
and U24762 (N_24762,N_24449,N_24474);
and U24763 (N_24763,N_24463,N_24401);
xnor U24764 (N_24764,N_24434,N_24567);
and U24765 (N_24765,N_24579,N_24430);
xnor U24766 (N_24766,N_24413,N_24542);
nand U24767 (N_24767,N_24519,N_24413);
nand U24768 (N_24768,N_24412,N_24578);
and U24769 (N_24769,N_24462,N_24466);
xor U24770 (N_24770,N_24590,N_24557);
or U24771 (N_24771,N_24583,N_24401);
nand U24772 (N_24772,N_24484,N_24572);
nor U24773 (N_24773,N_24424,N_24516);
and U24774 (N_24774,N_24428,N_24515);
nand U24775 (N_24775,N_24426,N_24546);
and U24776 (N_24776,N_24437,N_24532);
nand U24777 (N_24777,N_24430,N_24456);
or U24778 (N_24778,N_24411,N_24585);
nand U24779 (N_24779,N_24577,N_24592);
or U24780 (N_24780,N_24467,N_24468);
and U24781 (N_24781,N_24518,N_24555);
nand U24782 (N_24782,N_24423,N_24537);
or U24783 (N_24783,N_24429,N_24525);
xnor U24784 (N_24784,N_24433,N_24516);
xnor U24785 (N_24785,N_24557,N_24439);
or U24786 (N_24786,N_24456,N_24494);
xnor U24787 (N_24787,N_24515,N_24573);
xnor U24788 (N_24788,N_24514,N_24502);
and U24789 (N_24789,N_24467,N_24598);
xnor U24790 (N_24790,N_24410,N_24512);
nor U24791 (N_24791,N_24459,N_24439);
and U24792 (N_24792,N_24554,N_24448);
nor U24793 (N_24793,N_24472,N_24559);
and U24794 (N_24794,N_24484,N_24447);
nand U24795 (N_24795,N_24425,N_24512);
xor U24796 (N_24796,N_24477,N_24581);
and U24797 (N_24797,N_24448,N_24508);
nor U24798 (N_24798,N_24599,N_24421);
nor U24799 (N_24799,N_24590,N_24456);
or U24800 (N_24800,N_24675,N_24736);
nand U24801 (N_24801,N_24609,N_24717);
or U24802 (N_24802,N_24629,N_24769);
and U24803 (N_24803,N_24708,N_24718);
nor U24804 (N_24804,N_24678,N_24702);
nor U24805 (N_24805,N_24694,N_24787);
xor U24806 (N_24806,N_24658,N_24665);
nor U24807 (N_24807,N_24645,N_24650);
and U24808 (N_24808,N_24639,N_24620);
nand U24809 (N_24809,N_24605,N_24780);
nor U24810 (N_24810,N_24727,N_24669);
nor U24811 (N_24811,N_24604,N_24758);
nand U24812 (N_24812,N_24667,N_24796);
or U24813 (N_24813,N_24619,N_24764);
nand U24814 (N_24814,N_24630,N_24622);
nor U24815 (N_24815,N_24699,N_24679);
nor U24816 (N_24816,N_24797,N_24676);
nand U24817 (N_24817,N_24696,N_24773);
nand U24818 (N_24818,N_24747,N_24656);
nor U24819 (N_24819,N_24646,N_24766);
nor U24820 (N_24820,N_24648,N_24789);
or U24821 (N_24821,N_24625,N_24680);
or U24822 (N_24822,N_24759,N_24637);
nand U24823 (N_24823,N_24684,N_24690);
or U24824 (N_24824,N_24705,N_24738);
xnor U24825 (N_24825,N_24730,N_24716);
or U24826 (N_24826,N_24767,N_24654);
xnor U24827 (N_24827,N_24771,N_24725);
nand U24828 (N_24828,N_24757,N_24613);
and U24829 (N_24829,N_24781,N_24723);
or U24830 (N_24830,N_24616,N_24634);
or U24831 (N_24831,N_24704,N_24693);
nand U24832 (N_24832,N_24642,N_24799);
or U24833 (N_24833,N_24691,N_24701);
or U24834 (N_24834,N_24663,N_24776);
xor U24835 (N_24835,N_24710,N_24615);
or U24836 (N_24836,N_24724,N_24672);
or U24837 (N_24837,N_24611,N_24624);
xnor U24838 (N_24838,N_24778,N_24685);
or U24839 (N_24839,N_24794,N_24768);
nor U24840 (N_24840,N_24700,N_24608);
and U24841 (N_24841,N_24635,N_24782);
or U24842 (N_24842,N_24602,N_24770);
nor U24843 (N_24843,N_24741,N_24745);
nor U24844 (N_24844,N_24633,N_24688);
or U24845 (N_24845,N_24617,N_24784);
nand U24846 (N_24846,N_24640,N_24728);
or U24847 (N_24847,N_24600,N_24734);
and U24848 (N_24848,N_24673,N_24753);
xor U24849 (N_24849,N_24659,N_24737);
and U24850 (N_24850,N_24621,N_24732);
nor U24851 (N_24851,N_24618,N_24632);
and U24852 (N_24852,N_24682,N_24695);
nor U24853 (N_24853,N_24603,N_24711);
nand U24854 (N_24854,N_24733,N_24662);
nor U24855 (N_24855,N_24743,N_24779);
and U24856 (N_24856,N_24643,N_24692);
xor U24857 (N_24857,N_24783,N_24670);
nand U24858 (N_24858,N_24721,N_24775);
or U24859 (N_24859,N_24763,N_24698);
or U24860 (N_24860,N_24607,N_24677);
xor U24861 (N_24861,N_24792,N_24707);
xor U24862 (N_24862,N_24772,N_24644);
or U24863 (N_24863,N_24715,N_24668);
or U24864 (N_24864,N_24689,N_24748);
nand U24865 (N_24865,N_24740,N_24749);
nor U24866 (N_24866,N_24601,N_24636);
or U24867 (N_24867,N_24638,N_24674);
nor U24868 (N_24868,N_24720,N_24614);
and U24869 (N_24869,N_24765,N_24709);
nor U24870 (N_24870,N_24786,N_24641);
or U24871 (N_24871,N_24752,N_24790);
or U24872 (N_24872,N_24610,N_24687);
xor U24873 (N_24873,N_24798,N_24746);
or U24874 (N_24874,N_24647,N_24661);
nand U24875 (N_24875,N_24750,N_24731);
nor U24876 (N_24876,N_24651,N_24754);
or U24877 (N_24877,N_24657,N_24649);
or U24878 (N_24878,N_24664,N_24774);
or U24879 (N_24879,N_24795,N_24714);
nand U24880 (N_24880,N_24660,N_24742);
nand U24881 (N_24881,N_24606,N_24623);
nand U24882 (N_24882,N_24777,N_24626);
nand U24883 (N_24883,N_24719,N_24785);
or U24884 (N_24884,N_24653,N_24655);
or U24885 (N_24885,N_24760,N_24722);
xor U24886 (N_24886,N_24666,N_24726);
nand U24887 (N_24887,N_24683,N_24703);
and U24888 (N_24888,N_24735,N_24612);
nand U24889 (N_24889,N_24713,N_24652);
nand U24890 (N_24890,N_24791,N_24739);
nor U24891 (N_24891,N_24681,N_24706);
xnor U24892 (N_24892,N_24788,N_24628);
xnor U24893 (N_24893,N_24697,N_24762);
xor U24894 (N_24894,N_24756,N_24751);
xor U24895 (N_24895,N_24627,N_24631);
nor U24896 (N_24896,N_24671,N_24712);
xor U24897 (N_24897,N_24755,N_24744);
xor U24898 (N_24898,N_24793,N_24761);
nor U24899 (N_24899,N_24686,N_24729);
nor U24900 (N_24900,N_24792,N_24604);
and U24901 (N_24901,N_24716,N_24775);
and U24902 (N_24902,N_24738,N_24639);
xnor U24903 (N_24903,N_24756,N_24720);
or U24904 (N_24904,N_24616,N_24758);
nor U24905 (N_24905,N_24632,N_24757);
xnor U24906 (N_24906,N_24752,N_24725);
nor U24907 (N_24907,N_24619,N_24789);
xnor U24908 (N_24908,N_24706,N_24677);
xnor U24909 (N_24909,N_24746,N_24767);
xor U24910 (N_24910,N_24788,N_24779);
nor U24911 (N_24911,N_24610,N_24627);
and U24912 (N_24912,N_24674,N_24736);
and U24913 (N_24913,N_24739,N_24790);
and U24914 (N_24914,N_24686,N_24714);
or U24915 (N_24915,N_24715,N_24793);
and U24916 (N_24916,N_24636,N_24688);
nor U24917 (N_24917,N_24692,N_24623);
nor U24918 (N_24918,N_24764,N_24669);
or U24919 (N_24919,N_24623,N_24726);
xnor U24920 (N_24920,N_24614,N_24702);
nor U24921 (N_24921,N_24611,N_24750);
xnor U24922 (N_24922,N_24729,N_24652);
nor U24923 (N_24923,N_24615,N_24779);
nand U24924 (N_24924,N_24710,N_24676);
and U24925 (N_24925,N_24732,N_24719);
or U24926 (N_24926,N_24630,N_24716);
xnor U24927 (N_24927,N_24677,N_24698);
xor U24928 (N_24928,N_24676,N_24758);
or U24929 (N_24929,N_24686,N_24609);
and U24930 (N_24930,N_24606,N_24603);
xor U24931 (N_24931,N_24750,N_24697);
or U24932 (N_24932,N_24734,N_24691);
nor U24933 (N_24933,N_24634,N_24670);
or U24934 (N_24934,N_24606,N_24638);
xnor U24935 (N_24935,N_24659,N_24662);
xor U24936 (N_24936,N_24632,N_24660);
nand U24937 (N_24937,N_24684,N_24780);
or U24938 (N_24938,N_24718,N_24788);
or U24939 (N_24939,N_24675,N_24696);
and U24940 (N_24940,N_24713,N_24773);
nor U24941 (N_24941,N_24784,N_24730);
xnor U24942 (N_24942,N_24629,N_24654);
nand U24943 (N_24943,N_24760,N_24715);
nor U24944 (N_24944,N_24645,N_24632);
nor U24945 (N_24945,N_24712,N_24718);
and U24946 (N_24946,N_24678,N_24733);
and U24947 (N_24947,N_24629,N_24718);
and U24948 (N_24948,N_24760,N_24748);
and U24949 (N_24949,N_24722,N_24768);
and U24950 (N_24950,N_24761,N_24723);
and U24951 (N_24951,N_24770,N_24695);
nor U24952 (N_24952,N_24773,N_24692);
nand U24953 (N_24953,N_24663,N_24738);
or U24954 (N_24954,N_24618,N_24728);
and U24955 (N_24955,N_24659,N_24635);
nand U24956 (N_24956,N_24733,N_24716);
or U24957 (N_24957,N_24629,N_24724);
or U24958 (N_24958,N_24799,N_24646);
nand U24959 (N_24959,N_24736,N_24603);
nor U24960 (N_24960,N_24689,N_24745);
and U24961 (N_24961,N_24690,N_24605);
or U24962 (N_24962,N_24698,N_24783);
and U24963 (N_24963,N_24699,N_24737);
xor U24964 (N_24964,N_24710,N_24632);
nor U24965 (N_24965,N_24627,N_24783);
or U24966 (N_24966,N_24768,N_24744);
nor U24967 (N_24967,N_24784,N_24644);
and U24968 (N_24968,N_24773,N_24660);
nor U24969 (N_24969,N_24768,N_24793);
nor U24970 (N_24970,N_24616,N_24630);
or U24971 (N_24971,N_24631,N_24724);
xnor U24972 (N_24972,N_24769,N_24603);
nand U24973 (N_24973,N_24758,N_24679);
nor U24974 (N_24974,N_24770,N_24788);
nand U24975 (N_24975,N_24756,N_24635);
or U24976 (N_24976,N_24611,N_24672);
and U24977 (N_24977,N_24627,N_24747);
xnor U24978 (N_24978,N_24712,N_24675);
nand U24979 (N_24979,N_24651,N_24722);
nand U24980 (N_24980,N_24714,N_24767);
or U24981 (N_24981,N_24684,N_24696);
nand U24982 (N_24982,N_24758,N_24738);
or U24983 (N_24983,N_24627,N_24640);
or U24984 (N_24984,N_24677,N_24763);
xnor U24985 (N_24985,N_24633,N_24610);
nor U24986 (N_24986,N_24748,N_24717);
and U24987 (N_24987,N_24767,N_24743);
nand U24988 (N_24988,N_24775,N_24647);
nand U24989 (N_24989,N_24614,N_24664);
and U24990 (N_24990,N_24632,N_24779);
xnor U24991 (N_24991,N_24610,N_24609);
or U24992 (N_24992,N_24746,N_24653);
xnor U24993 (N_24993,N_24617,N_24753);
nand U24994 (N_24994,N_24778,N_24712);
nand U24995 (N_24995,N_24600,N_24775);
or U24996 (N_24996,N_24601,N_24706);
and U24997 (N_24997,N_24641,N_24770);
nor U24998 (N_24998,N_24666,N_24636);
and U24999 (N_24999,N_24756,N_24729);
xnor U25000 (N_25000,N_24946,N_24894);
nand U25001 (N_25001,N_24989,N_24925);
nor U25002 (N_25002,N_24817,N_24971);
or U25003 (N_25003,N_24911,N_24831);
nand U25004 (N_25004,N_24883,N_24953);
nand U25005 (N_25005,N_24900,N_24996);
or U25006 (N_25006,N_24871,N_24943);
or U25007 (N_25007,N_24874,N_24927);
nor U25008 (N_25008,N_24881,N_24800);
and U25009 (N_25009,N_24884,N_24885);
and U25010 (N_25010,N_24980,N_24917);
nor U25011 (N_25011,N_24896,N_24855);
xnor U25012 (N_25012,N_24934,N_24970);
nor U25013 (N_25013,N_24830,N_24928);
or U25014 (N_25014,N_24979,N_24918);
nand U25015 (N_25015,N_24833,N_24838);
xor U25016 (N_25016,N_24988,N_24818);
nand U25017 (N_25017,N_24923,N_24902);
nand U25018 (N_25018,N_24866,N_24876);
nor U25019 (N_25019,N_24933,N_24991);
nand U25020 (N_25020,N_24812,N_24997);
nor U25021 (N_25021,N_24870,N_24820);
nand U25022 (N_25022,N_24841,N_24805);
and U25023 (N_25023,N_24926,N_24921);
or U25024 (N_25024,N_24986,N_24810);
nor U25025 (N_25025,N_24813,N_24910);
nor U25026 (N_25026,N_24890,N_24882);
nand U25027 (N_25027,N_24898,N_24873);
xor U25028 (N_25028,N_24942,N_24967);
and U25029 (N_25029,N_24968,N_24856);
and U25030 (N_25030,N_24836,N_24857);
nor U25031 (N_25031,N_24877,N_24944);
and U25032 (N_25032,N_24957,N_24931);
nor U25033 (N_25033,N_24869,N_24982);
nor U25034 (N_25034,N_24956,N_24981);
nor U25035 (N_25035,N_24972,N_24941);
and U25036 (N_25036,N_24913,N_24978);
nand U25037 (N_25037,N_24845,N_24951);
nor U25038 (N_25038,N_24935,N_24827);
and U25039 (N_25039,N_24975,N_24875);
xnor U25040 (N_25040,N_24895,N_24985);
and U25041 (N_25041,N_24950,N_24815);
and U25042 (N_25042,N_24952,N_24889);
or U25043 (N_25043,N_24961,N_24822);
or U25044 (N_25044,N_24995,N_24906);
or U25045 (N_25045,N_24987,N_24872);
nand U25046 (N_25046,N_24990,N_24924);
xnor U25047 (N_25047,N_24919,N_24983);
and U25048 (N_25048,N_24843,N_24880);
nor U25049 (N_25049,N_24994,N_24998);
nor U25050 (N_25050,N_24832,N_24948);
xnor U25051 (N_25051,N_24835,N_24993);
nor U25052 (N_25052,N_24965,N_24816);
and U25053 (N_25053,N_24819,N_24806);
nand U25054 (N_25054,N_24809,N_24891);
and U25055 (N_25055,N_24825,N_24839);
nand U25056 (N_25056,N_24879,N_24920);
xnor U25057 (N_25057,N_24939,N_24984);
and U25058 (N_25058,N_24959,N_24958);
or U25059 (N_25059,N_24863,N_24848);
xnor U25060 (N_25060,N_24824,N_24846);
nand U25061 (N_25061,N_24887,N_24940);
and U25062 (N_25062,N_24909,N_24808);
and U25063 (N_25063,N_24938,N_24802);
or U25064 (N_25064,N_24821,N_24904);
xor U25065 (N_25065,N_24823,N_24865);
nor U25066 (N_25066,N_24828,N_24851);
xor U25067 (N_25067,N_24897,N_24974);
nor U25068 (N_25068,N_24912,N_24893);
xnor U25069 (N_25069,N_24852,N_24849);
and U25070 (N_25070,N_24969,N_24905);
nor U25071 (N_25071,N_24878,N_24963);
xor U25072 (N_25072,N_24907,N_24850);
or U25073 (N_25073,N_24842,N_24937);
nand U25074 (N_25074,N_24960,N_24964);
nor U25075 (N_25075,N_24914,N_24886);
nor U25076 (N_25076,N_24826,N_24908);
xnor U25077 (N_25077,N_24949,N_24837);
nor U25078 (N_25078,N_24804,N_24977);
nand U25079 (N_25079,N_24901,N_24962);
nor U25080 (N_25080,N_24888,N_24864);
and U25081 (N_25081,N_24999,N_24814);
and U25082 (N_25082,N_24922,N_24860);
nand U25083 (N_25083,N_24945,N_24966);
nor U25084 (N_25084,N_24955,N_24862);
nand U25085 (N_25085,N_24930,N_24947);
nand U25086 (N_25086,N_24801,N_24834);
and U25087 (N_25087,N_24932,N_24903);
and U25088 (N_25088,N_24992,N_24973);
nor U25089 (N_25089,N_24829,N_24854);
and U25090 (N_25090,N_24892,N_24811);
nor U25091 (N_25091,N_24853,N_24844);
nor U25092 (N_25092,N_24803,N_24954);
and U25093 (N_25093,N_24899,N_24840);
and U25094 (N_25094,N_24807,N_24915);
and U25095 (N_25095,N_24929,N_24861);
nor U25096 (N_25096,N_24976,N_24867);
nor U25097 (N_25097,N_24868,N_24847);
or U25098 (N_25098,N_24916,N_24858);
xnor U25099 (N_25099,N_24936,N_24859);
and U25100 (N_25100,N_24831,N_24958);
nand U25101 (N_25101,N_24936,N_24813);
or U25102 (N_25102,N_24910,N_24996);
nand U25103 (N_25103,N_24871,N_24917);
nand U25104 (N_25104,N_24972,N_24814);
and U25105 (N_25105,N_24932,N_24819);
nand U25106 (N_25106,N_24927,N_24969);
nand U25107 (N_25107,N_24957,N_24919);
nand U25108 (N_25108,N_24925,N_24931);
xor U25109 (N_25109,N_24899,N_24927);
or U25110 (N_25110,N_24806,N_24980);
and U25111 (N_25111,N_24947,N_24995);
or U25112 (N_25112,N_24839,N_24860);
xnor U25113 (N_25113,N_24883,N_24941);
or U25114 (N_25114,N_24963,N_24846);
or U25115 (N_25115,N_24853,N_24842);
nor U25116 (N_25116,N_24991,N_24997);
xor U25117 (N_25117,N_24902,N_24967);
nor U25118 (N_25118,N_24920,N_24896);
and U25119 (N_25119,N_24980,N_24849);
or U25120 (N_25120,N_24939,N_24952);
and U25121 (N_25121,N_24967,N_24809);
and U25122 (N_25122,N_24998,N_24806);
nor U25123 (N_25123,N_24803,N_24934);
and U25124 (N_25124,N_24904,N_24887);
nor U25125 (N_25125,N_24882,N_24848);
nor U25126 (N_25126,N_24928,N_24988);
nor U25127 (N_25127,N_24971,N_24901);
or U25128 (N_25128,N_24845,N_24892);
nand U25129 (N_25129,N_24846,N_24813);
and U25130 (N_25130,N_24862,N_24839);
nor U25131 (N_25131,N_24968,N_24889);
nand U25132 (N_25132,N_24942,N_24892);
nand U25133 (N_25133,N_24895,N_24807);
xor U25134 (N_25134,N_24972,N_24931);
and U25135 (N_25135,N_24974,N_24819);
and U25136 (N_25136,N_24890,N_24913);
or U25137 (N_25137,N_24851,N_24939);
xnor U25138 (N_25138,N_24803,N_24917);
xor U25139 (N_25139,N_24823,N_24885);
or U25140 (N_25140,N_24856,N_24925);
nand U25141 (N_25141,N_24981,N_24947);
xnor U25142 (N_25142,N_24877,N_24860);
nand U25143 (N_25143,N_24825,N_24904);
nand U25144 (N_25144,N_24879,N_24880);
nor U25145 (N_25145,N_24949,N_24955);
or U25146 (N_25146,N_24928,N_24804);
nor U25147 (N_25147,N_24967,N_24930);
xnor U25148 (N_25148,N_24923,N_24825);
xnor U25149 (N_25149,N_24945,N_24815);
or U25150 (N_25150,N_24856,N_24880);
nand U25151 (N_25151,N_24952,N_24995);
or U25152 (N_25152,N_24866,N_24919);
or U25153 (N_25153,N_24873,N_24978);
or U25154 (N_25154,N_24851,N_24920);
xnor U25155 (N_25155,N_24967,N_24859);
nor U25156 (N_25156,N_24903,N_24815);
xor U25157 (N_25157,N_24844,N_24984);
xnor U25158 (N_25158,N_24963,N_24805);
or U25159 (N_25159,N_24876,N_24893);
or U25160 (N_25160,N_24818,N_24926);
nor U25161 (N_25161,N_24915,N_24917);
and U25162 (N_25162,N_24886,N_24906);
and U25163 (N_25163,N_24808,N_24898);
nor U25164 (N_25164,N_24993,N_24981);
nor U25165 (N_25165,N_24941,N_24907);
xnor U25166 (N_25166,N_24939,N_24909);
or U25167 (N_25167,N_24924,N_24916);
or U25168 (N_25168,N_24808,N_24855);
nand U25169 (N_25169,N_24816,N_24927);
and U25170 (N_25170,N_24847,N_24938);
or U25171 (N_25171,N_24946,N_24943);
and U25172 (N_25172,N_24892,N_24999);
or U25173 (N_25173,N_24846,N_24949);
nor U25174 (N_25174,N_24981,N_24852);
nand U25175 (N_25175,N_24915,N_24850);
or U25176 (N_25176,N_24817,N_24925);
or U25177 (N_25177,N_24970,N_24946);
nor U25178 (N_25178,N_24953,N_24918);
nor U25179 (N_25179,N_24953,N_24969);
xor U25180 (N_25180,N_24800,N_24966);
or U25181 (N_25181,N_24814,N_24843);
nor U25182 (N_25182,N_24832,N_24856);
nand U25183 (N_25183,N_24908,N_24867);
or U25184 (N_25184,N_24827,N_24938);
and U25185 (N_25185,N_24854,N_24973);
or U25186 (N_25186,N_24979,N_24892);
nor U25187 (N_25187,N_24928,N_24862);
nand U25188 (N_25188,N_24919,N_24990);
or U25189 (N_25189,N_24881,N_24969);
nor U25190 (N_25190,N_24924,N_24873);
and U25191 (N_25191,N_24830,N_24847);
nor U25192 (N_25192,N_24963,N_24981);
or U25193 (N_25193,N_24856,N_24956);
nor U25194 (N_25194,N_24883,N_24903);
and U25195 (N_25195,N_24990,N_24922);
and U25196 (N_25196,N_24946,N_24876);
or U25197 (N_25197,N_24926,N_24827);
xor U25198 (N_25198,N_24840,N_24837);
or U25199 (N_25199,N_24863,N_24926);
or U25200 (N_25200,N_25028,N_25116);
xnor U25201 (N_25201,N_25166,N_25114);
nor U25202 (N_25202,N_25005,N_25135);
nand U25203 (N_25203,N_25027,N_25107);
nor U25204 (N_25204,N_25189,N_25025);
nor U25205 (N_25205,N_25173,N_25004);
nand U25206 (N_25206,N_25105,N_25043);
or U25207 (N_25207,N_25153,N_25077);
nand U25208 (N_25208,N_25119,N_25131);
and U25209 (N_25209,N_25164,N_25041);
or U25210 (N_25210,N_25083,N_25089);
or U25211 (N_25211,N_25023,N_25086);
and U25212 (N_25212,N_25084,N_25011);
or U25213 (N_25213,N_25049,N_25038);
or U25214 (N_25214,N_25087,N_25186);
and U25215 (N_25215,N_25016,N_25177);
and U25216 (N_25216,N_25017,N_25163);
nor U25217 (N_25217,N_25103,N_25062);
nand U25218 (N_25218,N_25156,N_25008);
nand U25219 (N_25219,N_25094,N_25014);
or U25220 (N_25220,N_25146,N_25054);
nand U25221 (N_25221,N_25154,N_25066);
nand U25222 (N_25222,N_25139,N_25098);
nand U25223 (N_25223,N_25081,N_25079);
and U25224 (N_25224,N_25015,N_25198);
nand U25225 (N_25225,N_25071,N_25165);
nand U25226 (N_25226,N_25144,N_25104);
and U25227 (N_25227,N_25151,N_25029);
nor U25228 (N_25228,N_25194,N_25145);
nor U25229 (N_25229,N_25031,N_25161);
nand U25230 (N_25230,N_25040,N_25174);
xor U25231 (N_25231,N_25178,N_25123);
nand U25232 (N_25232,N_25115,N_25090);
nand U25233 (N_25233,N_25170,N_25032);
or U25234 (N_25234,N_25117,N_25065);
and U25235 (N_25235,N_25188,N_25129);
xnor U25236 (N_25236,N_25196,N_25061);
nor U25237 (N_25237,N_25092,N_25120);
nor U25238 (N_25238,N_25073,N_25034);
or U25239 (N_25239,N_25074,N_25099);
nand U25240 (N_25240,N_25171,N_25030);
xnor U25241 (N_25241,N_25045,N_25007);
nor U25242 (N_25242,N_25091,N_25180);
nor U25243 (N_25243,N_25053,N_25158);
xnor U25244 (N_25244,N_25112,N_25001);
and U25245 (N_25245,N_25111,N_25149);
nand U25246 (N_25246,N_25072,N_25050);
xnor U25247 (N_25247,N_25124,N_25132);
and U25248 (N_25248,N_25024,N_25035);
xnor U25249 (N_25249,N_25052,N_25127);
nand U25250 (N_25250,N_25100,N_25182);
xnor U25251 (N_25251,N_25059,N_25152);
nand U25252 (N_25252,N_25068,N_25181);
nor U25253 (N_25253,N_25097,N_25192);
and U25254 (N_25254,N_25106,N_25133);
xor U25255 (N_25255,N_25010,N_25058);
nor U25256 (N_25256,N_25147,N_25009);
or U25257 (N_25257,N_25195,N_25018);
nand U25258 (N_25258,N_25126,N_25080);
and U25259 (N_25259,N_25051,N_25167);
or U25260 (N_25260,N_25187,N_25102);
xnor U25261 (N_25261,N_25155,N_25037);
or U25262 (N_25262,N_25006,N_25057);
or U25263 (N_25263,N_25002,N_25042);
or U25264 (N_25264,N_25064,N_25157);
xor U25265 (N_25265,N_25141,N_25121);
xnor U25266 (N_25266,N_25110,N_25136);
xnor U25267 (N_25267,N_25047,N_25193);
xor U25268 (N_25268,N_25137,N_25172);
and U25269 (N_25269,N_25113,N_25095);
nand U25270 (N_25270,N_25055,N_25046);
and U25271 (N_25271,N_25039,N_25075);
nor U25272 (N_25272,N_25159,N_25130);
xnor U25273 (N_25273,N_25160,N_25108);
and U25274 (N_25274,N_25020,N_25021);
xor U25275 (N_25275,N_25022,N_25128);
and U25276 (N_25276,N_25134,N_25122);
and U25277 (N_25277,N_25168,N_25013);
xnor U25278 (N_25278,N_25176,N_25197);
nor U25279 (N_25279,N_25076,N_25012);
xor U25280 (N_25280,N_25169,N_25143);
xnor U25281 (N_25281,N_25150,N_25142);
xnor U25282 (N_25282,N_25000,N_25162);
or U25283 (N_25283,N_25190,N_25138);
or U25284 (N_25284,N_25118,N_25175);
xor U25285 (N_25285,N_25096,N_25044);
xnor U25286 (N_25286,N_25060,N_25140);
nand U25287 (N_25287,N_25093,N_25125);
and U25288 (N_25288,N_25101,N_25191);
xnor U25289 (N_25289,N_25185,N_25088);
or U25290 (N_25290,N_25070,N_25063);
nor U25291 (N_25291,N_25003,N_25067);
and U25292 (N_25292,N_25033,N_25199);
nand U25293 (N_25293,N_25082,N_25056);
nand U25294 (N_25294,N_25026,N_25179);
xor U25295 (N_25295,N_25069,N_25036);
nand U25296 (N_25296,N_25078,N_25183);
xor U25297 (N_25297,N_25148,N_25085);
or U25298 (N_25298,N_25048,N_25184);
xnor U25299 (N_25299,N_25019,N_25109);
nor U25300 (N_25300,N_25045,N_25062);
nand U25301 (N_25301,N_25135,N_25114);
or U25302 (N_25302,N_25059,N_25197);
nor U25303 (N_25303,N_25158,N_25130);
xnor U25304 (N_25304,N_25096,N_25047);
xnor U25305 (N_25305,N_25142,N_25155);
and U25306 (N_25306,N_25092,N_25006);
and U25307 (N_25307,N_25096,N_25035);
xor U25308 (N_25308,N_25056,N_25025);
nand U25309 (N_25309,N_25075,N_25073);
or U25310 (N_25310,N_25032,N_25141);
nor U25311 (N_25311,N_25137,N_25148);
or U25312 (N_25312,N_25071,N_25119);
xnor U25313 (N_25313,N_25147,N_25027);
or U25314 (N_25314,N_25130,N_25055);
or U25315 (N_25315,N_25138,N_25186);
and U25316 (N_25316,N_25088,N_25146);
xor U25317 (N_25317,N_25021,N_25107);
nand U25318 (N_25318,N_25156,N_25018);
nor U25319 (N_25319,N_25115,N_25131);
xnor U25320 (N_25320,N_25168,N_25148);
or U25321 (N_25321,N_25033,N_25091);
or U25322 (N_25322,N_25084,N_25062);
nand U25323 (N_25323,N_25192,N_25003);
or U25324 (N_25324,N_25055,N_25135);
xnor U25325 (N_25325,N_25161,N_25041);
nand U25326 (N_25326,N_25071,N_25153);
nand U25327 (N_25327,N_25152,N_25119);
nand U25328 (N_25328,N_25116,N_25019);
and U25329 (N_25329,N_25186,N_25194);
and U25330 (N_25330,N_25182,N_25049);
and U25331 (N_25331,N_25016,N_25029);
nand U25332 (N_25332,N_25117,N_25093);
xor U25333 (N_25333,N_25137,N_25047);
and U25334 (N_25334,N_25093,N_25089);
xnor U25335 (N_25335,N_25085,N_25061);
nor U25336 (N_25336,N_25171,N_25166);
and U25337 (N_25337,N_25001,N_25152);
nor U25338 (N_25338,N_25021,N_25187);
nor U25339 (N_25339,N_25014,N_25190);
nand U25340 (N_25340,N_25181,N_25083);
nand U25341 (N_25341,N_25003,N_25094);
and U25342 (N_25342,N_25085,N_25078);
xor U25343 (N_25343,N_25052,N_25174);
and U25344 (N_25344,N_25147,N_25181);
or U25345 (N_25345,N_25144,N_25087);
nor U25346 (N_25346,N_25076,N_25066);
nor U25347 (N_25347,N_25035,N_25135);
or U25348 (N_25348,N_25081,N_25025);
nand U25349 (N_25349,N_25174,N_25118);
and U25350 (N_25350,N_25038,N_25172);
or U25351 (N_25351,N_25169,N_25179);
xor U25352 (N_25352,N_25133,N_25195);
nor U25353 (N_25353,N_25028,N_25180);
or U25354 (N_25354,N_25003,N_25182);
nand U25355 (N_25355,N_25068,N_25072);
nor U25356 (N_25356,N_25159,N_25027);
nand U25357 (N_25357,N_25035,N_25020);
xor U25358 (N_25358,N_25004,N_25177);
xor U25359 (N_25359,N_25150,N_25062);
or U25360 (N_25360,N_25088,N_25090);
and U25361 (N_25361,N_25121,N_25173);
xor U25362 (N_25362,N_25156,N_25127);
and U25363 (N_25363,N_25161,N_25162);
nand U25364 (N_25364,N_25044,N_25147);
or U25365 (N_25365,N_25173,N_25093);
or U25366 (N_25366,N_25003,N_25075);
and U25367 (N_25367,N_25161,N_25072);
or U25368 (N_25368,N_25124,N_25192);
xor U25369 (N_25369,N_25066,N_25102);
xnor U25370 (N_25370,N_25002,N_25085);
or U25371 (N_25371,N_25198,N_25036);
xor U25372 (N_25372,N_25033,N_25164);
nand U25373 (N_25373,N_25043,N_25158);
and U25374 (N_25374,N_25073,N_25113);
or U25375 (N_25375,N_25037,N_25071);
nor U25376 (N_25376,N_25171,N_25089);
nand U25377 (N_25377,N_25073,N_25067);
xor U25378 (N_25378,N_25054,N_25019);
nor U25379 (N_25379,N_25140,N_25168);
nand U25380 (N_25380,N_25142,N_25077);
nand U25381 (N_25381,N_25129,N_25013);
and U25382 (N_25382,N_25109,N_25065);
or U25383 (N_25383,N_25181,N_25187);
xor U25384 (N_25384,N_25098,N_25121);
nor U25385 (N_25385,N_25091,N_25165);
xor U25386 (N_25386,N_25109,N_25070);
nand U25387 (N_25387,N_25027,N_25165);
nand U25388 (N_25388,N_25070,N_25035);
and U25389 (N_25389,N_25018,N_25149);
and U25390 (N_25390,N_25091,N_25118);
xnor U25391 (N_25391,N_25145,N_25144);
and U25392 (N_25392,N_25159,N_25142);
xor U25393 (N_25393,N_25192,N_25151);
nand U25394 (N_25394,N_25124,N_25059);
xnor U25395 (N_25395,N_25005,N_25070);
nand U25396 (N_25396,N_25154,N_25068);
and U25397 (N_25397,N_25099,N_25012);
nor U25398 (N_25398,N_25008,N_25052);
nand U25399 (N_25399,N_25166,N_25191);
or U25400 (N_25400,N_25337,N_25281);
and U25401 (N_25401,N_25266,N_25320);
nor U25402 (N_25402,N_25251,N_25201);
nor U25403 (N_25403,N_25369,N_25319);
xor U25404 (N_25404,N_25203,N_25336);
nor U25405 (N_25405,N_25214,N_25398);
nand U25406 (N_25406,N_25298,N_25274);
or U25407 (N_25407,N_25240,N_25379);
and U25408 (N_25408,N_25211,N_25395);
nand U25409 (N_25409,N_25367,N_25239);
and U25410 (N_25410,N_25287,N_25272);
or U25411 (N_25411,N_25317,N_25318);
xor U25412 (N_25412,N_25200,N_25365);
and U25413 (N_25413,N_25223,N_25300);
nor U25414 (N_25414,N_25275,N_25321);
and U25415 (N_25415,N_25362,N_25227);
nand U25416 (N_25416,N_25270,N_25294);
nand U25417 (N_25417,N_25356,N_25390);
or U25418 (N_25418,N_25267,N_25210);
nand U25419 (N_25419,N_25208,N_25371);
or U25420 (N_25420,N_25396,N_25288);
xor U25421 (N_25421,N_25261,N_25224);
nand U25422 (N_25422,N_25231,N_25233);
nand U25423 (N_25423,N_25361,N_25343);
xor U25424 (N_25424,N_25380,N_25216);
and U25425 (N_25425,N_25333,N_25358);
or U25426 (N_25426,N_25256,N_25282);
and U25427 (N_25427,N_25363,N_25235);
nor U25428 (N_25428,N_25273,N_25276);
nor U25429 (N_25429,N_25241,N_25354);
nor U25430 (N_25430,N_25360,N_25340);
nand U25431 (N_25431,N_25234,N_25329);
and U25432 (N_25432,N_25378,N_25338);
nand U25433 (N_25433,N_25348,N_25301);
and U25434 (N_25434,N_25307,N_25387);
or U25435 (N_25435,N_25215,N_25204);
nand U25436 (N_25436,N_25246,N_25353);
xor U25437 (N_25437,N_25218,N_25255);
xnor U25438 (N_25438,N_25243,N_25334);
nand U25439 (N_25439,N_25264,N_25232);
xor U25440 (N_25440,N_25314,N_25389);
and U25441 (N_25441,N_25268,N_25278);
or U25442 (N_25442,N_25249,N_25346);
or U25443 (N_25443,N_25296,N_25399);
nand U25444 (N_25444,N_25219,N_25238);
nor U25445 (N_25445,N_25323,N_25258);
nand U25446 (N_25446,N_25308,N_25355);
nand U25447 (N_25447,N_25286,N_25388);
and U25448 (N_25448,N_25225,N_25289);
and U25449 (N_25449,N_25228,N_25366);
and U25450 (N_25450,N_25382,N_25259);
or U25451 (N_25451,N_25306,N_25383);
xor U25452 (N_25452,N_25217,N_25357);
nand U25453 (N_25453,N_25253,N_25325);
nor U25454 (N_25454,N_25309,N_25368);
xor U25455 (N_25455,N_25263,N_25326);
or U25456 (N_25456,N_25283,N_25248);
and U25457 (N_25457,N_25359,N_25345);
xor U25458 (N_25458,N_25302,N_25245);
nand U25459 (N_25459,N_25279,N_25271);
xor U25460 (N_25460,N_25242,N_25250);
and U25461 (N_25461,N_25364,N_25290);
nor U25462 (N_25462,N_25206,N_25322);
nand U25463 (N_25463,N_25324,N_25209);
xor U25464 (N_25464,N_25220,N_25376);
or U25465 (N_25465,N_25230,N_25384);
nor U25466 (N_25466,N_25375,N_25377);
nand U25467 (N_25467,N_25202,N_25339);
nand U25468 (N_25468,N_25292,N_25207);
or U25469 (N_25469,N_25293,N_25385);
or U25470 (N_25470,N_25386,N_25370);
and U25471 (N_25471,N_25374,N_25212);
xnor U25472 (N_25472,N_25265,N_25305);
xor U25473 (N_25473,N_25391,N_25229);
xor U25474 (N_25474,N_25311,N_25392);
or U25475 (N_25475,N_25303,N_25285);
or U25476 (N_25476,N_25394,N_25262);
nand U25477 (N_25477,N_25244,N_25269);
nor U25478 (N_25478,N_25299,N_25284);
nor U25479 (N_25479,N_25349,N_25277);
xnor U25480 (N_25480,N_25397,N_25291);
and U25481 (N_25481,N_25222,N_25236);
nor U25482 (N_25482,N_25205,N_25312);
nand U25483 (N_25483,N_25332,N_25342);
or U25484 (N_25484,N_25352,N_25330);
xor U25485 (N_25485,N_25328,N_25247);
or U25486 (N_25486,N_25213,N_25252);
or U25487 (N_25487,N_25310,N_25257);
xnor U25488 (N_25488,N_25260,N_25315);
nand U25489 (N_25489,N_25304,N_25341);
nand U25490 (N_25490,N_25344,N_25373);
xor U25491 (N_25491,N_25350,N_25335);
and U25492 (N_25492,N_25237,N_25316);
nor U25493 (N_25493,N_25313,N_25327);
or U25494 (N_25494,N_25297,N_25280);
or U25495 (N_25495,N_25331,N_25351);
nand U25496 (N_25496,N_25226,N_25295);
nand U25497 (N_25497,N_25372,N_25393);
and U25498 (N_25498,N_25221,N_25347);
nand U25499 (N_25499,N_25381,N_25254);
nor U25500 (N_25500,N_25283,N_25256);
and U25501 (N_25501,N_25333,N_25211);
xnor U25502 (N_25502,N_25269,N_25272);
nor U25503 (N_25503,N_25245,N_25256);
xnor U25504 (N_25504,N_25323,N_25375);
xnor U25505 (N_25505,N_25392,N_25278);
or U25506 (N_25506,N_25232,N_25253);
and U25507 (N_25507,N_25250,N_25213);
xor U25508 (N_25508,N_25356,N_25340);
nand U25509 (N_25509,N_25391,N_25217);
nor U25510 (N_25510,N_25214,N_25284);
and U25511 (N_25511,N_25265,N_25309);
nor U25512 (N_25512,N_25241,N_25281);
nand U25513 (N_25513,N_25366,N_25225);
nand U25514 (N_25514,N_25276,N_25315);
nor U25515 (N_25515,N_25333,N_25204);
nand U25516 (N_25516,N_25391,N_25395);
xnor U25517 (N_25517,N_25385,N_25325);
and U25518 (N_25518,N_25226,N_25301);
xor U25519 (N_25519,N_25367,N_25288);
nand U25520 (N_25520,N_25388,N_25325);
nand U25521 (N_25521,N_25265,N_25335);
nor U25522 (N_25522,N_25345,N_25395);
and U25523 (N_25523,N_25241,N_25377);
nor U25524 (N_25524,N_25369,N_25220);
nand U25525 (N_25525,N_25313,N_25345);
nor U25526 (N_25526,N_25299,N_25294);
or U25527 (N_25527,N_25316,N_25360);
xnor U25528 (N_25528,N_25357,N_25226);
xnor U25529 (N_25529,N_25244,N_25201);
and U25530 (N_25530,N_25358,N_25306);
nor U25531 (N_25531,N_25356,N_25244);
or U25532 (N_25532,N_25247,N_25388);
nor U25533 (N_25533,N_25306,N_25225);
and U25534 (N_25534,N_25344,N_25381);
xor U25535 (N_25535,N_25384,N_25293);
nor U25536 (N_25536,N_25250,N_25209);
nand U25537 (N_25537,N_25358,N_25210);
xor U25538 (N_25538,N_25265,N_25375);
and U25539 (N_25539,N_25259,N_25317);
or U25540 (N_25540,N_25361,N_25320);
and U25541 (N_25541,N_25272,N_25224);
or U25542 (N_25542,N_25318,N_25204);
xor U25543 (N_25543,N_25276,N_25201);
and U25544 (N_25544,N_25330,N_25204);
or U25545 (N_25545,N_25310,N_25350);
nand U25546 (N_25546,N_25206,N_25364);
nor U25547 (N_25547,N_25344,N_25302);
xor U25548 (N_25548,N_25386,N_25241);
nand U25549 (N_25549,N_25296,N_25325);
nand U25550 (N_25550,N_25218,N_25292);
nand U25551 (N_25551,N_25322,N_25390);
xor U25552 (N_25552,N_25363,N_25214);
xor U25553 (N_25553,N_25213,N_25356);
nor U25554 (N_25554,N_25255,N_25318);
or U25555 (N_25555,N_25305,N_25273);
nand U25556 (N_25556,N_25382,N_25200);
xnor U25557 (N_25557,N_25278,N_25366);
nor U25558 (N_25558,N_25391,N_25281);
and U25559 (N_25559,N_25313,N_25230);
nand U25560 (N_25560,N_25296,N_25393);
nand U25561 (N_25561,N_25371,N_25263);
or U25562 (N_25562,N_25307,N_25288);
and U25563 (N_25563,N_25234,N_25287);
xor U25564 (N_25564,N_25367,N_25345);
xnor U25565 (N_25565,N_25236,N_25392);
nor U25566 (N_25566,N_25281,N_25366);
and U25567 (N_25567,N_25320,N_25374);
nand U25568 (N_25568,N_25239,N_25345);
and U25569 (N_25569,N_25246,N_25283);
nand U25570 (N_25570,N_25295,N_25264);
xor U25571 (N_25571,N_25394,N_25393);
nor U25572 (N_25572,N_25390,N_25251);
or U25573 (N_25573,N_25208,N_25391);
or U25574 (N_25574,N_25254,N_25302);
nand U25575 (N_25575,N_25266,N_25335);
and U25576 (N_25576,N_25221,N_25376);
nor U25577 (N_25577,N_25277,N_25358);
nor U25578 (N_25578,N_25306,N_25211);
nand U25579 (N_25579,N_25259,N_25214);
or U25580 (N_25580,N_25394,N_25267);
nor U25581 (N_25581,N_25373,N_25303);
or U25582 (N_25582,N_25289,N_25286);
nand U25583 (N_25583,N_25223,N_25212);
nor U25584 (N_25584,N_25337,N_25376);
nand U25585 (N_25585,N_25271,N_25327);
and U25586 (N_25586,N_25343,N_25297);
nand U25587 (N_25587,N_25349,N_25387);
nor U25588 (N_25588,N_25334,N_25223);
xor U25589 (N_25589,N_25221,N_25343);
xnor U25590 (N_25590,N_25355,N_25259);
and U25591 (N_25591,N_25266,N_25211);
nor U25592 (N_25592,N_25200,N_25206);
nand U25593 (N_25593,N_25297,N_25365);
or U25594 (N_25594,N_25270,N_25203);
xnor U25595 (N_25595,N_25398,N_25365);
and U25596 (N_25596,N_25267,N_25232);
nor U25597 (N_25597,N_25265,N_25376);
or U25598 (N_25598,N_25284,N_25328);
or U25599 (N_25599,N_25231,N_25289);
xnor U25600 (N_25600,N_25411,N_25401);
nor U25601 (N_25601,N_25525,N_25439);
nand U25602 (N_25602,N_25574,N_25431);
nand U25603 (N_25603,N_25597,N_25562);
and U25604 (N_25604,N_25463,N_25555);
nand U25605 (N_25605,N_25424,N_25476);
xor U25606 (N_25606,N_25580,N_25488);
or U25607 (N_25607,N_25414,N_25451);
and U25608 (N_25608,N_25447,N_25455);
nand U25609 (N_25609,N_25446,N_25569);
xnor U25610 (N_25610,N_25575,N_25400);
xor U25611 (N_25611,N_25430,N_25436);
and U25612 (N_25612,N_25462,N_25497);
nor U25613 (N_25613,N_25478,N_25501);
nand U25614 (N_25614,N_25554,N_25568);
xor U25615 (N_25615,N_25523,N_25467);
and U25616 (N_25616,N_25520,N_25507);
and U25617 (N_25617,N_25524,N_25490);
xor U25618 (N_25618,N_25567,N_25543);
nand U25619 (N_25619,N_25416,N_25434);
and U25620 (N_25620,N_25548,N_25449);
and U25621 (N_25621,N_25561,N_25518);
and U25622 (N_25622,N_25421,N_25406);
nand U25623 (N_25623,N_25417,N_25563);
nor U25624 (N_25624,N_25502,N_25544);
and U25625 (N_25625,N_25445,N_25539);
or U25626 (N_25626,N_25547,N_25482);
nor U25627 (N_25627,N_25598,N_25465);
nand U25628 (N_25628,N_25587,N_25441);
nand U25629 (N_25629,N_25536,N_25504);
xor U25630 (N_25630,N_25402,N_25448);
nor U25631 (N_25631,N_25480,N_25531);
and U25632 (N_25632,N_25577,N_25459);
nand U25633 (N_25633,N_25556,N_25509);
xor U25634 (N_25634,N_25530,N_25566);
nand U25635 (N_25635,N_25572,N_25452);
xor U25636 (N_25636,N_25443,N_25422);
nand U25637 (N_25637,N_25475,N_25484);
or U25638 (N_25638,N_25412,N_25586);
xor U25639 (N_25639,N_25517,N_25512);
or U25640 (N_25640,N_25429,N_25468);
xor U25641 (N_25641,N_25408,N_25435);
and U25642 (N_25642,N_25466,N_25485);
nand U25643 (N_25643,N_25546,N_25426);
xnor U25644 (N_25644,N_25511,N_25407);
xnor U25645 (N_25645,N_25469,N_25550);
nand U25646 (N_25646,N_25535,N_25513);
nor U25647 (N_25647,N_25415,N_25489);
nand U25648 (N_25648,N_25405,N_25514);
nand U25649 (N_25649,N_25529,N_25481);
xnor U25650 (N_25650,N_25506,N_25519);
or U25651 (N_25651,N_25464,N_25522);
or U25652 (N_25652,N_25545,N_25599);
nor U25653 (N_25653,N_25591,N_25450);
nor U25654 (N_25654,N_25583,N_25585);
nor U25655 (N_25655,N_25570,N_25565);
nor U25656 (N_25656,N_25596,N_25413);
nor U25657 (N_25657,N_25487,N_25503);
and U25658 (N_25658,N_25582,N_25472);
and U25659 (N_25659,N_25534,N_25456);
nand U25660 (N_25660,N_25578,N_25494);
nor U25661 (N_25661,N_25594,N_25508);
nand U25662 (N_25662,N_25403,N_25595);
xnor U25663 (N_25663,N_25409,N_25540);
nor U25664 (N_25664,N_25526,N_25573);
xnor U25665 (N_25665,N_25495,N_25420);
nor U25666 (N_25666,N_25538,N_25593);
or U25667 (N_25667,N_25427,N_25440);
and U25668 (N_25668,N_25437,N_25558);
nor U25669 (N_25669,N_25527,N_25579);
xnor U25670 (N_25670,N_25552,N_25532);
nor U25671 (N_25671,N_25473,N_25438);
nor U25672 (N_25672,N_25590,N_25533);
or U25673 (N_25673,N_25584,N_25442);
and U25674 (N_25674,N_25454,N_25553);
xor U25675 (N_25675,N_25428,N_25588);
nand U25676 (N_25676,N_25521,N_25433);
and U25677 (N_25677,N_25474,N_25551);
nor U25678 (N_25678,N_25418,N_25589);
or U25679 (N_25679,N_25483,N_25516);
xnor U25680 (N_25680,N_25581,N_25479);
or U25681 (N_25681,N_25499,N_25492);
and U25682 (N_25682,N_25486,N_25457);
and U25683 (N_25683,N_25471,N_25425);
xnor U25684 (N_25684,N_25528,N_25461);
or U25685 (N_25685,N_25549,N_25432);
nor U25686 (N_25686,N_25559,N_25419);
or U25687 (N_25687,N_25477,N_25560);
and U25688 (N_25688,N_25470,N_25505);
xnor U25689 (N_25689,N_25423,N_25458);
nand U25690 (N_25690,N_25498,N_25541);
nor U25691 (N_25691,N_25557,N_25410);
xnor U25692 (N_25692,N_25510,N_25404);
or U25693 (N_25693,N_25571,N_25576);
and U25694 (N_25694,N_25592,N_25515);
and U25695 (N_25695,N_25564,N_25453);
nand U25696 (N_25696,N_25496,N_25444);
and U25697 (N_25697,N_25460,N_25500);
and U25698 (N_25698,N_25491,N_25537);
nand U25699 (N_25699,N_25542,N_25493);
and U25700 (N_25700,N_25441,N_25509);
xnor U25701 (N_25701,N_25436,N_25585);
nand U25702 (N_25702,N_25442,N_25420);
and U25703 (N_25703,N_25504,N_25440);
and U25704 (N_25704,N_25537,N_25439);
nand U25705 (N_25705,N_25445,N_25574);
xnor U25706 (N_25706,N_25425,N_25518);
and U25707 (N_25707,N_25582,N_25578);
xor U25708 (N_25708,N_25464,N_25547);
or U25709 (N_25709,N_25593,N_25433);
and U25710 (N_25710,N_25452,N_25489);
or U25711 (N_25711,N_25442,N_25492);
nor U25712 (N_25712,N_25476,N_25522);
or U25713 (N_25713,N_25474,N_25534);
nor U25714 (N_25714,N_25533,N_25570);
xnor U25715 (N_25715,N_25449,N_25434);
xnor U25716 (N_25716,N_25496,N_25467);
nor U25717 (N_25717,N_25474,N_25431);
nor U25718 (N_25718,N_25596,N_25491);
or U25719 (N_25719,N_25555,N_25572);
xor U25720 (N_25720,N_25581,N_25584);
xor U25721 (N_25721,N_25422,N_25414);
xnor U25722 (N_25722,N_25447,N_25443);
or U25723 (N_25723,N_25568,N_25480);
nor U25724 (N_25724,N_25471,N_25449);
xnor U25725 (N_25725,N_25458,N_25595);
or U25726 (N_25726,N_25551,N_25456);
nand U25727 (N_25727,N_25483,N_25459);
and U25728 (N_25728,N_25401,N_25529);
nor U25729 (N_25729,N_25477,N_25584);
and U25730 (N_25730,N_25549,N_25402);
and U25731 (N_25731,N_25511,N_25429);
nor U25732 (N_25732,N_25489,N_25520);
nand U25733 (N_25733,N_25556,N_25512);
or U25734 (N_25734,N_25495,N_25597);
or U25735 (N_25735,N_25574,N_25444);
and U25736 (N_25736,N_25417,N_25488);
xnor U25737 (N_25737,N_25547,N_25449);
or U25738 (N_25738,N_25497,N_25565);
nor U25739 (N_25739,N_25490,N_25494);
and U25740 (N_25740,N_25502,N_25572);
or U25741 (N_25741,N_25585,N_25437);
xor U25742 (N_25742,N_25506,N_25558);
nor U25743 (N_25743,N_25546,N_25544);
and U25744 (N_25744,N_25519,N_25591);
or U25745 (N_25745,N_25478,N_25462);
nand U25746 (N_25746,N_25568,N_25450);
xor U25747 (N_25747,N_25533,N_25483);
or U25748 (N_25748,N_25529,N_25445);
nor U25749 (N_25749,N_25563,N_25472);
nor U25750 (N_25750,N_25458,N_25412);
and U25751 (N_25751,N_25565,N_25543);
xnor U25752 (N_25752,N_25446,N_25572);
nor U25753 (N_25753,N_25521,N_25419);
nand U25754 (N_25754,N_25527,N_25482);
nor U25755 (N_25755,N_25432,N_25511);
xnor U25756 (N_25756,N_25457,N_25565);
nand U25757 (N_25757,N_25491,N_25444);
and U25758 (N_25758,N_25584,N_25456);
or U25759 (N_25759,N_25528,N_25542);
nor U25760 (N_25760,N_25419,N_25505);
nand U25761 (N_25761,N_25517,N_25531);
and U25762 (N_25762,N_25569,N_25545);
nor U25763 (N_25763,N_25467,N_25590);
xor U25764 (N_25764,N_25581,N_25579);
nand U25765 (N_25765,N_25529,N_25491);
nand U25766 (N_25766,N_25580,N_25508);
or U25767 (N_25767,N_25458,N_25590);
xnor U25768 (N_25768,N_25424,N_25490);
nor U25769 (N_25769,N_25538,N_25501);
xnor U25770 (N_25770,N_25424,N_25571);
and U25771 (N_25771,N_25484,N_25561);
xnor U25772 (N_25772,N_25533,N_25426);
nor U25773 (N_25773,N_25549,N_25476);
xnor U25774 (N_25774,N_25472,N_25574);
nand U25775 (N_25775,N_25423,N_25447);
nand U25776 (N_25776,N_25403,N_25542);
or U25777 (N_25777,N_25502,N_25521);
and U25778 (N_25778,N_25573,N_25595);
and U25779 (N_25779,N_25589,N_25425);
or U25780 (N_25780,N_25493,N_25575);
or U25781 (N_25781,N_25408,N_25406);
and U25782 (N_25782,N_25548,N_25483);
xnor U25783 (N_25783,N_25472,N_25560);
or U25784 (N_25784,N_25584,N_25458);
and U25785 (N_25785,N_25565,N_25510);
or U25786 (N_25786,N_25559,N_25525);
nor U25787 (N_25787,N_25491,N_25581);
nor U25788 (N_25788,N_25435,N_25466);
xnor U25789 (N_25789,N_25404,N_25494);
nand U25790 (N_25790,N_25469,N_25594);
and U25791 (N_25791,N_25528,N_25527);
nand U25792 (N_25792,N_25401,N_25456);
xor U25793 (N_25793,N_25555,N_25584);
nor U25794 (N_25794,N_25523,N_25580);
nor U25795 (N_25795,N_25599,N_25474);
and U25796 (N_25796,N_25486,N_25467);
and U25797 (N_25797,N_25412,N_25434);
xor U25798 (N_25798,N_25516,N_25578);
and U25799 (N_25799,N_25558,N_25436);
nor U25800 (N_25800,N_25600,N_25659);
nor U25801 (N_25801,N_25766,N_25710);
nand U25802 (N_25802,N_25789,N_25604);
or U25803 (N_25803,N_25756,N_25725);
nor U25804 (N_25804,N_25727,N_25745);
and U25805 (N_25805,N_25653,N_25774);
nand U25806 (N_25806,N_25788,N_25677);
xor U25807 (N_25807,N_25735,N_25690);
nand U25808 (N_25808,N_25631,N_25674);
nor U25809 (N_25809,N_25650,N_25623);
nand U25810 (N_25810,N_25684,N_25749);
nand U25811 (N_25811,N_25695,N_25737);
xor U25812 (N_25812,N_25634,N_25638);
or U25813 (N_25813,N_25668,N_25662);
nor U25814 (N_25814,N_25753,N_25757);
and U25815 (N_25815,N_25633,N_25602);
xnor U25816 (N_25816,N_25708,N_25765);
nand U25817 (N_25817,N_25670,N_25726);
or U25818 (N_25818,N_25799,N_25700);
or U25819 (N_25819,N_25618,N_25733);
or U25820 (N_25820,N_25741,N_25762);
nor U25821 (N_25821,N_25760,N_25794);
xor U25822 (N_25822,N_25642,N_25706);
nor U25823 (N_25823,N_25764,N_25782);
nand U25824 (N_25824,N_25730,N_25699);
and U25825 (N_25825,N_25791,N_25786);
or U25826 (N_25826,N_25603,N_25663);
or U25827 (N_25827,N_25629,N_25713);
nor U25828 (N_25828,N_25746,N_25728);
and U25829 (N_25829,N_25647,N_25665);
nor U25830 (N_25830,N_25759,N_25651);
and U25831 (N_25831,N_25722,N_25729);
or U25832 (N_25832,N_25754,N_25705);
xnor U25833 (N_25833,N_25793,N_25641);
nand U25834 (N_25834,N_25798,N_25687);
nand U25835 (N_25835,N_25654,N_25666);
nand U25836 (N_25836,N_25637,N_25776);
nand U25837 (N_25837,N_25620,N_25777);
nor U25838 (N_25838,N_25731,N_25681);
nand U25839 (N_25839,N_25775,N_25652);
nand U25840 (N_25840,N_25640,N_25770);
and U25841 (N_25841,N_25716,N_25625);
nor U25842 (N_25842,N_25704,N_25769);
nand U25843 (N_25843,N_25630,N_25692);
nand U25844 (N_25844,N_25748,N_25667);
nand U25845 (N_25845,N_25619,N_25648);
nor U25846 (N_25846,N_25673,N_25616);
nand U25847 (N_25847,N_25607,N_25610);
and U25848 (N_25848,N_25723,N_25701);
nand U25849 (N_25849,N_25715,N_25635);
and U25850 (N_25850,N_25658,N_25707);
or U25851 (N_25851,N_25724,N_25685);
nor U25852 (N_25852,N_25752,N_25732);
nand U25853 (N_25853,N_25747,N_25767);
nand U25854 (N_25854,N_25661,N_25780);
nor U25855 (N_25855,N_25790,N_25646);
nor U25856 (N_25856,N_25656,N_25622);
nor U25857 (N_25857,N_25721,N_25795);
nor U25858 (N_25858,N_25628,N_25691);
or U25859 (N_25859,N_25696,N_25643);
xor U25860 (N_25860,N_25783,N_25621);
nor U25861 (N_25861,N_25626,N_25739);
and U25862 (N_25862,N_25675,N_25645);
xor U25863 (N_25863,N_25614,N_25712);
xnor U25864 (N_25864,N_25763,N_25669);
nand U25865 (N_25865,N_25608,N_25719);
and U25866 (N_25866,N_25693,N_25718);
nor U25867 (N_25867,N_25717,N_25784);
and U25868 (N_25868,N_25711,N_25688);
nor U25869 (N_25869,N_25778,N_25649);
xnor U25870 (N_25870,N_25613,N_25671);
xor U25871 (N_25871,N_25639,N_25792);
xor U25872 (N_25872,N_25768,N_25697);
and U25873 (N_25873,N_25709,N_25787);
or U25874 (N_25874,N_25796,N_25609);
and U25875 (N_25875,N_25736,N_25627);
nand U25876 (N_25876,N_25664,N_25686);
nor U25877 (N_25877,N_25611,N_25772);
and U25878 (N_25878,N_25742,N_25612);
nor U25879 (N_25879,N_25676,N_25797);
xnor U25880 (N_25880,N_25657,N_25771);
nor U25881 (N_25881,N_25605,N_25624);
or U25882 (N_25882,N_25781,N_25655);
xor U25883 (N_25883,N_25702,N_25714);
or U25884 (N_25884,N_25751,N_25615);
and U25885 (N_25885,N_25678,N_25755);
nand U25886 (N_25886,N_25720,N_25703);
xnor U25887 (N_25887,N_25606,N_25758);
nor U25888 (N_25888,N_25689,N_25785);
nand U25889 (N_25889,N_25682,N_25761);
nand U25890 (N_25890,N_25636,N_25694);
and U25891 (N_25891,N_25601,N_25738);
xnor U25892 (N_25892,N_25779,N_25734);
nand U25893 (N_25893,N_25683,N_25672);
nand U25894 (N_25894,N_25750,N_25644);
or U25895 (N_25895,N_25744,N_25773);
xnor U25896 (N_25896,N_25698,N_25660);
nor U25897 (N_25897,N_25632,N_25679);
xnor U25898 (N_25898,N_25740,N_25743);
or U25899 (N_25899,N_25680,N_25617);
xnor U25900 (N_25900,N_25659,N_25601);
nor U25901 (N_25901,N_25749,N_25737);
nor U25902 (N_25902,N_25657,N_25649);
nor U25903 (N_25903,N_25772,N_25645);
xnor U25904 (N_25904,N_25750,N_25771);
or U25905 (N_25905,N_25768,N_25650);
and U25906 (N_25906,N_25620,N_25657);
nor U25907 (N_25907,N_25710,N_25611);
and U25908 (N_25908,N_25620,N_25769);
or U25909 (N_25909,N_25774,N_25609);
nor U25910 (N_25910,N_25769,N_25718);
nor U25911 (N_25911,N_25607,N_25795);
nor U25912 (N_25912,N_25788,N_25757);
xnor U25913 (N_25913,N_25600,N_25616);
nand U25914 (N_25914,N_25713,N_25760);
xor U25915 (N_25915,N_25637,N_25786);
and U25916 (N_25916,N_25699,N_25749);
xor U25917 (N_25917,N_25631,N_25727);
nor U25918 (N_25918,N_25659,N_25784);
or U25919 (N_25919,N_25749,N_25649);
nand U25920 (N_25920,N_25621,N_25758);
nand U25921 (N_25921,N_25720,N_25657);
and U25922 (N_25922,N_25637,N_25785);
nor U25923 (N_25923,N_25615,N_25742);
xnor U25924 (N_25924,N_25668,N_25658);
nor U25925 (N_25925,N_25753,N_25725);
nand U25926 (N_25926,N_25607,N_25676);
or U25927 (N_25927,N_25738,N_25765);
and U25928 (N_25928,N_25715,N_25720);
xnor U25929 (N_25929,N_25638,N_25729);
nor U25930 (N_25930,N_25603,N_25707);
nand U25931 (N_25931,N_25749,N_25725);
xor U25932 (N_25932,N_25773,N_25724);
or U25933 (N_25933,N_25755,N_25609);
nand U25934 (N_25934,N_25638,N_25747);
nor U25935 (N_25935,N_25752,N_25663);
or U25936 (N_25936,N_25631,N_25793);
or U25937 (N_25937,N_25612,N_25676);
nand U25938 (N_25938,N_25735,N_25604);
nor U25939 (N_25939,N_25707,N_25702);
nor U25940 (N_25940,N_25618,N_25633);
xor U25941 (N_25941,N_25739,N_25613);
nor U25942 (N_25942,N_25730,N_25708);
xnor U25943 (N_25943,N_25752,N_25781);
nor U25944 (N_25944,N_25660,N_25723);
nor U25945 (N_25945,N_25781,N_25641);
nand U25946 (N_25946,N_25782,N_25638);
xnor U25947 (N_25947,N_25685,N_25619);
nand U25948 (N_25948,N_25667,N_25636);
and U25949 (N_25949,N_25743,N_25616);
nor U25950 (N_25950,N_25687,N_25675);
nand U25951 (N_25951,N_25675,N_25600);
nand U25952 (N_25952,N_25607,N_25749);
or U25953 (N_25953,N_25684,N_25735);
and U25954 (N_25954,N_25763,N_25628);
and U25955 (N_25955,N_25646,N_25753);
or U25956 (N_25956,N_25733,N_25736);
nand U25957 (N_25957,N_25695,N_25611);
or U25958 (N_25958,N_25674,N_25645);
nand U25959 (N_25959,N_25715,N_25799);
or U25960 (N_25960,N_25769,N_25749);
xnor U25961 (N_25961,N_25711,N_25623);
nand U25962 (N_25962,N_25794,N_25778);
and U25963 (N_25963,N_25739,N_25618);
nand U25964 (N_25964,N_25751,N_25745);
xnor U25965 (N_25965,N_25619,N_25618);
nand U25966 (N_25966,N_25728,N_25675);
nand U25967 (N_25967,N_25738,N_25761);
xnor U25968 (N_25968,N_25659,N_25783);
and U25969 (N_25969,N_25607,N_25640);
nand U25970 (N_25970,N_25671,N_25644);
and U25971 (N_25971,N_25609,N_25637);
or U25972 (N_25972,N_25693,N_25639);
nand U25973 (N_25973,N_25689,N_25669);
xnor U25974 (N_25974,N_25654,N_25622);
nor U25975 (N_25975,N_25601,N_25792);
or U25976 (N_25976,N_25653,N_25725);
nor U25977 (N_25977,N_25702,N_25688);
nand U25978 (N_25978,N_25743,N_25639);
and U25979 (N_25979,N_25777,N_25657);
and U25980 (N_25980,N_25630,N_25678);
nand U25981 (N_25981,N_25762,N_25672);
xor U25982 (N_25982,N_25683,N_25783);
xor U25983 (N_25983,N_25689,N_25615);
nand U25984 (N_25984,N_25600,N_25718);
nor U25985 (N_25985,N_25788,N_25748);
or U25986 (N_25986,N_25690,N_25667);
nand U25987 (N_25987,N_25779,N_25703);
or U25988 (N_25988,N_25783,N_25635);
or U25989 (N_25989,N_25660,N_25606);
and U25990 (N_25990,N_25649,N_25618);
xnor U25991 (N_25991,N_25633,N_25707);
nand U25992 (N_25992,N_25684,N_25775);
nor U25993 (N_25993,N_25606,N_25782);
or U25994 (N_25994,N_25703,N_25795);
xnor U25995 (N_25995,N_25785,N_25697);
xor U25996 (N_25996,N_25695,N_25635);
and U25997 (N_25997,N_25712,N_25729);
or U25998 (N_25998,N_25762,N_25723);
xor U25999 (N_25999,N_25688,N_25685);
and U26000 (N_26000,N_25972,N_25948);
nor U26001 (N_26001,N_25907,N_25894);
nand U26002 (N_26002,N_25861,N_25831);
and U26003 (N_26003,N_25857,N_25875);
and U26004 (N_26004,N_25837,N_25947);
nand U26005 (N_26005,N_25812,N_25955);
nand U26006 (N_26006,N_25935,N_25844);
nand U26007 (N_26007,N_25827,N_25856);
nand U26008 (N_26008,N_25818,N_25928);
xor U26009 (N_26009,N_25978,N_25884);
or U26010 (N_26010,N_25999,N_25967);
xor U26011 (N_26011,N_25874,N_25880);
nand U26012 (N_26012,N_25905,N_25829);
xnor U26013 (N_26013,N_25866,N_25985);
nand U26014 (N_26014,N_25904,N_25939);
or U26015 (N_26015,N_25919,N_25817);
nand U26016 (N_26016,N_25819,N_25820);
nand U26017 (N_26017,N_25801,N_25941);
and U26018 (N_26018,N_25910,N_25879);
nor U26019 (N_26019,N_25852,N_25997);
nor U26020 (N_26020,N_25952,N_25876);
and U26021 (N_26021,N_25984,N_25983);
xnor U26022 (N_26022,N_25938,N_25925);
or U26023 (N_26023,N_25921,N_25990);
nand U26024 (N_26024,N_25949,N_25940);
nor U26025 (N_26025,N_25897,N_25891);
nor U26026 (N_26026,N_25864,N_25892);
nand U26027 (N_26027,N_25930,N_25973);
xor U26028 (N_26028,N_25834,N_25800);
and U26029 (N_26029,N_25975,N_25903);
nor U26030 (N_26030,N_25974,N_25873);
and U26031 (N_26031,N_25971,N_25946);
nand U26032 (N_26032,N_25806,N_25899);
and U26033 (N_26033,N_25863,N_25872);
nor U26034 (N_26034,N_25900,N_25993);
nand U26035 (N_26035,N_25957,N_25994);
and U26036 (N_26036,N_25916,N_25805);
and U26037 (N_26037,N_25840,N_25867);
nor U26038 (N_26038,N_25944,N_25987);
or U26039 (N_26039,N_25962,N_25917);
xnor U26040 (N_26040,N_25982,N_25803);
nand U26041 (N_26041,N_25881,N_25913);
and U26042 (N_26042,N_25860,N_25854);
nand U26043 (N_26043,N_25804,N_25869);
or U26044 (N_26044,N_25945,N_25963);
nand U26045 (N_26045,N_25835,N_25895);
or U26046 (N_26046,N_25981,N_25968);
nand U26047 (N_26047,N_25960,N_25950);
or U26048 (N_26048,N_25964,N_25845);
nor U26049 (N_26049,N_25901,N_25836);
nor U26050 (N_26050,N_25830,N_25826);
xnor U26051 (N_26051,N_25979,N_25932);
nor U26052 (N_26052,N_25885,N_25889);
or U26053 (N_26053,N_25802,N_25912);
nor U26054 (N_26054,N_25846,N_25886);
or U26055 (N_26055,N_25959,N_25943);
xor U26056 (N_26056,N_25998,N_25855);
and U26057 (N_26057,N_25893,N_25833);
and U26058 (N_26058,N_25936,N_25848);
and U26059 (N_26059,N_25850,N_25961);
nand U26060 (N_26060,N_25847,N_25953);
xnor U26061 (N_26061,N_25911,N_25989);
and U26062 (N_26062,N_25821,N_25858);
or U26063 (N_26063,N_25877,N_25976);
or U26064 (N_26064,N_25914,N_25988);
xnor U26065 (N_26065,N_25926,N_25839);
nor U26066 (N_26066,N_25832,N_25809);
and U26067 (N_26067,N_25843,N_25920);
nand U26068 (N_26068,N_25922,N_25842);
nor U26069 (N_26069,N_25813,N_25808);
and U26070 (N_26070,N_25966,N_25896);
nand U26071 (N_26071,N_25924,N_25906);
nor U26072 (N_26072,N_25824,N_25942);
nand U26073 (N_26073,N_25902,N_25853);
nor U26074 (N_26074,N_25986,N_25883);
or U26075 (N_26075,N_25882,N_25996);
nor U26076 (N_26076,N_25898,N_25927);
nand U26077 (N_26077,N_25908,N_25954);
and U26078 (N_26078,N_25825,N_25851);
nor U26079 (N_26079,N_25870,N_25977);
or U26080 (N_26080,N_25992,N_25965);
and U26081 (N_26081,N_25937,N_25991);
and U26082 (N_26082,N_25887,N_25995);
and U26083 (N_26083,N_25822,N_25807);
or U26084 (N_26084,N_25811,N_25823);
nand U26085 (N_26085,N_25909,N_25878);
or U26086 (N_26086,N_25828,N_25810);
nand U26087 (N_26087,N_25918,N_25888);
and U26088 (N_26088,N_25951,N_25865);
nor U26089 (N_26089,N_25929,N_25868);
or U26090 (N_26090,N_25956,N_25890);
and U26091 (N_26091,N_25969,N_25871);
nor U26092 (N_26092,N_25970,N_25859);
nand U26093 (N_26093,N_25862,N_25933);
nor U26094 (N_26094,N_25814,N_25815);
xnor U26095 (N_26095,N_25980,N_25838);
xor U26096 (N_26096,N_25816,N_25849);
nor U26097 (N_26097,N_25841,N_25923);
and U26098 (N_26098,N_25934,N_25915);
nand U26099 (N_26099,N_25931,N_25958);
xor U26100 (N_26100,N_25807,N_25921);
nor U26101 (N_26101,N_25862,N_25902);
or U26102 (N_26102,N_25825,N_25800);
and U26103 (N_26103,N_25999,N_25906);
or U26104 (N_26104,N_25800,N_25864);
xnor U26105 (N_26105,N_25983,N_25995);
or U26106 (N_26106,N_25946,N_25942);
and U26107 (N_26107,N_25890,N_25899);
nand U26108 (N_26108,N_25965,N_25932);
and U26109 (N_26109,N_25862,N_25842);
xor U26110 (N_26110,N_25979,N_25825);
xnor U26111 (N_26111,N_25994,N_25952);
and U26112 (N_26112,N_25929,N_25908);
and U26113 (N_26113,N_25882,N_25986);
nand U26114 (N_26114,N_25961,N_25848);
or U26115 (N_26115,N_25807,N_25814);
and U26116 (N_26116,N_25820,N_25806);
nor U26117 (N_26117,N_25978,N_25916);
nand U26118 (N_26118,N_25838,N_25998);
nor U26119 (N_26119,N_25929,N_25958);
nand U26120 (N_26120,N_25815,N_25839);
nand U26121 (N_26121,N_25884,N_25847);
xnor U26122 (N_26122,N_25835,N_25944);
and U26123 (N_26123,N_25864,N_25905);
or U26124 (N_26124,N_25932,N_25883);
nor U26125 (N_26125,N_25931,N_25864);
nor U26126 (N_26126,N_25872,N_25903);
or U26127 (N_26127,N_25936,N_25982);
or U26128 (N_26128,N_25991,N_25921);
xnor U26129 (N_26129,N_25955,N_25855);
nor U26130 (N_26130,N_25860,N_25924);
xnor U26131 (N_26131,N_25843,N_25959);
xnor U26132 (N_26132,N_25911,N_25858);
xor U26133 (N_26133,N_25894,N_25831);
and U26134 (N_26134,N_25993,N_25979);
nor U26135 (N_26135,N_25855,N_25858);
nor U26136 (N_26136,N_25958,N_25889);
nor U26137 (N_26137,N_25930,N_25901);
xnor U26138 (N_26138,N_25842,N_25930);
or U26139 (N_26139,N_25874,N_25906);
and U26140 (N_26140,N_25831,N_25953);
nand U26141 (N_26141,N_25976,N_25986);
nor U26142 (N_26142,N_25885,N_25966);
xnor U26143 (N_26143,N_25823,N_25966);
nor U26144 (N_26144,N_25840,N_25931);
nor U26145 (N_26145,N_25883,N_25865);
or U26146 (N_26146,N_25834,N_25930);
nor U26147 (N_26147,N_25945,N_25999);
nand U26148 (N_26148,N_25837,N_25959);
or U26149 (N_26149,N_25892,N_25802);
or U26150 (N_26150,N_25904,N_25959);
nor U26151 (N_26151,N_25869,N_25807);
xnor U26152 (N_26152,N_25841,N_25801);
or U26153 (N_26153,N_25821,N_25930);
nor U26154 (N_26154,N_25974,N_25981);
or U26155 (N_26155,N_25954,N_25906);
xor U26156 (N_26156,N_25828,N_25939);
nand U26157 (N_26157,N_25925,N_25833);
and U26158 (N_26158,N_25919,N_25991);
xnor U26159 (N_26159,N_25990,N_25930);
nor U26160 (N_26160,N_25802,N_25809);
and U26161 (N_26161,N_25845,N_25945);
and U26162 (N_26162,N_25887,N_25955);
xnor U26163 (N_26163,N_25890,N_25941);
and U26164 (N_26164,N_25993,N_25918);
xnor U26165 (N_26165,N_25835,N_25960);
or U26166 (N_26166,N_25815,N_25964);
and U26167 (N_26167,N_25902,N_25893);
and U26168 (N_26168,N_25996,N_25908);
or U26169 (N_26169,N_25837,N_25839);
or U26170 (N_26170,N_25932,N_25867);
nand U26171 (N_26171,N_25975,N_25977);
or U26172 (N_26172,N_25880,N_25970);
xor U26173 (N_26173,N_25899,N_25811);
and U26174 (N_26174,N_25989,N_25928);
nor U26175 (N_26175,N_25989,N_25942);
or U26176 (N_26176,N_25967,N_25833);
or U26177 (N_26177,N_25862,N_25964);
or U26178 (N_26178,N_25882,N_25958);
or U26179 (N_26179,N_25993,N_25864);
or U26180 (N_26180,N_25992,N_25961);
and U26181 (N_26181,N_25977,N_25824);
nand U26182 (N_26182,N_25893,N_25822);
nand U26183 (N_26183,N_25990,N_25950);
nand U26184 (N_26184,N_25851,N_25860);
nand U26185 (N_26185,N_25850,N_25860);
xnor U26186 (N_26186,N_25941,N_25875);
xor U26187 (N_26187,N_25972,N_25975);
nand U26188 (N_26188,N_25978,N_25819);
and U26189 (N_26189,N_25973,N_25855);
xnor U26190 (N_26190,N_25830,N_25864);
xnor U26191 (N_26191,N_25919,N_25825);
nand U26192 (N_26192,N_25924,N_25892);
nand U26193 (N_26193,N_25982,N_25897);
and U26194 (N_26194,N_25840,N_25964);
and U26195 (N_26195,N_25876,N_25961);
nor U26196 (N_26196,N_25953,N_25881);
nand U26197 (N_26197,N_25853,N_25999);
nand U26198 (N_26198,N_25972,N_25965);
or U26199 (N_26199,N_25897,N_25804);
or U26200 (N_26200,N_26134,N_26176);
nor U26201 (N_26201,N_26000,N_26180);
nor U26202 (N_26202,N_26058,N_26089);
xnor U26203 (N_26203,N_26175,N_26139);
nand U26204 (N_26204,N_26022,N_26094);
or U26205 (N_26205,N_26171,N_26132);
nor U26206 (N_26206,N_26034,N_26083);
nand U26207 (N_26207,N_26052,N_26152);
xnor U26208 (N_26208,N_26194,N_26010);
xnor U26209 (N_26209,N_26151,N_26140);
nor U26210 (N_26210,N_26019,N_26091);
nor U26211 (N_26211,N_26055,N_26046);
and U26212 (N_26212,N_26027,N_26100);
or U26213 (N_26213,N_26079,N_26068);
nor U26214 (N_26214,N_26125,N_26062);
nor U26215 (N_26215,N_26076,N_26072);
xnor U26216 (N_26216,N_26020,N_26098);
xnor U26217 (N_26217,N_26031,N_26166);
and U26218 (N_26218,N_26186,N_26084);
and U26219 (N_26219,N_26118,N_26016);
nand U26220 (N_26220,N_26156,N_26197);
or U26221 (N_26221,N_26012,N_26026);
or U26222 (N_26222,N_26102,N_26167);
xor U26223 (N_26223,N_26150,N_26008);
and U26224 (N_26224,N_26159,N_26173);
nor U26225 (N_26225,N_26169,N_26090);
and U26226 (N_26226,N_26121,N_26093);
or U26227 (N_26227,N_26196,N_26145);
nor U26228 (N_26228,N_26104,N_26047);
and U26229 (N_26229,N_26006,N_26028);
nand U26230 (N_26230,N_26048,N_26185);
nor U26231 (N_26231,N_26127,N_26191);
nand U26232 (N_26232,N_26192,N_26190);
nor U26233 (N_26233,N_26038,N_26074);
nor U26234 (N_26234,N_26099,N_26130);
nand U26235 (N_26235,N_26025,N_26164);
or U26236 (N_26236,N_26161,N_26040);
and U26237 (N_26237,N_26108,N_26182);
xnor U26238 (N_26238,N_26135,N_26071);
xor U26239 (N_26239,N_26122,N_26106);
nor U26240 (N_26240,N_26039,N_26033);
xor U26241 (N_26241,N_26177,N_26018);
or U26242 (N_26242,N_26195,N_26137);
xor U26243 (N_26243,N_26148,N_26172);
and U26244 (N_26244,N_26045,N_26075);
nor U26245 (N_26245,N_26157,N_26041);
xnor U26246 (N_26246,N_26111,N_26069);
or U26247 (N_26247,N_26126,N_26032);
nor U26248 (N_26248,N_26014,N_26184);
nor U26249 (N_26249,N_26149,N_26163);
nor U26250 (N_26250,N_26117,N_26054);
and U26251 (N_26251,N_26120,N_26154);
xor U26252 (N_26252,N_26059,N_26114);
or U26253 (N_26253,N_26086,N_26128);
or U26254 (N_26254,N_26035,N_26060);
nand U26255 (N_26255,N_26170,N_26065);
nor U26256 (N_26256,N_26049,N_26073);
xor U26257 (N_26257,N_26187,N_26042);
xor U26258 (N_26258,N_26110,N_26043);
or U26259 (N_26259,N_26015,N_26189);
or U26260 (N_26260,N_26005,N_26013);
xor U26261 (N_26261,N_26188,N_26051);
or U26262 (N_26262,N_26095,N_26179);
xnor U26263 (N_26263,N_26002,N_26142);
or U26264 (N_26264,N_26001,N_26107);
or U26265 (N_26265,N_26178,N_26160);
and U26266 (N_26266,N_26165,N_26168);
and U26267 (N_26267,N_26029,N_26081);
nand U26268 (N_26268,N_26153,N_26077);
nor U26269 (N_26269,N_26143,N_26063);
nor U26270 (N_26270,N_26085,N_26101);
nand U26271 (N_26271,N_26078,N_26003);
nor U26272 (N_26272,N_26183,N_26096);
nand U26273 (N_26273,N_26199,N_26080);
or U26274 (N_26274,N_26037,N_26082);
nand U26275 (N_26275,N_26129,N_26056);
nand U26276 (N_26276,N_26017,N_26158);
xnor U26277 (N_26277,N_26123,N_26133);
or U26278 (N_26278,N_26105,N_26144);
or U26279 (N_26279,N_26004,N_26024);
or U26280 (N_26280,N_26162,N_26193);
or U26281 (N_26281,N_26174,N_26147);
xnor U26282 (N_26282,N_26097,N_26141);
and U26283 (N_26283,N_26007,N_26064);
or U26284 (N_26284,N_26112,N_26011);
xor U26285 (N_26285,N_26087,N_26030);
xnor U26286 (N_26286,N_26103,N_26009);
and U26287 (N_26287,N_26131,N_26113);
nand U26288 (N_26288,N_26061,N_26181);
or U26289 (N_26289,N_26109,N_26116);
xor U26290 (N_26290,N_26146,N_26136);
nor U26291 (N_26291,N_26115,N_26138);
nor U26292 (N_26292,N_26198,N_26050);
nand U26293 (N_26293,N_26124,N_26092);
nor U26294 (N_26294,N_26070,N_26088);
nand U26295 (N_26295,N_26023,N_26053);
nor U26296 (N_26296,N_26057,N_26067);
nand U26297 (N_26297,N_26021,N_26119);
and U26298 (N_26298,N_26044,N_26036);
or U26299 (N_26299,N_26066,N_26155);
and U26300 (N_26300,N_26034,N_26013);
nor U26301 (N_26301,N_26185,N_26039);
nand U26302 (N_26302,N_26189,N_26160);
and U26303 (N_26303,N_26085,N_26105);
or U26304 (N_26304,N_26181,N_26103);
xnor U26305 (N_26305,N_26139,N_26099);
xnor U26306 (N_26306,N_26199,N_26003);
nor U26307 (N_26307,N_26038,N_26170);
nor U26308 (N_26308,N_26105,N_26080);
or U26309 (N_26309,N_26091,N_26094);
and U26310 (N_26310,N_26189,N_26029);
nand U26311 (N_26311,N_26056,N_26171);
or U26312 (N_26312,N_26095,N_26184);
nor U26313 (N_26313,N_26179,N_26101);
or U26314 (N_26314,N_26132,N_26107);
nand U26315 (N_26315,N_26120,N_26107);
nor U26316 (N_26316,N_26102,N_26012);
xnor U26317 (N_26317,N_26113,N_26050);
or U26318 (N_26318,N_26112,N_26051);
xor U26319 (N_26319,N_26123,N_26161);
or U26320 (N_26320,N_26018,N_26132);
xnor U26321 (N_26321,N_26090,N_26016);
nor U26322 (N_26322,N_26003,N_26039);
xnor U26323 (N_26323,N_26010,N_26165);
xnor U26324 (N_26324,N_26150,N_26065);
xnor U26325 (N_26325,N_26149,N_26160);
or U26326 (N_26326,N_26194,N_26136);
and U26327 (N_26327,N_26075,N_26027);
nor U26328 (N_26328,N_26089,N_26044);
nor U26329 (N_26329,N_26124,N_26055);
and U26330 (N_26330,N_26095,N_26041);
or U26331 (N_26331,N_26100,N_26157);
or U26332 (N_26332,N_26045,N_26179);
or U26333 (N_26333,N_26135,N_26199);
nand U26334 (N_26334,N_26009,N_26140);
nor U26335 (N_26335,N_26066,N_26011);
nand U26336 (N_26336,N_26007,N_26076);
nand U26337 (N_26337,N_26187,N_26112);
nand U26338 (N_26338,N_26129,N_26143);
nand U26339 (N_26339,N_26075,N_26074);
nor U26340 (N_26340,N_26062,N_26113);
nor U26341 (N_26341,N_26177,N_26136);
and U26342 (N_26342,N_26010,N_26183);
xnor U26343 (N_26343,N_26039,N_26115);
xnor U26344 (N_26344,N_26014,N_26082);
xnor U26345 (N_26345,N_26012,N_26166);
xnor U26346 (N_26346,N_26183,N_26013);
and U26347 (N_26347,N_26081,N_26041);
nor U26348 (N_26348,N_26143,N_26079);
or U26349 (N_26349,N_26015,N_26044);
nor U26350 (N_26350,N_26070,N_26011);
nor U26351 (N_26351,N_26069,N_26183);
xnor U26352 (N_26352,N_26180,N_26053);
and U26353 (N_26353,N_26023,N_26097);
nor U26354 (N_26354,N_26007,N_26093);
or U26355 (N_26355,N_26169,N_26029);
and U26356 (N_26356,N_26013,N_26016);
nor U26357 (N_26357,N_26149,N_26035);
nand U26358 (N_26358,N_26171,N_26133);
nand U26359 (N_26359,N_26156,N_26192);
nor U26360 (N_26360,N_26013,N_26075);
and U26361 (N_26361,N_26006,N_26179);
nor U26362 (N_26362,N_26164,N_26146);
or U26363 (N_26363,N_26009,N_26117);
nor U26364 (N_26364,N_26130,N_26019);
nor U26365 (N_26365,N_26038,N_26027);
or U26366 (N_26366,N_26023,N_26118);
or U26367 (N_26367,N_26013,N_26196);
and U26368 (N_26368,N_26170,N_26199);
and U26369 (N_26369,N_26149,N_26171);
and U26370 (N_26370,N_26156,N_26033);
and U26371 (N_26371,N_26039,N_26188);
or U26372 (N_26372,N_26104,N_26166);
xor U26373 (N_26373,N_26080,N_26148);
xor U26374 (N_26374,N_26170,N_26100);
or U26375 (N_26375,N_26179,N_26001);
or U26376 (N_26376,N_26171,N_26042);
nor U26377 (N_26377,N_26128,N_26079);
nor U26378 (N_26378,N_26174,N_26047);
nor U26379 (N_26379,N_26128,N_26199);
and U26380 (N_26380,N_26052,N_26061);
and U26381 (N_26381,N_26129,N_26030);
and U26382 (N_26382,N_26086,N_26096);
xor U26383 (N_26383,N_26193,N_26032);
and U26384 (N_26384,N_26102,N_26025);
xor U26385 (N_26385,N_26174,N_26136);
nor U26386 (N_26386,N_26174,N_26154);
and U26387 (N_26387,N_26199,N_26032);
and U26388 (N_26388,N_26073,N_26072);
nor U26389 (N_26389,N_26084,N_26023);
and U26390 (N_26390,N_26065,N_26154);
nor U26391 (N_26391,N_26150,N_26134);
and U26392 (N_26392,N_26157,N_26163);
or U26393 (N_26393,N_26081,N_26130);
or U26394 (N_26394,N_26193,N_26059);
xor U26395 (N_26395,N_26101,N_26111);
and U26396 (N_26396,N_26082,N_26126);
xor U26397 (N_26397,N_26065,N_26086);
and U26398 (N_26398,N_26128,N_26013);
or U26399 (N_26399,N_26150,N_26063);
xor U26400 (N_26400,N_26350,N_26310);
nand U26401 (N_26401,N_26294,N_26321);
xnor U26402 (N_26402,N_26317,N_26258);
nor U26403 (N_26403,N_26279,N_26335);
or U26404 (N_26404,N_26344,N_26233);
and U26405 (N_26405,N_26360,N_26222);
nand U26406 (N_26406,N_26251,N_26383);
and U26407 (N_26407,N_26303,N_26237);
and U26408 (N_26408,N_26220,N_26302);
and U26409 (N_26409,N_26327,N_26359);
and U26410 (N_26410,N_26299,N_26292);
or U26411 (N_26411,N_26297,N_26382);
nand U26412 (N_26412,N_26367,N_26380);
nand U26413 (N_26413,N_26241,N_26284);
and U26414 (N_26414,N_26267,N_26374);
nor U26415 (N_26415,N_26323,N_26266);
nor U26416 (N_26416,N_26261,N_26242);
nand U26417 (N_26417,N_26214,N_26260);
and U26418 (N_26418,N_26304,N_26391);
or U26419 (N_26419,N_26243,N_26217);
nand U26420 (N_26420,N_26291,N_26373);
and U26421 (N_26421,N_26215,N_26330);
nand U26422 (N_26422,N_26388,N_26309);
and U26423 (N_26423,N_26308,N_26311);
xor U26424 (N_26424,N_26329,N_26305);
nor U26425 (N_26425,N_26399,N_26244);
and U26426 (N_26426,N_26259,N_26378);
xor U26427 (N_26427,N_26226,N_26298);
nand U26428 (N_26428,N_26318,N_26338);
xnor U26429 (N_26429,N_26264,N_26315);
and U26430 (N_26430,N_26246,N_26366);
xnor U26431 (N_26431,N_26393,N_26219);
and U26432 (N_26432,N_26387,N_26397);
nand U26433 (N_26433,N_26232,N_26396);
xnor U26434 (N_26434,N_26265,N_26274);
nand U26435 (N_26435,N_26370,N_26349);
xnor U26436 (N_26436,N_26272,N_26293);
or U26437 (N_26437,N_26372,N_26342);
nand U26438 (N_26438,N_26336,N_26256);
nor U26439 (N_26439,N_26250,N_26202);
and U26440 (N_26440,N_26263,N_26351);
nand U26441 (N_26441,N_26249,N_26319);
nand U26442 (N_26442,N_26312,N_26296);
and U26443 (N_26443,N_26276,N_26239);
nor U26444 (N_26444,N_26283,N_26295);
and U26445 (N_26445,N_26270,N_26245);
or U26446 (N_26446,N_26314,N_26201);
nor U26447 (N_26447,N_26365,N_26255);
or U26448 (N_26448,N_26223,N_26271);
or U26449 (N_26449,N_26353,N_26326);
or U26450 (N_26450,N_26205,N_26213);
nand U26451 (N_26451,N_26355,N_26254);
xor U26452 (N_26452,N_26324,N_26231);
and U26453 (N_26453,N_26203,N_26225);
and U26454 (N_26454,N_26207,N_26262);
nand U26455 (N_26455,N_26313,N_26368);
or U26456 (N_26456,N_26362,N_26273);
nor U26457 (N_26457,N_26369,N_26381);
nor U26458 (N_26458,N_26307,N_26301);
xnor U26459 (N_26459,N_26257,N_26332);
nand U26460 (N_26460,N_26320,N_26281);
xnor U26461 (N_26461,N_26364,N_26227);
or U26462 (N_26462,N_26371,N_26376);
xnor U26463 (N_26463,N_26253,N_26287);
nor U26464 (N_26464,N_26218,N_26334);
and U26465 (N_26465,N_26200,N_26356);
nor U26466 (N_26466,N_26348,N_26210);
or U26467 (N_26467,N_26322,N_26390);
nor U26468 (N_26468,N_26386,N_26238);
xnor U26469 (N_26469,N_26275,N_26394);
and U26470 (N_26470,N_26288,N_26280);
nand U26471 (N_26471,N_26340,N_26343);
or U26472 (N_26472,N_26385,N_26268);
xor U26473 (N_26473,N_26247,N_26229);
xnor U26474 (N_26474,N_26300,N_26252);
nor U26475 (N_26475,N_26361,N_26224);
nand U26476 (N_26476,N_26289,N_26316);
or U26477 (N_26477,N_26206,N_26354);
and U26478 (N_26478,N_26337,N_26240);
nor U26479 (N_26479,N_26395,N_26375);
xnor U26480 (N_26480,N_26285,N_26346);
nand U26481 (N_26481,N_26333,N_26234);
xor U26482 (N_26482,N_26352,N_26212);
nor U26483 (N_26483,N_26392,N_26357);
and U26484 (N_26484,N_26384,N_26228);
nor U26485 (N_26485,N_26211,N_26277);
or U26486 (N_26486,N_26230,N_26236);
and U26487 (N_26487,N_26363,N_26286);
xnor U26488 (N_26488,N_26221,N_26379);
nand U26489 (N_26489,N_26278,N_26248);
and U26490 (N_26490,N_26398,N_26209);
or U26491 (N_26491,N_26269,N_26216);
and U26492 (N_26492,N_26235,N_26306);
or U26493 (N_26493,N_26204,N_26208);
nand U26494 (N_26494,N_26377,N_26331);
xnor U26495 (N_26495,N_26345,N_26341);
or U26496 (N_26496,N_26347,N_26389);
and U26497 (N_26497,N_26328,N_26339);
nor U26498 (N_26498,N_26290,N_26325);
nand U26499 (N_26499,N_26358,N_26282);
xnor U26500 (N_26500,N_26239,N_26371);
xor U26501 (N_26501,N_26353,N_26313);
and U26502 (N_26502,N_26238,N_26359);
nand U26503 (N_26503,N_26351,N_26244);
and U26504 (N_26504,N_26307,N_26280);
nand U26505 (N_26505,N_26237,N_26356);
nor U26506 (N_26506,N_26302,N_26269);
nand U26507 (N_26507,N_26366,N_26270);
xnor U26508 (N_26508,N_26243,N_26200);
xor U26509 (N_26509,N_26217,N_26230);
nand U26510 (N_26510,N_26358,N_26248);
nor U26511 (N_26511,N_26228,N_26236);
or U26512 (N_26512,N_26397,N_26287);
xnor U26513 (N_26513,N_26236,N_26399);
and U26514 (N_26514,N_26294,N_26348);
and U26515 (N_26515,N_26388,N_26379);
or U26516 (N_26516,N_26235,N_26356);
xnor U26517 (N_26517,N_26233,N_26210);
nand U26518 (N_26518,N_26361,N_26200);
and U26519 (N_26519,N_26224,N_26294);
or U26520 (N_26520,N_26293,N_26394);
nand U26521 (N_26521,N_26205,N_26238);
nand U26522 (N_26522,N_26230,N_26286);
nor U26523 (N_26523,N_26208,N_26212);
or U26524 (N_26524,N_26341,N_26337);
nor U26525 (N_26525,N_26275,N_26225);
xor U26526 (N_26526,N_26380,N_26273);
or U26527 (N_26527,N_26311,N_26380);
and U26528 (N_26528,N_26312,N_26289);
nand U26529 (N_26529,N_26340,N_26399);
or U26530 (N_26530,N_26343,N_26396);
nor U26531 (N_26531,N_26249,N_26362);
nor U26532 (N_26532,N_26332,N_26200);
xnor U26533 (N_26533,N_26368,N_26216);
and U26534 (N_26534,N_26395,N_26336);
nand U26535 (N_26535,N_26373,N_26374);
nand U26536 (N_26536,N_26374,N_26249);
xor U26537 (N_26537,N_26336,N_26372);
and U26538 (N_26538,N_26379,N_26317);
nand U26539 (N_26539,N_26334,N_26394);
and U26540 (N_26540,N_26269,N_26328);
xor U26541 (N_26541,N_26272,N_26370);
nor U26542 (N_26542,N_26231,N_26384);
nand U26543 (N_26543,N_26263,N_26341);
xnor U26544 (N_26544,N_26322,N_26255);
or U26545 (N_26545,N_26340,N_26254);
xnor U26546 (N_26546,N_26368,N_26294);
xor U26547 (N_26547,N_26350,N_26382);
xor U26548 (N_26548,N_26258,N_26304);
xor U26549 (N_26549,N_26229,N_26383);
and U26550 (N_26550,N_26341,N_26308);
xnor U26551 (N_26551,N_26284,N_26205);
and U26552 (N_26552,N_26326,N_26394);
nand U26553 (N_26553,N_26290,N_26333);
and U26554 (N_26554,N_26326,N_26286);
or U26555 (N_26555,N_26234,N_26355);
and U26556 (N_26556,N_26285,N_26396);
nor U26557 (N_26557,N_26253,N_26364);
xor U26558 (N_26558,N_26365,N_26277);
xor U26559 (N_26559,N_26234,N_26325);
nand U26560 (N_26560,N_26347,N_26280);
or U26561 (N_26561,N_26203,N_26370);
or U26562 (N_26562,N_26364,N_26219);
or U26563 (N_26563,N_26360,N_26303);
nand U26564 (N_26564,N_26210,N_26279);
and U26565 (N_26565,N_26340,N_26398);
xor U26566 (N_26566,N_26238,N_26316);
and U26567 (N_26567,N_26207,N_26394);
xor U26568 (N_26568,N_26313,N_26328);
or U26569 (N_26569,N_26332,N_26370);
nor U26570 (N_26570,N_26282,N_26296);
xnor U26571 (N_26571,N_26376,N_26241);
or U26572 (N_26572,N_26394,N_26320);
and U26573 (N_26573,N_26383,N_26235);
or U26574 (N_26574,N_26365,N_26328);
and U26575 (N_26575,N_26320,N_26362);
nand U26576 (N_26576,N_26277,N_26212);
and U26577 (N_26577,N_26378,N_26384);
or U26578 (N_26578,N_26330,N_26305);
and U26579 (N_26579,N_26348,N_26277);
nor U26580 (N_26580,N_26302,N_26213);
nand U26581 (N_26581,N_26374,N_26318);
nor U26582 (N_26582,N_26283,N_26332);
or U26583 (N_26583,N_26325,N_26373);
nand U26584 (N_26584,N_26254,N_26215);
nand U26585 (N_26585,N_26332,N_26362);
nor U26586 (N_26586,N_26378,N_26310);
nand U26587 (N_26587,N_26398,N_26213);
nor U26588 (N_26588,N_26315,N_26268);
nand U26589 (N_26589,N_26389,N_26326);
or U26590 (N_26590,N_26328,N_26292);
nand U26591 (N_26591,N_26232,N_26329);
or U26592 (N_26592,N_26312,N_26233);
nor U26593 (N_26593,N_26237,N_26377);
nand U26594 (N_26594,N_26261,N_26237);
and U26595 (N_26595,N_26255,N_26274);
nand U26596 (N_26596,N_26203,N_26358);
or U26597 (N_26597,N_26203,N_26264);
nor U26598 (N_26598,N_26333,N_26279);
xnor U26599 (N_26599,N_26314,N_26340);
nand U26600 (N_26600,N_26400,N_26558);
nand U26601 (N_26601,N_26472,N_26473);
or U26602 (N_26602,N_26403,N_26542);
and U26603 (N_26603,N_26545,N_26439);
nand U26604 (N_26604,N_26499,N_26429);
and U26605 (N_26605,N_26547,N_26583);
nand U26606 (N_26606,N_26581,N_26511);
xnor U26607 (N_26607,N_26577,N_26526);
xor U26608 (N_26608,N_26584,N_26458);
or U26609 (N_26609,N_26470,N_26559);
and U26610 (N_26610,N_26405,N_26446);
or U26611 (N_26611,N_26563,N_26460);
nor U26612 (N_26612,N_26505,N_26415);
or U26613 (N_26613,N_26543,N_26532);
nand U26614 (N_26614,N_26561,N_26567);
or U26615 (N_26615,N_26548,N_26442);
xnor U26616 (N_26616,N_26433,N_26503);
nand U26617 (N_26617,N_26578,N_26535);
nand U26618 (N_26618,N_26564,N_26410);
nand U26619 (N_26619,N_26518,N_26420);
nor U26620 (N_26620,N_26438,N_26588);
xor U26621 (N_26621,N_26457,N_26557);
xor U26622 (N_26622,N_26521,N_26502);
or U26623 (N_26623,N_26407,N_26412);
nand U26624 (N_26624,N_26556,N_26476);
or U26625 (N_26625,N_26538,N_26540);
or U26626 (N_26626,N_26527,N_26454);
or U26627 (N_26627,N_26534,N_26597);
and U26628 (N_26628,N_26552,N_26435);
and U26629 (N_26629,N_26553,N_26569);
and U26630 (N_26630,N_26571,N_26546);
nand U26631 (N_26631,N_26479,N_26582);
or U26632 (N_26632,N_26555,N_26523);
or U26633 (N_26633,N_26531,N_26414);
nor U26634 (N_26634,N_26507,N_26508);
or U26635 (N_26635,N_26536,N_26506);
nand U26636 (N_26636,N_26539,N_26444);
and U26637 (N_26637,N_26486,N_26464);
nor U26638 (N_26638,N_26504,N_26490);
and U26639 (N_26639,N_26431,N_26576);
xnor U26640 (N_26640,N_26537,N_26560);
xor U26641 (N_26641,N_26580,N_26425);
or U26642 (N_26642,N_26519,N_26474);
or U26643 (N_26643,N_26497,N_26402);
or U26644 (N_26644,N_26598,N_26409);
nor U26645 (N_26645,N_26517,N_26418);
xor U26646 (N_26646,N_26530,N_26411);
nor U26647 (N_26647,N_26516,N_26453);
and U26648 (N_26648,N_26466,N_26417);
nor U26649 (N_26649,N_26436,N_26572);
nor U26650 (N_26650,N_26467,N_26512);
nor U26651 (N_26651,N_26586,N_26492);
nand U26652 (N_26652,N_26449,N_26595);
nand U26653 (N_26653,N_26599,N_26533);
and U26654 (N_26654,N_26522,N_26437);
nor U26655 (N_26655,N_26591,N_26477);
xnor U26656 (N_26656,N_26524,N_26424);
and U26657 (N_26657,N_26423,N_26450);
or U26658 (N_26658,N_26408,N_26549);
xnor U26659 (N_26659,N_26525,N_26445);
xnor U26660 (N_26660,N_26481,N_26565);
nor U26661 (N_26661,N_26587,N_26488);
xor U26662 (N_26662,N_26432,N_26513);
xor U26663 (N_26663,N_26416,N_26422);
xnor U26664 (N_26664,N_26554,N_26495);
nor U26665 (N_26665,N_26509,N_26455);
or U26666 (N_26666,N_26514,N_26461);
nand U26667 (N_26667,N_26551,N_26448);
xor U26668 (N_26668,N_26462,N_26568);
nor U26669 (N_26669,N_26478,N_26575);
nor U26670 (N_26670,N_26480,N_26501);
nor U26671 (N_26671,N_26494,N_26421);
and U26672 (N_26672,N_26456,N_26441);
and U26673 (N_26673,N_26440,N_26471);
nand U26674 (N_26674,N_26529,N_26404);
nand U26675 (N_26675,N_26596,N_26427);
xnor U26676 (N_26676,N_26528,N_26475);
nand U26677 (N_26677,N_26574,N_26585);
xnor U26678 (N_26678,N_26493,N_26566);
or U26679 (N_26679,N_26594,N_26510);
and U26680 (N_26680,N_26491,N_26443);
xor U26681 (N_26681,N_26434,N_26484);
or U26682 (N_26682,N_26589,N_26592);
or U26683 (N_26683,N_26496,N_26544);
nor U26684 (N_26684,N_26428,N_26426);
xor U26685 (N_26685,N_26520,N_26489);
or U26686 (N_26686,N_26485,N_26593);
and U26687 (N_26687,N_26482,N_26570);
and U26688 (N_26688,N_26498,N_26430);
or U26689 (N_26689,N_26573,N_26451);
xnor U26690 (N_26690,N_26465,N_26401);
and U26691 (N_26691,N_26579,N_26468);
nand U26692 (N_26692,N_26541,N_26515);
and U26693 (N_26693,N_26419,N_26413);
and U26694 (N_26694,N_26590,N_26562);
nor U26695 (N_26695,N_26487,N_26550);
nor U26696 (N_26696,N_26447,N_26406);
xor U26697 (N_26697,N_26500,N_26452);
nand U26698 (N_26698,N_26459,N_26469);
nor U26699 (N_26699,N_26483,N_26463);
nor U26700 (N_26700,N_26592,N_26597);
xnor U26701 (N_26701,N_26441,N_26561);
or U26702 (N_26702,N_26453,N_26405);
or U26703 (N_26703,N_26518,N_26544);
nor U26704 (N_26704,N_26575,N_26494);
and U26705 (N_26705,N_26508,N_26439);
or U26706 (N_26706,N_26556,N_26550);
nand U26707 (N_26707,N_26526,N_26555);
xor U26708 (N_26708,N_26439,N_26529);
or U26709 (N_26709,N_26429,N_26589);
and U26710 (N_26710,N_26588,N_26426);
nor U26711 (N_26711,N_26529,N_26599);
or U26712 (N_26712,N_26499,N_26524);
and U26713 (N_26713,N_26562,N_26540);
nand U26714 (N_26714,N_26548,N_26424);
nor U26715 (N_26715,N_26572,N_26467);
or U26716 (N_26716,N_26539,N_26537);
xor U26717 (N_26717,N_26554,N_26453);
nor U26718 (N_26718,N_26441,N_26471);
xor U26719 (N_26719,N_26519,N_26522);
or U26720 (N_26720,N_26482,N_26589);
and U26721 (N_26721,N_26481,N_26486);
nand U26722 (N_26722,N_26442,N_26422);
or U26723 (N_26723,N_26591,N_26519);
nor U26724 (N_26724,N_26483,N_26512);
and U26725 (N_26725,N_26591,N_26502);
nand U26726 (N_26726,N_26424,N_26595);
and U26727 (N_26727,N_26449,N_26550);
nand U26728 (N_26728,N_26519,N_26492);
or U26729 (N_26729,N_26549,N_26422);
nand U26730 (N_26730,N_26461,N_26433);
nor U26731 (N_26731,N_26598,N_26568);
nor U26732 (N_26732,N_26578,N_26406);
nand U26733 (N_26733,N_26557,N_26438);
nor U26734 (N_26734,N_26572,N_26457);
nor U26735 (N_26735,N_26466,N_26522);
nand U26736 (N_26736,N_26492,N_26506);
nand U26737 (N_26737,N_26485,N_26595);
nand U26738 (N_26738,N_26537,N_26407);
xor U26739 (N_26739,N_26548,N_26428);
nor U26740 (N_26740,N_26416,N_26576);
nand U26741 (N_26741,N_26502,N_26490);
and U26742 (N_26742,N_26508,N_26411);
xnor U26743 (N_26743,N_26525,N_26419);
xor U26744 (N_26744,N_26461,N_26572);
xnor U26745 (N_26745,N_26495,N_26417);
or U26746 (N_26746,N_26491,N_26532);
xor U26747 (N_26747,N_26524,N_26531);
nand U26748 (N_26748,N_26545,N_26418);
nor U26749 (N_26749,N_26578,N_26425);
or U26750 (N_26750,N_26515,N_26463);
or U26751 (N_26751,N_26551,N_26565);
nand U26752 (N_26752,N_26531,N_26460);
or U26753 (N_26753,N_26541,N_26559);
xor U26754 (N_26754,N_26476,N_26566);
nor U26755 (N_26755,N_26474,N_26403);
nor U26756 (N_26756,N_26542,N_26500);
or U26757 (N_26757,N_26461,N_26415);
and U26758 (N_26758,N_26593,N_26580);
xnor U26759 (N_26759,N_26572,N_26488);
nor U26760 (N_26760,N_26508,N_26529);
nor U26761 (N_26761,N_26590,N_26469);
nor U26762 (N_26762,N_26509,N_26595);
xor U26763 (N_26763,N_26473,N_26402);
and U26764 (N_26764,N_26430,N_26548);
or U26765 (N_26765,N_26423,N_26429);
and U26766 (N_26766,N_26461,N_26540);
nand U26767 (N_26767,N_26488,N_26556);
and U26768 (N_26768,N_26489,N_26417);
or U26769 (N_26769,N_26440,N_26573);
and U26770 (N_26770,N_26401,N_26565);
nor U26771 (N_26771,N_26469,N_26451);
nand U26772 (N_26772,N_26419,N_26454);
nor U26773 (N_26773,N_26529,N_26580);
nor U26774 (N_26774,N_26441,N_26403);
and U26775 (N_26775,N_26426,N_26422);
nor U26776 (N_26776,N_26581,N_26548);
or U26777 (N_26777,N_26505,N_26525);
xnor U26778 (N_26778,N_26443,N_26542);
nand U26779 (N_26779,N_26463,N_26573);
xor U26780 (N_26780,N_26589,N_26583);
xor U26781 (N_26781,N_26516,N_26529);
or U26782 (N_26782,N_26444,N_26400);
and U26783 (N_26783,N_26410,N_26485);
xor U26784 (N_26784,N_26459,N_26436);
xnor U26785 (N_26785,N_26409,N_26487);
xor U26786 (N_26786,N_26508,N_26559);
nor U26787 (N_26787,N_26435,N_26404);
nor U26788 (N_26788,N_26493,N_26507);
xnor U26789 (N_26789,N_26485,N_26421);
and U26790 (N_26790,N_26470,N_26456);
nor U26791 (N_26791,N_26447,N_26439);
xnor U26792 (N_26792,N_26578,N_26552);
or U26793 (N_26793,N_26452,N_26476);
nand U26794 (N_26794,N_26489,N_26453);
nand U26795 (N_26795,N_26484,N_26511);
or U26796 (N_26796,N_26527,N_26538);
xnor U26797 (N_26797,N_26545,N_26483);
nand U26798 (N_26798,N_26453,N_26437);
nor U26799 (N_26799,N_26587,N_26589);
nand U26800 (N_26800,N_26615,N_26799);
and U26801 (N_26801,N_26654,N_26675);
or U26802 (N_26802,N_26606,N_26769);
xor U26803 (N_26803,N_26762,N_26611);
and U26804 (N_26804,N_26635,N_26692);
and U26805 (N_26805,N_26610,N_26684);
xor U26806 (N_26806,N_26625,N_26763);
nand U26807 (N_26807,N_26639,N_26704);
nor U26808 (N_26808,N_26748,N_26766);
nor U26809 (N_26809,N_26712,N_26780);
xor U26810 (N_26810,N_26656,N_26691);
xor U26811 (N_26811,N_26680,N_26666);
nand U26812 (N_26812,N_26727,N_26785);
nor U26813 (N_26813,N_26758,N_26767);
or U26814 (N_26814,N_26796,N_26641);
and U26815 (N_26815,N_26753,N_26792);
and U26816 (N_26816,N_26690,N_26781);
nor U26817 (N_26817,N_26761,N_26744);
nor U26818 (N_26818,N_26798,N_26613);
and U26819 (N_26819,N_26677,N_26775);
and U26820 (N_26820,N_26765,N_26633);
nor U26821 (N_26821,N_26681,N_26661);
or U26822 (N_26822,N_26617,N_26784);
or U26823 (N_26823,N_26730,N_26673);
nor U26824 (N_26824,N_26795,N_26788);
nor U26825 (N_26825,N_26721,N_26787);
xor U26826 (N_26826,N_26772,N_26738);
and U26827 (N_26827,N_26618,N_26671);
or U26828 (N_26828,N_26773,N_26733);
nand U26829 (N_26829,N_26755,N_26621);
xnor U26830 (N_26830,N_26698,N_26764);
nand U26831 (N_26831,N_26628,N_26734);
xor U26832 (N_26832,N_26664,N_26634);
nor U26833 (N_26833,N_26644,N_26689);
nor U26834 (N_26834,N_26728,N_26693);
or U26835 (N_26835,N_26720,N_26695);
or U26836 (N_26836,N_26778,N_26756);
nor U26837 (N_26837,N_26601,N_26687);
and U26838 (N_26838,N_26776,N_26623);
nor U26839 (N_26839,N_26736,N_26669);
and U26840 (N_26840,N_26667,N_26746);
or U26841 (N_26841,N_26682,N_26713);
xor U26842 (N_26842,N_26794,N_26790);
nor U26843 (N_26843,N_26760,N_26739);
and U26844 (N_26844,N_26652,N_26616);
and U26845 (N_26845,N_26686,N_26632);
nand U26846 (N_26846,N_26797,N_26724);
nand U26847 (N_26847,N_26685,N_26731);
nand U26848 (N_26848,N_26650,N_26705);
or U26849 (N_26849,N_26636,N_26709);
or U26850 (N_26850,N_26782,N_26768);
and U26851 (N_26851,N_26646,N_26607);
or U26852 (N_26852,N_26626,N_26688);
xnor U26853 (N_26853,N_26743,N_26662);
xor U26854 (N_26854,N_26609,N_26624);
nand U26855 (N_26855,N_26751,N_26694);
or U26856 (N_26856,N_26678,N_26676);
nand U26857 (N_26857,N_26683,N_26608);
and U26858 (N_26858,N_26726,N_26770);
or U26859 (N_26859,N_26714,N_26679);
nand U26860 (N_26860,N_26722,N_26707);
and U26861 (N_26861,N_26672,N_26702);
nand U26862 (N_26862,N_26620,N_26789);
or U26863 (N_26863,N_26774,N_26779);
nor U26864 (N_26864,N_26631,N_26604);
and U26865 (N_26865,N_26710,N_26791);
nand U26866 (N_26866,N_26700,N_26729);
and U26867 (N_26867,N_26600,N_26670);
nor U26868 (N_26868,N_26655,N_26706);
nor U26869 (N_26869,N_26629,N_26786);
xor U26870 (N_26870,N_26660,N_26605);
or U26871 (N_26871,N_26750,N_26752);
and U26872 (N_26872,N_26640,N_26732);
or U26873 (N_26873,N_26674,N_26708);
nand U26874 (N_26874,N_26668,N_26659);
or U26875 (N_26875,N_26663,N_26719);
and U26876 (N_26876,N_26737,N_26699);
and U26877 (N_26877,N_26645,N_26749);
or U26878 (N_26878,N_26715,N_26703);
or U26879 (N_26879,N_26658,N_26793);
xnor U26880 (N_26880,N_26651,N_26657);
nor U26881 (N_26881,N_26711,N_26602);
xnor U26882 (N_26882,N_26742,N_26638);
nand U26883 (N_26883,N_26637,N_26647);
and U26884 (N_26884,N_26701,N_26757);
or U26885 (N_26885,N_26783,N_26740);
nor U26886 (N_26886,N_26653,N_26745);
or U26887 (N_26887,N_26665,N_26747);
and U26888 (N_26888,N_26627,N_26643);
or U26889 (N_26889,N_26697,N_26642);
or U26890 (N_26890,N_26696,N_26735);
and U26891 (N_26891,N_26619,N_26716);
nor U26892 (N_26892,N_26648,N_26718);
and U26893 (N_26893,N_26622,N_26754);
xnor U26894 (N_26894,N_26630,N_26725);
xnor U26895 (N_26895,N_26612,N_26717);
xnor U26896 (N_26896,N_26759,N_26777);
xor U26897 (N_26897,N_26741,N_26723);
or U26898 (N_26898,N_26603,N_26649);
nor U26899 (N_26899,N_26614,N_26771);
and U26900 (N_26900,N_26748,N_26772);
xor U26901 (N_26901,N_26753,N_26693);
nor U26902 (N_26902,N_26680,N_26708);
nor U26903 (N_26903,N_26776,N_26789);
nand U26904 (N_26904,N_26706,N_26766);
nor U26905 (N_26905,N_26747,N_26794);
nand U26906 (N_26906,N_26740,N_26743);
nor U26907 (N_26907,N_26736,N_26617);
nand U26908 (N_26908,N_26614,N_26716);
or U26909 (N_26909,N_26670,N_26718);
nand U26910 (N_26910,N_26772,N_26737);
nor U26911 (N_26911,N_26638,N_26741);
nand U26912 (N_26912,N_26693,N_26716);
nand U26913 (N_26913,N_26614,N_26786);
or U26914 (N_26914,N_26746,N_26771);
and U26915 (N_26915,N_26681,N_26644);
xnor U26916 (N_26916,N_26682,N_26794);
and U26917 (N_26917,N_26797,N_26652);
or U26918 (N_26918,N_26657,N_26762);
or U26919 (N_26919,N_26608,N_26708);
nand U26920 (N_26920,N_26757,N_26666);
xnor U26921 (N_26921,N_26674,N_26618);
nand U26922 (N_26922,N_26635,N_26697);
or U26923 (N_26923,N_26710,N_26746);
nand U26924 (N_26924,N_26714,N_26707);
xnor U26925 (N_26925,N_26737,N_26749);
and U26926 (N_26926,N_26620,N_26786);
and U26927 (N_26927,N_26759,N_26771);
nor U26928 (N_26928,N_26706,N_26763);
nor U26929 (N_26929,N_26782,N_26648);
xnor U26930 (N_26930,N_26607,N_26790);
or U26931 (N_26931,N_26765,N_26735);
nand U26932 (N_26932,N_26690,N_26656);
xnor U26933 (N_26933,N_26775,N_26616);
or U26934 (N_26934,N_26763,N_26675);
or U26935 (N_26935,N_26693,N_26600);
nor U26936 (N_26936,N_26672,N_26684);
xor U26937 (N_26937,N_26792,N_26790);
or U26938 (N_26938,N_26715,N_26651);
or U26939 (N_26939,N_26760,N_26729);
or U26940 (N_26940,N_26723,N_26750);
and U26941 (N_26941,N_26757,N_26650);
nand U26942 (N_26942,N_26721,N_26740);
nor U26943 (N_26943,N_26722,N_26669);
nand U26944 (N_26944,N_26663,N_26678);
or U26945 (N_26945,N_26621,N_26667);
and U26946 (N_26946,N_26601,N_26699);
xor U26947 (N_26947,N_26631,N_26747);
or U26948 (N_26948,N_26751,N_26774);
xor U26949 (N_26949,N_26730,N_26684);
nor U26950 (N_26950,N_26775,N_26780);
nand U26951 (N_26951,N_26779,N_26621);
and U26952 (N_26952,N_26757,N_26649);
and U26953 (N_26953,N_26600,N_26749);
nor U26954 (N_26954,N_26703,N_26725);
xnor U26955 (N_26955,N_26637,N_26741);
xnor U26956 (N_26956,N_26740,N_26724);
and U26957 (N_26957,N_26700,N_26756);
and U26958 (N_26958,N_26664,N_26656);
or U26959 (N_26959,N_26670,N_26710);
nor U26960 (N_26960,N_26605,N_26628);
xor U26961 (N_26961,N_26640,N_26744);
xor U26962 (N_26962,N_26641,N_26700);
and U26963 (N_26963,N_26640,N_26634);
or U26964 (N_26964,N_26734,N_26736);
xnor U26965 (N_26965,N_26668,N_26794);
and U26966 (N_26966,N_26701,N_26716);
nor U26967 (N_26967,N_26732,N_26743);
xor U26968 (N_26968,N_26617,N_26793);
and U26969 (N_26969,N_26727,N_26746);
xor U26970 (N_26970,N_26667,N_26799);
and U26971 (N_26971,N_26797,N_26662);
or U26972 (N_26972,N_26790,N_26780);
and U26973 (N_26973,N_26789,N_26613);
or U26974 (N_26974,N_26670,N_26675);
nand U26975 (N_26975,N_26740,N_26681);
xor U26976 (N_26976,N_26656,N_26759);
nand U26977 (N_26977,N_26775,N_26744);
xnor U26978 (N_26978,N_26648,N_26756);
nand U26979 (N_26979,N_26721,N_26760);
xnor U26980 (N_26980,N_26644,N_26622);
nand U26981 (N_26981,N_26654,N_26788);
and U26982 (N_26982,N_26658,N_26774);
nor U26983 (N_26983,N_26647,N_26617);
xor U26984 (N_26984,N_26616,N_26624);
nor U26985 (N_26985,N_26701,N_26752);
nor U26986 (N_26986,N_26701,N_26736);
nand U26987 (N_26987,N_26752,N_26782);
and U26988 (N_26988,N_26634,N_26711);
nor U26989 (N_26989,N_26734,N_26710);
and U26990 (N_26990,N_26605,N_26629);
nand U26991 (N_26991,N_26610,N_26737);
nor U26992 (N_26992,N_26740,N_26629);
or U26993 (N_26993,N_26633,N_26764);
or U26994 (N_26994,N_26637,N_26791);
or U26995 (N_26995,N_26600,N_26770);
xnor U26996 (N_26996,N_26716,N_26658);
nor U26997 (N_26997,N_26797,N_26639);
nor U26998 (N_26998,N_26712,N_26725);
and U26999 (N_26999,N_26767,N_26760);
and U27000 (N_27000,N_26820,N_26854);
or U27001 (N_27001,N_26981,N_26895);
and U27002 (N_27002,N_26857,N_26961);
nor U27003 (N_27003,N_26993,N_26996);
nand U27004 (N_27004,N_26874,N_26827);
or U27005 (N_27005,N_26889,N_26964);
or U27006 (N_27006,N_26836,N_26811);
and U27007 (N_27007,N_26896,N_26858);
and U27008 (N_27008,N_26882,N_26939);
nand U27009 (N_27009,N_26872,N_26891);
nor U27010 (N_27010,N_26990,N_26830);
or U27011 (N_27011,N_26831,N_26944);
or U27012 (N_27012,N_26845,N_26800);
nor U27013 (N_27013,N_26812,N_26869);
xor U27014 (N_27014,N_26992,N_26978);
or U27015 (N_27015,N_26974,N_26899);
or U27016 (N_27016,N_26938,N_26833);
xor U27017 (N_27017,N_26849,N_26824);
or U27018 (N_27018,N_26839,N_26890);
nand U27019 (N_27019,N_26953,N_26893);
nand U27020 (N_27020,N_26852,N_26848);
nand U27021 (N_27021,N_26828,N_26955);
or U27022 (N_27022,N_26968,N_26966);
or U27023 (N_27023,N_26832,N_26884);
xor U27024 (N_27024,N_26888,N_26919);
and U27025 (N_27025,N_26900,N_26958);
nor U27026 (N_27026,N_26924,N_26904);
or U27027 (N_27027,N_26875,N_26954);
xnor U27028 (N_27028,N_26868,N_26998);
nand U27029 (N_27029,N_26829,N_26844);
or U27030 (N_27030,N_26945,N_26862);
and U27031 (N_27031,N_26816,N_26851);
and U27032 (N_27032,N_26999,N_26801);
nor U27033 (N_27033,N_26806,N_26894);
nor U27034 (N_27034,N_26907,N_26947);
and U27035 (N_27035,N_26949,N_26963);
nor U27036 (N_27036,N_26918,N_26980);
xor U27037 (N_27037,N_26805,N_26972);
or U27038 (N_27038,N_26864,N_26835);
xnor U27039 (N_27039,N_26903,N_26809);
nand U27040 (N_27040,N_26914,N_26948);
nor U27041 (N_27041,N_26901,N_26883);
and U27042 (N_27042,N_26892,N_26970);
and U27043 (N_27043,N_26840,N_26923);
and U27044 (N_27044,N_26834,N_26908);
and U27045 (N_27045,N_26881,N_26979);
or U27046 (N_27046,N_26937,N_26917);
nor U27047 (N_27047,N_26973,N_26988);
nand U27048 (N_27048,N_26926,N_26930);
or U27049 (N_27049,N_26865,N_26913);
xnor U27050 (N_27050,N_26847,N_26879);
or U27051 (N_27051,N_26905,N_26826);
nor U27052 (N_27052,N_26962,N_26977);
nand U27053 (N_27053,N_26986,N_26985);
nand U27054 (N_27054,N_26956,N_26860);
xor U27055 (N_27055,N_26936,N_26843);
xor U27056 (N_27056,N_26817,N_26871);
nand U27057 (N_27057,N_26821,N_26969);
nor U27058 (N_27058,N_26942,N_26957);
nand U27059 (N_27059,N_26912,N_26976);
and U27060 (N_27060,N_26850,N_26971);
xor U27061 (N_27061,N_26982,N_26935);
or U27062 (N_27062,N_26995,N_26898);
xnor U27063 (N_27063,N_26994,N_26989);
xnor U27064 (N_27064,N_26846,N_26873);
nor U27065 (N_27065,N_26943,N_26842);
nor U27066 (N_27066,N_26837,N_26886);
and U27067 (N_27067,N_26838,N_26960);
and U27068 (N_27068,N_26921,N_26802);
nand U27069 (N_27069,N_26859,N_26822);
nand U27070 (N_27070,N_26853,N_26819);
nor U27071 (N_27071,N_26877,N_26876);
nand U27072 (N_27072,N_26929,N_26878);
nor U27073 (N_27073,N_26967,N_26940);
xnor U27074 (N_27074,N_26915,N_26810);
and U27075 (N_27075,N_26856,N_26870);
and U27076 (N_27076,N_26928,N_26931);
or U27077 (N_27077,N_26902,N_26861);
and U27078 (N_27078,N_26946,N_26991);
xor U27079 (N_27079,N_26867,N_26823);
nand U27080 (N_27080,N_26803,N_26959);
and U27081 (N_27081,N_26841,N_26927);
and U27082 (N_27082,N_26950,N_26932);
or U27083 (N_27083,N_26813,N_26952);
or U27084 (N_27084,N_26825,N_26909);
and U27085 (N_27085,N_26983,N_26965);
and U27086 (N_27086,N_26987,N_26897);
nand U27087 (N_27087,N_26911,N_26951);
xnor U27088 (N_27088,N_26887,N_26934);
and U27089 (N_27089,N_26975,N_26815);
nand U27090 (N_27090,N_26941,N_26925);
or U27091 (N_27091,N_26880,N_26920);
xor U27092 (N_27092,N_26814,N_26855);
and U27093 (N_27093,N_26863,N_26922);
nor U27094 (N_27094,N_26997,N_26910);
or U27095 (N_27095,N_26916,N_26804);
or U27096 (N_27096,N_26818,N_26807);
nand U27097 (N_27097,N_26906,N_26866);
xor U27098 (N_27098,N_26885,N_26933);
nand U27099 (N_27099,N_26808,N_26984);
nor U27100 (N_27100,N_26970,N_26837);
xor U27101 (N_27101,N_26997,N_26883);
or U27102 (N_27102,N_26844,N_26835);
and U27103 (N_27103,N_26876,N_26810);
xnor U27104 (N_27104,N_26953,N_26867);
nand U27105 (N_27105,N_26831,N_26907);
nand U27106 (N_27106,N_26873,N_26927);
nor U27107 (N_27107,N_26806,N_26929);
nor U27108 (N_27108,N_26947,N_26972);
nor U27109 (N_27109,N_26883,N_26985);
xnor U27110 (N_27110,N_26880,N_26835);
or U27111 (N_27111,N_26845,N_26815);
nor U27112 (N_27112,N_26928,N_26980);
or U27113 (N_27113,N_26989,N_26858);
nor U27114 (N_27114,N_26935,N_26863);
or U27115 (N_27115,N_26921,N_26880);
nand U27116 (N_27116,N_26878,N_26837);
xnor U27117 (N_27117,N_26971,N_26987);
nand U27118 (N_27118,N_26982,N_26953);
and U27119 (N_27119,N_26978,N_26820);
nor U27120 (N_27120,N_26951,N_26812);
and U27121 (N_27121,N_26880,N_26970);
or U27122 (N_27122,N_26964,N_26894);
xnor U27123 (N_27123,N_26970,N_26985);
nor U27124 (N_27124,N_26979,N_26874);
nor U27125 (N_27125,N_26876,N_26893);
xnor U27126 (N_27126,N_26904,N_26940);
or U27127 (N_27127,N_26953,N_26989);
nand U27128 (N_27128,N_26987,N_26830);
xnor U27129 (N_27129,N_26876,N_26872);
or U27130 (N_27130,N_26946,N_26949);
xor U27131 (N_27131,N_26844,N_26823);
nor U27132 (N_27132,N_26814,N_26942);
and U27133 (N_27133,N_26855,N_26947);
or U27134 (N_27134,N_26902,N_26899);
xor U27135 (N_27135,N_26903,N_26801);
and U27136 (N_27136,N_26889,N_26852);
nor U27137 (N_27137,N_26819,N_26966);
nor U27138 (N_27138,N_26844,N_26898);
and U27139 (N_27139,N_26896,N_26848);
and U27140 (N_27140,N_26937,N_26812);
and U27141 (N_27141,N_26943,N_26927);
xor U27142 (N_27142,N_26960,N_26948);
nand U27143 (N_27143,N_26861,N_26986);
nand U27144 (N_27144,N_26979,N_26946);
or U27145 (N_27145,N_26924,N_26844);
xnor U27146 (N_27146,N_26891,N_26895);
nand U27147 (N_27147,N_26857,N_26898);
nor U27148 (N_27148,N_26916,N_26833);
or U27149 (N_27149,N_26964,N_26838);
xnor U27150 (N_27150,N_26988,N_26819);
and U27151 (N_27151,N_26999,N_26851);
nand U27152 (N_27152,N_26992,N_26982);
and U27153 (N_27153,N_26983,N_26905);
nand U27154 (N_27154,N_26953,N_26814);
and U27155 (N_27155,N_26900,N_26816);
and U27156 (N_27156,N_26824,N_26809);
or U27157 (N_27157,N_26877,N_26976);
and U27158 (N_27158,N_26826,N_26943);
and U27159 (N_27159,N_26985,N_26967);
nand U27160 (N_27160,N_26808,N_26974);
or U27161 (N_27161,N_26891,N_26940);
or U27162 (N_27162,N_26866,N_26969);
nor U27163 (N_27163,N_26921,N_26996);
nand U27164 (N_27164,N_26867,N_26815);
xor U27165 (N_27165,N_26837,N_26861);
or U27166 (N_27166,N_26939,N_26827);
and U27167 (N_27167,N_26916,N_26948);
nand U27168 (N_27168,N_26803,N_26833);
and U27169 (N_27169,N_26955,N_26981);
or U27170 (N_27170,N_26887,N_26918);
and U27171 (N_27171,N_26811,N_26904);
and U27172 (N_27172,N_26952,N_26964);
and U27173 (N_27173,N_26915,N_26835);
or U27174 (N_27174,N_26863,N_26908);
nor U27175 (N_27175,N_26985,N_26963);
xnor U27176 (N_27176,N_26906,N_26828);
xor U27177 (N_27177,N_26843,N_26812);
and U27178 (N_27178,N_26907,N_26825);
nand U27179 (N_27179,N_26826,N_26819);
or U27180 (N_27180,N_26956,N_26847);
xor U27181 (N_27181,N_26977,N_26975);
or U27182 (N_27182,N_26885,N_26982);
nor U27183 (N_27183,N_26809,N_26946);
and U27184 (N_27184,N_26926,N_26855);
nand U27185 (N_27185,N_26817,N_26828);
xnor U27186 (N_27186,N_26940,N_26966);
or U27187 (N_27187,N_26811,N_26848);
xnor U27188 (N_27188,N_26996,N_26899);
nor U27189 (N_27189,N_26904,N_26886);
or U27190 (N_27190,N_26847,N_26936);
nor U27191 (N_27191,N_26953,N_26956);
nand U27192 (N_27192,N_26884,N_26952);
or U27193 (N_27193,N_26801,N_26812);
and U27194 (N_27194,N_26905,N_26932);
or U27195 (N_27195,N_26854,N_26909);
and U27196 (N_27196,N_26898,N_26975);
or U27197 (N_27197,N_26949,N_26973);
nor U27198 (N_27198,N_26800,N_26984);
nor U27199 (N_27199,N_26848,N_26952);
xnor U27200 (N_27200,N_27105,N_27190);
and U27201 (N_27201,N_27171,N_27043);
or U27202 (N_27202,N_27081,N_27066);
and U27203 (N_27203,N_27017,N_27189);
or U27204 (N_27204,N_27070,N_27113);
nor U27205 (N_27205,N_27160,N_27022);
or U27206 (N_27206,N_27136,N_27085);
or U27207 (N_27207,N_27013,N_27187);
and U27208 (N_27208,N_27041,N_27087);
or U27209 (N_27209,N_27166,N_27122);
xor U27210 (N_27210,N_27064,N_27094);
nand U27211 (N_27211,N_27121,N_27026);
and U27212 (N_27212,N_27052,N_27021);
xor U27213 (N_27213,N_27132,N_27069);
and U27214 (N_27214,N_27089,N_27147);
nor U27215 (N_27215,N_27126,N_27019);
nand U27216 (N_27216,N_27175,N_27120);
nor U27217 (N_27217,N_27169,N_27141);
nor U27218 (N_27218,N_27037,N_27006);
or U27219 (N_27219,N_27130,N_27191);
and U27220 (N_27220,N_27199,N_27174);
nand U27221 (N_27221,N_27049,N_27086);
or U27222 (N_27222,N_27040,N_27134);
or U27223 (N_27223,N_27117,N_27046);
or U27224 (N_27224,N_27153,N_27124);
nand U27225 (N_27225,N_27036,N_27010);
and U27226 (N_27226,N_27050,N_27196);
nand U27227 (N_27227,N_27033,N_27186);
or U27228 (N_27228,N_27084,N_27009);
nor U27229 (N_27229,N_27073,N_27032);
or U27230 (N_27230,N_27107,N_27020);
nand U27231 (N_27231,N_27044,N_27163);
nand U27232 (N_27232,N_27156,N_27159);
or U27233 (N_27233,N_27148,N_27127);
or U27234 (N_27234,N_27014,N_27146);
nor U27235 (N_27235,N_27027,N_27045);
and U27236 (N_27236,N_27076,N_27091);
nor U27237 (N_27237,N_27170,N_27092);
and U27238 (N_27238,N_27179,N_27158);
or U27239 (N_27239,N_27011,N_27038);
nand U27240 (N_27240,N_27077,N_27133);
or U27241 (N_27241,N_27003,N_27035);
or U27242 (N_27242,N_27135,N_27001);
and U27243 (N_27243,N_27071,N_27031);
nand U27244 (N_27244,N_27154,N_27048);
xnor U27245 (N_27245,N_27181,N_27079);
nor U27246 (N_27246,N_27051,N_27164);
xnor U27247 (N_27247,N_27062,N_27194);
xnor U27248 (N_27248,N_27161,N_27099);
nor U27249 (N_27249,N_27007,N_27144);
and U27250 (N_27250,N_27123,N_27162);
or U27251 (N_27251,N_27053,N_27184);
xnor U27252 (N_27252,N_27042,N_27197);
nor U27253 (N_27253,N_27063,N_27104);
and U27254 (N_27254,N_27178,N_27072);
nor U27255 (N_27255,N_27112,N_27074);
nand U27256 (N_27256,N_27145,N_27155);
nand U27257 (N_27257,N_27028,N_27188);
or U27258 (N_27258,N_27097,N_27056);
nor U27259 (N_27259,N_27143,N_27109);
or U27260 (N_27260,N_27125,N_27150);
or U27261 (N_27261,N_27030,N_27012);
or U27262 (N_27262,N_27088,N_27152);
or U27263 (N_27263,N_27068,N_27131);
nor U27264 (N_27264,N_27103,N_27114);
xnor U27265 (N_27265,N_27142,N_27098);
nand U27266 (N_27266,N_27065,N_27168);
nor U27267 (N_27267,N_27128,N_27096);
or U27268 (N_27268,N_27139,N_27039);
or U27269 (N_27269,N_27080,N_27111);
nor U27270 (N_27270,N_27185,N_27167);
nor U27271 (N_27271,N_27024,N_27034);
xnor U27272 (N_27272,N_27182,N_27172);
and U27273 (N_27273,N_27100,N_27023);
nand U27274 (N_27274,N_27008,N_27078);
nand U27275 (N_27275,N_27059,N_27093);
and U27276 (N_27276,N_27005,N_27176);
nand U27277 (N_27277,N_27180,N_27018);
or U27278 (N_27278,N_27151,N_27106);
and U27279 (N_27279,N_27137,N_27192);
xnor U27280 (N_27280,N_27057,N_27075);
nand U27281 (N_27281,N_27198,N_27067);
xnor U27282 (N_27282,N_27102,N_27054);
or U27283 (N_27283,N_27082,N_27101);
or U27284 (N_27284,N_27025,N_27119);
xnor U27285 (N_27285,N_27110,N_27061);
and U27286 (N_27286,N_27193,N_27004);
nand U27287 (N_27287,N_27195,N_27016);
or U27288 (N_27288,N_27047,N_27118);
or U27289 (N_27289,N_27000,N_27173);
xor U27290 (N_27290,N_27090,N_27095);
nand U27291 (N_27291,N_27140,N_27083);
or U27292 (N_27292,N_27177,N_27157);
nor U27293 (N_27293,N_27165,N_27029);
nand U27294 (N_27294,N_27058,N_27116);
or U27295 (N_27295,N_27002,N_27183);
and U27296 (N_27296,N_27055,N_27015);
xnor U27297 (N_27297,N_27060,N_27108);
or U27298 (N_27298,N_27115,N_27138);
or U27299 (N_27299,N_27129,N_27149);
xnor U27300 (N_27300,N_27082,N_27159);
and U27301 (N_27301,N_27080,N_27161);
xor U27302 (N_27302,N_27045,N_27037);
and U27303 (N_27303,N_27161,N_27179);
nor U27304 (N_27304,N_27081,N_27183);
xnor U27305 (N_27305,N_27090,N_27058);
xor U27306 (N_27306,N_27055,N_27103);
and U27307 (N_27307,N_27040,N_27096);
xor U27308 (N_27308,N_27186,N_27018);
nand U27309 (N_27309,N_27050,N_27049);
or U27310 (N_27310,N_27061,N_27001);
nor U27311 (N_27311,N_27192,N_27092);
and U27312 (N_27312,N_27053,N_27103);
nand U27313 (N_27313,N_27001,N_27199);
nand U27314 (N_27314,N_27009,N_27087);
nand U27315 (N_27315,N_27147,N_27063);
xor U27316 (N_27316,N_27153,N_27005);
nor U27317 (N_27317,N_27050,N_27038);
nor U27318 (N_27318,N_27157,N_27054);
or U27319 (N_27319,N_27119,N_27030);
nor U27320 (N_27320,N_27068,N_27090);
and U27321 (N_27321,N_27140,N_27147);
and U27322 (N_27322,N_27003,N_27010);
nor U27323 (N_27323,N_27003,N_27114);
and U27324 (N_27324,N_27198,N_27147);
xor U27325 (N_27325,N_27107,N_27110);
xor U27326 (N_27326,N_27085,N_27082);
and U27327 (N_27327,N_27139,N_27055);
and U27328 (N_27328,N_27076,N_27065);
or U27329 (N_27329,N_27104,N_27133);
nor U27330 (N_27330,N_27045,N_27024);
and U27331 (N_27331,N_27175,N_27188);
and U27332 (N_27332,N_27162,N_27036);
or U27333 (N_27333,N_27070,N_27025);
and U27334 (N_27334,N_27048,N_27070);
nor U27335 (N_27335,N_27028,N_27081);
and U27336 (N_27336,N_27152,N_27177);
nand U27337 (N_27337,N_27016,N_27005);
or U27338 (N_27338,N_27010,N_27163);
nor U27339 (N_27339,N_27065,N_27156);
nor U27340 (N_27340,N_27018,N_27083);
nand U27341 (N_27341,N_27197,N_27151);
xnor U27342 (N_27342,N_27181,N_27178);
or U27343 (N_27343,N_27149,N_27104);
nand U27344 (N_27344,N_27051,N_27109);
nor U27345 (N_27345,N_27068,N_27159);
nor U27346 (N_27346,N_27124,N_27008);
nand U27347 (N_27347,N_27111,N_27015);
or U27348 (N_27348,N_27078,N_27053);
nand U27349 (N_27349,N_27138,N_27108);
and U27350 (N_27350,N_27012,N_27176);
and U27351 (N_27351,N_27018,N_27151);
nand U27352 (N_27352,N_27156,N_27178);
or U27353 (N_27353,N_27161,N_27081);
and U27354 (N_27354,N_27147,N_27072);
nand U27355 (N_27355,N_27069,N_27023);
and U27356 (N_27356,N_27079,N_27029);
or U27357 (N_27357,N_27062,N_27005);
xor U27358 (N_27358,N_27023,N_27077);
nand U27359 (N_27359,N_27041,N_27117);
xor U27360 (N_27360,N_27153,N_27171);
nand U27361 (N_27361,N_27032,N_27138);
and U27362 (N_27362,N_27193,N_27088);
or U27363 (N_27363,N_27004,N_27034);
nand U27364 (N_27364,N_27104,N_27050);
and U27365 (N_27365,N_27071,N_27023);
nor U27366 (N_27366,N_27103,N_27195);
nand U27367 (N_27367,N_27150,N_27035);
xnor U27368 (N_27368,N_27190,N_27070);
nand U27369 (N_27369,N_27194,N_27115);
nor U27370 (N_27370,N_27085,N_27010);
nor U27371 (N_27371,N_27068,N_27013);
and U27372 (N_27372,N_27135,N_27031);
and U27373 (N_27373,N_27104,N_27056);
xor U27374 (N_27374,N_27156,N_27106);
and U27375 (N_27375,N_27181,N_27179);
nand U27376 (N_27376,N_27161,N_27033);
nand U27377 (N_27377,N_27062,N_27198);
or U27378 (N_27378,N_27079,N_27171);
nand U27379 (N_27379,N_27127,N_27015);
nor U27380 (N_27380,N_27003,N_27161);
xnor U27381 (N_27381,N_27182,N_27103);
xor U27382 (N_27382,N_27059,N_27008);
nor U27383 (N_27383,N_27028,N_27132);
or U27384 (N_27384,N_27040,N_27131);
nor U27385 (N_27385,N_27130,N_27157);
and U27386 (N_27386,N_27099,N_27019);
and U27387 (N_27387,N_27068,N_27133);
nor U27388 (N_27388,N_27025,N_27082);
or U27389 (N_27389,N_27196,N_27076);
and U27390 (N_27390,N_27013,N_27098);
xor U27391 (N_27391,N_27026,N_27137);
and U27392 (N_27392,N_27141,N_27002);
nor U27393 (N_27393,N_27060,N_27096);
and U27394 (N_27394,N_27092,N_27059);
and U27395 (N_27395,N_27130,N_27071);
and U27396 (N_27396,N_27104,N_27123);
nor U27397 (N_27397,N_27042,N_27142);
nand U27398 (N_27398,N_27138,N_27079);
nand U27399 (N_27399,N_27191,N_27013);
nor U27400 (N_27400,N_27346,N_27258);
nor U27401 (N_27401,N_27380,N_27291);
or U27402 (N_27402,N_27230,N_27370);
or U27403 (N_27403,N_27302,N_27266);
nor U27404 (N_27404,N_27221,N_27259);
nand U27405 (N_27405,N_27364,N_27326);
or U27406 (N_27406,N_27375,N_27392);
or U27407 (N_27407,N_27287,N_27212);
and U27408 (N_27408,N_27286,N_27357);
nor U27409 (N_27409,N_27306,N_27332);
or U27410 (N_27410,N_27308,N_27237);
or U27411 (N_27411,N_27272,N_27398);
nor U27412 (N_27412,N_27253,N_27394);
nand U27413 (N_27413,N_27310,N_27391);
nand U27414 (N_27414,N_27340,N_27356);
xnor U27415 (N_27415,N_27211,N_27361);
nand U27416 (N_27416,N_27251,N_27264);
nand U27417 (N_27417,N_27240,N_27355);
xor U27418 (N_27418,N_27319,N_27265);
and U27419 (N_27419,N_27373,N_27307);
and U27420 (N_27420,N_27204,N_27331);
and U27421 (N_27421,N_27383,N_27389);
or U27422 (N_27422,N_27213,N_27231);
nand U27423 (N_27423,N_27284,N_27312);
xor U27424 (N_27424,N_27320,N_27246);
and U27425 (N_27425,N_27330,N_27371);
and U27426 (N_27426,N_27256,N_27268);
nor U27427 (N_27427,N_27233,N_27245);
nor U27428 (N_27428,N_27374,N_27229);
or U27429 (N_27429,N_27208,N_27317);
nand U27430 (N_27430,N_27384,N_27271);
nand U27431 (N_27431,N_27338,N_27219);
nand U27432 (N_27432,N_27366,N_27323);
or U27433 (N_27433,N_27283,N_27359);
and U27434 (N_27434,N_27292,N_27378);
nand U27435 (N_27435,N_27296,N_27209);
nor U27436 (N_27436,N_27289,N_27234);
nor U27437 (N_27437,N_27224,N_27305);
nand U27438 (N_27438,N_27393,N_27311);
nand U27439 (N_27439,N_27248,N_27262);
or U27440 (N_27440,N_27313,N_27299);
xnor U27441 (N_27441,N_27318,N_27387);
and U27442 (N_27442,N_27277,N_27236);
xor U27443 (N_27443,N_27200,N_27205);
or U27444 (N_27444,N_27328,N_27218);
xnor U27445 (N_27445,N_27395,N_27341);
nand U27446 (N_27446,N_27261,N_27396);
nor U27447 (N_27447,N_27379,N_27363);
nand U27448 (N_27448,N_27222,N_27358);
nor U27449 (N_27449,N_27390,N_27282);
or U27450 (N_27450,N_27257,N_27327);
xnor U27451 (N_27451,N_27267,N_27397);
xor U27452 (N_27452,N_27334,N_27314);
nand U27453 (N_27453,N_27281,N_27207);
nand U27454 (N_27454,N_27269,N_27254);
xnor U27455 (N_27455,N_27322,N_27369);
or U27456 (N_27456,N_27298,N_27349);
xnor U27457 (N_27457,N_27350,N_27273);
or U27458 (N_27458,N_27223,N_27270);
and U27459 (N_27459,N_27290,N_27352);
nand U27460 (N_27460,N_27335,N_27376);
nor U27461 (N_27461,N_27216,N_27227);
nor U27462 (N_27462,N_27316,N_27381);
nor U27463 (N_27463,N_27343,N_27278);
nor U27464 (N_27464,N_27324,N_27339);
or U27465 (N_27465,N_27276,N_27220);
nand U27466 (N_27466,N_27372,N_27347);
nor U27467 (N_27467,N_27241,N_27354);
nor U27468 (N_27468,N_27368,N_27280);
and U27469 (N_27469,N_27301,N_27274);
or U27470 (N_27470,N_27238,N_27351);
and U27471 (N_27471,N_27365,N_27250);
or U27472 (N_27472,N_27303,N_27247);
xor U27473 (N_27473,N_27342,N_27336);
and U27474 (N_27474,N_27226,N_27242);
and U27475 (N_27475,N_27285,N_27295);
xor U27476 (N_27476,N_27377,N_27249);
nand U27477 (N_27477,N_27386,N_27360);
nand U27478 (N_27478,N_27388,N_27367);
and U27479 (N_27479,N_27203,N_27337);
and U27480 (N_27480,N_27348,N_27293);
nand U27481 (N_27481,N_27345,N_27225);
or U27482 (N_27482,N_27252,N_27304);
nor U27483 (N_27483,N_27329,N_27325);
xnor U27484 (N_27484,N_27215,N_27244);
or U27485 (N_27485,N_27279,N_27217);
and U27486 (N_27486,N_27300,N_27232);
and U27487 (N_27487,N_27255,N_27362);
xor U27488 (N_27488,N_27206,N_27275);
nand U27489 (N_27489,N_27353,N_27294);
and U27490 (N_27490,N_27297,N_27333);
or U27491 (N_27491,N_27263,N_27288);
and U27492 (N_27492,N_27239,N_27309);
or U27493 (N_27493,N_27214,N_27235);
nor U27494 (N_27494,N_27321,N_27210);
nor U27495 (N_27495,N_27243,N_27344);
nor U27496 (N_27496,N_27399,N_27228);
nand U27497 (N_27497,N_27260,N_27385);
nor U27498 (N_27498,N_27202,N_27382);
nand U27499 (N_27499,N_27315,N_27201);
nand U27500 (N_27500,N_27394,N_27373);
nand U27501 (N_27501,N_27269,N_27209);
nor U27502 (N_27502,N_27255,N_27366);
nor U27503 (N_27503,N_27292,N_27228);
and U27504 (N_27504,N_27212,N_27291);
and U27505 (N_27505,N_27247,N_27316);
or U27506 (N_27506,N_27320,N_27283);
nand U27507 (N_27507,N_27382,N_27272);
or U27508 (N_27508,N_27368,N_27348);
nor U27509 (N_27509,N_27224,N_27228);
xor U27510 (N_27510,N_27282,N_27302);
xnor U27511 (N_27511,N_27248,N_27282);
xnor U27512 (N_27512,N_27216,N_27374);
nand U27513 (N_27513,N_27286,N_27233);
nor U27514 (N_27514,N_27349,N_27217);
or U27515 (N_27515,N_27279,N_27275);
nor U27516 (N_27516,N_27361,N_27378);
and U27517 (N_27517,N_27390,N_27298);
or U27518 (N_27518,N_27256,N_27322);
nor U27519 (N_27519,N_27276,N_27376);
and U27520 (N_27520,N_27363,N_27250);
xor U27521 (N_27521,N_27394,N_27365);
xnor U27522 (N_27522,N_27373,N_27296);
or U27523 (N_27523,N_27335,N_27398);
nor U27524 (N_27524,N_27218,N_27248);
nand U27525 (N_27525,N_27349,N_27314);
xnor U27526 (N_27526,N_27220,N_27234);
or U27527 (N_27527,N_27321,N_27267);
nand U27528 (N_27528,N_27305,N_27233);
nor U27529 (N_27529,N_27234,N_27232);
xor U27530 (N_27530,N_27234,N_27266);
xnor U27531 (N_27531,N_27291,N_27202);
nand U27532 (N_27532,N_27363,N_27386);
xnor U27533 (N_27533,N_27342,N_27329);
xnor U27534 (N_27534,N_27343,N_27391);
and U27535 (N_27535,N_27222,N_27279);
nor U27536 (N_27536,N_27269,N_27393);
or U27537 (N_27537,N_27279,N_27372);
or U27538 (N_27538,N_27240,N_27366);
or U27539 (N_27539,N_27301,N_27235);
nor U27540 (N_27540,N_27209,N_27223);
nand U27541 (N_27541,N_27367,N_27390);
nand U27542 (N_27542,N_27210,N_27298);
and U27543 (N_27543,N_27363,N_27278);
and U27544 (N_27544,N_27368,N_27302);
and U27545 (N_27545,N_27259,N_27385);
nor U27546 (N_27546,N_27231,N_27261);
xor U27547 (N_27547,N_27354,N_27300);
nor U27548 (N_27548,N_27260,N_27357);
nor U27549 (N_27549,N_27364,N_27268);
xor U27550 (N_27550,N_27286,N_27300);
nand U27551 (N_27551,N_27288,N_27253);
or U27552 (N_27552,N_27274,N_27349);
xnor U27553 (N_27553,N_27399,N_27333);
nor U27554 (N_27554,N_27263,N_27246);
and U27555 (N_27555,N_27330,N_27254);
xor U27556 (N_27556,N_27241,N_27222);
nor U27557 (N_27557,N_27264,N_27385);
xor U27558 (N_27558,N_27369,N_27319);
xnor U27559 (N_27559,N_27204,N_27371);
nor U27560 (N_27560,N_27228,N_27211);
nor U27561 (N_27561,N_27207,N_27392);
nor U27562 (N_27562,N_27321,N_27202);
or U27563 (N_27563,N_27287,N_27336);
nand U27564 (N_27564,N_27270,N_27368);
or U27565 (N_27565,N_27288,N_27218);
and U27566 (N_27566,N_27333,N_27382);
and U27567 (N_27567,N_27335,N_27353);
and U27568 (N_27568,N_27345,N_27330);
or U27569 (N_27569,N_27306,N_27288);
nor U27570 (N_27570,N_27308,N_27356);
or U27571 (N_27571,N_27356,N_27358);
and U27572 (N_27572,N_27398,N_27399);
and U27573 (N_27573,N_27388,N_27255);
nand U27574 (N_27574,N_27268,N_27360);
xor U27575 (N_27575,N_27256,N_27301);
and U27576 (N_27576,N_27230,N_27366);
nor U27577 (N_27577,N_27340,N_27223);
or U27578 (N_27578,N_27302,N_27219);
and U27579 (N_27579,N_27399,N_27224);
and U27580 (N_27580,N_27277,N_27313);
and U27581 (N_27581,N_27239,N_27227);
or U27582 (N_27582,N_27230,N_27240);
xnor U27583 (N_27583,N_27271,N_27257);
or U27584 (N_27584,N_27283,N_27355);
and U27585 (N_27585,N_27230,N_27286);
and U27586 (N_27586,N_27232,N_27288);
nor U27587 (N_27587,N_27225,N_27235);
and U27588 (N_27588,N_27233,N_27274);
nor U27589 (N_27589,N_27270,N_27391);
nand U27590 (N_27590,N_27295,N_27345);
and U27591 (N_27591,N_27286,N_27322);
nor U27592 (N_27592,N_27251,N_27337);
xor U27593 (N_27593,N_27293,N_27346);
and U27594 (N_27594,N_27392,N_27282);
and U27595 (N_27595,N_27295,N_27294);
or U27596 (N_27596,N_27327,N_27204);
and U27597 (N_27597,N_27225,N_27351);
nand U27598 (N_27598,N_27303,N_27381);
nor U27599 (N_27599,N_27335,N_27319);
nor U27600 (N_27600,N_27493,N_27587);
and U27601 (N_27601,N_27456,N_27409);
xor U27602 (N_27602,N_27460,N_27418);
and U27603 (N_27603,N_27511,N_27439);
and U27604 (N_27604,N_27518,N_27457);
nor U27605 (N_27605,N_27470,N_27589);
nor U27606 (N_27606,N_27403,N_27554);
or U27607 (N_27607,N_27442,N_27578);
nand U27608 (N_27608,N_27410,N_27400);
nand U27609 (N_27609,N_27421,N_27451);
or U27610 (N_27610,N_27429,N_27523);
and U27611 (N_27611,N_27454,N_27441);
xor U27612 (N_27612,N_27501,N_27513);
or U27613 (N_27613,N_27596,N_27468);
nor U27614 (N_27614,N_27407,N_27562);
or U27615 (N_27615,N_27595,N_27541);
nor U27616 (N_27616,N_27434,N_27514);
nor U27617 (N_27617,N_27526,N_27411);
and U27618 (N_27618,N_27505,N_27425);
or U27619 (N_27619,N_27423,N_27565);
nand U27620 (N_27620,N_27569,N_27459);
nor U27621 (N_27621,N_27545,N_27450);
nand U27622 (N_27622,N_27559,N_27427);
nor U27623 (N_27623,N_27424,N_27496);
nor U27624 (N_27624,N_27521,N_27416);
or U27625 (N_27625,N_27534,N_27476);
xnor U27626 (N_27626,N_27506,N_27447);
nand U27627 (N_27627,N_27499,N_27431);
and U27628 (N_27628,N_27548,N_27568);
xnor U27629 (N_27629,N_27445,N_27500);
xnor U27630 (N_27630,N_27404,N_27527);
xnor U27631 (N_27631,N_27497,N_27485);
nand U27632 (N_27632,N_27469,N_27529);
xnor U27633 (N_27633,N_27494,N_27530);
nand U27634 (N_27634,N_27560,N_27449);
or U27635 (N_27635,N_27571,N_27519);
nor U27636 (N_27636,N_27579,N_27414);
nor U27637 (N_27637,N_27401,N_27440);
or U27638 (N_27638,N_27558,N_27502);
nor U27639 (N_27639,N_27550,N_27438);
or U27640 (N_27640,N_27553,N_27586);
and U27641 (N_27641,N_27581,N_27446);
nor U27642 (N_27642,N_27417,N_27477);
xor U27643 (N_27643,N_27516,N_27537);
xor U27644 (N_27644,N_27535,N_27444);
xnor U27645 (N_27645,N_27566,N_27539);
or U27646 (N_27646,N_27585,N_27563);
or U27647 (N_27647,N_27413,N_27588);
or U27648 (N_27648,N_27488,N_27492);
nand U27649 (N_27649,N_27561,N_27582);
and U27650 (N_27650,N_27556,N_27590);
nand U27651 (N_27651,N_27528,N_27532);
and U27652 (N_27652,N_27593,N_27551);
and U27653 (N_27653,N_27402,N_27510);
nor U27654 (N_27654,N_27557,N_27515);
nand U27655 (N_27655,N_27584,N_27508);
nand U27656 (N_27656,N_27484,N_27599);
nor U27657 (N_27657,N_27422,N_27448);
or U27658 (N_27658,N_27426,N_27463);
nand U27659 (N_27659,N_27504,N_27509);
nand U27660 (N_27660,N_27486,N_27475);
xor U27661 (N_27661,N_27577,N_27572);
nand U27662 (N_27662,N_27435,N_27428);
nor U27663 (N_27663,N_27462,N_27544);
nand U27664 (N_27664,N_27415,N_27533);
xor U27665 (N_27665,N_27574,N_27443);
nand U27666 (N_27666,N_27594,N_27531);
nor U27667 (N_27667,N_27583,N_27473);
nor U27668 (N_27668,N_27481,N_27471);
xnor U27669 (N_27669,N_27461,N_27495);
nand U27670 (N_27670,N_27549,N_27430);
nand U27671 (N_27671,N_27580,N_27592);
and U27672 (N_27672,N_27525,N_27503);
nor U27673 (N_27673,N_27546,N_27487);
nand U27674 (N_27674,N_27408,N_27412);
xor U27675 (N_27675,N_27507,N_27540);
nor U27676 (N_27676,N_27405,N_27598);
and U27677 (N_27677,N_27489,N_27479);
xnor U27678 (N_27678,N_27591,N_27474);
nand U27679 (N_27679,N_27472,N_27543);
and U27680 (N_27680,N_27547,N_27522);
nor U27681 (N_27681,N_27524,N_27455);
nand U27682 (N_27682,N_27573,N_27490);
or U27683 (N_27683,N_27466,N_27482);
nor U27684 (N_27684,N_27419,N_27576);
nand U27685 (N_27685,N_27564,N_27437);
nor U27686 (N_27686,N_27555,N_27552);
nand U27687 (N_27687,N_27480,N_27491);
or U27688 (N_27688,N_27433,N_27536);
nor U27689 (N_27689,N_27465,N_27542);
nand U27690 (N_27690,N_27452,N_27597);
xnor U27691 (N_27691,N_27453,N_27567);
xor U27692 (N_27692,N_27420,N_27570);
nand U27693 (N_27693,N_27512,N_27432);
or U27694 (N_27694,N_27406,N_27538);
and U27695 (N_27695,N_27464,N_27458);
nor U27696 (N_27696,N_27478,N_27436);
nor U27697 (N_27697,N_27498,N_27517);
nand U27698 (N_27698,N_27483,N_27575);
xnor U27699 (N_27699,N_27520,N_27467);
or U27700 (N_27700,N_27547,N_27519);
and U27701 (N_27701,N_27473,N_27454);
nor U27702 (N_27702,N_27403,N_27494);
nand U27703 (N_27703,N_27540,N_27590);
xnor U27704 (N_27704,N_27442,N_27498);
and U27705 (N_27705,N_27448,N_27450);
nand U27706 (N_27706,N_27587,N_27557);
and U27707 (N_27707,N_27570,N_27497);
and U27708 (N_27708,N_27453,N_27562);
nor U27709 (N_27709,N_27475,N_27401);
and U27710 (N_27710,N_27493,N_27444);
and U27711 (N_27711,N_27508,N_27518);
or U27712 (N_27712,N_27578,N_27443);
nand U27713 (N_27713,N_27428,N_27599);
and U27714 (N_27714,N_27507,N_27461);
or U27715 (N_27715,N_27485,N_27576);
or U27716 (N_27716,N_27468,N_27500);
and U27717 (N_27717,N_27580,N_27420);
and U27718 (N_27718,N_27418,N_27405);
nand U27719 (N_27719,N_27508,N_27430);
nor U27720 (N_27720,N_27534,N_27438);
or U27721 (N_27721,N_27403,N_27411);
nand U27722 (N_27722,N_27439,N_27492);
nand U27723 (N_27723,N_27522,N_27471);
nand U27724 (N_27724,N_27418,N_27593);
nand U27725 (N_27725,N_27476,N_27426);
nand U27726 (N_27726,N_27523,N_27417);
nor U27727 (N_27727,N_27474,N_27490);
nand U27728 (N_27728,N_27469,N_27539);
xnor U27729 (N_27729,N_27473,N_27432);
nand U27730 (N_27730,N_27435,N_27529);
nand U27731 (N_27731,N_27527,N_27571);
xnor U27732 (N_27732,N_27453,N_27530);
nand U27733 (N_27733,N_27448,N_27534);
or U27734 (N_27734,N_27407,N_27442);
xor U27735 (N_27735,N_27581,N_27428);
nand U27736 (N_27736,N_27581,N_27538);
and U27737 (N_27737,N_27507,N_27576);
nand U27738 (N_27738,N_27459,N_27590);
and U27739 (N_27739,N_27431,N_27586);
xor U27740 (N_27740,N_27513,N_27499);
nand U27741 (N_27741,N_27463,N_27408);
nand U27742 (N_27742,N_27416,N_27503);
or U27743 (N_27743,N_27403,N_27476);
xnor U27744 (N_27744,N_27594,N_27556);
and U27745 (N_27745,N_27428,N_27533);
and U27746 (N_27746,N_27510,N_27565);
nor U27747 (N_27747,N_27518,N_27510);
and U27748 (N_27748,N_27559,N_27546);
and U27749 (N_27749,N_27564,N_27476);
and U27750 (N_27750,N_27520,N_27538);
or U27751 (N_27751,N_27480,N_27426);
nand U27752 (N_27752,N_27487,N_27413);
xnor U27753 (N_27753,N_27500,N_27548);
nor U27754 (N_27754,N_27577,N_27509);
nor U27755 (N_27755,N_27534,N_27539);
or U27756 (N_27756,N_27544,N_27590);
nand U27757 (N_27757,N_27473,N_27522);
nand U27758 (N_27758,N_27512,N_27517);
xnor U27759 (N_27759,N_27576,N_27400);
and U27760 (N_27760,N_27462,N_27513);
nor U27761 (N_27761,N_27578,N_27514);
nor U27762 (N_27762,N_27505,N_27570);
nor U27763 (N_27763,N_27495,N_27439);
xnor U27764 (N_27764,N_27490,N_27592);
and U27765 (N_27765,N_27595,N_27550);
or U27766 (N_27766,N_27467,N_27493);
nand U27767 (N_27767,N_27411,N_27487);
or U27768 (N_27768,N_27403,N_27505);
or U27769 (N_27769,N_27447,N_27454);
and U27770 (N_27770,N_27444,N_27551);
nor U27771 (N_27771,N_27549,N_27408);
and U27772 (N_27772,N_27508,N_27495);
and U27773 (N_27773,N_27412,N_27585);
and U27774 (N_27774,N_27571,N_27452);
nor U27775 (N_27775,N_27573,N_27459);
nor U27776 (N_27776,N_27559,N_27575);
or U27777 (N_27777,N_27582,N_27522);
or U27778 (N_27778,N_27472,N_27588);
and U27779 (N_27779,N_27587,N_27548);
or U27780 (N_27780,N_27445,N_27569);
or U27781 (N_27781,N_27545,N_27410);
xor U27782 (N_27782,N_27520,N_27401);
or U27783 (N_27783,N_27469,N_27461);
nand U27784 (N_27784,N_27494,N_27523);
or U27785 (N_27785,N_27559,N_27416);
or U27786 (N_27786,N_27446,N_27594);
or U27787 (N_27787,N_27463,N_27526);
or U27788 (N_27788,N_27403,N_27564);
or U27789 (N_27789,N_27465,N_27472);
and U27790 (N_27790,N_27533,N_27571);
nor U27791 (N_27791,N_27556,N_27510);
nor U27792 (N_27792,N_27447,N_27496);
nor U27793 (N_27793,N_27439,N_27456);
nor U27794 (N_27794,N_27489,N_27487);
nand U27795 (N_27795,N_27511,N_27469);
or U27796 (N_27796,N_27456,N_27424);
nor U27797 (N_27797,N_27517,N_27531);
or U27798 (N_27798,N_27513,N_27406);
and U27799 (N_27799,N_27480,N_27418);
nor U27800 (N_27800,N_27647,N_27659);
and U27801 (N_27801,N_27654,N_27762);
or U27802 (N_27802,N_27635,N_27711);
nor U27803 (N_27803,N_27718,N_27642);
nand U27804 (N_27804,N_27777,N_27629);
and U27805 (N_27805,N_27799,N_27617);
xnor U27806 (N_27806,N_27724,N_27779);
xnor U27807 (N_27807,N_27712,N_27767);
nand U27808 (N_27808,N_27685,N_27672);
xor U27809 (N_27809,N_27790,N_27774);
nor U27810 (N_27810,N_27632,N_27671);
or U27811 (N_27811,N_27795,N_27722);
nand U27812 (N_27812,N_27730,N_27726);
or U27813 (N_27813,N_27689,N_27785);
and U27814 (N_27814,N_27792,N_27789);
nand U27815 (N_27815,N_27612,N_27710);
xnor U27816 (N_27816,N_27641,N_27747);
and U27817 (N_27817,N_27615,N_27706);
nor U27818 (N_27818,N_27739,N_27748);
nand U27819 (N_27819,N_27791,N_27663);
nor U27820 (N_27820,N_27648,N_27652);
and U27821 (N_27821,N_27613,N_27657);
or U27822 (N_27822,N_27668,N_27787);
and U27823 (N_27823,N_27796,N_27660);
xor U27824 (N_27824,N_27743,N_27776);
or U27825 (N_27825,N_27728,N_27793);
xor U27826 (N_27826,N_27770,N_27670);
xnor U27827 (N_27827,N_27610,N_27696);
and U27828 (N_27828,N_27764,N_27715);
and U27829 (N_27829,N_27650,N_27622);
or U27830 (N_27830,N_27666,N_27752);
xnor U27831 (N_27831,N_27639,N_27757);
nand U27832 (N_27832,N_27771,N_27619);
or U27833 (N_27833,N_27631,N_27608);
and U27834 (N_27834,N_27611,N_27769);
xor U27835 (N_27835,N_27678,N_27602);
nand U27836 (N_27836,N_27624,N_27798);
or U27837 (N_27837,N_27614,N_27758);
and U27838 (N_27838,N_27754,N_27716);
and U27839 (N_27839,N_27677,N_27753);
and U27840 (N_27840,N_27725,N_27731);
nand U27841 (N_27841,N_27623,N_27662);
xor U27842 (N_27842,N_27675,N_27765);
or U27843 (N_27843,N_27603,N_27797);
nor U27844 (N_27844,N_27626,N_27708);
nand U27845 (N_27845,N_27698,N_27640);
and U27846 (N_27846,N_27750,N_27607);
nor U27847 (N_27847,N_27692,N_27719);
xnor U27848 (N_27848,N_27699,N_27656);
and U27849 (N_27849,N_27628,N_27618);
nand U27850 (N_27850,N_27676,N_27609);
xor U27851 (N_27851,N_27749,N_27649);
and U27852 (N_27852,N_27600,N_27697);
xor U27853 (N_27853,N_27721,N_27633);
and U27854 (N_27854,N_27646,N_27653);
nor U27855 (N_27855,N_27700,N_27766);
or U27856 (N_27856,N_27738,N_27773);
xnor U27857 (N_27857,N_27784,N_27736);
nand U27858 (N_27858,N_27705,N_27788);
or U27859 (N_27859,N_27780,N_27745);
nor U27860 (N_27860,N_27794,N_27768);
and U27861 (N_27861,N_27664,N_27683);
and U27862 (N_27862,N_27667,N_27778);
or U27863 (N_27863,N_27606,N_27687);
nor U27864 (N_27864,N_27604,N_27634);
xor U27865 (N_27865,N_27720,N_27638);
or U27866 (N_27866,N_27694,N_27704);
xnor U27867 (N_27867,N_27709,N_27695);
and U27868 (N_27868,N_27686,N_27605);
nand U27869 (N_27869,N_27760,N_27786);
or U27870 (N_27870,N_27701,N_27717);
xnor U27871 (N_27871,N_27636,N_27681);
xor U27872 (N_27872,N_27682,N_27742);
nor U27873 (N_27873,N_27755,N_27684);
xor U27874 (N_27874,N_27658,N_27688);
or U27875 (N_27875,N_27673,N_27645);
nand U27876 (N_27876,N_27772,N_27703);
or U27877 (N_27877,N_27729,N_27637);
or U27878 (N_27878,N_27775,N_27669);
or U27879 (N_27879,N_27643,N_27734);
and U27880 (N_27880,N_27713,N_27782);
and U27881 (N_27881,N_27644,N_27620);
nor U27882 (N_27882,N_27630,N_27665);
or U27883 (N_27883,N_27763,N_27714);
and U27884 (N_27884,N_27746,N_27621);
and U27885 (N_27885,N_27783,N_27616);
xnor U27886 (N_27886,N_27751,N_27691);
nor U27887 (N_27887,N_27727,N_27723);
or U27888 (N_27888,N_27693,N_27759);
or U27889 (N_27889,N_27679,N_27661);
nand U27890 (N_27890,N_27651,N_27737);
nand U27891 (N_27891,N_27741,N_27761);
xnor U27892 (N_27892,N_27601,N_27655);
xor U27893 (N_27893,N_27625,N_27733);
nand U27894 (N_27894,N_27756,N_27735);
nor U27895 (N_27895,N_27740,N_27674);
nand U27896 (N_27896,N_27744,N_27702);
nand U27897 (N_27897,N_27680,N_27690);
xor U27898 (N_27898,N_27707,N_27732);
or U27899 (N_27899,N_27627,N_27781);
and U27900 (N_27900,N_27728,N_27697);
and U27901 (N_27901,N_27772,N_27608);
nand U27902 (N_27902,N_27721,N_27706);
xor U27903 (N_27903,N_27749,N_27795);
xnor U27904 (N_27904,N_27639,N_27640);
or U27905 (N_27905,N_27697,N_27746);
and U27906 (N_27906,N_27621,N_27699);
or U27907 (N_27907,N_27632,N_27661);
nor U27908 (N_27908,N_27798,N_27631);
nand U27909 (N_27909,N_27765,N_27697);
nor U27910 (N_27910,N_27631,N_27725);
nor U27911 (N_27911,N_27606,N_27627);
xor U27912 (N_27912,N_27634,N_27691);
nand U27913 (N_27913,N_27768,N_27732);
and U27914 (N_27914,N_27694,N_27760);
xor U27915 (N_27915,N_27773,N_27684);
or U27916 (N_27916,N_27715,N_27738);
xnor U27917 (N_27917,N_27656,N_27745);
and U27918 (N_27918,N_27649,N_27689);
xor U27919 (N_27919,N_27664,N_27712);
nor U27920 (N_27920,N_27772,N_27731);
or U27921 (N_27921,N_27704,N_27777);
and U27922 (N_27922,N_27628,N_27659);
nand U27923 (N_27923,N_27743,N_27689);
or U27924 (N_27924,N_27658,N_27728);
and U27925 (N_27925,N_27635,N_27644);
or U27926 (N_27926,N_27641,N_27762);
xor U27927 (N_27927,N_27651,N_27769);
nand U27928 (N_27928,N_27600,N_27776);
nand U27929 (N_27929,N_27643,N_27743);
or U27930 (N_27930,N_27698,N_27650);
nor U27931 (N_27931,N_27738,N_27697);
and U27932 (N_27932,N_27654,N_27617);
xnor U27933 (N_27933,N_27672,N_27721);
nand U27934 (N_27934,N_27627,N_27706);
and U27935 (N_27935,N_27632,N_27748);
nand U27936 (N_27936,N_27682,N_27741);
nand U27937 (N_27937,N_27722,N_27623);
nor U27938 (N_27938,N_27651,N_27790);
nand U27939 (N_27939,N_27782,N_27666);
nand U27940 (N_27940,N_27644,N_27610);
nand U27941 (N_27941,N_27669,N_27634);
and U27942 (N_27942,N_27732,N_27735);
nand U27943 (N_27943,N_27744,N_27628);
nand U27944 (N_27944,N_27761,N_27680);
nor U27945 (N_27945,N_27769,N_27706);
nand U27946 (N_27946,N_27779,N_27736);
xnor U27947 (N_27947,N_27741,N_27667);
nor U27948 (N_27948,N_27799,N_27633);
nor U27949 (N_27949,N_27730,N_27666);
xnor U27950 (N_27950,N_27648,N_27685);
nand U27951 (N_27951,N_27752,N_27734);
and U27952 (N_27952,N_27649,N_27731);
or U27953 (N_27953,N_27712,N_27635);
xnor U27954 (N_27954,N_27668,N_27770);
nand U27955 (N_27955,N_27677,N_27604);
nand U27956 (N_27956,N_27609,N_27660);
or U27957 (N_27957,N_27614,N_27711);
and U27958 (N_27958,N_27614,N_27608);
nand U27959 (N_27959,N_27781,N_27713);
xor U27960 (N_27960,N_27771,N_27625);
xor U27961 (N_27961,N_27686,N_27706);
or U27962 (N_27962,N_27725,N_27616);
xor U27963 (N_27963,N_27751,N_27612);
xnor U27964 (N_27964,N_27708,N_27722);
nand U27965 (N_27965,N_27758,N_27645);
nor U27966 (N_27966,N_27600,N_27696);
and U27967 (N_27967,N_27667,N_27712);
and U27968 (N_27968,N_27655,N_27610);
nand U27969 (N_27969,N_27648,N_27748);
xnor U27970 (N_27970,N_27673,N_27630);
and U27971 (N_27971,N_27717,N_27698);
nor U27972 (N_27972,N_27705,N_27744);
and U27973 (N_27973,N_27710,N_27753);
and U27974 (N_27974,N_27706,N_27670);
nand U27975 (N_27975,N_27652,N_27729);
xnor U27976 (N_27976,N_27706,N_27687);
nor U27977 (N_27977,N_27664,N_27632);
or U27978 (N_27978,N_27694,N_27648);
or U27979 (N_27979,N_27630,N_27797);
xor U27980 (N_27980,N_27615,N_27786);
xnor U27981 (N_27981,N_27774,N_27635);
nand U27982 (N_27982,N_27774,N_27797);
nor U27983 (N_27983,N_27730,N_27629);
or U27984 (N_27984,N_27670,N_27645);
nor U27985 (N_27985,N_27693,N_27617);
or U27986 (N_27986,N_27646,N_27679);
and U27987 (N_27987,N_27727,N_27670);
nand U27988 (N_27988,N_27649,N_27764);
nor U27989 (N_27989,N_27705,N_27761);
nand U27990 (N_27990,N_27776,N_27795);
nor U27991 (N_27991,N_27719,N_27614);
xnor U27992 (N_27992,N_27700,N_27701);
or U27993 (N_27993,N_27745,N_27701);
nand U27994 (N_27994,N_27688,N_27703);
nor U27995 (N_27995,N_27688,N_27648);
nand U27996 (N_27996,N_27617,N_27765);
nor U27997 (N_27997,N_27600,N_27623);
nand U27998 (N_27998,N_27622,N_27786);
or U27999 (N_27999,N_27698,N_27758);
nor U28000 (N_28000,N_27956,N_27802);
nand U28001 (N_28001,N_27930,N_27894);
nand U28002 (N_28002,N_27887,N_27916);
nor U28003 (N_28003,N_27948,N_27908);
or U28004 (N_28004,N_27852,N_27839);
nor U28005 (N_28005,N_27922,N_27947);
nor U28006 (N_28006,N_27877,N_27935);
xor U28007 (N_28007,N_27964,N_27957);
xor U28008 (N_28008,N_27832,N_27861);
and U28009 (N_28009,N_27933,N_27962);
or U28010 (N_28010,N_27958,N_27815);
nor U28011 (N_28011,N_27854,N_27872);
or U28012 (N_28012,N_27803,N_27897);
nor U28013 (N_28013,N_27899,N_27939);
or U28014 (N_28014,N_27886,N_27848);
xor U28015 (N_28015,N_27972,N_27955);
and U28016 (N_28016,N_27924,N_27992);
or U28017 (N_28017,N_27889,N_27902);
nor U28018 (N_28018,N_27813,N_27904);
xnor U28019 (N_28019,N_27912,N_27966);
nor U28020 (N_28020,N_27943,N_27817);
and U28021 (N_28021,N_27995,N_27806);
or U28022 (N_28022,N_27827,N_27835);
or U28023 (N_28023,N_27941,N_27884);
nor U28024 (N_28024,N_27856,N_27867);
xor U28025 (N_28025,N_27984,N_27860);
nor U28026 (N_28026,N_27853,N_27976);
and U28027 (N_28027,N_27847,N_27882);
and U28028 (N_28028,N_27844,N_27828);
xor U28029 (N_28029,N_27951,N_27927);
or U28030 (N_28030,N_27991,N_27918);
and U28031 (N_28031,N_27859,N_27881);
nor U28032 (N_28032,N_27879,N_27906);
or U28033 (N_28033,N_27961,N_27915);
or U28034 (N_28034,N_27807,N_27934);
nand U28035 (N_28035,N_27804,N_27925);
and U28036 (N_28036,N_27805,N_27843);
or U28037 (N_28037,N_27893,N_27871);
or U28038 (N_28038,N_27836,N_27980);
nand U28039 (N_28039,N_27910,N_27842);
and U28040 (N_28040,N_27949,N_27896);
or U28041 (N_28041,N_27946,N_27826);
nand U28042 (N_28042,N_27845,N_27870);
and U28043 (N_28043,N_27875,N_27833);
or U28044 (N_28044,N_27923,N_27811);
or U28045 (N_28045,N_27900,N_27869);
or U28046 (N_28046,N_27953,N_27849);
or U28047 (N_28047,N_27998,N_27876);
nor U28048 (N_28048,N_27862,N_27830);
xnor U28049 (N_28049,N_27824,N_27858);
xor U28050 (N_28050,N_27829,N_27838);
xnor U28051 (N_28051,N_27960,N_27969);
and U28052 (N_28052,N_27954,N_27865);
or U28053 (N_28053,N_27970,N_27978);
xnor U28054 (N_28054,N_27928,N_27952);
nand U28055 (N_28055,N_27973,N_27901);
or U28056 (N_28056,N_27816,N_27909);
nor U28057 (N_28057,N_27979,N_27937);
nor U28058 (N_28058,N_27890,N_27857);
nand U28059 (N_28059,N_27866,N_27989);
and U28060 (N_28060,N_27841,N_27938);
and U28061 (N_28061,N_27840,N_27959);
nor U28062 (N_28062,N_27987,N_27965);
nand U28063 (N_28063,N_27968,N_27885);
and U28064 (N_28064,N_27967,N_27950);
and U28065 (N_28065,N_27974,N_27850);
nor U28066 (N_28066,N_27990,N_27888);
nor U28067 (N_28067,N_27810,N_27863);
or U28068 (N_28068,N_27883,N_27999);
or U28069 (N_28069,N_27821,N_27920);
xnor U28070 (N_28070,N_27864,N_27808);
nor U28071 (N_28071,N_27818,N_27994);
nor U28072 (N_28072,N_27825,N_27820);
nor U28073 (N_28073,N_27809,N_27873);
nand U28074 (N_28074,N_27814,N_27891);
nand U28075 (N_28075,N_27993,N_27905);
xnor U28076 (N_28076,N_27919,N_27988);
or U28077 (N_28077,N_27819,N_27831);
nor U28078 (N_28078,N_27801,N_27936);
or U28079 (N_28079,N_27812,N_27985);
xnor U28080 (N_28080,N_27855,N_27982);
or U28081 (N_28081,N_27975,N_27926);
and U28082 (N_28082,N_27944,N_27878);
xnor U28083 (N_28083,N_27868,N_27846);
xor U28084 (N_28084,N_27917,N_27921);
xor U28085 (N_28085,N_27895,N_27945);
nand U28086 (N_28086,N_27822,N_27851);
nor U28087 (N_28087,N_27932,N_27834);
nand U28088 (N_28088,N_27997,N_27963);
xnor U28089 (N_28089,N_27986,N_27903);
nor U28090 (N_28090,N_27940,N_27914);
nand U28091 (N_28091,N_27977,N_27800);
or U28092 (N_28092,N_27874,N_27898);
nand U28093 (N_28093,N_27911,N_27837);
xor U28094 (N_28094,N_27983,N_27892);
xnor U28095 (N_28095,N_27942,N_27823);
nand U28096 (N_28096,N_27929,N_27971);
nor U28097 (N_28097,N_27880,N_27907);
and U28098 (N_28098,N_27981,N_27996);
xnor U28099 (N_28099,N_27931,N_27913);
nand U28100 (N_28100,N_27969,N_27995);
xor U28101 (N_28101,N_27959,N_27969);
or U28102 (N_28102,N_27852,N_27871);
and U28103 (N_28103,N_27803,N_27891);
xnor U28104 (N_28104,N_27963,N_27814);
or U28105 (N_28105,N_27939,N_27928);
or U28106 (N_28106,N_27922,N_27928);
xor U28107 (N_28107,N_27839,N_27801);
nor U28108 (N_28108,N_27889,N_27867);
nand U28109 (N_28109,N_27986,N_27828);
nor U28110 (N_28110,N_27818,N_27844);
xor U28111 (N_28111,N_27993,N_27828);
or U28112 (N_28112,N_27864,N_27815);
or U28113 (N_28113,N_27914,N_27988);
and U28114 (N_28114,N_27938,N_27989);
xor U28115 (N_28115,N_27973,N_27946);
and U28116 (N_28116,N_27970,N_27820);
nand U28117 (N_28117,N_27979,N_27982);
nand U28118 (N_28118,N_27947,N_27835);
and U28119 (N_28119,N_27861,N_27839);
xor U28120 (N_28120,N_27948,N_27893);
or U28121 (N_28121,N_27894,N_27925);
xnor U28122 (N_28122,N_27913,N_27927);
or U28123 (N_28123,N_27874,N_27948);
and U28124 (N_28124,N_27988,N_27941);
nor U28125 (N_28125,N_27829,N_27840);
nor U28126 (N_28126,N_27933,N_27877);
xor U28127 (N_28127,N_27936,N_27876);
and U28128 (N_28128,N_27815,N_27896);
or U28129 (N_28129,N_27962,N_27983);
or U28130 (N_28130,N_27960,N_27879);
xnor U28131 (N_28131,N_27999,N_27856);
nand U28132 (N_28132,N_27961,N_27834);
and U28133 (N_28133,N_27980,N_27944);
nand U28134 (N_28134,N_27913,N_27827);
or U28135 (N_28135,N_27879,N_27988);
or U28136 (N_28136,N_27998,N_27878);
nand U28137 (N_28137,N_27948,N_27800);
xor U28138 (N_28138,N_27930,N_27812);
xnor U28139 (N_28139,N_27987,N_27875);
or U28140 (N_28140,N_27861,N_27835);
or U28141 (N_28141,N_27930,N_27822);
or U28142 (N_28142,N_27997,N_27986);
xnor U28143 (N_28143,N_27987,N_27859);
xor U28144 (N_28144,N_27956,N_27970);
and U28145 (N_28145,N_27855,N_27968);
and U28146 (N_28146,N_27901,N_27958);
or U28147 (N_28147,N_27834,N_27919);
or U28148 (N_28148,N_27982,N_27984);
and U28149 (N_28149,N_27905,N_27916);
or U28150 (N_28150,N_27901,N_27994);
xnor U28151 (N_28151,N_27882,N_27987);
nor U28152 (N_28152,N_27979,N_27904);
nor U28153 (N_28153,N_27967,N_27854);
or U28154 (N_28154,N_27871,N_27806);
xor U28155 (N_28155,N_27928,N_27938);
nor U28156 (N_28156,N_27931,N_27838);
or U28157 (N_28157,N_27806,N_27853);
xor U28158 (N_28158,N_27983,N_27910);
nand U28159 (N_28159,N_27966,N_27990);
and U28160 (N_28160,N_27901,N_27921);
nor U28161 (N_28161,N_27813,N_27909);
or U28162 (N_28162,N_27904,N_27831);
nor U28163 (N_28163,N_27916,N_27974);
or U28164 (N_28164,N_27884,N_27838);
and U28165 (N_28165,N_27964,N_27860);
xnor U28166 (N_28166,N_27925,N_27959);
or U28167 (N_28167,N_27942,N_27835);
nand U28168 (N_28168,N_27844,N_27951);
xor U28169 (N_28169,N_27953,N_27842);
and U28170 (N_28170,N_27873,N_27967);
and U28171 (N_28171,N_27816,N_27863);
or U28172 (N_28172,N_27851,N_27812);
nor U28173 (N_28173,N_27886,N_27817);
nand U28174 (N_28174,N_27949,N_27862);
xor U28175 (N_28175,N_27836,N_27822);
or U28176 (N_28176,N_27860,N_27903);
and U28177 (N_28177,N_27925,N_27949);
nand U28178 (N_28178,N_27835,N_27967);
nor U28179 (N_28179,N_27902,N_27995);
and U28180 (N_28180,N_27817,N_27908);
and U28181 (N_28181,N_27977,N_27850);
nor U28182 (N_28182,N_27897,N_27856);
nand U28183 (N_28183,N_27881,N_27902);
and U28184 (N_28184,N_27933,N_27863);
nand U28185 (N_28185,N_27869,N_27951);
nand U28186 (N_28186,N_27997,N_27983);
and U28187 (N_28187,N_27860,N_27934);
and U28188 (N_28188,N_27918,N_27965);
or U28189 (N_28189,N_27886,N_27805);
nor U28190 (N_28190,N_27845,N_27976);
xor U28191 (N_28191,N_27906,N_27820);
and U28192 (N_28192,N_27811,N_27849);
or U28193 (N_28193,N_27983,N_27904);
xnor U28194 (N_28194,N_27835,N_27915);
xor U28195 (N_28195,N_27878,N_27920);
nor U28196 (N_28196,N_27938,N_27963);
and U28197 (N_28197,N_27914,N_27998);
xor U28198 (N_28198,N_27859,N_27812);
nor U28199 (N_28199,N_27908,N_27826);
nand U28200 (N_28200,N_28075,N_28110);
nor U28201 (N_28201,N_28166,N_28141);
or U28202 (N_28202,N_28108,N_28043);
xnor U28203 (N_28203,N_28015,N_28102);
or U28204 (N_28204,N_28100,N_28098);
nand U28205 (N_28205,N_28135,N_28091);
nand U28206 (N_28206,N_28073,N_28169);
xnor U28207 (N_28207,N_28033,N_28105);
nand U28208 (N_28208,N_28037,N_28142);
or U28209 (N_28209,N_28176,N_28183);
or U28210 (N_28210,N_28174,N_28190);
and U28211 (N_28211,N_28162,N_28045);
nand U28212 (N_28212,N_28197,N_28074);
and U28213 (N_28213,N_28002,N_28010);
and U28214 (N_28214,N_28158,N_28023);
nand U28215 (N_28215,N_28006,N_28021);
xor U28216 (N_28216,N_28035,N_28184);
and U28217 (N_28217,N_28181,N_28192);
nor U28218 (N_28218,N_28124,N_28149);
or U28219 (N_28219,N_28012,N_28125);
and U28220 (N_28220,N_28078,N_28143);
nor U28221 (N_28221,N_28063,N_28112);
or U28222 (N_28222,N_28147,N_28089);
or U28223 (N_28223,N_28080,N_28048);
or U28224 (N_28224,N_28022,N_28069);
and U28225 (N_28225,N_28017,N_28072);
or U28226 (N_28226,N_28189,N_28032);
nand U28227 (N_28227,N_28177,N_28107);
nand U28228 (N_28228,N_28179,N_28085);
and U28229 (N_28229,N_28016,N_28011);
or U28230 (N_28230,N_28101,N_28053);
and U28231 (N_28231,N_28175,N_28103);
nor U28232 (N_28232,N_28027,N_28131);
xnor U28233 (N_28233,N_28092,N_28150);
nand U28234 (N_28234,N_28173,N_28165);
nand U28235 (N_28235,N_28159,N_28128);
xnor U28236 (N_28236,N_28090,N_28029);
or U28237 (N_28237,N_28066,N_28031);
and U28238 (N_28238,N_28121,N_28084);
nor U28239 (N_28239,N_28172,N_28062);
nor U28240 (N_28240,N_28134,N_28161);
xor U28241 (N_28241,N_28140,N_28148);
or U28242 (N_28242,N_28038,N_28046);
nand U28243 (N_28243,N_28019,N_28094);
xnor U28244 (N_28244,N_28160,N_28057);
or U28245 (N_28245,N_28061,N_28186);
and U28246 (N_28246,N_28138,N_28130);
nor U28247 (N_28247,N_28146,N_28115);
and U28248 (N_28248,N_28157,N_28077);
or U28249 (N_28249,N_28058,N_28060);
nor U28250 (N_28250,N_28003,N_28154);
nand U28251 (N_28251,N_28195,N_28026);
or U28252 (N_28252,N_28117,N_28139);
and U28253 (N_28253,N_28034,N_28056);
nand U28254 (N_28254,N_28054,N_28164);
nand U28255 (N_28255,N_28178,N_28059);
nor U28256 (N_28256,N_28133,N_28096);
xnor U28257 (N_28257,N_28009,N_28024);
nand U28258 (N_28258,N_28137,N_28086);
or U28259 (N_28259,N_28049,N_28004);
or U28260 (N_28260,N_28007,N_28151);
or U28261 (N_28261,N_28114,N_28047);
xnor U28262 (N_28262,N_28129,N_28081);
nand U28263 (N_28263,N_28155,N_28180);
or U28264 (N_28264,N_28118,N_28093);
nand U28265 (N_28265,N_28144,N_28005);
or U28266 (N_28266,N_28187,N_28167);
nor U28267 (N_28267,N_28122,N_28042);
nand U28268 (N_28268,N_28170,N_28095);
xor U28269 (N_28269,N_28132,N_28194);
nor U28270 (N_28270,N_28126,N_28099);
and U28271 (N_28271,N_28040,N_28065);
and U28272 (N_28272,N_28052,N_28050);
nand U28273 (N_28273,N_28156,N_28018);
nor U28274 (N_28274,N_28008,N_28044);
nand U28275 (N_28275,N_28185,N_28028);
or U28276 (N_28276,N_28113,N_28000);
nor U28277 (N_28277,N_28083,N_28088);
nand U28278 (N_28278,N_28193,N_28111);
nand U28279 (N_28279,N_28136,N_28152);
or U28280 (N_28280,N_28039,N_28163);
and U28281 (N_28281,N_28087,N_28116);
or U28282 (N_28282,N_28001,N_28051);
nand U28283 (N_28283,N_28182,N_28041);
or U28284 (N_28284,N_28068,N_28030);
nor U28285 (N_28285,N_28196,N_28104);
xnor U28286 (N_28286,N_28123,N_28082);
xor U28287 (N_28287,N_28199,N_28071);
xor U28288 (N_28288,N_28064,N_28036);
nand U28289 (N_28289,N_28097,N_28020);
nor U28290 (N_28290,N_28191,N_28013);
xnor U28291 (N_28291,N_28109,N_28067);
or U28292 (N_28292,N_28127,N_28076);
xor U28293 (N_28293,N_28120,N_28198);
nand U28294 (N_28294,N_28106,N_28153);
and U28295 (N_28295,N_28119,N_28014);
nand U28296 (N_28296,N_28025,N_28079);
nor U28297 (N_28297,N_28055,N_28171);
xnor U28298 (N_28298,N_28168,N_28070);
or U28299 (N_28299,N_28188,N_28145);
or U28300 (N_28300,N_28117,N_28060);
nor U28301 (N_28301,N_28174,N_28175);
xnor U28302 (N_28302,N_28029,N_28071);
nor U28303 (N_28303,N_28034,N_28122);
or U28304 (N_28304,N_28043,N_28005);
xnor U28305 (N_28305,N_28131,N_28019);
xor U28306 (N_28306,N_28191,N_28060);
xor U28307 (N_28307,N_28120,N_28134);
nor U28308 (N_28308,N_28196,N_28167);
or U28309 (N_28309,N_28087,N_28192);
or U28310 (N_28310,N_28033,N_28022);
or U28311 (N_28311,N_28064,N_28148);
nor U28312 (N_28312,N_28178,N_28177);
nor U28313 (N_28313,N_28092,N_28194);
xor U28314 (N_28314,N_28116,N_28189);
and U28315 (N_28315,N_28055,N_28197);
and U28316 (N_28316,N_28067,N_28011);
and U28317 (N_28317,N_28069,N_28100);
and U28318 (N_28318,N_28088,N_28179);
nand U28319 (N_28319,N_28186,N_28054);
and U28320 (N_28320,N_28182,N_28030);
xnor U28321 (N_28321,N_28031,N_28005);
and U28322 (N_28322,N_28100,N_28153);
nor U28323 (N_28323,N_28092,N_28044);
xor U28324 (N_28324,N_28179,N_28130);
xnor U28325 (N_28325,N_28110,N_28169);
nor U28326 (N_28326,N_28042,N_28000);
and U28327 (N_28327,N_28032,N_28060);
xnor U28328 (N_28328,N_28164,N_28046);
nor U28329 (N_28329,N_28192,N_28016);
xor U28330 (N_28330,N_28131,N_28125);
and U28331 (N_28331,N_28099,N_28046);
or U28332 (N_28332,N_28032,N_28066);
nor U28333 (N_28333,N_28160,N_28137);
nand U28334 (N_28334,N_28170,N_28085);
and U28335 (N_28335,N_28111,N_28123);
nand U28336 (N_28336,N_28006,N_28111);
or U28337 (N_28337,N_28161,N_28020);
or U28338 (N_28338,N_28126,N_28149);
nor U28339 (N_28339,N_28048,N_28041);
nor U28340 (N_28340,N_28109,N_28192);
or U28341 (N_28341,N_28109,N_28164);
nor U28342 (N_28342,N_28170,N_28005);
xor U28343 (N_28343,N_28150,N_28164);
nor U28344 (N_28344,N_28158,N_28118);
xnor U28345 (N_28345,N_28141,N_28010);
and U28346 (N_28346,N_28054,N_28197);
nand U28347 (N_28347,N_28153,N_28198);
or U28348 (N_28348,N_28193,N_28030);
or U28349 (N_28349,N_28097,N_28023);
or U28350 (N_28350,N_28167,N_28083);
nor U28351 (N_28351,N_28042,N_28025);
or U28352 (N_28352,N_28189,N_28136);
and U28353 (N_28353,N_28074,N_28123);
and U28354 (N_28354,N_28016,N_28134);
nand U28355 (N_28355,N_28132,N_28087);
nor U28356 (N_28356,N_28180,N_28162);
nor U28357 (N_28357,N_28048,N_28185);
xor U28358 (N_28358,N_28018,N_28122);
nand U28359 (N_28359,N_28181,N_28130);
xnor U28360 (N_28360,N_28048,N_28164);
xor U28361 (N_28361,N_28032,N_28199);
and U28362 (N_28362,N_28033,N_28081);
nand U28363 (N_28363,N_28082,N_28059);
or U28364 (N_28364,N_28044,N_28180);
xnor U28365 (N_28365,N_28019,N_28027);
nor U28366 (N_28366,N_28182,N_28199);
nor U28367 (N_28367,N_28108,N_28152);
nor U28368 (N_28368,N_28093,N_28010);
or U28369 (N_28369,N_28013,N_28176);
xor U28370 (N_28370,N_28102,N_28055);
nand U28371 (N_28371,N_28196,N_28136);
or U28372 (N_28372,N_28001,N_28141);
xnor U28373 (N_28373,N_28199,N_28181);
nor U28374 (N_28374,N_28010,N_28048);
or U28375 (N_28375,N_28034,N_28028);
nor U28376 (N_28376,N_28110,N_28151);
and U28377 (N_28377,N_28191,N_28113);
and U28378 (N_28378,N_28047,N_28076);
or U28379 (N_28379,N_28180,N_28149);
xor U28380 (N_28380,N_28062,N_28022);
or U28381 (N_28381,N_28020,N_28140);
nor U28382 (N_28382,N_28147,N_28155);
nand U28383 (N_28383,N_28198,N_28131);
nand U28384 (N_28384,N_28062,N_28019);
and U28385 (N_28385,N_28175,N_28189);
nor U28386 (N_28386,N_28095,N_28071);
or U28387 (N_28387,N_28088,N_28023);
and U28388 (N_28388,N_28063,N_28001);
nor U28389 (N_28389,N_28032,N_28009);
nand U28390 (N_28390,N_28163,N_28173);
nand U28391 (N_28391,N_28048,N_28062);
nor U28392 (N_28392,N_28014,N_28101);
and U28393 (N_28393,N_28145,N_28115);
nor U28394 (N_28394,N_28099,N_28158);
nor U28395 (N_28395,N_28123,N_28196);
xor U28396 (N_28396,N_28194,N_28020);
nand U28397 (N_28397,N_28011,N_28162);
and U28398 (N_28398,N_28121,N_28052);
and U28399 (N_28399,N_28020,N_28050);
and U28400 (N_28400,N_28354,N_28216);
nand U28401 (N_28401,N_28374,N_28367);
and U28402 (N_28402,N_28304,N_28246);
or U28403 (N_28403,N_28315,N_28231);
and U28404 (N_28404,N_28218,N_28344);
nand U28405 (N_28405,N_28392,N_28361);
xnor U28406 (N_28406,N_28395,N_28225);
xor U28407 (N_28407,N_28261,N_28278);
nand U28408 (N_28408,N_28250,N_28251);
or U28409 (N_28409,N_28248,N_28378);
nor U28410 (N_28410,N_28204,N_28329);
or U28411 (N_28411,N_28317,N_28272);
nor U28412 (N_28412,N_28215,N_28287);
nand U28413 (N_28413,N_28305,N_28267);
nor U28414 (N_28414,N_28381,N_28312);
and U28415 (N_28415,N_28235,N_28295);
or U28416 (N_28416,N_28323,N_28290);
nand U28417 (N_28417,N_28343,N_28217);
xor U28418 (N_28418,N_28281,N_28228);
xor U28419 (N_28419,N_28286,N_28206);
nor U28420 (N_28420,N_28283,N_28234);
or U28421 (N_28421,N_28226,N_28256);
or U28422 (N_28422,N_28365,N_28252);
nand U28423 (N_28423,N_28334,N_28389);
xor U28424 (N_28424,N_28316,N_28385);
xor U28425 (N_28425,N_28351,N_28306);
or U28426 (N_28426,N_28280,N_28349);
nor U28427 (N_28427,N_28275,N_28296);
xor U28428 (N_28428,N_28284,N_28239);
nor U28429 (N_28429,N_28331,N_28253);
xnor U28430 (N_28430,N_28375,N_28314);
nand U28431 (N_28431,N_28237,N_28242);
and U28432 (N_28432,N_28310,N_28363);
nand U28433 (N_28433,N_28222,N_28373);
nand U28434 (N_28434,N_28386,N_28266);
xnor U28435 (N_28435,N_28370,N_28391);
nand U28436 (N_28436,N_28247,N_28353);
or U28437 (N_28437,N_28200,N_28350);
or U28438 (N_28438,N_28233,N_28293);
xor U28439 (N_28439,N_28236,N_28338);
nand U28440 (N_28440,N_28227,N_28270);
nor U28441 (N_28441,N_28336,N_28399);
nand U28442 (N_28442,N_28273,N_28264);
nor U28443 (N_28443,N_28262,N_28357);
nand U28444 (N_28444,N_28319,N_28372);
nor U28445 (N_28445,N_28297,N_28397);
nor U28446 (N_28446,N_28309,N_28318);
xnor U28447 (N_28447,N_28209,N_28355);
or U28448 (N_28448,N_28269,N_28330);
nor U28449 (N_28449,N_28211,N_28327);
or U28450 (N_28450,N_28207,N_28324);
nand U28451 (N_28451,N_28332,N_28241);
or U28452 (N_28452,N_28255,N_28277);
or U28453 (N_28453,N_28288,N_28282);
or U28454 (N_28454,N_28383,N_28307);
nand U28455 (N_28455,N_28291,N_28202);
or U28456 (N_28456,N_28366,N_28232);
and U28457 (N_28457,N_28380,N_28294);
or U28458 (N_28458,N_28249,N_28276);
nand U28459 (N_28459,N_28258,N_28360);
nand U28460 (N_28460,N_28348,N_28302);
or U28461 (N_28461,N_28292,N_28208);
nor U28462 (N_28462,N_28342,N_28274);
nor U28463 (N_28463,N_28326,N_28285);
nand U28464 (N_28464,N_28201,N_28322);
xnor U28465 (N_28465,N_28393,N_28333);
or U28466 (N_28466,N_28203,N_28337);
or U28467 (N_28467,N_28303,N_28238);
and U28468 (N_28468,N_28388,N_28394);
and U28469 (N_28469,N_28346,N_28219);
and U28470 (N_28470,N_28213,N_28221);
nand U28471 (N_28471,N_28358,N_28223);
nand U28472 (N_28472,N_28244,N_28260);
nor U28473 (N_28473,N_28268,N_28390);
nand U28474 (N_28474,N_28259,N_28359);
xnor U28475 (N_28475,N_28254,N_28263);
nor U28476 (N_28476,N_28210,N_28311);
nor U28477 (N_28477,N_28300,N_28279);
nor U28478 (N_28478,N_28387,N_28205);
nand U28479 (N_28479,N_28313,N_28376);
nor U28480 (N_28480,N_28325,N_28214);
or U28481 (N_28481,N_28289,N_28328);
and U28482 (N_28482,N_28298,N_28362);
nor U28483 (N_28483,N_28398,N_28308);
or U28484 (N_28484,N_28224,N_28379);
nand U28485 (N_28485,N_28341,N_28320);
nor U28486 (N_28486,N_28335,N_28369);
xor U28487 (N_28487,N_28301,N_28245);
or U28488 (N_28488,N_28265,N_28371);
nand U28489 (N_28489,N_28271,N_28340);
and U28490 (N_28490,N_28339,N_28229);
nand U28491 (N_28491,N_28382,N_28377);
and U28492 (N_28492,N_28347,N_28364);
nand U28493 (N_28493,N_28230,N_28243);
and U28494 (N_28494,N_28356,N_28257);
nand U28495 (N_28495,N_28212,N_28220);
and U28496 (N_28496,N_28345,N_28321);
nor U28497 (N_28497,N_28352,N_28396);
nand U28498 (N_28498,N_28368,N_28299);
or U28499 (N_28499,N_28240,N_28384);
nor U28500 (N_28500,N_28338,N_28203);
nor U28501 (N_28501,N_28255,N_28399);
or U28502 (N_28502,N_28357,N_28206);
xor U28503 (N_28503,N_28399,N_28252);
nor U28504 (N_28504,N_28351,N_28319);
and U28505 (N_28505,N_28222,N_28205);
and U28506 (N_28506,N_28310,N_28221);
or U28507 (N_28507,N_28239,N_28283);
or U28508 (N_28508,N_28200,N_28260);
nor U28509 (N_28509,N_28222,N_28301);
xnor U28510 (N_28510,N_28357,N_28362);
xor U28511 (N_28511,N_28265,N_28330);
and U28512 (N_28512,N_28262,N_28222);
or U28513 (N_28513,N_28333,N_28326);
nor U28514 (N_28514,N_28371,N_28282);
and U28515 (N_28515,N_28349,N_28285);
xor U28516 (N_28516,N_28299,N_28330);
nor U28517 (N_28517,N_28353,N_28214);
or U28518 (N_28518,N_28219,N_28324);
and U28519 (N_28519,N_28259,N_28340);
nor U28520 (N_28520,N_28200,N_28267);
or U28521 (N_28521,N_28331,N_28393);
nor U28522 (N_28522,N_28362,N_28324);
and U28523 (N_28523,N_28379,N_28289);
nand U28524 (N_28524,N_28219,N_28236);
nand U28525 (N_28525,N_28338,N_28344);
xor U28526 (N_28526,N_28224,N_28385);
and U28527 (N_28527,N_28377,N_28356);
nand U28528 (N_28528,N_28346,N_28325);
and U28529 (N_28529,N_28358,N_28231);
xor U28530 (N_28530,N_28381,N_28215);
nor U28531 (N_28531,N_28333,N_28214);
nand U28532 (N_28532,N_28249,N_28373);
nand U28533 (N_28533,N_28384,N_28329);
or U28534 (N_28534,N_28247,N_28388);
nor U28535 (N_28535,N_28358,N_28314);
nor U28536 (N_28536,N_28227,N_28382);
or U28537 (N_28537,N_28313,N_28317);
or U28538 (N_28538,N_28362,N_28398);
nand U28539 (N_28539,N_28354,N_28219);
nor U28540 (N_28540,N_28372,N_28359);
or U28541 (N_28541,N_28383,N_28331);
nor U28542 (N_28542,N_28344,N_28271);
or U28543 (N_28543,N_28392,N_28362);
nand U28544 (N_28544,N_28333,N_28216);
xor U28545 (N_28545,N_28218,N_28331);
nand U28546 (N_28546,N_28343,N_28204);
or U28547 (N_28547,N_28381,N_28255);
and U28548 (N_28548,N_28384,N_28211);
xor U28549 (N_28549,N_28337,N_28273);
nand U28550 (N_28550,N_28335,N_28216);
xor U28551 (N_28551,N_28292,N_28228);
nand U28552 (N_28552,N_28366,N_28367);
nand U28553 (N_28553,N_28361,N_28214);
nor U28554 (N_28554,N_28202,N_28263);
or U28555 (N_28555,N_28363,N_28260);
nand U28556 (N_28556,N_28325,N_28202);
and U28557 (N_28557,N_28290,N_28201);
and U28558 (N_28558,N_28233,N_28248);
nand U28559 (N_28559,N_28295,N_28268);
xnor U28560 (N_28560,N_28238,N_28257);
xor U28561 (N_28561,N_28399,N_28223);
and U28562 (N_28562,N_28310,N_28245);
or U28563 (N_28563,N_28367,N_28318);
or U28564 (N_28564,N_28201,N_28312);
xnor U28565 (N_28565,N_28278,N_28240);
nor U28566 (N_28566,N_28339,N_28313);
nor U28567 (N_28567,N_28321,N_28272);
or U28568 (N_28568,N_28205,N_28265);
nor U28569 (N_28569,N_28343,N_28340);
or U28570 (N_28570,N_28238,N_28219);
or U28571 (N_28571,N_28222,N_28238);
nand U28572 (N_28572,N_28206,N_28392);
or U28573 (N_28573,N_28216,N_28282);
and U28574 (N_28574,N_28257,N_28280);
and U28575 (N_28575,N_28386,N_28293);
nand U28576 (N_28576,N_28364,N_28299);
and U28577 (N_28577,N_28245,N_28267);
nor U28578 (N_28578,N_28341,N_28286);
or U28579 (N_28579,N_28370,N_28376);
nand U28580 (N_28580,N_28269,N_28331);
xor U28581 (N_28581,N_28338,N_28290);
nor U28582 (N_28582,N_28387,N_28382);
xnor U28583 (N_28583,N_28254,N_28230);
or U28584 (N_28584,N_28228,N_28345);
nor U28585 (N_28585,N_28249,N_28314);
and U28586 (N_28586,N_28206,N_28350);
or U28587 (N_28587,N_28281,N_28343);
and U28588 (N_28588,N_28254,N_28272);
and U28589 (N_28589,N_28370,N_28221);
xnor U28590 (N_28590,N_28315,N_28369);
nor U28591 (N_28591,N_28342,N_28269);
xnor U28592 (N_28592,N_28215,N_28208);
or U28593 (N_28593,N_28324,N_28266);
and U28594 (N_28594,N_28206,N_28245);
or U28595 (N_28595,N_28304,N_28309);
xor U28596 (N_28596,N_28320,N_28338);
or U28597 (N_28597,N_28243,N_28370);
nand U28598 (N_28598,N_28318,N_28210);
nand U28599 (N_28599,N_28319,N_28285);
nand U28600 (N_28600,N_28406,N_28574);
or U28601 (N_28601,N_28421,N_28502);
or U28602 (N_28602,N_28419,N_28469);
xor U28603 (N_28603,N_28577,N_28534);
nor U28604 (N_28604,N_28438,N_28448);
or U28605 (N_28605,N_28560,N_28578);
nor U28606 (N_28606,N_28441,N_28517);
and U28607 (N_28607,N_28532,N_28556);
nor U28608 (N_28608,N_28597,N_28535);
nand U28609 (N_28609,N_28423,N_28417);
or U28610 (N_28610,N_28473,N_28480);
xnor U28611 (N_28611,N_28458,N_28564);
and U28612 (N_28612,N_28568,N_28450);
xnor U28613 (N_28613,N_28401,N_28414);
and U28614 (N_28614,N_28454,N_28452);
nor U28615 (N_28615,N_28554,N_28595);
and U28616 (N_28616,N_28413,N_28569);
xnor U28617 (N_28617,N_28516,N_28487);
or U28618 (N_28618,N_28466,N_28529);
and U28619 (N_28619,N_28429,N_28476);
or U28620 (N_28620,N_28507,N_28445);
xor U28621 (N_28621,N_28494,N_28424);
nor U28622 (N_28622,N_28579,N_28477);
nand U28623 (N_28623,N_28462,N_28582);
nand U28624 (N_28624,N_28489,N_28474);
nor U28625 (N_28625,N_28433,N_28530);
nor U28626 (N_28626,N_28425,N_28478);
nor U28627 (N_28627,N_28519,N_28485);
xnor U28628 (N_28628,N_28408,N_28580);
nor U28629 (N_28629,N_28453,N_28594);
nand U28630 (N_28630,N_28447,N_28404);
or U28631 (N_28631,N_28465,N_28513);
nand U28632 (N_28632,N_28443,N_28427);
or U28633 (N_28633,N_28528,N_28537);
nand U28634 (N_28634,N_28540,N_28542);
nand U28635 (N_28635,N_28451,N_28561);
or U28636 (N_28636,N_28486,N_28590);
nand U28637 (N_28637,N_28434,N_28576);
or U28638 (N_28638,N_28488,N_28432);
nand U28639 (N_28639,N_28500,N_28479);
and U28640 (N_28640,N_28572,N_28400);
and U28641 (N_28641,N_28503,N_28536);
or U28642 (N_28642,N_28546,N_28410);
and U28643 (N_28643,N_28555,N_28459);
or U28644 (N_28644,N_28440,N_28557);
nand U28645 (N_28645,N_28570,N_28598);
nand U28646 (N_28646,N_28539,N_28435);
nand U28647 (N_28647,N_28510,N_28599);
and U28648 (N_28648,N_28405,N_28456);
nor U28649 (N_28649,N_28509,N_28495);
and U28650 (N_28650,N_28596,N_28512);
nand U28651 (N_28651,N_28523,N_28437);
xnor U28652 (N_28652,N_28520,N_28531);
xor U28653 (N_28653,N_28407,N_28589);
or U28654 (N_28654,N_28481,N_28547);
xnor U28655 (N_28655,N_28563,N_28403);
nor U28656 (N_28656,N_28552,N_28455);
or U28657 (N_28657,N_28591,N_28499);
nand U28658 (N_28658,N_28412,N_28428);
nand U28659 (N_28659,N_28550,N_28583);
nand U28660 (N_28660,N_28467,N_28492);
nand U28661 (N_28661,N_28426,N_28463);
nand U28662 (N_28662,N_28566,N_28562);
xor U28663 (N_28663,N_28498,N_28411);
xnor U28664 (N_28664,N_28504,N_28586);
and U28665 (N_28665,N_28422,N_28418);
or U28666 (N_28666,N_28436,N_28431);
and U28667 (N_28667,N_28565,N_28468);
xnor U28668 (N_28668,N_28548,N_28558);
or U28669 (N_28669,N_28420,N_28416);
or U28670 (N_28670,N_28439,N_28430);
xnor U28671 (N_28671,N_28541,N_28484);
nand U28672 (N_28672,N_28515,N_28573);
nand U28673 (N_28673,N_28442,N_28559);
xnor U28674 (N_28674,N_28457,N_28446);
nand U28675 (N_28675,N_28514,N_28444);
nand U28676 (N_28676,N_28508,N_28490);
nor U28677 (N_28677,N_28475,N_28415);
xnor U28678 (N_28678,N_28482,N_28491);
nor U28679 (N_28679,N_28472,N_28409);
nand U28680 (N_28680,N_28501,N_28533);
and U28681 (N_28681,N_28551,N_28575);
or U28682 (N_28682,N_28549,N_28581);
nor U28683 (N_28683,N_28493,N_28553);
nand U28684 (N_28684,N_28571,N_28585);
nand U28685 (N_28685,N_28593,N_28471);
nand U28686 (N_28686,N_28588,N_28567);
nand U28687 (N_28687,N_28527,N_28506);
and U28688 (N_28688,N_28522,N_28470);
nand U28689 (N_28689,N_28449,N_28483);
xnor U28690 (N_28690,N_28526,N_28518);
xnor U28691 (N_28691,N_28464,N_28543);
nor U28692 (N_28692,N_28505,N_28402);
xnor U28693 (N_28693,N_28511,N_28460);
nor U28694 (N_28694,N_28496,N_28538);
or U28695 (N_28695,N_28497,N_28544);
xnor U28696 (N_28696,N_28461,N_28525);
xnor U28697 (N_28697,N_28584,N_28521);
xor U28698 (N_28698,N_28592,N_28524);
xor U28699 (N_28699,N_28545,N_28587);
nor U28700 (N_28700,N_28445,N_28500);
nor U28701 (N_28701,N_28457,N_28498);
nand U28702 (N_28702,N_28461,N_28535);
xor U28703 (N_28703,N_28520,N_28480);
and U28704 (N_28704,N_28570,N_28546);
xor U28705 (N_28705,N_28582,N_28459);
or U28706 (N_28706,N_28408,N_28423);
xnor U28707 (N_28707,N_28455,N_28458);
nor U28708 (N_28708,N_28523,N_28403);
or U28709 (N_28709,N_28538,N_28495);
nor U28710 (N_28710,N_28442,N_28510);
xor U28711 (N_28711,N_28434,N_28413);
nand U28712 (N_28712,N_28490,N_28579);
and U28713 (N_28713,N_28506,N_28409);
nor U28714 (N_28714,N_28409,N_28583);
xnor U28715 (N_28715,N_28492,N_28563);
xor U28716 (N_28716,N_28559,N_28584);
nand U28717 (N_28717,N_28578,N_28554);
and U28718 (N_28718,N_28477,N_28434);
nor U28719 (N_28719,N_28474,N_28505);
nand U28720 (N_28720,N_28411,N_28566);
and U28721 (N_28721,N_28468,N_28533);
or U28722 (N_28722,N_28521,N_28495);
and U28723 (N_28723,N_28485,N_28509);
xor U28724 (N_28724,N_28473,N_28560);
or U28725 (N_28725,N_28560,N_28597);
nand U28726 (N_28726,N_28438,N_28581);
and U28727 (N_28727,N_28438,N_28538);
nor U28728 (N_28728,N_28527,N_28588);
and U28729 (N_28729,N_28501,N_28475);
and U28730 (N_28730,N_28519,N_28525);
and U28731 (N_28731,N_28466,N_28472);
xor U28732 (N_28732,N_28469,N_28480);
and U28733 (N_28733,N_28412,N_28564);
nor U28734 (N_28734,N_28543,N_28559);
nor U28735 (N_28735,N_28549,N_28478);
nand U28736 (N_28736,N_28528,N_28471);
and U28737 (N_28737,N_28488,N_28505);
xor U28738 (N_28738,N_28476,N_28427);
or U28739 (N_28739,N_28599,N_28541);
and U28740 (N_28740,N_28460,N_28412);
or U28741 (N_28741,N_28496,N_28514);
nor U28742 (N_28742,N_28593,N_28505);
nor U28743 (N_28743,N_28554,N_28460);
or U28744 (N_28744,N_28577,N_28432);
nand U28745 (N_28745,N_28427,N_28428);
or U28746 (N_28746,N_28462,N_28506);
or U28747 (N_28747,N_28489,N_28485);
and U28748 (N_28748,N_28495,N_28591);
or U28749 (N_28749,N_28548,N_28568);
or U28750 (N_28750,N_28590,N_28404);
xnor U28751 (N_28751,N_28534,N_28540);
xor U28752 (N_28752,N_28440,N_28564);
and U28753 (N_28753,N_28577,N_28560);
and U28754 (N_28754,N_28418,N_28486);
nor U28755 (N_28755,N_28515,N_28578);
nand U28756 (N_28756,N_28558,N_28480);
or U28757 (N_28757,N_28561,N_28586);
nand U28758 (N_28758,N_28560,N_28434);
nor U28759 (N_28759,N_28523,N_28521);
and U28760 (N_28760,N_28409,N_28400);
xor U28761 (N_28761,N_28472,N_28511);
nor U28762 (N_28762,N_28517,N_28429);
or U28763 (N_28763,N_28511,N_28430);
and U28764 (N_28764,N_28489,N_28437);
xnor U28765 (N_28765,N_28500,N_28545);
nor U28766 (N_28766,N_28475,N_28592);
nor U28767 (N_28767,N_28448,N_28468);
xnor U28768 (N_28768,N_28551,N_28427);
and U28769 (N_28769,N_28423,N_28449);
and U28770 (N_28770,N_28541,N_28512);
and U28771 (N_28771,N_28510,N_28525);
and U28772 (N_28772,N_28412,N_28462);
nand U28773 (N_28773,N_28537,N_28546);
or U28774 (N_28774,N_28542,N_28442);
nor U28775 (N_28775,N_28422,N_28518);
and U28776 (N_28776,N_28410,N_28521);
or U28777 (N_28777,N_28587,N_28436);
or U28778 (N_28778,N_28476,N_28521);
nor U28779 (N_28779,N_28463,N_28571);
and U28780 (N_28780,N_28480,N_28564);
nand U28781 (N_28781,N_28595,N_28416);
xor U28782 (N_28782,N_28536,N_28549);
or U28783 (N_28783,N_28492,N_28460);
nand U28784 (N_28784,N_28444,N_28567);
and U28785 (N_28785,N_28579,N_28408);
nor U28786 (N_28786,N_28490,N_28551);
nand U28787 (N_28787,N_28540,N_28479);
nor U28788 (N_28788,N_28402,N_28511);
or U28789 (N_28789,N_28460,N_28587);
and U28790 (N_28790,N_28580,N_28563);
nand U28791 (N_28791,N_28534,N_28421);
and U28792 (N_28792,N_28487,N_28436);
or U28793 (N_28793,N_28444,N_28427);
and U28794 (N_28794,N_28511,N_28593);
nor U28795 (N_28795,N_28584,N_28536);
xnor U28796 (N_28796,N_28451,N_28418);
and U28797 (N_28797,N_28426,N_28421);
xnor U28798 (N_28798,N_28447,N_28505);
and U28799 (N_28799,N_28492,N_28438);
xor U28800 (N_28800,N_28622,N_28778);
xnor U28801 (N_28801,N_28736,N_28627);
or U28802 (N_28802,N_28725,N_28638);
and U28803 (N_28803,N_28619,N_28766);
xnor U28804 (N_28804,N_28623,N_28641);
or U28805 (N_28805,N_28695,N_28747);
and U28806 (N_28806,N_28709,N_28728);
xnor U28807 (N_28807,N_28737,N_28755);
or U28808 (N_28808,N_28752,N_28779);
and U28809 (N_28809,N_28681,N_28714);
or U28810 (N_28810,N_28765,N_28699);
or U28811 (N_28811,N_28793,N_28629);
or U28812 (N_28812,N_28648,N_28729);
or U28813 (N_28813,N_28609,N_28723);
nor U28814 (N_28814,N_28760,N_28684);
xnor U28815 (N_28815,N_28751,N_28688);
or U28816 (N_28816,N_28618,N_28746);
xnor U28817 (N_28817,N_28745,N_28621);
and U28818 (N_28818,N_28718,N_28740);
nor U28819 (N_28819,N_28664,N_28775);
xnor U28820 (N_28820,N_28739,N_28724);
xor U28821 (N_28821,N_28617,N_28726);
and U28822 (N_28822,N_28659,N_28764);
xor U28823 (N_28823,N_28717,N_28720);
or U28824 (N_28824,N_28744,N_28611);
nand U28825 (N_28825,N_28690,N_28692);
or U28826 (N_28826,N_28615,N_28646);
xnor U28827 (N_28827,N_28706,N_28784);
or U28828 (N_28828,N_28620,N_28781);
xor U28829 (N_28829,N_28730,N_28658);
nor U28830 (N_28830,N_28603,N_28691);
or U28831 (N_28831,N_28694,N_28696);
nor U28832 (N_28832,N_28742,N_28642);
nor U28833 (N_28833,N_28614,N_28647);
xnor U28834 (N_28834,N_28639,N_28708);
or U28835 (N_28835,N_28673,N_28705);
and U28836 (N_28836,N_28634,N_28763);
nand U28837 (N_28837,N_28758,N_28657);
or U28838 (N_28838,N_28776,N_28704);
and U28839 (N_28839,N_28677,N_28749);
and U28840 (N_28840,N_28660,N_28687);
or U28841 (N_28841,N_28796,N_28722);
nand U28842 (N_28842,N_28783,N_28713);
or U28843 (N_28843,N_28667,N_28732);
nor U28844 (N_28844,N_28773,N_28640);
xnor U28845 (N_28845,N_28743,N_28750);
nor U28846 (N_28846,N_28666,N_28731);
xnor U28847 (N_28847,N_28649,N_28719);
nand U28848 (N_28848,N_28693,N_28756);
or U28849 (N_28849,N_28636,N_28741);
nand U28850 (N_28850,N_28715,N_28735);
and U28851 (N_28851,N_28768,N_28786);
xnor U28852 (N_28852,N_28600,N_28761);
and U28853 (N_28853,N_28656,N_28676);
nor U28854 (N_28854,N_28748,N_28663);
xnor U28855 (N_28855,N_28734,N_28661);
or U28856 (N_28856,N_28601,N_28613);
nor U28857 (N_28857,N_28702,N_28669);
or U28858 (N_28858,N_28716,N_28630);
nor U28859 (N_28859,N_28602,N_28655);
nand U28860 (N_28860,N_28777,N_28799);
xnor U28861 (N_28861,N_28754,N_28697);
nor U28862 (N_28862,N_28665,N_28712);
or U28863 (N_28863,N_28662,N_28653);
nor U28864 (N_28864,N_28678,N_28707);
nand U28865 (N_28865,N_28635,N_28733);
or U28866 (N_28866,N_28605,N_28645);
or U28867 (N_28867,N_28797,N_28604);
nand U28868 (N_28868,N_28628,N_28683);
xor U28869 (N_28869,N_28789,N_28685);
nor U28870 (N_28870,N_28769,N_28791);
nand U28871 (N_28871,N_28782,N_28686);
nand U28872 (N_28872,N_28795,N_28610);
nand U28873 (N_28873,N_28637,N_28790);
or U28874 (N_28874,N_28626,N_28767);
xnor U28875 (N_28875,N_28727,N_28780);
nand U28876 (N_28876,N_28700,N_28703);
or U28877 (N_28877,N_28682,N_28757);
and U28878 (N_28878,N_28633,N_28785);
xor U28879 (N_28879,N_28631,N_28625);
nor U28880 (N_28880,N_28643,N_28794);
nor U28881 (N_28881,N_28710,N_28632);
nor U28882 (N_28882,N_28674,N_28770);
or U28883 (N_28883,N_28650,N_28608);
xnor U28884 (N_28884,N_28672,N_28753);
xnor U28885 (N_28885,N_28644,N_28624);
nand U28886 (N_28886,N_28668,N_28607);
or U28887 (N_28887,N_28701,N_28798);
xnor U28888 (N_28888,N_28652,N_28721);
and U28889 (N_28889,N_28675,N_28689);
nand U28890 (N_28890,N_28759,N_28612);
or U28891 (N_28891,N_28774,N_28654);
xor U28892 (N_28892,N_28738,N_28762);
nand U28893 (N_28893,N_28670,N_28698);
xnor U28894 (N_28894,N_28711,N_28616);
nand U28895 (N_28895,N_28787,N_28772);
and U28896 (N_28896,N_28788,N_28680);
nor U28897 (N_28897,N_28771,N_28679);
xnor U28898 (N_28898,N_28606,N_28671);
and U28899 (N_28899,N_28651,N_28792);
nand U28900 (N_28900,N_28663,N_28712);
xnor U28901 (N_28901,N_28772,N_28744);
or U28902 (N_28902,N_28738,N_28682);
and U28903 (N_28903,N_28746,N_28794);
or U28904 (N_28904,N_28649,N_28634);
or U28905 (N_28905,N_28669,N_28716);
or U28906 (N_28906,N_28649,N_28687);
nor U28907 (N_28907,N_28641,N_28664);
nand U28908 (N_28908,N_28682,N_28717);
xnor U28909 (N_28909,N_28769,N_28792);
or U28910 (N_28910,N_28614,N_28693);
xnor U28911 (N_28911,N_28729,N_28756);
nand U28912 (N_28912,N_28660,N_28621);
xnor U28913 (N_28913,N_28700,N_28623);
nand U28914 (N_28914,N_28751,N_28740);
xnor U28915 (N_28915,N_28661,N_28610);
and U28916 (N_28916,N_28696,N_28771);
or U28917 (N_28917,N_28707,N_28684);
xor U28918 (N_28918,N_28619,N_28778);
xor U28919 (N_28919,N_28774,N_28662);
or U28920 (N_28920,N_28650,N_28739);
or U28921 (N_28921,N_28635,N_28716);
xnor U28922 (N_28922,N_28680,N_28704);
or U28923 (N_28923,N_28667,N_28682);
and U28924 (N_28924,N_28618,N_28645);
or U28925 (N_28925,N_28626,N_28712);
xor U28926 (N_28926,N_28672,N_28734);
and U28927 (N_28927,N_28706,N_28727);
nand U28928 (N_28928,N_28713,N_28750);
nor U28929 (N_28929,N_28745,N_28700);
nor U28930 (N_28930,N_28631,N_28746);
and U28931 (N_28931,N_28663,N_28625);
or U28932 (N_28932,N_28631,N_28784);
xnor U28933 (N_28933,N_28726,N_28779);
and U28934 (N_28934,N_28715,N_28774);
nor U28935 (N_28935,N_28653,N_28691);
nand U28936 (N_28936,N_28679,N_28783);
nand U28937 (N_28937,N_28785,N_28646);
and U28938 (N_28938,N_28687,N_28731);
xnor U28939 (N_28939,N_28682,N_28654);
nor U28940 (N_28940,N_28759,N_28651);
nand U28941 (N_28941,N_28772,N_28616);
xor U28942 (N_28942,N_28796,N_28771);
or U28943 (N_28943,N_28672,N_28790);
nand U28944 (N_28944,N_28643,N_28756);
xnor U28945 (N_28945,N_28700,N_28722);
nor U28946 (N_28946,N_28739,N_28779);
nand U28947 (N_28947,N_28695,N_28740);
xnor U28948 (N_28948,N_28665,N_28670);
nand U28949 (N_28949,N_28729,N_28616);
nand U28950 (N_28950,N_28795,N_28727);
nand U28951 (N_28951,N_28743,N_28644);
nor U28952 (N_28952,N_28691,N_28761);
nor U28953 (N_28953,N_28649,N_28691);
nor U28954 (N_28954,N_28690,N_28795);
xnor U28955 (N_28955,N_28626,N_28765);
and U28956 (N_28956,N_28746,N_28669);
or U28957 (N_28957,N_28741,N_28663);
xor U28958 (N_28958,N_28756,N_28610);
xor U28959 (N_28959,N_28655,N_28727);
nor U28960 (N_28960,N_28679,N_28646);
nand U28961 (N_28961,N_28705,N_28648);
nand U28962 (N_28962,N_28612,N_28668);
nand U28963 (N_28963,N_28770,N_28621);
nand U28964 (N_28964,N_28698,N_28778);
nor U28965 (N_28965,N_28788,N_28710);
and U28966 (N_28966,N_28693,N_28752);
nor U28967 (N_28967,N_28645,N_28721);
or U28968 (N_28968,N_28734,N_28623);
nand U28969 (N_28969,N_28722,N_28711);
nand U28970 (N_28970,N_28793,N_28683);
nand U28971 (N_28971,N_28736,N_28758);
nor U28972 (N_28972,N_28645,N_28789);
and U28973 (N_28973,N_28664,N_28620);
xnor U28974 (N_28974,N_28774,N_28771);
nand U28975 (N_28975,N_28622,N_28761);
and U28976 (N_28976,N_28708,N_28705);
or U28977 (N_28977,N_28791,N_28678);
nand U28978 (N_28978,N_28601,N_28752);
or U28979 (N_28979,N_28795,N_28688);
and U28980 (N_28980,N_28729,N_28798);
nor U28981 (N_28981,N_28656,N_28784);
xor U28982 (N_28982,N_28769,N_28759);
nand U28983 (N_28983,N_28763,N_28626);
xnor U28984 (N_28984,N_28726,N_28667);
or U28985 (N_28985,N_28619,N_28753);
or U28986 (N_28986,N_28700,N_28737);
and U28987 (N_28987,N_28602,N_28719);
nand U28988 (N_28988,N_28673,N_28655);
and U28989 (N_28989,N_28744,N_28790);
nand U28990 (N_28990,N_28763,N_28664);
nor U28991 (N_28991,N_28692,N_28749);
xnor U28992 (N_28992,N_28677,N_28709);
and U28993 (N_28993,N_28781,N_28738);
xnor U28994 (N_28994,N_28757,N_28633);
xor U28995 (N_28995,N_28616,N_28683);
xnor U28996 (N_28996,N_28697,N_28673);
and U28997 (N_28997,N_28713,N_28632);
xor U28998 (N_28998,N_28608,N_28729);
or U28999 (N_28999,N_28761,N_28660);
nand U29000 (N_29000,N_28875,N_28973);
nand U29001 (N_29001,N_28901,N_28820);
nand U29002 (N_29002,N_28997,N_28924);
xnor U29003 (N_29003,N_28862,N_28891);
or U29004 (N_29004,N_28941,N_28839);
xnor U29005 (N_29005,N_28966,N_28970);
nand U29006 (N_29006,N_28876,N_28934);
and U29007 (N_29007,N_28958,N_28967);
and U29008 (N_29008,N_28965,N_28897);
nand U29009 (N_29009,N_28841,N_28860);
and U29010 (N_29010,N_28998,N_28883);
nand U29011 (N_29011,N_28822,N_28936);
nor U29012 (N_29012,N_28816,N_28939);
xnor U29013 (N_29013,N_28912,N_28851);
nor U29014 (N_29014,N_28834,N_28995);
nand U29015 (N_29015,N_28856,N_28903);
nor U29016 (N_29016,N_28978,N_28893);
or U29017 (N_29017,N_28949,N_28923);
nand U29018 (N_29018,N_28869,N_28831);
and U29019 (N_29019,N_28850,N_28858);
or U29020 (N_29020,N_28947,N_28867);
nand U29021 (N_29021,N_28945,N_28805);
and U29022 (N_29022,N_28999,N_28910);
or U29023 (N_29023,N_28873,N_28812);
xor U29024 (N_29024,N_28938,N_28960);
nand U29025 (N_29025,N_28896,N_28884);
and U29026 (N_29026,N_28919,N_28861);
xor U29027 (N_29027,N_28830,N_28943);
or U29028 (N_29028,N_28866,N_28927);
xor U29029 (N_29029,N_28928,N_28962);
xnor U29030 (N_29030,N_28881,N_28833);
or U29031 (N_29031,N_28979,N_28977);
nand U29032 (N_29032,N_28802,N_28926);
xor U29033 (N_29033,N_28853,N_28889);
or U29034 (N_29034,N_28852,N_28991);
xor U29035 (N_29035,N_28905,N_28818);
and U29036 (N_29036,N_28929,N_28863);
xnor U29037 (N_29037,N_28952,N_28922);
and U29038 (N_29038,N_28835,N_28809);
or U29039 (N_29039,N_28844,N_28990);
xor U29040 (N_29040,N_28933,N_28838);
and U29041 (N_29041,N_28921,N_28932);
nand U29042 (N_29042,N_28864,N_28909);
xor U29043 (N_29043,N_28840,N_28857);
nand U29044 (N_29044,N_28946,N_28971);
xor U29045 (N_29045,N_28810,N_28907);
or U29046 (N_29046,N_28984,N_28827);
nand U29047 (N_29047,N_28837,N_28983);
or U29048 (N_29048,N_28871,N_28976);
xor U29049 (N_29049,N_28887,N_28982);
and U29050 (N_29050,N_28894,N_28854);
and U29051 (N_29051,N_28968,N_28944);
and U29052 (N_29052,N_28955,N_28888);
nor U29053 (N_29053,N_28845,N_28828);
and U29054 (N_29054,N_28956,N_28898);
nand U29055 (N_29055,N_28975,N_28855);
or U29056 (N_29056,N_28974,N_28980);
or U29057 (N_29057,N_28957,N_28914);
nand U29058 (N_29058,N_28806,N_28951);
and U29059 (N_29059,N_28925,N_28950);
or U29060 (N_29060,N_28846,N_28814);
nand U29061 (N_29061,N_28913,N_28961);
nor U29062 (N_29062,N_28904,N_28915);
nor U29063 (N_29063,N_28801,N_28972);
and U29064 (N_29064,N_28849,N_28868);
or U29065 (N_29065,N_28807,N_28821);
and U29066 (N_29066,N_28892,N_28880);
or U29067 (N_29067,N_28832,N_28902);
or U29068 (N_29068,N_28900,N_28917);
nor U29069 (N_29069,N_28877,N_28813);
or U29070 (N_29070,N_28935,N_28992);
or U29071 (N_29071,N_28899,N_28890);
or U29072 (N_29072,N_28916,N_28920);
nand U29073 (N_29073,N_28959,N_28940);
and U29074 (N_29074,N_28870,N_28836);
and U29075 (N_29075,N_28826,N_28963);
and U29076 (N_29076,N_28969,N_28815);
nand U29077 (N_29077,N_28865,N_28829);
nor U29078 (N_29078,N_28993,N_28989);
and U29079 (N_29079,N_28886,N_28874);
nor U29080 (N_29080,N_28811,N_28817);
xor U29081 (N_29081,N_28872,N_28819);
and U29082 (N_29082,N_28859,N_28808);
and U29083 (N_29083,N_28842,N_28885);
xor U29084 (N_29084,N_28882,N_28986);
nand U29085 (N_29085,N_28803,N_28964);
nor U29086 (N_29086,N_28848,N_28800);
nor U29087 (N_29087,N_28823,N_28906);
or U29088 (N_29088,N_28994,N_28911);
and U29089 (N_29089,N_28981,N_28987);
nand U29090 (N_29090,N_28918,N_28954);
nor U29091 (N_29091,N_28985,N_28847);
or U29092 (N_29092,N_28996,N_28878);
nor U29093 (N_29093,N_28908,N_28804);
xor U29094 (N_29094,N_28942,N_28824);
nand U29095 (N_29095,N_28937,N_28879);
and U29096 (N_29096,N_28953,N_28895);
xor U29097 (N_29097,N_28948,N_28931);
xnor U29098 (N_29098,N_28988,N_28843);
or U29099 (N_29099,N_28930,N_28825);
xnor U29100 (N_29100,N_28840,N_28864);
nand U29101 (N_29101,N_28957,N_28926);
nand U29102 (N_29102,N_28997,N_28899);
and U29103 (N_29103,N_28959,N_28840);
nand U29104 (N_29104,N_28948,N_28945);
nor U29105 (N_29105,N_28880,N_28825);
nand U29106 (N_29106,N_28847,N_28885);
nand U29107 (N_29107,N_28810,N_28899);
nand U29108 (N_29108,N_28969,N_28949);
nand U29109 (N_29109,N_28818,N_28911);
and U29110 (N_29110,N_28961,N_28981);
nor U29111 (N_29111,N_28889,N_28816);
xnor U29112 (N_29112,N_28951,N_28903);
nor U29113 (N_29113,N_28929,N_28961);
or U29114 (N_29114,N_28909,N_28987);
or U29115 (N_29115,N_28997,N_28803);
nor U29116 (N_29116,N_28808,N_28928);
or U29117 (N_29117,N_28864,N_28813);
nand U29118 (N_29118,N_28956,N_28810);
nand U29119 (N_29119,N_28800,N_28957);
nor U29120 (N_29120,N_28850,N_28986);
and U29121 (N_29121,N_28883,N_28949);
nand U29122 (N_29122,N_28815,N_28992);
xnor U29123 (N_29123,N_28954,N_28830);
or U29124 (N_29124,N_28883,N_28981);
nor U29125 (N_29125,N_28938,N_28956);
xnor U29126 (N_29126,N_28823,N_28942);
nand U29127 (N_29127,N_28898,N_28957);
nand U29128 (N_29128,N_28803,N_28914);
and U29129 (N_29129,N_28996,N_28923);
and U29130 (N_29130,N_28926,N_28833);
nor U29131 (N_29131,N_28891,N_28879);
nor U29132 (N_29132,N_28848,N_28842);
xor U29133 (N_29133,N_28955,N_28833);
and U29134 (N_29134,N_28909,N_28859);
nor U29135 (N_29135,N_28890,N_28984);
nor U29136 (N_29136,N_28867,N_28990);
or U29137 (N_29137,N_28834,N_28897);
nor U29138 (N_29138,N_28957,N_28925);
nor U29139 (N_29139,N_28990,N_28843);
nand U29140 (N_29140,N_28849,N_28981);
or U29141 (N_29141,N_28923,N_28887);
and U29142 (N_29142,N_28886,N_28805);
and U29143 (N_29143,N_28855,N_28817);
nand U29144 (N_29144,N_28963,N_28997);
or U29145 (N_29145,N_28891,N_28989);
nor U29146 (N_29146,N_28888,N_28852);
xor U29147 (N_29147,N_28899,N_28878);
nor U29148 (N_29148,N_28849,N_28835);
nand U29149 (N_29149,N_28805,N_28807);
or U29150 (N_29150,N_28891,N_28888);
or U29151 (N_29151,N_28839,N_28955);
nand U29152 (N_29152,N_28866,N_28847);
or U29153 (N_29153,N_28802,N_28821);
xnor U29154 (N_29154,N_28980,N_28926);
or U29155 (N_29155,N_28901,N_28824);
nor U29156 (N_29156,N_28854,N_28903);
nor U29157 (N_29157,N_28853,N_28982);
nand U29158 (N_29158,N_28888,N_28910);
and U29159 (N_29159,N_28819,N_28937);
and U29160 (N_29160,N_28896,N_28939);
xnor U29161 (N_29161,N_28838,N_28951);
or U29162 (N_29162,N_28906,N_28963);
nor U29163 (N_29163,N_28801,N_28846);
nand U29164 (N_29164,N_28914,N_28981);
xnor U29165 (N_29165,N_28961,N_28854);
nand U29166 (N_29166,N_28841,N_28994);
nand U29167 (N_29167,N_28933,N_28980);
nor U29168 (N_29168,N_28835,N_28967);
nor U29169 (N_29169,N_28848,N_28956);
and U29170 (N_29170,N_28949,N_28928);
xor U29171 (N_29171,N_28932,N_28950);
nand U29172 (N_29172,N_28956,N_28833);
xor U29173 (N_29173,N_28832,N_28947);
xor U29174 (N_29174,N_28901,N_28987);
xnor U29175 (N_29175,N_28920,N_28863);
or U29176 (N_29176,N_28849,N_28983);
and U29177 (N_29177,N_28831,N_28822);
nand U29178 (N_29178,N_28904,N_28858);
nor U29179 (N_29179,N_28851,N_28804);
nor U29180 (N_29180,N_28988,N_28994);
nand U29181 (N_29181,N_28831,N_28964);
nor U29182 (N_29182,N_28895,N_28983);
xnor U29183 (N_29183,N_28988,N_28815);
nor U29184 (N_29184,N_28803,N_28936);
nand U29185 (N_29185,N_28829,N_28860);
or U29186 (N_29186,N_28950,N_28989);
or U29187 (N_29187,N_28898,N_28851);
and U29188 (N_29188,N_28831,N_28887);
and U29189 (N_29189,N_28999,N_28811);
and U29190 (N_29190,N_28937,N_28913);
or U29191 (N_29191,N_28836,N_28893);
and U29192 (N_29192,N_28949,N_28919);
and U29193 (N_29193,N_28956,N_28949);
xor U29194 (N_29194,N_28881,N_28936);
or U29195 (N_29195,N_28900,N_28999);
or U29196 (N_29196,N_28980,N_28840);
nor U29197 (N_29197,N_28968,N_28908);
nor U29198 (N_29198,N_28866,N_28815);
and U29199 (N_29199,N_28945,N_28853);
nor U29200 (N_29200,N_29066,N_29186);
xor U29201 (N_29201,N_29086,N_29172);
xnor U29202 (N_29202,N_29149,N_29037);
xnor U29203 (N_29203,N_29015,N_29072);
xnor U29204 (N_29204,N_29009,N_29089);
or U29205 (N_29205,N_29139,N_29063);
or U29206 (N_29206,N_29061,N_29169);
nor U29207 (N_29207,N_29095,N_29020);
and U29208 (N_29208,N_29116,N_29023);
nand U29209 (N_29209,N_29014,N_29173);
nand U29210 (N_29210,N_29058,N_29168);
or U29211 (N_29211,N_29003,N_29096);
xnor U29212 (N_29212,N_29145,N_29043);
nor U29213 (N_29213,N_29137,N_29171);
nor U29214 (N_29214,N_29107,N_29065);
or U29215 (N_29215,N_29097,N_29144);
nor U29216 (N_29216,N_29184,N_29188);
or U29217 (N_29217,N_29038,N_29024);
or U29218 (N_29218,N_29099,N_29152);
nand U29219 (N_29219,N_29178,N_29133);
xor U29220 (N_29220,N_29123,N_29019);
nand U29221 (N_29221,N_29028,N_29102);
nand U29222 (N_29222,N_29070,N_29104);
nor U29223 (N_29223,N_29074,N_29045);
or U29224 (N_29224,N_29068,N_29193);
and U29225 (N_29225,N_29039,N_29140);
xor U29226 (N_29226,N_29001,N_29055);
nor U29227 (N_29227,N_29151,N_29120);
xor U29228 (N_29228,N_29180,N_29067);
and U29229 (N_29229,N_29077,N_29141);
nand U29230 (N_29230,N_29108,N_29013);
nand U29231 (N_29231,N_29158,N_29159);
xor U29232 (N_29232,N_29117,N_29142);
and U29233 (N_29233,N_29008,N_29010);
nand U29234 (N_29234,N_29194,N_29165);
nor U29235 (N_29235,N_29143,N_29093);
xnor U29236 (N_29236,N_29044,N_29121);
and U29237 (N_29237,N_29082,N_29189);
xnor U29238 (N_29238,N_29146,N_29154);
and U29239 (N_29239,N_29128,N_29012);
nor U29240 (N_29240,N_29053,N_29118);
or U29241 (N_29241,N_29105,N_29134);
nand U29242 (N_29242,N_29198,N_29035);
xor U29243 (N_29243,N_29100,N_29113);
or U29244 (N_29244,N_29106,N_29056);
and U29245 (N_29245,N_29185,N_29170);
nor U29246 (N_29246,N_29148,N_29109);
nor U29247 (N_29247,N_29060,N_29050);
or U29248 (N_29248,N_29125,N_29174);
or U29249 (N_29249,N_29182,N_29018);
xnor U29250 (N_29250,N_29085,N_29195);
or U29251 (N_29251,N_29101,N_29087);
or U29252 (N_29252,N_29111,N_29092);
nor U29253 (N_29253,N_29042,N_29199);
nand U29254 (N_29254,N_29062,N_29187);
and U29255 (N_29255,N_29091,N_29163);
or U29256 (N_29256,N_29026,N_29021);
nand U29257 (N_29257,N_29156,N_29005);
or U29258 (N_29258,N_29197,N_29132);
or U29259 (N_29259,N_29176,N_29022);
xnor U29260 (N_29260,N_29006,N_29078);
and U29261 (N_29261,N_29049,N_29161);
or U29262 (N_29262,N_29080,N_29179);
nand U29263 (N_29263,N_29160,N_29071);
xor U29264 (N_29264,N_29033,N_29183);
or U29265 (N_29265,N_29131,N_29057);
xor U29266 (N_29266,N_29094,N_29027);
xor U29267 (N_29267,N_29054,N_29147);
and U29268 (N_29268,N_29048,N_29150);
nor U29269 (N_29269,N_29047,N_29129);
nand U29270 (N_29270,N_29127,N_29059);
or U29271 (N_29271,N_29052,N_29103);
or U29272 (N_29272,N_29088,N_29031);
nand U29273 (N_29273,N_29190,N_29196);
nand U29274 (N_29274,N_29075,N_29112);
and U29275 (N_29275,N_29136,N_29076);
nor U29276 (N_29276,N_29032,N_29017);
and U29277 (N_29277,N_29046,N_29034);
nor U29278 (N_29278,N_29029,N_29162);
and U29279 (N_29279,N_29051,N_29177);
or U29280 (N_29280,N_29084,N_29167);
xor U29281 (N_29281,N_29079,N_29114);
and U29282 (N_29282,N_29122,N_29040);
nor U29283 (N_29283,N_29004,N_29157);
nor U29284 (N_29284,N_29191,N_29090);
or U29285 (N_29285,N_29025,N_29124);
nor U29286 (N_29286,N_29166,N_29000);
and U29287 (N_29287,N_29064,N_29011);
nand U29288 (N_29288,N_29036,N_29135);
and U29289 (N_29289,N_29130,N_29164);
or U29290 (N_29290,N_29138,N_29153);
and U29291 (N_29291,N_29119,N_29115);
xnor U29292 (N_29292,N_29098,N_29083);
xnor U29293 (N_29293,N_29030,N_29002);
nand U29294 (N_29294,N_29073,N_29016);
nand U29295 (N_29295,N_29175,N_29181);
xor U29296 (N_29296,N_29007,N_29041);
xnor U29297 (N_29297,N_29110,N_29069);
or U29298 (N_29298,N_29081,N_29126);
and U29299 (N_29299,N_29192,N_29155);
and U29300 (N_29300,N_29169,N_29130);
and U29301 (N_29301,N_29106,N_29080);
nand U29302 (N_29302,N_29118,N_29085);
nand U29303 (N_29303,N_29155,N_29007);
or U29304 (N_29304,N_29034,N_29195);
or U29305 (N_29305,N_29152,N_29145);
nor U29306 (N_29306,N_29069,N_29038);
nor U29307 (N_29307,N_29143,N_29115);
xor U29308 (N_29308,N_29158,N_29133);
xor U29309 (N_29309,N_29032,N_29073);
and U29310 (N_29310,N_29041,N_29080);
nor U29311 (N_29311,N_29181,N_29185);
or U29312 (N_29312,N_29011,N_29124);
nand U29313 (N_29313,N_29004,N_29117);
or U29314 (N_29314,N_29157,N_29074);
nand U29315 (N_29315,N_29019,N_29074);
xnor U29316 (N_29316,N_29091,N_29166);
nand U29317 (N_29317,N_29172,N_29057);
or U29318 (N_29318,N_29018,N_29080);
nand U29319 (N_29319,N_29116,N_29082);
and U29320 (N_29320,N_29097,N_29043);
nand U29321 (N_29321,N_29126,N_29059);
xnor U29322 (N_29322,N_29157,N_29021);
nand U29323 (N_29323,N_29195,N_29078);
xor U29324 (N_29324,N_29062,N_29080);
or U29325 (N_29325,N_29038,N_29057);
nor U29326 (N_29326,N_29049,N_29085);
and U29327 (N_29327,N_29165,N_29021);
xor U29328 (N_29328,N_29011,N_29013);
or U29329 (N_29329,N_29129,N_29172);
xor U29330 (N_29330,N_29041,N_29097);
xnor U29331 (N_29331,N_29091,N_29098);
and U29332 (N_29332,N_29136,N_29122);
nand U29333 (N_29333,N_29109,N_29105);
or U29334 (N_29334,N_29050,N_29023);
xor U29335 (N_29335,N_29092,N_29167);
and U29336 (N_29336,N_29089,N_29150);
and U29337 (N_29337,N_29173,N_29065);
xor U29338 (N_29338,N_29044,N_29067);
xor U29339 (N_29339,N_29147,N_29112);
or U29340 (N_29340,N_29167,N_29130);
or U29341 (N_29341,N_29042,N_29084);
xnor U29342 (N_29342,N_29011,N_29079);
nor U29343 (N_29343,N_29182,N_29067);
nand U29344 (N_29344,N_29014,N_29065);
and U29345 (N_29345,N_29035,N_29049);
nand U29346 (N_29346,N_29167,N_29024);
xor U29347 (N_29347,N_29139,N_29099);
xor U29348 (N_29348,N_29038,N_29124);
and U29349 (N_29349,N_29196,N_29166);
nor U29350 (N_29350,N_29132,N_29195);
and U29351 (N_29351,N_29187,N_29148);
nand U29352 (N_29352,N_29149,N_29169);
nor U29353 (N_29353,N_29045,N_29065);
xnor U29354 (N_29354,N_29168,N_29043);
or U29355 (N_29355,N_29164,N_29049);
nor U29356 (N_29356,N_29024,N_29075);
nand U29357 (N_29357,N_29122,N_29147);
nor U29358 (N_29358,N_29018,N_29191);
or U29359 (N_29359,N_29014,N_29001);
nor U29360 (N_29360,N_29028,N_29100);
xnor U29361 (N_29361,N_29183,N_29073);
or U29362 (N_29362,N_29025,N_29131);
or U29363 (N_29363,N_29041,N_29087);
nor U29364 (N_29364,N_29142,N_29182);
or U29365 (N_29365,N_29157,N_29029);
nand U29366 (N_29366,N_29156,N_29049);
and U29367 (N_29367,N_29089,N_29066);
xor U29368 (N_29368,N_29152,N_29139);
nor U29369 (N_29369,N_29030,N_29051);
xor U29370 (N_29370,N_29016,N_29010);
xnor U29371 (N_29371,N_29143,N_29007);
xor U29372 (N_29372,N_29172,N_29025);
and U29373 (N_29373,N_29075,N_29091);
xnor U29374 (N_29374,N_29103,N_29019);
and U29375 (N_29375,N_29041,N_29135);
nor U29376 (N_29376,N_29129,N_29093);
and U29377 (N_29377,N_29006,N_29011);
or U29378 (N_29378,N_29114,N_29002);
xor U29379 (N_29379,N_29198,N_29171);
nand U29380 (N_29380,N_29054,N_29039);
nor U29381 (N_29381,N_29039,N_29180);
xor U29382 (N_29382,N_29128,N_29115);
nand U29383 (N_29383,N_29046,N_29056);
or U29384 (N_29384,N_29012,N_29032);
and U29385 (N_29385,N_29024,N_29008);
nor U29386 (N_29386,N_29175,N_29048);
or U29387 (N_29387,N_29146,N_29102);
and U29388 (N_29388,N_29135,N_29165);
or U29389 (N_29389,N_29003,N_29071);
nand U29390 (N_29390,N_29190,N_29176);
nor U29391 (N_29391,N_29011,N_29021);
or U29392 (N_29392,N_29003,N_29128);
nand U29393 (N_29393,N_29109,N_29188);
nand U29394 (N_29394,N_29030,N_29064);
nor U29395 (N_29395,N_29082,N_29055);
and U29396 (N_29396,N_29194,N_29130);
and U29397 (N_29397,N_29199,N_29013);
nand U29398 (N_29398,N_29191,N_29138);
and U29399 (N_29399,N_29086,N_29116);
nor U29400 (N_29400,N_29213,N_29335);
nand U29401 (N_29401,N_29275,N_29389);
nand U29402 (N_29402,N_29274,N_29298);
xor U29403 (N_29403,N_29272,N_29289);
and U29404 (N_29404,N_29259,N_29229);
nor U29405 (N_29405,N_29283,N_29236);
xor U29406 (N_29406,N_29203,N_29214);
or U29407 (N_29407,N_29384,N_29367);
xor U29408 (N_29408,N_29372,N_29294);
or U29409 (N_29409,N_29306,N_29363);
and U29410 (N_29410,N_29221,N_29260);
nor U29411 (N_29411,N_29304,N_29208);
or U29412 (N_29412,N_29357,N_29356);
xnor U29413 (N_29413,N_29264,N_29212);
and U29414 (N_29414,N_29330,N_29353);
and U29415 (N_29415,N_29354,N_29303);
nor U29416 (N_29416,N_29322,N_29237);
nor U29417 (N_29417,N_29318,N_29320);
or U29418 (N_29418,N_29247,N_29355);
nand U29419 (N_29419,N_29211,N_29364);
xor U29420 (N_29420,N_29215,N_29328);
nand U29421 (N_29421,N_29383,N_29325);
xor U29422 (N_29422,N_29233,N_29269);
nand U29423 (N_29423,N_29337,N_29348);
xnor U29424 (N_29424,N_29216,N_29299);
nand U29425 (N_29425,N_29387,N_29321);
or U29426 (N_29426,N_29234,N_29346);
xor U29427 (N_29427,N_29315,N_29377);
xor U29428 (N_29428,N_29368,N_29201);
xor U29429 (N_29429,N_29376,N_29378);
or U29430 (N_29430,N_29265,N_29380);
and U29431 (N_29431,N_29398,N_29246);
nand U29432 (N_29432,N_29279,N_29266);
xnor U29433 (N_29433,N_29358,N_29295);
and U29434 (N_29434,N_29277,N_29336);
or U29435 (N_29435,N_29273,N_29256);
or U29436 (N_29436,N_29316,N_29224);
and U29437 (N_29437,N_29390,N_29204);
and U29438 (N_29438,N_29352,N_29301);
xor U29439 (N_29439,N_29385,N_29267);
nand U29440 (N_29440,N_29243,N_29228);
or U29441 (N_29441,N_29312,N_29332);
nand U29442 (N_29442,N_29305,N_29381);
or U29443 (N_29443,N_29382,N_29231);
nor U29444 (N_29444,N_29349,N_29341);
or U29445 (N_29445,N_29252,N_29386);
and U29446 (N_29446,N_29327,N_29226);
and U29447 (N_29447,N_29338,N_29317);
nand U29448 (N_29448,N_29209,N_29206);
xor U29449 (N_29449,N_29244,N_29388);
nand U29450 (N_29450,N_29296,N_29326);
xor U29451 (N_29451,N_29223,N_29324);
xor U29452 (N_29452,N_29205,N_29248);
and U29453 (N_29453,N_29302,N_29251);
xor U29454 (N_29454,N_29263,N_29290);
nor U29455 (N_29455,N_29394,N_29292);
nand U29456 (N_29456,N_29278,N_29255);
nand U29457 (N_29457,N_29309,N_29369);
or U29458 (N_29458,N_29361,N_29242);
nand U29459 (N_29459,N_29210,N_29297);
nor U29460 (N_29460,N_29281,N_29391);
nand U29461 (N_29461,N_29362,N_29399);
or U29462 (N_29462,N_29240,N_29287);
or U29463 (N_29463,N_29241,N_29339);
xnor U29464 (N_29464,N_29350,N_29220);
xor U29465 (N_29465,N_29397,N_29284);
or U29466 (N_29466,N_29261,N_29254);
nor U29467 (N_29467,N_29323,N_29313);
nand U29468 (N_29468,N_29239,N_29351);
xor U29469 (N_29469,N_29342,N_29393);
and U29470 (N_29470,N_29365,N_29217);
nor U29471 (N_29471,N_29291,N_29340);
or U29472 (N_29472,N_29202,N_29396);
xnor U29473 (N_29473,N_29373,N_29329);
and U29474 (N_29474,N_29276,N_29285);
xor U29475 (N_29475,N_29311,N_29257);
xor U29476 (N_29476,N_29250,N_29200);
nand U29477 (N_29477,N_29343,N_29379);
or U29478 (N_29478,N_29307,N_29227);
nand U29479 (N_29479,N_29258,N_29345);
nand U29480 (N_29480,N_29218,N_29319);
xor U29481 (N_29481,N_29366,N_29262);
nand U29482 (N_29482,N_29310,N_29268);
nor U29483 (N_29483,N_29371,N_29334);
and U29484 (N_29484,N_29225,N_29207);
and U29485 (N_29485,N_29286,N_29395);
nor U29486 (N_29486,N_29331,N_29374);
or U29487 (N_29487,N_29300,N_29232);
and U29488 (N_29488,N_29271,N_29293);
or U29489 (N_29489,N_29360,N_29375);
nor U29490 (N_29490,N_29314,N_29359);
or U29491 (N_29491,N_29280,N_29238);
nor U29492 (N_29492,N_29245,N_29253);
xnor U29493 (N_29493,N_29235,N_29347);
xnor U29494 (N_29494,N_29230,N_29282);
or U29495 (N_29495,N_29344,N_29249);
or U29496 (N_29496,N_29222,N_29270);
xnor U29497 (N_29497,N_29288,N_29333);
nor U29498 (N_29498,N_29392,N_29370);
nand U29499 (N_29499,N_29308,N_29219);
nor U29500 (N_29500,N_29387,N_29271);
nand U29501 (N_29501,N_29232,N_29307);
xor U29502 (N_29502,N_29282,N_29288);
nor U29503 (N_29503,N_29337,N_29275);
xor U29504 (N_29504,N_29318,N_29359);
xor U29505 (N_29505,N_29219,N_29248);
or U29506 (N_29506,N_29399,N_29326);
or U29507 (N_29507,N_29295,N_29309);
nor U29508 (N_29508,N_29358,N_29213);
nor U29509 (N_29509,N_29239,N_29394);
nor U29510 (N_29510,N_29305,N_29320);
nor U29511 (N_29511,N_29240,N_29319);
nand U29512 (N_29512,N_29303,N_29224);
nand U29513 (N_29513,N_29224,N_29332);
nor U29514 (N_29514,N_29242,N_29230);
or U29515 (N_29515,N_29269,N_29354);
nand U29516 (N_29516,N_29260,N_29344);
and U29517 (N_29517,N_29377,N_29264);
nor U29518 (N_29518,N_29381,N_29219);
xnor U29519 (N_29519,N_29272,N_29240);
nor U29520 (N_29520,N_29391,N_29372);
nor U29521 (N_29521,N_29239,N_29358);
nand U29522 (N_29522,N_29213,N_29227);
xnor U29523 (N_29523,N_29311,N_29371);
xnor U29524 (N_29524,N_29298,N_29318);
nand U29525 (N_29525,N_29217,N_29373);
nor U29526 (N_29526,N_29264,N_29350);
xnor U29527 (N_29527,N_29206,N_29287);
nor U29528 (N_29528,N_29226,N_29297);
nor U29529 (N_29529,N_29390,N_29371);
or U29530 (N_29530,N_29269,N_29363);
nand U29531 (N_29531,N_29337,N_29389);
nor U29532 (N_29532,N_29371,N_29233);
xor U29533 (N_29533,N_29277,N_29270);
nor U29534 (N_29534,N_29390,N_29255);
nand U29535 (N_29535,N_29290,N_29316);
nand U29536 (N_29536,N_29294,N_29304);
nand U29537 (N_29537,N_29383,N_29353);
or U29538 (N_29538,N_29204,N_29397);
xor U29539 (N_29539,N_29314,N_29240);
nand U29540 (N_29540,N_29226,N_29363);
or U29541 (N_29541,N_29209,N_29352);
nor U29542 (N_29542,N_29208,N_29378);
or U29543 (N_29543,N_29289,N_29383);
or U29544 (N_29544,N_29257,N_29252);
nand U29545 (N_29545,N_29263,N_29226);
nand U29546 (N_29546,N_29351,N_29287);
xor U29547 (N_29547,N_29351,N_29325);
nor U29548 (N_29548,N_29227,N_29216);
xnor U29549 (N_29549,N_29318,N_29385);
xnor U29550 (N_29550,N_29354,N_29205);
xor U29551 (N_29551,N_29268,N_29227);
nor U29552 (N_29552,N_29350,N_29354);
nor U29553 (N_29553,N_29308,N_29253);
or U29554 (N_29554,N_29365,N_29361);
nand U29555 (N_29555,N_29239,N_29234);
nand U29556 (N_29556,N_29369,N_29227);
nor U29557 (N_29557,N_29283,N_29373);
nand U29558 (N_29558,N_29247,N_29236);
or U29559 (N_29559,N_29219,N_29241);
or U29560 (N_29560,N_29266,N_29296);
xor U29561 (N_29561,N_29205,N_29388);
nand U29562 (N_29562,N_29332,N_29391);
nor U29563 (N_29563,N_29378,N_29334);
nand U29564 (N_29564,N_29240,N_29325);
xnor U29565 (N_29565,N_29336,N_29248);
xor U29566 (N_29566,N_29380,N_29374);
nor U29567 (N_29567,N_29217,N_29238);
nor U29568 (N_29568,N_29237,N_29394);
xor U29569 (N_29569,N_29281,N_29315);
nor U29570 (N_29570,N_29216,N_29246);
nand U29571 (N_29571,N_29318,N_29214);
or U29572 (N_29572,N_29391,N_29228);
nand U29573 (N_29573,N_29230,N_29323);
nor U29574 (N_29574,N_29299,N_29253);
xnor U29575 (N_29575,N_29213,N_29268);
xor U29576 (N_29576,N_29367,N_29323);
and U29577 (N_29577,N_29223,N_29311);
nand U29578 (N_29578,N_29326,N_29209);
xnor U29579 (N_29579,N_29361,N_29314);
nand U29580 (N_29580,N_29253,N_29267);
and U29581 (N_29581,N_29265,N_29260);
or U29582 (N_29582,N_29316,N_29350);
nand U29583 (N_29583,N_29335,N_29271);
or U29584 (N_29584,N_29227,N_29357);
or U29585 (N_29585,N_29371,N_29315);
nand U29586 (N_29586,N_29382,N_29243);
or U29587 (N_29587,N_29276,N_29399);
nand U29588 (N_29588,N_29292,N_29246);
nor U29589 (N_29589,N_29281,N_29390);
or U29590 (N_29590,N_29268,N_29338);
xnor U29591 (N_29591,N_29315,N_29277);
and U29592 (N_29592,N_29239,N_29390);
and U29593 (N_29593,N_29298,N_29371);
nand U29594 (N_29594,N_29306,N_29329);
or U29595 (N_29595,N_29249,N_29273);
nand U29596 (N_29596,N_29222,N_29350);
or U29597 (N_29597,N_29333,N_29272);
xor U29598 (N_29598,N_29266,N_29355);
and U29599 (N_29599,N_29249,N_29335);
xnor U29600 (N_29600,N_29458,N_29493);
nor U29601 (N_29601,N_29405,N_29462);
nand U29602 (N_29602,N_29571,N_29543);
or U29603 (N_29603,N_29526,N_29419);
nand U29604 (N_29604,N_29408,N_29410);
or U29605 (N_29605,N_29556,N_29426);
and U29606 (N_29606,N_29551,N_29586);
or U29607 (N_29607,N_29402,N_29530);
nand U29608 (N_29608,N_29446,N_29504);
nor U29609 (N_29609,N_29572,N_29502);
nor U29610 (N_29610,N_29582,N_29562);
nor U29611 (N_29611,N_29533,N_29517);
or U29612 (N_29612,N_29557,N_29550);
nor U29613 (N_29613,N_29421,N_29461);
xor U29614 (N_29614,N_29574,N_29479);
nor U29615 (N_29615,N_29460,N_29455);
or U29616 (N_29616,N_29538,N_29429);
or U29617 (N_29617,N_29569,N_29514);
or U29618 (N_29618,N_29585,N_29523);
and U29619 (N_29619,N_29593,N_29555);
nand U29620 (N_29620,N_29487,N_29436);
nor U29621 (N_29621,N_29466,N_29590);
and U29622 (N_29622,N_29537,N_29409);
nor U29623 (N_29623,N_29521,N_29563);
and U29624 (N_29624,N_29529,N_29592);
or U29625 (N_29625,N_29503,N_29411);
and U29626 (N_29626,N_29528,N_29474);
or U29627 (N_29627,N_29469,N_29577);
and U29628 (N_29628,N_29565,N_29475);
nand U29629 (N_29629,N_29495,N_29415);
and U29630 (N_29630,N_29536,N_29486);
nand U29631 (N_29631,N_29518,N_29567);
or U29632 (N_29632,N_29481,N_29471);
and U29633 (N_29633,N_29463,N_29428);
and U29634 (N_29634,N_29473,N_29568);
or U29635 (N_29635,N_29512,N_29454);
nor U29636 (N_29636,N_29406,N_29488);
and U29637 (N_29637,N_29423,N_29413);
xor U29638 (N_29638,N_29499,N_29430);
xor U29639 (N_29639,N_29456,N_29440);
xnor U29640 (N_29640,N_29452,N_29407);
nand U29641 (N_29641,N_29534,N_29507);
or U29642 (N_29642,N_29575,N_29438);
nand U29643 (N_29643,N_29589,N_29525);
xor U29644 (N_29644,N_29595,N_29418);
nor U29645 (N_29645,N_29596,N_29524);
or U29646 (N_29646,N_29432,N_29477);
xor U29647 (N_29647,N_29468,N_29578);
xnor U29648 (N_29648,N_29435,N_29439);
and U29649 (N_29649,N_29480,N_29425);
nor U29650 (N_29650,N_29494,N_29449);
nor U29651 (N_29651,N_29464,N_29588);
or U29652 (N_29652,N_29444,N_29580);
nand U29653 (N_29653,N_29545,N_29403);
xnor U29654 (N_29654,N_29506,N_29583);
or U29655 (N_29655,N_29520,N_29519);
nand U29656 (N_29656,N_29431,N_29482);
and U29657 (N_29657,N_29422,N_29470);
nor U29658 (N_29658,N_29465,N_29535);
xor U29659 (N_29659,N_29433,N_29416);
or U29660 (N_29660,N_29424,N_29496);
or U29661 (N_29661,N_29478,N_29591);
and U29662 (N_29662,N_29453,N_29576);
nor U29663 (N_29663,N_29544,N_29400);
or U29664 (N_29664,N_29467,N_29579);
and U29665 (N_29665,N_29552,N_29427);
nor U29666 (N_29666,N_29548,N_29566);
nor U29667 (N_29667,N_29509,N_29492);
nand U29668 (N_29668,N_29501,N_29527);
xnor U29669 (N_29669,N_29450,N_29522);
nand U29670 (N_29670,N_29597,N_29558);
or U29671 (N_29671,N_29559,N_29542);
nand U29672 (N_29672,N_29570,N_29511);
nand U29673 (N_29673,N_29434,N_29485);
and U29674 (N_29674,N_29553,N_29573);
and U29675 (N_29675,N_29546,N_29457);
nor U29676 (N_29676,N_29515,N_29516);
nand U29677 (N_29677,N_29564,N_29447);
and U29678 (N_29678,N_29505,N_29476);
xnor U29679 (N_29679,N_29500,N_29484);
and U29680 (N_29680,N_29451,N_29560);
nand U29681 (N_29681,N_29541,N_29532);
and U29682 (N_29682,N_29412,N_29510);
or U29683 (N_29683,N_29490,N_29539);
and U29684 (N_29684,N_29549,N_29584);
xnor U29685 (N_29685,N_29581,N_29459);
or U29686 (N_29686,N_29513,N_29448);
nand U29687 (N_29687,N_29442,N_29443);
nor U29688 (N_29688,N_29598,N_29404);
or U29689 (N_29689,N_29561,N_29547);
xnor U29690 (N_29690,N_29498,N_29472);
or U29691 (N_29691,N_29437,N_29489);
or U29692 (N_29692,N_29417,N_29401);
nor U29693 (N_29693,N_29554,N_29594);
or U29694 (N_29694,N_29599,N_29414);
nor U29695 (N_29695,N_29420,N_29531);
or U29696 (N_29696,N_29540,N_29441);
or U29697 (N_29697,N_29508,N_29483);
nor U29698 (N_29698,N_29491,N_29445);
nand U29699 (N_29699,N_29587,N_29497);
nand U29700 (N_29700,N_29427,N_29523);
or U29701 (N_29701,N_29533,N_29488);
xnor U29702 (N_29702,N_29537,N_29447);
nand U29703 (N_29703,N_29454,N_29590);
xor U29704 (N_29704,N_29509,N_29453);
or U29705 (N_29705,N_29592,N_29479);
xnor U29706 (N_29706,N_29587,N_29477);
xnor U29707 (N_29707,N_29505,N_29525);
and U29708 (N_29708,N_29556,N_29547);
nand U29709 (N_29709,N_29570,N_29466);
nand U29710 (N_29710,N_29588,N_29412);
xor U29711 (N_29711,N_29531,N_29568);
xnor U29712 (N_29712,N_29535,N_29493);
nor U29713 (N_29713,N_29412,N_29503);
and U29714 (N_29714,N_29576,N_29546);
xnor U29715 (N_29715,N_29510,N_29518);
nand U29716 (N_29716,N_29520,N_29521);
or U29717 (N_29717,N_29416,N_29422);
xor U29718 (N_29718,N_29520,N_29514);
nor U29719 (N_29719,N_29582,N_29523);
nand U29720 (N_29720,N_29409,N_29467);
xnor U29721 (N_29721,N_29416,N_29548);
and U29722 (N_29722,N_29502,N_29462);
xnor U29723 (N_29723,N_29476,N_29454);
nand U29724 (N_29724,N_29443,N_29532);
or U29725 (N_29725,N_29419,N_29536);
nand U29726 (N_29726,N_29435,N_29454);
and U29727 (N_29727,N_29414,N_29498);
nor U29728 (N_29728,N_29448,N_29430);
and U29729 (N_29729,N_29438,N_29498);
and U29730 (N_29730,N_29500,N_29571);
and U29731 (N_29731,N_29582,N_29571);
and U29732 (N_29732,N_29483,N_29518);
or U29733 (N_29733,N_29519,N_29413);
nand U29734 (N_29734,N_29467,N_29400);
nor U29735 (N_29735,N_29566,N_29488);
or U29736 (N_29736,N_29442,N_29535);
xnor U29737 (N_29737,N_29512,N_29435);
nor U29738 (N_29738,N_29474,N_29410);
nand U29739 (N_29739,N_29510,N_29478);
xor U29740 (N_29740,N_29482,N_29484);
or U29741 (N_29741,N_29413,N_29404);
and U29742 (N_29742,N_29540,N_29503);
nand U29743 (N_29743,N_29498,N_29445);
or U29744 (N_29744,N_29419,N_29493);
nor U29745 (N_29745,N_29439,N_29500);
nor U29746 (N_29746,N_29410,N_29576);
nand U29747 (N_29747,N_29471,N_29433);
or U29748 (N_29748,N_29546,N_29575);
xnor U29749 (N_29749,N_29567,N_29495);
and U29750 (N_29750,N_29450,N_29587);
nor U29751 (N_29751,N_29559,N_29422);
nor U29752 (N_29752,N_29519,N_29471);
and U29753 (N_29753,N_29554,N_29491);
or U29754 (N_29754,N_29474,N_29590);
or U29755 (N_29755,N_29456,N_29482);
xnor U29756 (N_29756,N_29488,N_29499);
and U29757 (N_29757,N_29552,N_29423);
nand U29758 (N_29758,N_29548,N_29452);
and U29759 (N_29759,N_29455,N_29451);
and U29760 (N_29760,N_29421,N_29482);
xnor U29761 (N_29761,N_29528,N_29524);
or U29762 (N_29762,N_29407,N_29494);
nand U29763 (N_29763,N_29583,N_29519);
xor U29764 (N_29764,N_29413,N_29498);
nand U29765 (N_29765,N_29541,N_29409);
xor U29766 (N_29766,N_29559,N_29557);
nand U29767 (N_29767,N_29591,N_29524);
and U29768 (N_29768,N_29557,N_29537);
nor U29769 (N_29769,N_29466,N_29554);
nor U29770 (N_29770,N_29513,N_29556);
nor U29771 (N_29771,N_29524,N_29413);
xor U29772 (N_29772,N_29440,N_29454);
xor U29773 (N_29773,N_29437,N_29494);
or U29774 (N_29774,N_29405,N_29499);
or U29775 (N_29775,N_29456,N_29539);
or U29776 (N_29776,N_29499,N_29536);
nor U29777 (N_29777,N_29424,N_29581);
or U29778 (N_29778,N_29455,N_29494);
xor U29779 (N_29779,N_29435,N_29526);
or U29780 (N_29780,N_29404,N_29472);
and U29781 (N_29781,N_29425,N_29534);
or U29782 (N_29782,N_29557,N_29530);
nor U29783 (N_29783,N_29529,N_29426);
and U29784 (N_29784,N_29492,N_29486);
or U29785 (N_29785,N_29495,N_29528);
nand U29786 (N_29786,N_29560,N_29561);
and U29787 (N_29787,N_29444,N_29512);
and U29788 (N_29788,N_29457,N_29469);
nand U29789 (N_29789,N_29477,N_29580);
nor U29790 (N_29790,N_29477,N_29407);
and U29791 (N_29791,N_29443,N_29475);
xor U29792 (N_29792,N_29521,N_29447);
xor U29793 (N_29793,N_29581,N_29432);
or U29794 (N_29794,N_29553,N_29501);
nand U29795 (N_29795,N_29531,N_29503);
xnor U29796 (N_29796,N_29432,N_29500);
xor U29797 (N_29797,N_29443,N_29458);
nand U29798 (N_29798,N_29434,N_29444);
nor U29799 (N_29799,N_29557,N_29463);
or U29800 (N_29800,N_29721,N_29787);
nor U29801 (N_29801,N_29651,N_29785);
or U29802 (N_29802,N_29636,N_29676);
nor U29803 (N_29803,N_29729,N_29699);
nand U29804 (N_29804,N_29748,N_29642);
and U29805 (N_29805,N_29774,N_29775);
xor U29806 (N_29806,N_29627,N_29616);
nor U29807 (N_29807,N_29684,N_29706);
and U29808 (N_29808,N_29796,N_29660);
or U29809 (N_29809,N_29694,N_29618);
and U29810 (N_29810,N_29714,N_29662);
nor U29811 (N_29811,N_29665,N_29621);
nor U29812 (N_29812,N_29711,N_29666);
or U29813 (N_29813,N_29615,N_29794);
or U29814 (N_29814,N_29623,N_29613);
or U29815 (N_29815,N_29743,N_29768);
nand U29816 (N_29816,N_29739,N_29722);
and U29817 (N_29817,N_29709,N_29674);
or U29818 (N_29818,N_29737,N_29695);
or U29819 (N_29819,N_29663,N_29780);
and U29820 (N_29820,N_29776,N_29765);
nor U29821 (N_29821,N_29608,N_29769);
nand U29822 (N_29822,N_29773,N_29688);
or U29823 (N_29823,N_29726,N_29647);
xor U29824 (N_29824,N_29679,N_29798);
nand U29825 (N_29825,N_29777,N_29669);
nor U29826 (N_29826,N_29718,N_29710);
nor U29827 (N_29827,N_29734,N_29788);
and U29828 (N_29828,N_29650,N_29609);
or U29829 (N_29829,N_29719,N_29640);
and U29830 (N_29830,N_29746,N_29781);
nor U29831 (N_29831,N_29644,N_29703);
or U29832 (N_29832,N_29759,N_29753);
nor U29833 (N_29833,N_29762,N_29620);
xnor U29834 (N_29834,N_29659,N_29655);
and U29835 (N_29835,N_29637,N_29723);
and U29836 (N_29836,N_29632,N_29680);
or U29837 (N_29837,N_29678,N_29728);
nor U29838 (N_29838,N_29742,N_29603);
nand U29839 (N_29839,N_29772,N_29630);
nand U29840 (N_29840,N_29735,N_29779);
xnor U29841 (N_29841,N_29664,N_29646);
nor U29842 (N_29842,N_29605,N_29799);
nor U29843 (N_29843,N_29629,N_29732);
xor U29844 (N_29844,N_29658,N_29771);
or U29845 (N_29845,N_29782,N_29705);
or U29846 (N_29846,N_29764,N_29653);
and U29847 (N_29847,N_29625,N_29745);
nand U29848 (N_29848,N_29791,N_29795);
xor U29849 (N_29849,N_29724,N_29626);
xor U29850 (N_29850,N_29789,N_29715);
or U29851 (N_29851,N_29740,N_29687);
xnor U29852 (N_29852,N_29610,N_29778);
and U29853 (N_29853,N_29634,N_29786);
nor U29854 (N_29854,N_29704,N_29619);
xor U29855 (N_29855,N_29631,N_29741);
and U29856 (N_29856,N_29783,N_29792);
nand U29857 (N_29857,N_29677,N_29793);
nand U29858 (N_29858,N_29693,N_29763);
and U29859 (N_29859,N_29717,N_29602);
nand U29860 (N_29860,N_29600,N_29738);
nand U29861 (N_29861,N_29643,N_29720);
and U29862 (N_29862,N_29766,N_29749);
xor U29863 (N_29863,N_29635,N_29667);
nor U29864 (N_29864,N_29639,N_29790);
nand U29865 (N_29865,N_29784,N_29601);
nand U29866 (N_29866,N_29713,N_29606);
or U29867 (N_29867,N_29654,N_29611);
nor U29868 (N_29868,N_29645,N_29657);
nand U29869 (N_29869,N_29731,N_29638);
or U29870 (N_29870,N_29641,N_29733);
or U29871 (N_29871,N_29698,N_29708);
or U29872 (N_29872,N_29624,N_29770);
or U29873 (N_29873,N_29673,N_29712);
and U29874 (N_29874,N_29716,N_29672);
and U29875 (N_29875,N_29685,N_29661);
and U29876 (N_29876,N_29755,N_29683);
or U29877 (N_29877,N_29707,N_29752);
or U29878 (N_29878,N_29689,N_29736);
and U29879 (N_29879,N_29700,N_29686);
nor U29880 (N_29880,N_29690,N_29670);
xor U29881 (N_29881,N_29758,N_29696);
xor U29882 (N_29882,N_29730,N_29604);
nand U29883 (N_29883,N_29668,N_29747);
or U29884 (N_29884,N_29751,N_29628);
xor U29885 (N_29885,N_29607,N_29725);
or U29886 (N_29886,N_29682,N_29744);
or U29887 (N_29887,N_29649,N_29691);
or U29888 (N_29888,N_29692,N_29675);
nor U29889 (N_29889,N_29701,N_29633);
or U29890 (N_29890,N_29617,N_29756);
and U29891 (N_29891,N_29681,N_29648);
or U29892 (N_29892,N_29614,N_29767);
xnor U29893 (N_29893,N_29656,N_29761);
xor U29894 (N_29894,N_29671,N_29612);
or U29895 (N_29895,N_29760,N_29754);
or U29896 (N_29896,N_29702,N_29697);
and U29897 (N_29897,N_29757,N_29727);
xnor U29898 (N_29898,N_29622,N_29750);
and U29899 (N_29899,N_29652,N_29797);
xor U29900 (N_29900,N_29790,N_29671);
and U29901 (N_29901,N_29676,N_29644);
nand U29902 (N_29902,N_29765,N_29746);
or U29903 (N_29903,N_29758,N_29757);
nor U29904 (N_29904,N_29657,N_29792);
xnor U29905 (N_29905,N_29687,N_29647);
xor U29906 (N_29906,N_29711,N_29614);
xor U29907 (N_29907,N_29692,N_29777);
and U29908 (N_29908,N_29671,N_29601);
or U29909 (N_29909,N_29627,N_29788);
and U29910 (N_29910,N_29779,N_29644);
or U29911 (N_29911,N_29641,N_29702);
nor U29912 (N_29912,N_29676,N_29764);
nand U29913 (N_29913,N_29629,N_29719);
or U29914 (N_29914,N_29634,N_29728);
and U29915 (N_29915,N_29772,N_29624);
or U29916 (N_29916,N_29636,N_29628);
nand U29917 (N_29917,N_29633,N_29741);
nand U29918 (N_29918,N_29644,N_29777);
or U29919 (N_29919,N_29607,N_29645);
xor U29920 (N_29920,N_29738,N_29668);
nor U29921 (N_29921,N_29741,N_29610);
or U29922 (N_29922,N_29632,N_29736);
nor U29923 (N_29923,N_29686,N_29640);
and U29924 (N_29924,N_29713,N_29783);
xnor U29925 (N_29925,N_29673,N_29691);
and U29926 (N_29926,N_29758,N_29775);
nand U29927 (N_29927,N_29786,N_29749);
and U29928 (N_29928,N_29738,N_29633);
xnor U29929 (N_29929,N_29754,N_29669);
nor U29930 (N_29930,N_29780,N_29721);
xnor U29931 (N_29931,N_29710,N_29698);
or U29932 (N_29932,N_29703,N_29735);
nor U29933 (N_29933,N_29633,N_29789);
xnor U29934 (N_29934,N_29652,N_29765);
xor U29935 (N_29935,N_29764,N_29757);
or U29936 (N_29936,N_29651,N_29677);
and U29937 (N_29937,N_29719,N_29657);
or U29938 (N_29938,N_29615,N_29763);
nor U29939 (N_29939,N_29733,N_29655);
xor U29940 (N_29940,N_29705,N_29652);
nand U29941 (N_29941,N_29750,N_29774);
and U29942 (N_29942,N_29617,N_29689);
and U29943 (N_29943,N_29751,N_29633);
xnor U29944 (N_29944,N_29732,N_29759);
or U29945 (N_29945,N_29724,N_29677);
and U29946 (N_29946,N_29643,N_29614);
or U29947 (N_29947,N_29604,N_29685);
nor U29948 (N_29948,N_29670,N_29668);
nor U29949 (N_29949,N_29693,N_29714);
xnor U29950 (N_29950,N_29639,N_29750);
or U29951 (N_29951,N_29762,N_29790);
nor U29952 (N_29952,N_29777,N_29694);
nand U29953 (N_29953,N_29690,N_29641);
xor U29954 (N_29954,N_29661,N_29756);
nor U29955 (N_29955,N_29632,N_29690);
nand U29956 (N_29956,N_29759,N_29645);
or U29957 (N_29957,N_29752,N_29775);
xnor U29958 (N_29958,N_29630,N_29778);
nand U29959 (N_29959,N_29762,N_29768);
and U29960 (N_29960,N_29685,N_29683);
nand U29961 (N_29961,N_29738,N_29678);
or U29962 (N_29962,N_29691,N_29618);
and U29963 (N_29963,N_29797,N_29769);
and U29964 (N_29964,N_29768,N_29610);
xnor U29965 (N_29965,N_29610,N_29651);
and U29966 (N_29966,N_29602,N_29657);
or U29967 (N_29967,N_29721,N_29744);
xor U29968 (N_29968,N_29685,N_29777);
xor U29969 (N_29969,N_29735,N_29666);
or U29970 (N_29970,N_29744,N_29722);
nand U29971 (N_29971,N_29604,N_29615);
nand U29972 (N_29972,N_29638,N_29626);
nor U29973 (N_29973,N_29641,N_29630);
or U29974 (N_29974,N_29662,N_29784);
nor U29975 (N_29975,N_29702,N_29615);
or U29976 (N_29976,N_29632,N_29639);
nor U29977 (N_29977,N_29701,N_29759);
xor U29978 (N_29978,N_29797,N_29641);
or U29979 (N_29979,N_29755,N_29752);
xnor U29980 (N_29980,N_29711,N_29639);
or U29981 (N_29981,N_29659,N_29730);
and U29982 (N_29982,N_29630,N_29656);
nor U29983 (N_29983,N_29656,N_29606);
xnor U29984 (N_29984,N_29722,N_29611);
and U29985 (N_29985,N_29635,N_29639);
and U29986 (N_29986,N_29761,N_29745);
xor U29987 (N_29987,N_29721,N_29606);
nor U29988 (N_29988,N_29728,N_29791);
and U29989 (N_29989,N_29714,N_29635);
or U29990 (N_29990,N_29783,N_29680);
nand U29991 (N_29991,N_29754,N_29788);
and U29992 (N_29992,N_29665,N_29716);
nor U29993 (N_29993,N_29705,N_29664);
and U29994 (N_29994,N_29682,N_29619);
nand U29995 (N_29995,N_29795,N_29713);
and U29996 (N_29996,N_29678,N_29626);
or U29997 (N_29997,N_29767,N_29797);
nor U29998 (N_29998,N_29783,N_29681);
nand U29999 (N_29999,N_29698,N_29643);
nor UO_0 (O_0,N_29970,N_29894);
and UO_1 (O_1,N_29892,N_29932);
xor UO_2 (O_2,N_29985,N_29919);
xnor UO_3 (O_3,N_29931,N_29975);
and UO_4 (O_4,N_29935,N_29829);
or UO_5 (O_5,N_29902,N_29821);
xor UO_6 (O_6,N_29890,N_29838);
xor UO_7 (O_7,N_29895,N_29836);
and UO_8 (O_8,N_29904,N_29860);
nor UO_9 (O_9,N_29954,N_29965);
xor UO_10 (O_10,N_29880,N_29847);
xor UO_11 (O_11,N_29943,N_29853);
nand UO_12 (O_12,N_29807,N_29855);
or UO_13 (O_13,N_29955,N_29837);
or UO_14 (O_14,N_29842,N_29827);
and UO_15 (O_15,N_29803,N_29924);
nand UO_16 (O_16,N_29898,N_29800);
xor UO_17 (O_17,N_29804,N_29858);
or UO_18 (O_18,N_29964,N_29945);
nand UO_19 (O_19,N_29967,N_29949);
xnor UO_20 (O_20,N_29813,N_29960);
nor UO_21 (O_21,N_29977,N_29899);
and UO_22 (O_22,N_29962,N_29887);
nor UO_23 (O_23,N_29815,N_29879);
nor UO_24 (O_24,N_29885,N_29817);
and UO_25 (O_25,N_29849,N_29979);
and UO_26 (O_26,N_29997,N_29802);
nor UO_27 (O_27,N_29988,N_29835);
and UO_28 (O_28,N_29917,N_29848);
nor UO_29 (O_29,N_29995,N_29882);
xor UO_30 (O_30,N_29875,N_29929);
nor UO_31 (O_31,N_29822,N_29870);
and UO_32 (O_32,N_29959,N_29814);
nor UO_33 (O_33,N_29994,N_29871);
or UO_34 (O_34,N_29972,N_29812);
nor UO_35 (O_35,N_29884,N_29891);
nand UO_36 (O_36,N_29819,N_29856);
nor UO_37 (O_37,N_29886,N_29996);
and UO_38 (O_38,N_29916,N_29841);
or UO_39 (O_39,N_29862,N_29991);
and UO_40 (O_40,N_29944,N_29881);
and UO_41 (O_41,N_29947,N_29930);
nor UO_42 (O_42,N_29986,N_29911);
and UO_43 (O_43,N_29914,N_29978);
nand UO_44 (O_44,N_29820,N_29832);
or UO_45 (O_45,N_29920,N_29983);
or UO_46 (O_46,N_29874,N_29901);
nor UO_47 (O_47,N_29867,N_29981);
xor UO_48 (O_48,N_29912,N_29951);
xor UO_49 (O_49,N_29888,N_29844);
or UO_50 (O_50,N_29834,N_29926);
and UO_51 (O_51,N_29907,N_29825);
xor UO_52 (O_52,N_29843,N_29968);
and UO_53 (O_53,N_29811,N_29942);
or UO_54 (O_54,N_29941,N_29966);
or UO_55 (O_55,N_29897,N_29877);
or UO_56 (O_56,N_29805,N_29846);
and UO_57 (O_57,N_29845,N_29974);
nand UO_58 (O_58,N_29989,N_29973);
and UO_59 (O_59,N_29958,N_29937);
or UO_60 (O_60,N_29938,N_29831);
or UO_61 (O_61,N_29992,N_29946);
and UO_62 (O_62,N_29953,N_29840);
xor UO_63 (O_63,N_29810,N_29861);
nor UO_64 (O_64,N_29873,N_29915);
or UO_65 (O_65,N_29950,N_29852);
or UO_66 (O_66,N_29956,N_29854);
or UO_67 (O_67,N_29934,N_29823);
xor UO_68 (O_68,N_29833,N_29906);
nand UO_69 (O_69,N_29830,N_29921);
xnor UO_70 (O_70,N_29976,N_29936);
or UO_71 (O_71,N_29922,N_29857);
nor UO_72 (O_72,N_29866,N_29824);
nand UO_73 (O_73,N_29828,N_29982);
and UO_74 (O_74,N_29993,N_29903);
and UO_75 (O_75,N_29969,N_29948);
and UO_76 (O_76,N_29961,N_29933);
nor UO_77 (O_77,N_29883,N_29865);
and UO_78 (O_78,N_29918,N_29851);
xor UO_79 (O_79,N_29963,N_29927);
nor UO_80 (O_80,N_29984,N_29806);
or UO_81 (O_81,N_29987,N_29900);
nor UO_82 (O_82,N_29925,N_29878);
or UO_83 (O_83,N_29952,N_29971);
nand UO_84 (O_84,N_29940,N_29896);
nor UO_85 (O_85,N_29859,N_29998);
nand UO_86 (O_86,N_29893,N_29872);
or UO_87 (O_87,N_29909,N_29850);
nand UO_88 (O_88,N_29801,N_29869);
or UO_89 (O_89,N_29816,N_29913);
and UO_90 (O_90,N_29957,N_29868);
nand UO_91 (O_91,N_29864,N_29910);
nor UO_92 (O_92,N_29863,N_29839);
nor UO_93 (O_93,N_29939,N_29908);
xnor UO_94 (O_94,N_29808,N_29889);
nor UO_95 (O_95,N_29990,N_29980);
and UO_96 (O_96,N_29818,N_29923);
or UO_97 (O_97,N_29928,N_29999);
and UO_98 (O_98,N_29826,N_29876);
and UO_99 (O_99,N_29809,N_29905);
nand UO_100 (O_100,N_29948,N_29921);
and UO_101 (O_101,N_29800,N_29858);
and UO_102 (O_102,N_29865,N_29978);
xnor UO_103 (O_103,N_29909,N_29845);
xnor UO_104 (O_104,N_29911,N_29889);
nor UO_105 (O_105,N_29868,N_29952);
nor UO_106 (O_106,N_29815,N_29812);
nor UO_107 (O_107,N_29935,N_29884);
nand UO_108 (O_108,N_29912,N_29811);
or UO_109 (O_109,N_29873,N_29947);
nand UO_110 (O_110,N_29815,N_29921);
or UO_111 (O_111,N_29946,N_29832);
nor UO_112 (O_112,N_29907,N_29917);
and UO_113 (O_113,N_29951,N_29978);
nand UO_114 (O_114,N_29810,N_29811);
xor UO_115 (O_115,N_29965,N_29867);
nand UO_116 (O_116,N_29935,N_29881);
xor UO_117 (O_117,N_29961,N_29949);
and UO_118 (O_118,N_29977,N_29921);
or UO_119 (O_119,N_29894,N_29932);
nand UO_120 (O_120,N_29872,N_29976);
nor UO_121 (O_121,N_29923,N_29892);
or UO_122 (O_122,N_29995,N_29905);
nand UO_123 (O_123,N_29852,N_29908);
and UO_124 (O_124,N_29958,N_29817);
xnor UO_125 (O_125,N_29830,N_29891);
nor UO_126 (O_126,N_29914,N_29923);
nor UO_127 (O_127,N_29901,N_29832);
or UO_128 (O_128,N_29815,N_29810);
or UO_129 (O_129,N_29963,N_29945);
xnor UO_130 (O_130,N_29930,N_29946);
nand UO_131 (O_131,N_29902,N_29932);
nand UO_132 (O_132,N_29950,N_29837);
nor UO_133 (O_133,N_29936,N_29888);
xor UO_134 (O_134,N_29878,N_29855);
xor UO_135 (O_135,N_29817,N_29821);
xnor UO_136 (O_136,N_29875,N_29818);
nor UO_137 (O_137,N_29970,N_29841);
nor UO_138 (O_138,N_29978,N_29902);
nand UO_139 (O_139,N_29915,N_29842);
xor UO_140 (O_140,N_29875,N_29802);
or UO_141 (O_141,N_29811,N_29922);
nand UO_142 (O_142,N_29942,N_29890);
and UO_143 (O_143,N_29911,N_29979);
nor UO_144 (O_144,N_29825,N_29984);
nor UO_145 (O_145,N_29873,N_29874);
nand UO_146 (O_146,N_29979,N_29956);
nor UO_147 (O_147,N_29947,N_29863);
nor UO_148 (O_148,N_29856,N_29837);
nor UO_149 (O_149,N_29892,N_29827);
nand UO_150 (O_150,N_29919,N_29838);
and UO_151 (O_151,N_29981,N_29919);
xor UO_152 (O_152,N_29897,N_29934);
xor UO_153 (O_153,N_29833,N_29940);
and UO_154 (O_154,N_29960,N_29811);
or UO_155 (O_155,N_29875,N_29838);
and UO_156 (O_156,N_29937,N_29991);
xor UO_157 (O_157,N_29812,N_29944);
and UO_158 (O_158,N_29922,N_29868);
xnor UO_159 (O_159,N_29892,N_29822);
or UO_160 (O_160,N_29948,N_29943);
nand UO_161 (O_161,N_29946,N_29909);
nor UO_162 (O_162,N_29910,N_29895);
and UO_163 (O_163,N_29949,N_29835);
xor UO_164 (O_164,N_29949,N_29887);
and UO_165 (O_165,N_29821,N_29923);
and UO_166 (O_166,N_29835,N_29959);
and UO_167 (O_167,N_29908,N_29897);
nor UO_168 (O_168,N_29823,N_29916);
xor UO_169 (O_169,N_29802,N_29886);
nand UO_170 (O_170,N_29897,N_29826);
xor UO_171 (O_171,N_29922,N_29813);
nand UO_172 (O_172,N_29841,N_29971);
nand UO_173 (O_173,N_29846,N_29949);
nor UO_174 (O_174,N_29991,N_29951);
or UO_175 (O_175,N_29818,N_29995);
nor UO_176 (O_176,N_29962,N_29912);
nor UO_177 (O_177,N_29972,N_29805);
and UO_178 (O_178,N_29832,N_29856);
or UO_179 (O_179,N_29929,N_29812);
and UO_180 (O_180,N_29978,N_29931);
and UO_181 (O_181,N_29969,N_29900);
nand UO_182 (O_182,N_29892,N_29802);
nand UO_183 (O_183,N_29879,N_29817);
nor UO_184 (O_184,N_29955,N_29951);
xor UO_185 (O_185,N_29979,N_29873);
nor UO_186 (O_186,N_29910,N_29901);
nor UO_187 (O_187,N_29928,N_29831);
xor UO_188 (O_188,N_29888,N_29804);
and UO_189 (O_189,N_29887,N_29834);
xnor UO_190 (O_190,N_29871,N_29895);
and UO_191 (O_191,N_29859,N_29962);
nor UO_192 (O_192,N_29934,N_29893);
or UO_193 (O_193,N_29813,N_29857);
or UO_194 (O_194,N_29919,N_29835);
or UO_195 (O_195,N_29883,N_29817);
or UO_196 (O_196,N_29986,N_29942);
xnor UO_197 (O_197,N_29982,N_29807);
xor UO_198 (O_198,N_29890,N_29937);
nand UO_199 (O_199,N_29916,N_29835);
nand UO_200 (O_200,N_29901,N_29802);
xor UO_201 (O_201,N_29867,N_29956);
nand UO_202 (O_202,N_29805,N_29858);
nor UO_203 (O_203,N_29846,N_29834);
or UO_204 (O_204,N_29940,N_29834);
xor UO_205 (O_205,N_29865,N_29809);
nand UO_206 (O_206,N_29833,N_29907);
and UO_207 (O_207,N_29918,N_29919);
and UO_208 (O_208,N_29955,N_29944);
nand UO_209 (O_209,N_29800,N_29863);
or UO_210 (O_210,N_29909,N_29977);
and UO_211 (O_211,N_29903,N_29864);
nor UO_212 (O_212,N_29934,N_29840);
nor UO_213 (O_213,N_29863,N_29949);
or UO_214 (O_214,N_29859,N_29847);
nor UO_215 (O_215,N_29827,N_29824);
nor UO_216 (O_216,N_29947,N_29855);
or UO_217 (O_217,N_29974,N_29862);
xor UO_218 (O_218,N_29927,N_29887);
xnor UO_219 (O_219,N_29897,N_29947);
xnor UO_220 (O_220,N_29891,N_29992);
xnor UO_221 (O_221,N_29963,N_29859);
xnor UO_222 (O_222,N_29939,N_29878);
nand UO_223 (O_223,N_29959,N_29978);
or UO_224 (O_224,N_29913,N_29985);
xor UO_225 (O_225,N_29860,N_29828);
xnor UO_226 (O_226,N_29815,N_29973);
and UO_227 (O_227,N_29935,N_29942);
xor UO_228 (O_228,N_29978,N_29929);
and UO_229 (O_229,N_29965,N_29932);
xor UO_230 (O_230,N_29922,N_29828);
or UO_231 (O_231,N_29928,N_29841);
nand UO_232 (O_232,N_29804,N_29808);
nor UO_233 (O_233,N_29998,N_29802);
nor UO_234 (O_234,N_29885,N_29879);
nand UO_235 (O_235,N_29869,N_29947);
nor UO_236 (O_236,N_29861,N_29864);
nand UO_237 (O_237,N_29893,N_29989);
nor UO_238 (O_238,N_29905,N_29900);
xor UO_239 (O_239,N_29822,N_29986);
and UO_240 (O_240,N_29980,N_29907);
xnor UO_241 (O_241,N_29872,N_29911);
or UO_242 (O_242,N_29969,N_29805);
or UO_243 (O_243,N_29800,N_29970);
nor UO_244 (O_244,N_29925,N_29980);
or UO_245 (O_245,N_29811,N_29839);
nor UO_246 (O_246,N_29923,N_29901);
nand UO_247 (O_247,N_29812,N_29862);
and UO_248 (O_248,N_29982,N_29891);
or UO_249 (O_249,N_29883,N_29826);
or UO_250 (O_250,N_29848,N_29899);
nand UO_251 (O_251,N_29807,N_29837);
nand UO_252 (O_252,N_29848,N_29960);
nor UO_253 (O_253,N_29970,N_29921);
nand UO_254 (O_254,N_29843,N_29975);
or UO_255 (O_255,N_29985,N_29855);
and UO_256 (O_256,N_29801,N_29889);
nand UO_257 (O_257,N_29959,N_29904);
nor UO_258 (O_258,N_29806,N_29914);
nand UO_259 (O_259,N_29947,N_29883);
or UO_260 (O_260,N_29926,N_29839);
xor UO_261 (O_261,N_29801,N_29822);
and UO_262 (O_262,N_29947,N_29820);
xnor UO_263 (O_263,N_29908,N_29933);
and UO_264 (O_264,N_29836,N_29875);
xnor UO_265 (O_265,N_29884,N_29833);
or UO_266 (O_266,N_29894,N_29823);
or UO_267 (O_267,N_29904,N_29842);
nor UO_268 (O_268,N_29936,N_29811);
and UO_269 (O_269,N_29998,N_29895);
xor UO_270 (O_270,N_29988,N_29906);
xnor UO_271 (O_271,N_29876,N_29984);
and UO_272 (O_272,N_29857,N_29898);
nand UO_273 (O_273,N_29872,N_29941);
nand UO_274 (O_274,N_29871,N_29897);
and UO_275 (O_275,N_29936,N_29922);
xnor UO_276 (O_276,N_29895,N_29946);
xor UO_277 (O_277,N_29820,N_29899);
nand UO_278 (O_278,N_29861,N_29989);
and UO_279 (O_279,N_29835,N_29821);
nor UO_280 (O_280,N_29959,N_29988);
xnor UO_281 (O_281,N_29851,N_29871);
or UO_282 (O_282,N_29904,N_29810);
or UO_283 (O_283,N_29918,N_29939);
xnor UO_284 (O_284,N_29979,N_29917);
and UO_285 (O_285,N_29810,N_29812);
nor UO_286 (O_286,N_29882,N_29894);
and UO_287 (O_287,N_29839,N_29962);
nor UO_288 (O_288,N_29813,N_29953);
and UO_289 (O_289,N_29847,N_29900);
xor UO_290 (O_290,N_29937,N_29827);
nand UO_291 (O_291,N_29917,N_29883);
xor UO_292 (O_292,N_29968,N_29929);
xnor UO_293 (O_293,N_29899,N_29866);
nand UO_294 (O_294,N_29985,N_29963);
xnor UO_295 (O_295,N_29828,N_29822);
or UO_296 (O_296,N_29868,N_29850);
and UO_297 (O_297,N_29819,N_29941);
nor UO_298 (O_298,N_29978,N_29987);
or UO_299 (O_299,N_29885,N_29946);
nand UO_300 (O_300,N_29865,N_29841);
nor UO_301 (O_301,N_29980,N_29831);
nor UO_302 (O_302,N_29978,N_29934);
nand UO_303 (O_303,N_29866,N_29943);
xor UO_304 (O_304,N_29946,N_29875);
and UO_305 (O_305,N_29915,N_29864);
and UO_306 (O_306,N_29883,N_29823);
or UO_307 (O_307,N_29847,N_29841);
xnor UO_308 (O_308,N_29878,N_29813);
and UO_309 (O_309,N_29894,N_29851);
xor UO_310 (O_310,N_29961,N_29983);
or UO_311 (O_311,N_29806,N_29970);
and UO_312 (O_312,N_29881,N_29816);
and UO_313 (O_313,N_29849,N_29997);
and UO_314 (O_314,N_29965,N_29953);
nand UO_315 (O_315,N_29894,N_29892);
xor UO_316 (O_316,N_29870,N_29986);
and UO_317 (O_317,N_29823,N_29851);
nand UO_318 (O_318,N_29905,N_29810);
xnor UO_319 (O_319,N_29973,N_29926);
or UO_320 (O_320,N_29847,N_29889);
or UO_321 (O_321,N_29841,N_29903);
nor UO_322 (O_322,N_29834,N_29938);
nor UO_323 (O_323,N_29892,N_29909);
xor UO_324 (O_324,N_29940,N_29906);
nor UO_325 (O_325,N_29996,N_29952);
and UO_326 (O_326,N_29883,N_29837);
xor UO_327 (O_327,N_29854,N_29802);
nor UO_328 (O_328,N_29914,N_29814);
nand UO_329 (O_329,N_29973,N_29925);
or UO_330 (O_330,N_29890,N_29846);
nand UO_331 (O_331,N_29898,N_29961);
xor UO_332 (O_332,N_29880,N_29825);
nand UO_333 (O_333,N_29832,N_29862);
nand UO_334 (O_334,N_29946,N_29824);
and UO_335 (O_335,N_29806,N_29816);
xnor UO_336 (O_336,N_29875,N_29863);
and UO_337 (O_337,N_29861,N_29924);
xnor UO_338 (O_338,N_29800,N_29900);
xnor UO_339 (O_339,N_29916,N_29906);
and UO_340 (O_340,N_29974,N_29987);
and UO_341 (O_341,N_29901,N_29879);
or UO_342 (O_342,N_29842,N_29891);
xor UO_343 (O_343,N_29948,N_29813);
and UO_344 (O_344,N_29821,N_29803);
xnor UO_345 (O_345,N_29925,N_29993);
and UO_346 (O_346,N_29961,N_29882);
nand UO_347 (O_347,N_29877,N_29923);
nor UO_348 (O_348,N_29921,N_29873);
xor UO_349 (O_349,N_29856,N_29927);
and UO_350 (O_350,N_29824,N_29978);
and UO_351 (O_351,N_29865,N_29830);
nand UO_352 (O_352,N_29833,N_29912);
xnor UO_353 (O_353,N_29827,N_29803);
nand UO_354 (O_354,N_29832,N_29981);
and UO_355 (O_355,N_29884,N_29981);
and UO_356 (O_356,N_29805,N_29864);
nor UO_357 (O_357,N_29858,N_29911);
xor UO_358 (O_358,N_29847,N_29803);
nand UO_359 (O_359,N_29917,N_29985);
nand UO_360 (O_360,N_29935,N_29962);
or UO_361 (O_361,N_29808,N_29870);
xnor UO_362 (O_362,N_29947,N_29928);
nand UO_363 (O_363,N_29917,N_29970);
nand UO_364 (O_364,N_29950,N_29874);
nor UO_365 (O_365,N_29919,N_29994);
or UO_366 (O_366,N_29969,N_29814);
nor UO_367 (O_367,N_29950,N_29967);
xnor UO_368 (O_368,N_29984,N_29830);
or UO_369 (O_369,N_29986,N_29854);
and UO_370 (O_370,N_29977,N_29820);
or UO_371 (O_371,N_29928,N_29984);
nor UO_372 (O_372,N_29937,N_29996);
and UO_373 (O_373,N_29875,N_29877);
xnor UO_374 (O_374,N_29813,N_29927);
or UO_375 (O_375,N_29985,N_29984);
xnor UO_376 (O_376,N_29865,N_29826);
or UO_377 (O_377,N_29865,N_29900);
nor UO_378 (O_378,N_29994,N_29985);
nand UO_379 (O_379,N_29910,N_29830);
nor UO_380 (O_380,N_29965,N_29821);
nor UO_381 (O_381,N_29842,N_29929);
or UO_382 (O_382,N_29810,N_29813);
nand UO_383 (O_383,N_29979,N_29879);
nor UO_384 (O_384,N_29836,N_29987);
and UO_385 (O_385,N_29961,N_29901);
xnor UO_386 (O_386,N_29875,N_29813);
nand UO_387 (O_387,N_29889,N_29806);
or UO_388 (O_388,N_29961,N_29967);
or UO_389 (O_389,N_29958,N_29922);
nand UO_390 (O_390,N_29907,N_29894);
nand UO_391 (O_391,N_29878,N_29891);
xnor UO_392 (O_392,N_29894,N_29936);
nor UO_393 (O_393,N_29982,N_29835);
or UO_394 (O_394,N_29926,N_29884);
nor UO_395 (O_395,N_29972,N_29801);
xnor UO_396 (O_396,N_29924,N_29862);
and UO_397 (O_397,N_29853,N_29807);
nor UO_398 (O_398,N_29893,N_29882);
or UO_399 (O_399,N_29854,N_29865);
xor UO_400 (O_400,N_29990,N_29816);
nand UO_401 (O_401,N_29868,N_29960);
nand UO_402 (O_402,N_29924,N_29882);
xor UO_403 (O_403,N_29931,N_29965);
nand UO_404 (O_404,N_29876,N_29884);
nand UO_405 (O_405,N_29984,N_29946);
or UO_406 (O_406,N_29969,N_29945);
nor UO_407 (O_407,N_29897,N_29894);
nand UO_408 (O_408,N_29918,N_29966);
nor UO_409 (O_409,N_29847,N_29804);
nand UO_410 (O_410,N_29944,N_29800);
nor UO_411 (O_411,N_29930,N_29945);
and UO_412 (O_412,N_29974,N_29926);
and UO_413 (O_413,N_29924,N_29934);
nand UO_414 (O_414,N_29969,N_29917);
or UO_415 (O_415,N_29848,N_29882);
or UO_416 (O_416,N_29891,N_29831);
or UO_417 (O_417,N_29870,N_29915);
nor UO_418 (O_418,N_29817,N_29980);
nor UO_419 (O_419,N_29827,N_29959);
nor UO_420 (O_420,N_29986,N_29846);
xor UO_421 (O_421,N_29994,N_29935);
and UO_422 (O_422,N_29801,N_29936);
xnor UO_423 (O_423,N_29910,N_29918);
nor UO_424 (O_424,N_29866,N_29873);
and UO_425 (O_425,N_29944,N_29861);
and UO_426 (O_426,N_29801,N_29857);
and UO_427 (O_427,N_29987,N_29952);
and UO_428 (O_428,N_29948,N_29853);
and UO_429 (O_429,N_29941,N_29976);
nand UO_430 (O_430,N_29849,N_29933);
nand UO_431 (O_431,N_29920,N_29948);
xor UO_432 (O_432,N_29873,N_29970);
nand UO_433 (O_433,N_29970,N_29834);
and UO_434 (O_434,N_29961,N_29973);
nand UO_435 (O_435,N_29949,N_29910);
xor UO_436 (O_436,N_29852,N_29823);
or UO_437 (O_437,N_29919,N_29905);
xor UO_438 (O_438,N_29828,N_29928);
and UO_439 (O_439,N_29990,N_29962);
and UO_440 (O_440,N_29978,N_29933);
or UO_441 (O_441,N_29897,N_29984);
nor UO_442 (O_442,N_29893,N_29880);
and UO_443 (O_443,N_29814,N_29906);
xor UO_444 (O_444,N_29961,N_29813);
nor UO_445 (O_445,N_29817,N_29948);
or UO_446 (O_446,N_29895,N_29881);
and UO_447 (O_447,N_29817,N_29880);
nor UO_448 (O_448,N_29813,N_29898);
nor UO_449 (O_449,N_29929,N_29957);
nand UO_450 (O_450,N_29872,N_29852);
and UO_451 (O_451,N_29800,N_29812);
nand UO_452 (O_452,N_29921,N_29946);
and UO_453 (O_453,N_29801,N_29834);
xnor UO_454 (O_454,N_29955,N_29851);
and UO_455 (O_455,N_29983,N_29936);
and UO_456 (O_456,N_29967,N_29975);
xor UO_457 (O_457,N_29818,N_29904);
or UO_458 (O_458,N_29863,N_29841);
and UO_459 (O_459,N_29993,N_29937);
or UO_460 (O_460,N_29942,N_29857);
xnor UO_461 (O_461,N_29824,N_29932);
nor UO_462 (O_462,N_29847,N_29969);
nand UO_463 (O_463,N_29959,N_29963);
and UO_464 (O_464,N_29989,N_29913);
or UO_465 (O_465,N_29971,N_29977);
and UO_466 (O_466,N_29994,N_29848);
and UO_467 (O_467,N_29846,N_29867);
and UO_468 (O_468,N_29815,N_29924);
nor UO_469 (O_469,N_29947,N_29953);
nor UO_470 (O_470,N_29895,N_29807);
nand UO_471 (O_471,N_29873,N_29903);
or UO_472 (O_472,N_29802,N_29983);
nand UO_473 (O_473,N_29810,N_29921);
xor UO_474 (O_474,N_29943,N_29900);
xnor UO_475 (O_475,N_29895,N_29947);
nor UO_476 (O_476,N_29817,N_29842);
and UO_477 (O_477,N_29874,N_29946);
nand UO_478 (O_478,N_29976,N_29836);
nand UO_479 (O_479,N_29878,N_29958);
nor UO_480 (O_480,N_29814,N_29980);
nand UO_481 (O_481,N_29920,N_29918);
xor UO_482 (O_482,N_29811,N_29956);
nand UO_483 (O_483,N_29875,N_29979);
nand UO_484 (O_484,N_29888,N_29984);
and UO_485 (O_485,N_29934,N_29895);
and UO_486 (O_486,N_29877,N_29872);
or UO_487 (O_487,N_29817,N_29833);
nand UO_488 (O_488,N_29853,N_29800);
or UO_489 (O_489,N_29904,N_29824);
xor UO_490 (O_490,N_29863,N_29884);
or UO_491 (O_491,N_29961,N_29987);
nand UO_492 (O_492,N_29967,N_29994);
nor UO_493 (O_493,N_29844,N_29885);
and UO_494 (O_494,N_29879,N_29906);
or UO_495 (O_495,N_29990,N_29848);
nand UO_496 (O_496,N_29888,N_29865);
xnor UO_497 (O_497,N_29984,N_29913);
nor UO_498 (O_498,N_29867,N_29949);
nor UO_499 (O_499,N_29983,N_29832);
xor UO_500 (O_500,N_29916,N_29836);
xor UO_501 (O_501,N_29847,N_29891);
xnor UO_502 (O_502,N_29892,N_29999);
nor UO_503 (O_503,N_29929,N_29913);
or UO_504 (O_504,N_29999,N_29877);
and UO_505 (O_505,N_29977,N_29839);
xor UO_506 (O_506,N_29878,N_29935);
xnor UO_507 (O_507,N_29873,N_29837);
and UO_508 (O_508,N_29979,N_29961);
nand UO_509 (O_509,N_29999,N_29899);
or UO_510 (O_510,N_29808,N_29969);
or UO_511 (O_511,N_29818,N_29909);
xor UO_512 (O_512,N_29872,N_29814);
nor UO_513 (O_513,N_29899,N_29918);
nor UO_514 (O_514,N_29866,N_29858);
and UO_515 (O_515,N_29980,N_29838);
nor UO_516 (O_516,N_29959,N_29948);
xor UO_517 (O_517,N_29952,N_29890);
nand UO_518 (O_518,N_29933,N_29905);
and UO_519 (O_519,N_29972,N_29974);
and UO_520 (O_520,N_29824,N_29942);
nor UO_521 (O_521,N_29952,N_29948);
xnor UO_522 (O_522,N_29816,N_29991);
nand UO_523 (O_523,N_29894,N_29972);
nor UO_524 (O_524,N_29851,N_29990);
nor UO_525 (O_525,N_29974,N_29847);
nand UO_526 (O_526,N_29857,N_29996);
xor UO_527 (O_527,N_29857,N_29893);
xor UO_528 (O_528,N_29915,N_29923);
or UO_529 (O_529,N_29874,N_29976);
xor UO_530 (O_530,N_29814,N_29870);
xnor UO_531 (O_531,N_29817,N_29900);
nand UO_532 (O_532,N_29937,N_29826);
nor UO_533 (O_533,N_29919,N_29849);
nor UO_534 (O_534,N_29972,N_29879);
nor UO_535 (O_535,N_29806,N_29834);
or UO_536 (O_536,N_29905,N_29985);
or UO_537 (O_537,N_29963,N_29949);
nor UO_538 (O_538,N_29929,N_29947);
nand UO_539 (O_539,N_29888,N_29961);
nor UO_540 (O_540,N_29873,N_29954);
xor UO_541 (O_541,N_29859,N_29823);
nand UO_542 (O_542,N_29942,N_29895);
xor UO_543 (O_543,N_29922,N_29893);
nand UO_544 (O_544,N_29973,N_29826);
xnor UO_545 (O_545,N_29989,N_29948);
xnor UO_546 (O_546,N_29914,N_29927);
and UO_547 (O_547,N_29880,N_29981);
nand UO_548 (O_548,N_29935,N_29919);
nand UO_549 (O_549,N_29985,N_29803);
and UO_550 (O_550,N_29897,N_29974);
or UO_551 (O_551,N_29820,N_29881);
nand UO_552 (O_552,N_29959,N_29832);
xor UO_553 (O_553,N_29883,N_29849);
nor UO_554 (O_554,N_29971,N_29871);
and UO_555 (O_555,N_29956,N_29946);
and UO_556 (O_556,N_29951,N_29980);
and UO_557 (O_557,N_29992,N_29812);
nor UO_558 (O_558,N_29813,N_29984);
and UO_559 (O_559,N_29801,N_29849);
nor UO_560 (O_560,N_29975,N_29851);
nor UO_561 (O_561,N_29843,N_29909);
nand UO_562 (O_562,N_29988,N_29928);
and UO_563 (O_563,N_29929,N_29839);
or UO_564 (O_564,N_29870,N_29868);
and UO_565 (O_565,N_29825,N_29939);
xnor UO_566 (O_566,N_29878,N_29837);
xor UO_567 (O_567,N_29822,N_29965);
nor UO_568 (O_568,N_29993,N_29902);
xor UO_569 (O_569,N_29849,N_29927);
or UO_570 (O_570,N_29888,N_29915);
and UO_571 (O_571,N_29818,N_29997);
nor UO_572 (O_572,N_29802,N_29945);
xnor UO_573 (O_573,N_29897,N_29813);
or UO_574 (O_574,N_29894,N_29959);
or UO_575 (O_575,N_29936,N_29859);
xor UO_576 (O_576,N_29857,N_29817);
or UO_577 (O_577,N_29834,N_29830);
or UO_578 (O_578,N_29961,N_29812);
and UO_579 (O_579,N_29874,N_29909);
and UO_580 (O_580,N_29941,N_29999);
xnor UO_581 (O_581,N_29850,N_29996);
xor UO_582 (O_582,N_29904,N_29929);
or UO_583 (O_583,N_29852,N_29848);
nor UO_584 (O_584,N_29840,N_29800);
xor UO_585 (O_585,N_29800,N_29816);
xnor UO_586 (O_586,N_29836,N_29889);
nand UO_587 (O_587,N_29823,N_29872);
nand UO_588 (O_588,N_29943,N_29858);
or UO_589 (O_589,N_29821,N_29820);
nand UO_590 (O_590,N_29901,N_29842);
nor UO_591 (O_591,N_29950,N_29858);
nor UO_592 (O_592,N_29909,N_29978);
and UO_593 (O_593,N_29847,N_29927);
nand UO_594 (O_594,N_29844,N_29950);
and UO_595 (O_595,N_29846,N_29816);
nand UO_596 (O_596,N_29917,N_29857);
or UO_597 (O_597,N_29996,N_29888);
or UO_598 (O_598,N_29935,N_29894);
and UO_599 (O_599,N_29986,N_29951);
or UO_600 (O_600,N_29860,N_29928);
nor UO_601 (O_601,N_29842,N_29852);
nor UO_602 (O_602,N_29878,N_29957);
nand UO_603 (O_603,N_29921,N_29863);
nand UO_604 (O_604,N_29889,N_29913);
xnor UO_605 (O_605,N_29897,N_29836);
and UO_606 (O_606,N_29886,N_29986);
or UO_607 (O_607,N_29805,N_29874);
xnor UO_608 (O_608,N_29856,N_29877);
or UO_609 (O_609,N_29992,N_29818);
and UO_610 (O_610,N_29813,N_29860);
or UO_611 (O_611,N_29804,N_29829);
and UO_612 (O_612,N_29870,N_29931);
nand UO_613 (O_613,N_29861,N_29827);
nor UO_614 (O_614,N_29953,N_29848);
nor UO_615 (O_615,N_29973,N_29938);
nor UO_616 (O_616,N_29991,N_29924);
and UO_617 (O_617,N_29875,N_29974);
nor UO_618 (O_618,N_29998,N_29864);
nand UO_619 (O_619,N_29963,N_29962);
nand UO_620 (O_620,N_29905,N_29941);
nor UO_621 (O_621,N_29960,N_29842);
nand UO_622 (O_622,N_29984,N_29822);
or UO_623 (O_623,N_29944,N_29884);
or UO_624 (O_624,N_29826,N_29825);
or UO_625 (O_625,N_29903,N_29874);
or UO_626 (O_626,N_29937,N_29825);
or UO_627 (O_627,N_29892,N_29926);
or UO_628 (O_628,N_29890,N_29814);
and UO_629 (O_629,N_29943,N_29857);
nor UO_630 (O_630,N_29928,N_29863);
or UO_631 (O_631,N_29861,N_29970);
xnor UO_632 (O_632,N_29848,N_29958);
or UO_633 (O_633,N_29868,N_29892);
nand UO_634 (O_634,N_29905,N_29981);
and UO_635 (O_635,N_29928,N_29968);
and UO_636 (O_636,N_29979,N_29883);
or UO_637 (O_637,N_29912,N_29856);
and UO_638 (O_638,N_29982,N_29929);
nor UO_639 (O_639,N_29933,N_29922);
xor UO_640 (O_640,N_29976,N_29998);
nand UO_641 (O_641,N_29975,N_29990);
or UO_642 (O_642,N_29820,N_29945);
or UO_643 (O_643,N_29825,N_29947);
and UO_644 (O_644,N_29899,N_29902);
xor UO_645 (O_645,N_29866,N_29805);
and UO_646 (O_646,N_29853,N_29848);
nand UO_647 (O_647,N_29839,N_29937);
nand UO_648 (O_648,N_29909,N_29920);
nor UO_649 (O_649,N_29951,N_29809);
nor UO_650 (O_650,N_29981,N_29887);
or UO_651 (O_651,N_29839,N_29865);
xor UO_652 (O_652,N_29812,N_29983);
and UO_653 (O_653,N_29858,N_29856);
nand UO_654 (O_654,N_29893,N_29958);
and UO_655 (O_655,N_29893,N_29898);
nand UO_656 (O_656,N_29974,N_29970);
and UO_657 (O_657,N_29844,N_29808);
nand UO_658 (O_658,N_29982,N_29976);
nor UO_659 (O_659,N_29957,N_29926);
and UO_660 (O_660,N_29909,N_29817);
nor UO_661 (O_661,N_29892,N_29815);
nand UO_662 (O_662,N_29999,N_29874);
or UO_663 (O_663,N_29965,N_29829);
nand UO_664 (O_664,N_29823,N_29919);
nor UO_665 (O_665,N_29846,N_29979);
and UO_666 (O_666,N_29842,N_29908);
nand UO_667 (O_667,N_29980,N_29941);
and UO_668 (O_668,N_29996,N_29848);
or UO_669 (O_669,N_29888,N_29848);
and UO_670 (O_670,N_29864,N_29956);
or UO_671 (O_671,N_29894,N_29842);
xor UO_672 (O_672,N_29922,N_29965);
nand UO_673 (O_673,N_29859,N_29992);
nand UO_674 (O_674,N_29959,N_29952);
nor UO_675 (O_675,N_29864,N_29964);
or UO_676 (O_676,N_29946,N_29998);
nand UO_677 (O_677,N_29801,N_29924);
xor UO_678 (O_678,N_29819,N_29854);
and UO_679 (O_679,N_29899,N_29881);
or UO_680 (O_680,N_29860,N_29941);
and UO_681 (O_681,N_29858,N_29854);
or UO_682 (O_682,N_29818,N_29849);
nand UO_683 (O_683,N_29959,N_29925);
nand UO_684 (O_684,N_29807,N_29850);
nor UO_685 (O_685,N_29875,N_29895);
and UO_686 (O_686,N_29982,N_29939);
or UO_687 (O_687,N_29850,N_29849);
nor UO_688 (O_688,N_29961,N_29926);
nor UO_689 (O_689,N_29835,N_29849);
xnor UO_690 (O_690,N_29879,N_29853);
nand UO_691 (O_691,N_29933,N_29871);
xnor UO_692 (O_692,N_29849,N_29871);
or UO_693 (O_693,N_29884,N_29807);
nor UO_694 (O_694,N_29912,N_29993);
and UO_695 (O_695,N_29803,N_29842);
nor UO_696 (O_696,N_29896,N_29886);
or UO_697 (O_697,N_29860,N_29949);
and UO_698 (O_698,N_29940,N_29961);
or UO_699 (O_699,N_29833,N_29910);
nand UO_700 (O_700,N_29839,N_29828);
nor UO_701 (O_701,N_29986,N_29818);
nor UO_702 (O_702,N_29936,N_29826);
and UO_703 (O_703,N_29906,N_29819);
or UO_704 (O_704,N_29893,N_29903);
or UO_705 (O_705,N_29939,N_29932);
nand UO_706 (O_706,N_29877,N_29802);
and UO_707 (O_707,N_29972,N_29883);
or UO_708 (O_708,N_29987,N_29909);
and UO_709 (O_709,N_29868,N_29928);
nor UO_710 (O_710,N_29970,N_29804);
nor UO_711 (O_711,N_29977,N_29881);
nand UO_712 (O_712,N_29937,N_29928);
xnor UO_713 (O_713,N_29904,N_29952);
xnor UO_714 (O_714,N_29845,N_29897);
nand UO_715 (O_715,N_29929,N_29948);
nor UO_716 (O_716,N_29848,N_29952);
and UO_717 (O_717,N_29950,N_29991);
nor UO_718 (O_718,N_29902,N_29914);
and UO_719 (O_719,N_29986,N_29804);
xor UO_720 (O_720,N_29898,N_29871);
and UO_721 (O_721,N_29881,N_29951);
nand UO_722 (O_722,N_29996,N_29879);
and UO_723 (O_723,N_29804,N_29863);
nor UO_724 (O_724,N_29861,N_29888);
nand UO_725 (O_725,N_29954,N_29993);
nor UO_726 (O_726,N_29816,N_29930);
nand UO_727 (O_727,N_29906,N_29899);
and UO_728 (O_728,N_29879,N_29880);
nor UO_729 (O_729,N_29870,N_29945);
nand UO_730 (O_730,N_29824,N_29808);
nor UO_731 (O_731,N_29923,N_29908);
or UO_732 (O_732,N_29889,N_29825);
and UO_733 (O_733,N_29813,N_29942);
xor UO_734 (O_734,N_29995,N_29843);
and UO_735 (O_735,N_29947,N_29916);
xnor UO_736 (O_736,N_29886,N_29932);
and UO_737 (O_737,N_29809,N_29820);
nand UO_738 (O_738,N_29940,N_29801);
xnor UO_739 (O_739,N_29896,N_29801);
nor UO_740 (O_740,N_29982,N_29842);
nor UO_741 (O_741,N_29877,N_29977);
nand UO_742 (O_742,N_29852,N_29859);
xor UO_743 (O_743,N_29968,N_29901);
and UO_744 (O_744,N_29967,N_29859);
or UO_745 (O_745,N_29967,N_29952);
nand UO_746 (O_746,N_29880,N_29821);
or UO_747 (O_747,N_29957,N_29970);
nor UO_748 (O_748,N_29915,N_29835);
nand UO_749 (O_749,N_29816,N_29933);
and UO_750 (O_750,N_29903,N_29908);
nand UO_751 (O_751,N_29895,N_29909);
nand UO_752 (O_752,N_29803,N_29820);
nand UO_753 (O_753,N_29916,N_29813);
xor UO_754 (O_754,N_29951,N_29889);
xor UO_755 (O_755,N_29891,N_29833);
or UO_756 (O_756,N_29811,N_29906);
or UO_757 (O_757,N_29964,N_29972);
xnor UO_758 (O_758,N_29939,N_29973);
or UO_759 (O_759,N_29950,N_29824);
nand UO_760 (O_760,N_29889,N_29870);
xnor UO_761 (O_761,N_29958,N_29960);
or UO_762 (O_762,N_29810,N_29825);
xnor UO_763 (O_763,N_29908,N_29959);
and UO_764 (O_764,N_29824,N_29896);
nor UO_765 (O_765,N_29965,N_29814);
nand UO_766 (O_766,N_29898,N_29944);
and UO_767 (O_767,N_29984,N_29960);
and UO_768 (O_768,N_29883,N_29950);
xnor UO_769 (O_769,N_29878,N_29897);
and UO_770 (O_770,N_29909,N_29854);
or UO_771 (O_771,N_29905,N_29989);
nor UO_772 (O_772,N_29836,N_29820);
nor UO_773 (O_773,N_29807,N_29902);
nand UO_774 (O_774,N_29945,N_29914);
xor UO_775 (O_775,N_29926,N_29843);
nand UO_776 (O_776,N_29977,N_29967);
and UO_777 (O_777,N_29850,N_29898);
xor UO_778 (O_778,N_29932,N_29968);
nor UO_779 (O_779,N_29873,N_29989);
nor UO_780 (O_780,N_29828,N_29955);
or UO_781 (O_781,N_29966,N_29990);
or UO_782 (O_782,N_29889,N_29831);
or UO_783 (O_783,N_29921,N_29897);
and UO_784 (O_784,N_29868,N_29946);
xor UO_785 (O_785,N_29982,N_29846);
nand UO_786 (O_786,N_29815,N_29932);
xor UO_787 (O_787,N_29906,N_29989);
xnor UO_788 (O_788,N_29914,N_29817);
and UO_789 (O_789,N_29947,N_29956);
or UO_790 (O_790,N_29909,N_29835);
nand UO_791 (O_791,N_29998,N_29961);
nor UO_792 (O_792,N_29827,N_29891);
xnor UO_793 (O_793,N_29862,N_29916);
and UO_794 (O_794,N_29818,N_29945);
or UO_795 (O_795,N_29853,N_29854);
and UO_796 (O_796,N_29963,N_29941);
nor UO_797 (O_797,N_29915,N_29899);
or UO_798 (O_798,N_29800,N_29927);
nand UO_799 (O_799,N_29938,N_29874);
nand UO_800 (O_800,N_29956,N_29903);
nor UO_801 (O_801,N_29818,N_29955);
nand UO_802 (O_802,N_29974,N_29912);
nand UO_803 (O_803,N_29818,N_29937);
or UO_804 (O_804,N_29882,N_29846);
nor UO_805 (O_805,N_29824,N_29877);
nand UO_806 (O_806,N_29982,N_29849);
nand UO_807 (O_807,N_29895,N_29984);
nand UO_808 (O_808,N_29940,N_29845);
and UO_809 (O_809,N_29830,N_29831);
nor UO_810 (O_810,N_29834,N_29982);
xor UO_811 (O_811,N_29931,N_29970);
nor UO_812 (O_812,N_29903,N_29872);
xnor UO_813 (O_813,N_29806,N_29960);
xor UO_814 (O_814,N_29916,N_29816);
or UO_815 (O_815,N_29813,N_29800);
or UO_816 (O_816,N_29871,N_29920);
nand UO_817 (O_817,N_29979,N_29923);
nor UO_818 (O_818,N_29986,N_29812);
nand UO_819 (O_819,N_29816,N_29902);
nand UO_820 (O_820,N_29920,N_29965);
nand UO_821 (O_821,N_29843,N_29816);
nor UO_822 (O_822,N_29820,N_29819);
or UO_823 (O_823,N_29929,N_29951);
or UO_824 (O_824,N_29967,N_29922);
nand UO_825 (O_825,N_29954,N_29811);
xor UO_826 (O_826,N_29899,N_29838);
and UO_827 (O_827,N_29985,N_29966);
nor UO_828 (O_828,N_29802,N_29811);
xnor UO_829 (O_829,N_29882,N_29927);
nand UO_830 (O_830,N_29852,N_29917);
or UO_831 (O_831,N_29995,N_29945);
nand UO_832 (O_832,N_29819,N_29972);
xnor UO_833 (O_833,N_29806,N_29908);
and UO_834 (O_834,N_29823,N_29902);
nor UO_835 (O_835,N_29971,N_29942);
nand UO_836 (O_836,N_29874,N_29889);
nor UO_837 (O_837,N_29944,N_29832);
and UO_838 (O_838,N_29845,N_29907);
xor UO_839 (O_839,N_29928,N_29924);
xnor UO_840 (O_840,N_29941,N_29832);
or UO_841 (O_841,N_29909,N_29939);
and UO_842 (O_842,N_29839,N_29964);
nor UO_843 (O_843,N_29980,N_29806);
nor UO_844 (O_844,N_29937,N_29920);
nor UO_845 (O_845,N_29846,N_29939);
nand UO_846 (O_846,N_29878,N_29989);
xnor UO_847 (O_847,N_29965,N_29894);
and UO_848 (O_848,N_29994,N_29869);
and UO_849 (O_849,N_29819,N_29957);
or UO_850 (O_850,N_29836,N_29938);
and UO_851 (O_851,N_29951,N_29840);
xnor UO_852 (O_852,N_29967,N_29809);
nor UO_853 (O_853,N_29848,N_29870);
xnor UO_854 (O_854,N_29926,N_29952);
xor UO_855 (O_855,N_29918,N_29837);
xnor UO_856 (O_856,N_29838,N_29813);
xnor UO_857 (O_857,N_29999,N_29875);
xor UO_858 (O_858,N_29854,N_29833);
xnor UO_859 (O_859,N_29960,N_29951);
nand UO_860 (O_860,N_29891,N_29851);
or UO_861 (O_861,N_29892,N_29958);
nor UO_862 (O_862,N_29905,N_29866);
nand UO_863 (O_863,N_29832,N_29879);
nor UO_864 (O_864,N_29870,N_29852);
nor UO_865 (O_865,N_29990,N_29934);
and UO_866 (O_866,N_29883,N_29852);
and UO_867 (O_867,N_29808,N_29919);
or UO_868 (O_868,N_29860,N_29903);
nor UO_869 (O_869,N_29840,N_29892);
nor UO_870 (O_870,N_29942,N_29867);
nor UO_871 (O_871,N_29944,N_29975);
and UO_872 (O_872,N_29844,N_29930);
and UO_873 (O_873,N_29830,N_29844);
or UO_874 (O_874,N_29844,N_29845);
and UO_875 (O_875,N_29885,N_29857);
or UO_876 (O_876,N_29824,N_29829);
xnor UO_877 (O_877,N_29976,N_29833);
xnor UO_878 (O_878,N_29867,N_29947);
and UO_879 (O_879,N_29885,N_29852);
and UO_880 (O_880,N_29885,N_29993);
and UO_881 (O_881,N_29857,N_29829);
nor UO_882 (O_882,N_29888,N_29972);
or UO_883 (O_883,N_29902,N_29893);
or UO_884 (O_884,N_29868,N_29804);
and UO_885 (O_885,N_29890,N_29842);
xor UO_886 (O_886,N_29977,N_29837);
xor UO_887 (O_887,N_29976,N_29837);
or UO_888 (O_888,N_29868,N_29896);
nand UO_889 (O_889,N_29891,N_29839);
nor UO_890 (O_890,N_29946,N_29817);
nand UO_891 (O_891,N_29998,N_29813);
nand UO_892 (O_892,N_29881,N_29972);
and UO_893 (O_893,N_29931,N_29972);
or UO_894 (O_894,N_29875,N_29864);
xnor UO_895 (O_895,N_29960,N_29872);
or UO_896 (O_896,N_29971,N_29813);
or UO_897 (O_897,N_29800,N_29857);
nor UO_898 (O_898,N_29888,N_29927);
nand UO_899 (O_899,N_29929,N_29967);
and UO_900 (O_900,N_29951,N_29931);
or UO_901 (O_901,N_29955,N_29889);
xor UO_902 (O_902,N_29862,N_29996);
xnor UO_903 (O_903,N_29827,N_29988);
nand UO_904 (O_904,N_29841,N_29891);
nand UO_905 (O_905,N_29856,N_29980);
or UO_906 (O_906,N_29911,N_29919);
nor UO_907 (O_907,N_29826,N_29814);
nor UO_908 (O_908,N_29960,N_29818);
nand UO_909 (O_909,N_29832,N_29891);
nand UO_910 (O_910,N_29862,N_29836);
and UO_911 (O_911,N_29951,N_29831);
xor UO_912 (O_912,N_29941,N_29967);
and UO_913 (O_913,N_29920,N_29894);
or UO_914 (O_914,N_29939,N_29984);
xnor UO_915 (O_915,N_29959,N_29872);
xor UO_916 (O_916,N_29833,N_29815);
or UO_917 (O_917,N_29898,N_29900);
xor UO_918 (O_918,N_29999,N_29922);
xor UO_919 (O_919,N_29950,N_29906);
xor UO_920 (O_920,N_29934,N_29941);
xor UO_921 (O_921,N_29873,N_29940);
nor UO_922 (O_922,N_29833,N_29918);
and UO_923 (O_923,N_29911,N_29906);
nand UO_924 (O_924,N_29956,N_29917);
nor UO_925 (O_925,N_29931,N_29876);
and UO_926 (O_926,N_29806,N_29969);
nor UO_927 (O_927,N_29917,N_29999);
and UO_928 (O_928,N_29826,N_29823);
and UO_929 (O_929,N_29985,N_29830);
and UO_930 (O_930,N_29916,N_29994);
or UO_931 (O_931,N_29881,N_29845);
and UO_932 (O_932,N_29990,N_29830);
nor UO_933 (O_933,N_29954,N_29921);
nor UO_934 (O_934,N_29823,N_29874);
or UO_935 (O_935,N_29844,N_29919);
or UO_936 (O_936,N_29936,N_29955);
xor UO_937 (O_937,N_29890,N_29992);
or UO_938 (O_938,N_29862,N_29856);
nor UO_939 (O_939,N_29974,N_29803);
nand UO_940 (O_940,N_29843,N_29973);
and UO_941 (O_941,N_29881,N_29828);
xor UO_942 (O_942,N_29951,N_29879);
and UO_943 (O_943,N_29922,N_29902);
nor UO_944 (O_944,N_29813,N_29896);
nand UO_945 (O_945,N_29899,N_29809);
xor UO_946 (O_946,N_29843,N_29951);
nand UO_947 (O_947,N_29922,N_29920);
nor UO_948 (O_948,N_29802,N_29955);
and UO_949 (O_949,N_29856,N_29955);
nor UO_950 (O_950,N_29873,N_29896);
nor UO_951 (O_951,N_29827,N_29820);
or UO_952 (O_952,N_29970,N_29825);
xor UO_953 (O_953,N_29848,N_29854);
and UO_954 (O_954,N_29833,N_29963);
xnor UO_955 (O_955,N_29839,N_29948);
nor UO_956 (O_956,N_29934,N_29872);
nor UO_957 (O_957,N_29945,N_29976);
xor UO_958 (O_958,N_29979,N_29855);
xor UO_959 (O_959,N_29915,N_29971);
and UO_960 (O_960,N_29969,N_29954);
nor UO_961 (O_961,N_29960,N_29910);
xnor UO_962 (O_962,N_29878,N_29819);
or UO_963 (O_963,N_29805,N_29837);
nand UO_964 (O_964,N_29921,N_29885);
nor UO_965 (O_965,N_29870,N_29871);
nand UO_966 (O_966,N_29936,N_29855);
nor UO_967 (O_967,N_29802,N_29804);
nand UO_968 (O_968,N_29879,N_29921);
or UO_969 (O_969,N_29929,N_29818);
or UO_970 (O_970,N_29898,N_29845);
nand UO_971 (O_971,N_29852,N_29815);
and UO_972 (O_972,N_29945,N_29908);
nor UO_973 (O_973,N_29934,N_29869);
or UO_974 (O_974,N_29823,N_29870);
nand UO_975 (O_975,N_29841,N_29868);
nand UO_976 (O_976,N_29821,N_29857);
nand UO_977 (O_977,N_29850,N_29876);
nand UO_978 (O_978,N_29870,N_29981);
nand UO_979 (O_979,N_29917,N_29866);
nand UO_980 (O_980,N_29872,N_29947);
and UO_981 (O_981,N_29982,N_29869);
xor UO_982 (O_982,N_29901,N_29878);
nand UO_983 (O_983,N_29927,N_29805);
nand UO_984 (O_984,N_29838,N_29997);
and UO_985 (O_985,N_29817,N_29981);
nand UO_986 (O_986,N_29991,N_29931);
xnor UO_987 (O_987,N_29834,N_29955);
or UO_988 (O_988,N_29856,N_29982);
nor UO_989 (O_989,N_29998,N_29831);
xor UO_990 (O_990,N_29932,N_29946);
and UO_991 (O_991,N_29856,N_29820);
xnor UO_992 (O_992,N_29855,N_29860);
nor UO_993 (O_993,N_29864,N_29819);
or UO_994 (O_994,N_29961,N_29854);
nand UO_995 (O_995,N_29958,N_29870);
and UO_996 (O_996,N_29959,N_29810);
and UO_997 (O_997,N_29921,N_29931);
and UO_998 (O_998,N_29854,N_29996);
nand UO_999 (O_999,N_29898,N_29978);
and UO_1000 (O_1000,N_29911,N_29829);
and UO_1001 (O_1001,N_29931,N_29896);
xnor UO_1002 (O_1002,N_29813,N_29990);
xor UO_1003 (O_1003,N_29945,N_29922);
or UO_1004 (O_1004,N_29993,N_29964);
nand UO_1005 (O_1005,N_29812,N_29844);
nor UO_1006 (O_1006,N_29989,N_29966);
nand UO_1007 (O_1007,N_29961,N_29950);
nand UO_1008 (O_1008,N_29837,N_29994);
xnor UO_1009 (O_1009,N_29830,N_29997);
or UO_1010 (O_1010,N_29880,N_29976);
nor UO_1011 (O_1011,N_29818,N_29857);
xnor UO_1012 (O_1012,N_29991,N_29836);
or UO_1013 (O_1013,N_29810,N_29908);
xnor UO_1014 (O_1014,N_29889,N_29949);
nor UO_1015 (O_1015,N_29944,N_29924);
or UO_1016 (O_1016,N_29866,N_29837);
and UO_1017 (O_1017,N_29921,N_29866);
and UO_1018 (O_1018,N_29970,N_29892);
or UO_1019 (O_1019,N_29920,N_29907);
nand UO_1020 (O_1020,N_29953,N_29992);
and UO_1021 (O_1021,N_29980,N_29839);
or UO_1022 (O_1022,N_29914,N_29842);
nand UO_1023 (O_1023,N_29819,N_29920);
or UO_1024 (O_1024,N_29938,N_29994);
or UO_1025 (O_1025,N_29914,N_29895);
xor UO_1026 (O_1026,N_29954,N_29972);
and UO_1027 (O_1027,N_29999,N_29881);
nand UO_1028 (O_1028,N_29858,N_29974);
nor UO_1029 (O_1029,N_29879,N_29871);
nor UO_1030 (O_1030,N_29969,N_29801);
nand UO_1031 (O_1031,N_29934,N_29833);
and UO_1032 (O_1032,N_29902,N_29982);
xnor UO_1033 (O_1033,N_29933,N_29925);
or UO_1034 (O_1034,N_29923,N_29900);
nor UO_1035 (O_1035,N_29952,N_29986);
xor UO_1036 (O_1036,N_29824,N_29867);
nand UO_1037 (O_1037,N_29999,N_29884);
nor UO_1038 (O_1038,N_29880,N_29873);
xor UO_1039 (O_1039,N_29990,N_29999);
or UO_1040 (O_1040,N_29828,N_29888);
and UO_1041 (O_1041,N_29878,N_29922);
nand UO_1042 (O_1042,N_29932,N_29926);
and UO_1043 (O_1043,N_29921,N_29940);
and UO_1044 (O_1044,N_29829,N_29927);
and UO_1045 (O_1045,N_29873,N_29805);
nand UO_1046 (O_1046,N_29819,N_29965);
nor UO_1047 (O_1047,N_29878,N_29984);
nand UO_1048 (O_1048,N_29918,N_29887);
or UO_1049 (O_1049,N_29885,N_29904);
nor UO_1050 (O_1050,N_29958,N_29843);
or UO_1051 (O_1051,N_29844,N_29814);
and UO_1052 (O_1052,N_29951,N_29952);
nor UO_1053 (O_1053,N_29900,N_29874);
and UO_1054 (O_1054,N_29959,N_29984);
or UO_1055 (O_1055,N_29946,N_29966);
nor UO_1056 (O_1056,N_29847,N_29812);
or UO_1057 (O_1057,N_29907,N_29971);
and UO_1058 (O_1058,N_29888,N_29886);
and UO_1059 (O_1059,N_29918,N_29806);
nor UO_1060 (O_1060,N_29862,N_29952);
nand UO_1061 (O_1061,N_29939,N_29950);
or UO_1062 (O_1062,N_29909,N_29974);
and UO_1063 (O_1063,N_29863,N_29918);
or UO_1064 (O_1064,N_29893,N_29936);
and UO_1065 (O_1065,N_29816,N_29859);
nand UO_1066 (O_1066,N_29822,N_29890);
and UO_1067 (O_1067,N_29905,N_29996);
and UO_1068 (O_1068,N_29928,N_29809);
and UO_1069 (O_1069,N_29932,N_29976);
or UO_1070 (O_1070,N_29958,N_29938);
and UO_1071 (O_1071,N_29876,N_29934);
or UO_1072 (O_1072,N_29812,N_29853);
xnor UO_1073 (O_1073,N_29873,N_29820);
xnor UO_1074 (O_1074,N_29956,N_29916);
and UO_1075 (O_1075,N_29855,N_29982);
nand UO_1076 (O_1076,N_29830,N_29992);
nand UO_1077 (O_1077,N_29980,N_29819);
xnor UO_1078 (O_1078,N_29940,N_29988);
xnor UO_1079 (O_1079,N_29934,N_29800);
and UO_1080 (O_1080,N_29873,N_29815);
or UO_1081 (O_1081,N_29890,N_29819);
or UO_1082 (O_1082,N_29888,N_29945);
or UO_1083 (O_1083,N_29990,N_29955);
and UO_1084 (O_1084,N_29821,N_29848);
or UO_1085 (O_1085,N_29970,N_29870);
and UO_1086 (O_1086,N_29935,N_29893);
and UO_1087 (O_1087,N_29815,N_29884);
xnor UO_1088 (O_1088,N_29868,N_29980);
nor UO_1089 (O_1089,N_29869,N_29893);
or UO_1090 (O_1090,N_29943,N_29936);
xor UO_1091 (O_1091,N_29888,N_29834);
xnor UO_1092 (O_1092,N_29935,N_29924);
nand UO_1093 (O_1093,N_29912,N_29829);
nor UO_1094 (O_1094,N_29817,N_29983);
or UO_1095 (O_1095,N_29981,N_29922);
and UO_1096 (O_1096,N_29869,N_29847);
nor UO_1097 (O_1097,N_29837,N_29857);
nand UO_1098 (O_1098,N_29826,N_29955);
xnor UO_1099 (O_1099,N_29853,N_29843);
and UO_1100 (O_1100,N_29831,N_29853);
nand UO_1101 (O_1101,N_29993,N_29894);
nor UO_1102 (O_1102,N_29878,N_29867);
nand UO_1103 (O_1103,N_29883,N_29953);
xnor UO_1104 (O_1104,N_29958,N_29881);
nand UO_1105 (O_1105,N_29843,N_29937);
or UO_1106 (O_1106,N_29860,N_29818);
nor UO_1107 (O_1107,N_29931,N_29987);
or UO_1108 (O_1108,N_29955,N_29989);
nand UO_1109 (O_1109,N_29996,N_29967);
and UO_1110 (O_1110,N_29926,N_29825);
nor UO_1111 (O_1111,N_29884,N_29872);
nor UO_1112 (O_1112,N_29802,N_29991);
nor UO_1113 (O_1113,N_29954,N_29805);
nor UO_1114 (O_1114,N_29948,N_29939);
nor UO_1115 (O_1115,N_29891,N_29922);
nor UO_1116 (O_1116,N_29906,N_29895);
and UO_1117 (O_1117,N_29835,N_29936);
xor UO_1118 (O_1118,N_29957,N_29827);
nor UO_1119 (O_1119,N_29809,N_29962);
xnor UO_1120 (O_1120,N_29866,N_29959);
nand UO_1121 (O_1121,N_29900,N_29853);
nand UO_1122 (O_1122,N_29866,N_29999);
nor UO_1123 (O_1123,N_29884,N_29913);
xnor UO_1124 (O_1124,N_29905,N_29946);
and UO_1125 (O_1125,N_29860,N_29878);
and UO_1126 (O_1126,N_29890,N_29816);
nor UO_1127 (O_1127,N_29956,N_29872);
xnor UO_1128 (O_1128,N_29811,N_29940);
nor UO_1129 (O_1129,N_29873,N_29910);
nand UO_1130 (O_1130,N_29833,N_29954);
or UO_1131 (O_1131,N_29908,N_29911);
nor UO_1132 (O_1132,N_29843,N_29992);
or UO_1133 (O_1133,N_29933,N_29819);
and UO_1134 (O_1134,N_29990,N_29821);
nor UO_1135 (O_1135,N_29970,N_29896);
and UO_1136 (O_1136,N_29883,N_29931);
nor UO_1137 (O_1137,N_29803,N_29919);
xor UO_1138 (O_1138,N_29865,N_29966);
nor UO_1139 (O_1139,N_29924,N_29912);
or UO_1140 (O_1140,N_29829,N_29850);
and UO_1141 (O_1141,N_29899,N_29804);
nand UO_1142 (O_1142,N_29955,N_29833);
nand UO_1143 (O_1143,N_29956,N_29815);
xnor UO_1144 (O_1144,N_29816,N_29883);
xnor UO_1145 (O_1145,N_29841,N_29925);
or UO_1146 (O_1146,N_29938,N_29878);
nand UO_1147 (O_1147,N_29813,N_29899);
or UO_1148 (O_1148,N_29949,N_29929);
or UO_1149 (O_1149,N_29985,N_29847);
or UO_1150 (O_1150,N_29839,N_29921);
nand UO_1151 (O_1151,N_29908,N_29862);
nand UO_1152 (O_1152,N_29953,N_29924);
or UO_1153 (O_1153,N_29913,N_29862);
or UO_1154 (O_1154,N_29950,N_29830);
and UO_1155 (O_1155,N_29987,N_29833);
xnor UO_1156 (O_1156,N_29963,N_29908);
or UO_1157 (O_1157,N_29982,N_29885);
xnor UO_1158 (O_1158,N_29909,N_29984);
xor UO_1159 (O_1159,N_29940,N_29909);
or UO_1160 (O_1160,N_29999,N_29968);
nand UO_1161 (O_1161,N_29997,N_29908);
and UO_1162 (O_1162,N_29801,N_29879);
nand UO_1163 (O_1163,N_29825,N_29808);
xor UO_1164 (O_1164,N_29926,N_29945);
or UO_1165 (O_1165,N_29817,N_29944);
xor UO_1166 (O_1166,N_29863,N_29963);
and UO_1167 (O_1167,N_29913,N_29858);
and UO_1168 (O_1168,N_29896,N_29854);
or UO_1169 (O_1169,N_29858,N_29926);
xnor UO_1170 (O_1170,N_29914,N_29982);
or UO_1171 (O_1171,N_29908,N_29905);
xor UO_1172 (O_1172,N_29887,N_29811);
nand UO_1173 (O_1173,N_29881,N_29863);
or UO_1174 (O_1174,N_29952,N_29839);
nor UO_1175 (O_1175,N_29886,N_29830);
nor UO_1176 (O_1176,N_29892,N_29900);
and UO_1177 (O_1177,N_29918,N_29877);
nand UO_1178 (O_1178,N_29832,N_29883);
or UO_1179 (O_1179,N_29946,N_29977);
nand UO_1180 (O_1180,N_29849,N_29978);
and UO_1181 (O_1181,N_29821,N_29945);
xor UO_1182 (O_1182,N_29940,N_29969);
or UO_1183 (O_1183,N_29803,N_29920);
nor UO_1184 (O_1184,N_29876,N_29999);
nor UO_1185 (O_1185,N_29917,N_29926);
nand UO_1186 (O_1186,N_29835,N_29888);
xor UO_1187 (O_1187,N_29868,N_29948);
nor UO_1188 (O_1188,N_29938,N_29853);
and UO_1189 (O_1189,N_29872,N_29928);
and UO_1190 (O_1190,N_29933,N_29927);
or UO_1191 (O_1191,N_29939,N_29876);
or UO_1192 (O_1192,N_29835,N_29856);
nor UO_1193 (O_1193,N_29970,N_29856);
or UO_1194 (O_1194,N_29930,N_29963);
nand UO_1195 (O_1195,N_29818,N_29855);
or UO_1196 (O_1196,N_29897,N_29989);
xor UO_1197 (O_1197,N_29967,N_29937);
or UO_1198 (O_1198,N_29835,N_29862);
nand UO_1199 (O_1199,N_29831,N_29837);
and UO_1200 (O_1200,N_29916,N_29943);
nor UO_1201 (O_1201,N_29956,N_29935);
nor UO_1202 (O_1202,N_29915,N_29853);
and UO_1203 (O_1203,N_29880,N_29840);
and UO_1204 (O_1204,N_29804,N_29949);
nand UO_1205 (O_1205,N_29817,N_29941);
nand UO_1206 (O_1206,N_29904,N_29966);
nor UO_1207 (O_1207,N_29803,N_29913);
nor UO_1208 (O_1208,N_29940,N_29962);
nor UO_1209 (O_1209,N_29828,N_29890);
nand UO_1210 (O_1210,N_29942,N_29801);
nor UO_1211 (O_1211,N_29943,N_29903);
nor UO_1212 (O_1212,N_29809,N_29886);
xnor UO_1213 (O_1213,N_29869,N_29865);
or UO_1214 (O_1214,N_29966,N_29978);
and UO_1215 (O_1215,N_29983,N_29960);
nand UO_1216 (O_1216,N_29805,N_29940);
xnor UO_1217 (O_1217,N_29903,N_29811);
xnor UO_1218 (O_1218,N_29952,N_29896);
nor UO_1219 (O_1219,N_29957,N_29840);
or UO_1220 (O_1220,N_29818,N_29953);
and UO_1221 (O_1221,N_29841,N_29938);
xnor UO_1222 (O_1222,N_29914,N_29950);
or UO_1223 (O_1223,N_29932,N_29903);
xnor UO_1224 (O_1224,N_29980,N_29813);
nand UO_1225 (O_1225,N_29972,N_29833);
nand UO_1226 (O_1226,N_29972,N_29800);
and UO_1227 (O_1227,N_29986,N_29943);
xnor UO_1228 (O_1228,N_29864,N_29850);
or UO_1229 (O_1229,N_29806,N_29957);
nand UO_1230 (O_1230,N_29931,N_29984);
or UO_1231 (O_1231,N_29830,N_29976);
nand UO_1232 (O_1232,N_29944,N_29996);
or UO_1233 (O_1233,N_29825,N_29997);
and UO_1234 (O_1234,N_29828,N_29975);
nand UO_1235 (O_1235,N_29944,N_29905);
or UO_1236 (O_1236,N_29940,N_29957);
nand UO_1237 (O_1237,N_29942,N_29951);
and UO_1238 (O_1238,N_29821,N_29886);
nand UO_1239 (O_1239,N_29843,N_29871);
xor UO_1240 (O_1240,N_29812,N_29859);
nor UO_1241 (O_1241,N_29836,N_29990);
nand UO_1242 (O_1242,N_29839,N_29853);
xor UO_1243 (O_1243,N_29835,N_29813);
and UO_1244 (O_1244,N_29982,N_29935);
nand UO_1245 (O_1245,N_29871,N_29948);
nand UO_1246 (O_1246,N_29981,N_29958);
nand UO_1247 (O_1247,N_29879,N_29809);
nand UO_1248 (O_1248,N_29906,N_29840);
or UO_1249 (O_1249,N_29809,N_29903);
nand UO_1250 (O_1250,N_29885,N_29805);
xor UO_1251 (O_1251,N_29841,N_29840);
or UO_1252 (O_1252,N_29875,N_29911);
or UO_1253 (O_1253,N_29874,N_29923);
xor UO_1254 (O_1254,N_29997,N_29918);
nor UO_1255 (O_1255,N_29837,N_29882);
xnor UO_1256 (O_1256,N_29964,N_29854);
nand UO_1257 (O_1257,N_29961,N_29853);
nor UO_1258 (O_1258,N_29833,N_29812);
nand UO_1259 (O_1259,N_29851,N_29970);
xor UO_1260 (O_1260,N_29817,N_29905);
and UO_1261 (O_1261,N_29895,N_29822);
nor UO_1262 (O_1262,N_29841,N_29873);
and UO_1263 (O_1263,N_29966,N_29919);
nand UO_1264 (O_1264,N_29928,N_29834);
or UO_1265 (O_1265,N_29809,N_29868);
and UO_1266 (O_1266,N_29833,N_29911);
or UO_1267 (O_1267,N_29961,N_29931);
nand UO_1268 (O_1268,N_29808,N_29987);
or UO_1269 (O_1269,N_29818,N_29958);
or UO_1270 (O_1270,N_29974,N_29883);
nor UO_1271 (O_1271,N_29870,N_29888);
or UO_1272 (O_1272,N_29912,N_29961);
xnor UO_1273 (O_1273,N_29805,N_29998);
nor UO_1274 (O_1274,N_29952,N_29918);
or UO_1275 (O_1275,N_29901,N_29905);
nand UO_1276 (O_1276,N_29945,N_29853);
or UO_1277 (O_1277,N_29850,N_29882);
nand UO_1278 (O_1278,N_29935,N_29807);
nand UO_1279 (O_1279,N_29886,N_29982);
or UO_1280 (O_1280,N_29930,N_29843);
nand UO_1281 (O_1281,N_29867,N_29881);
nand UO_1282 (O_1282,N_29805,N_29882);
nor UO_1283 (O_1283,N_29984,N_29837);
nand UO_1284 (O_1284,N_29887,N_29862);
or UO_1285 (O_1285,N_29954,N_29819);
and UO_1286 (O_1286,N_29975,N_29852);
nand UO_1287 (O_1287,N_29993,N_29909);
and UO_1288 (O_1288,N_29973,N_29850);
or UO_1289 (O_1289,N_29814,N_29854);
and UO_1290 (O_1290,N_29830,N_29955);
and UO_1291 (O_1291,N_29912,N_29823);
nand UO_1292 (O_1292,N_29879,N_29949);
nand UO_1293 (O_1293,N_29845,N_29840);
nor UO_1294 (O_1294,N_29953,N_29946);
or UO_1295 (O_1295,N_29871,N_29914);
nand UO_1296 (O_1296,N_29993,N_29953);
nor UO_1297 (O_1297,N_29872,N_29929);
or UO_1298 (O_1298,N_29834,N_29807);
xnor UO_1299 (O_1299,N_29912,N_29943);
and UO_1300 (O_1300,N_29897,N_29967);
xnor UO_1301 (O_1301,N_29831,N_29933);
or UO_1302 (O_1302,N_29850,N_29828);
and UO_1303 (O_1303,N_29871,N_29992);
nor UO_1304 (O_1304,N_29927,N_29921);
xnor UO_1305 (O_1305,N_29894,N_29889);
nand UO_1306 (O_1306,N_29829,N_29876);
nor UO_1307 (O_1307,N_29818,N_29807);
nor UO_1308 (O_1308,N_29874,N_29955);
and UO_1309 (O_1309,N_29904,N_29928);
xnor UO_1310 (O_1310,N_29871,N_29972);
nor UO_1311 (O_1311,N_29830,N_29852);
nand UO_1312 (O_1312,N_29892,N_29879);
or UO_1313 (O_1313,N_29998,N_29847);
and UO_1314 (O_1314,N_29982,N_29997);
nand UO_1315 (O_1315,N_29834,N_29883);
or UO_1316 (O_1316,N_29896,N_29976);
nand UO_1317 (O_1317,N_29849,N_29989);
or UO_1318 (O_1318,N_29878,N_29987);
or UO_1319 (O_1319,N_29943,N_29944);
nor UO_1320 (O_1320,N_29862,N_29940);
or UO_1321 (O_1321,N_29848,N_29906);
nor UO_1322 (O_1322,N_29988,N_29853);
or UO_1323 (O_1323,N_29978,N_29873);
nor UO_1324 (O_1324,N_29821,N_29836);
or UO_1325 (O_1325,N_29919,N_29836);
nand UO_1326 (O_1326,N_29834,N_29954);
nor UO_1327 (O_1327,N_29976,N_29881);
or UO_1328 (O_1328,N_29921,N_29816);
or UO_1329 (O_1329,N_29959,N_29911);
nor UO_1330 (O_1330,N_29874,N_29920);
or UO_1331 (O_1331,N_29840,N_29833);
or UO_1332 (O_1332,N_29929,N_29923);
xor UO_1333 (O_1333,N_29848,N_29857);
nor UO_1334 (O_1334,N_29985,N_29950);
and UO_1335 (O_1335,N_29824,N_29873);
or UO_1336 (O_1336,N_29925,N_29961);
and UO_1337 (O_1337,N_29807,N_29829);
or UO_1338 (O_1338,N_29832,N_29878);
and UO_1339 (O_1339,N_29849,N_29894);
xnor UO_1340 (O_1340,N_29845,N_29904);
xor UO_1341 (O_1341,N_29843,N_29809);
and UO_1342 (O_1342,N_29887,N_29890);
and UO_1343 (O_1343,N_29948,N_29914);
nand UO_1344 (O_1344,N_29962,N_29911);
and UO_1345 (O_1345,N_29933,N_29900);
xor UO_1346 (O_1346,N_29912,N_29861);
or UO_1347 (O_1347,N_29803,N_29945);
or UO_1348 (O_1348,N_29859,N_29952);
nor UO_1349 (O_1349,N_29978,N_29938);
and UO_1350 (O_1350,N_29954,N_29916);
and UO_1351 (O_1351,N_29919,N_29928);
or UO_1352 (O_1352,N_29817,N_29989);
nor UO_1353 (O_1353,N_29982,N_29857);
or UO_1354 (O_1354,N_29983,N_29996);
and UO_1355 (O_1355,N_29805,N_29986);
xnor UO_1356 (O_1356,N_29865,N_29941);
nand UO_1357 (O_1357,N_29907,N_29965);
nor UO_1358 (O_1358,N_29995,N_29851);
and UO_1359 (O_1359,N_29983,N_29969);
nor UO_1360 (O_1360,N_29822,N_29829);
nor UO_1361 (O_1361,N_29877,N_29903);
xnor UO_1362 (O_1362,N_29951,N_29907);
and UO_1363 (O_1363,N_29950,N_29965);
and UO_1364 (O_1364,N_29970,N_29986);
nor UO_1365 (O_1365,N_29808,N_29998);
nor UO_1366 (O_1366,N_29864,N_29973);
or UO_1367 (O_1367,N_29932,N_29896);
xor UO_1368 (O_1368,N_29872,N_29813);
or UO_1369 (O_1369,N_29885,N_29869);
and UO_1370 (O_1370,N_29828,N_29974);
nor UO_1371 (O_1371,N_29837,N_29906);
nand UO_1372 (O_1372,N_29990,N_29823);
nor UO_1373 (O_1373,N_29859,N_29979);
and UO_1374 (O_1374,N_29853,N_29830);
or UO_1375 (O_1375,N_29832,N_29903);
nor UO_1376 (O_1376,N_29815,N_29960);
nand UO_1377 (O_1377,N_29918,N_29895);
and UO_1378 (O_1378,N_29839,N_29908);
nand UO_1379 (O_1379,N_29841,N_29983);
nor UO_1380 (O_1380,N_29919,N_29906);
nor UO_1381 (O_1381,N_29868,N_29965);
or UO_1382 (O_1382,N_29925,N_29944);
nor UO_1383 (O_1383,N_29981,N_29960);
and UO_1384 (O_1384,N_29845,N_29972);
xor UO_1385 (O_1385,N_29855,N_29869);
and UO_1386 (O_1386,N_29935,N_29908);
nor UO_1387 (O_1387,N_29885,N_29989);
xor UO_1388 (O_1388,N_29955,N_29880);
and UO_1389 (O_1389,N_29838,N_29896);
and UO_1390 (O_1390,N_29850,N_29942);
or UO_1391 (O_1391,N_29861,N_29951);
nand UO_1392 (O_1392,N_29962,N_29925);
and UO_1393 (O_1393,N_29855,N_29988);
and UO_1394 (O_1394,N_29824,N_29854);
and UO_1395 (O_1395,N_29965,N_29901);
nor UO_1396 (O_1396,N_29964,N_29915);
nor UO_1397 (O_1397,N_29859,N_29966);
and UO_1398 (O_1398,N_29966,N_29982);
nand UO_1399 (O_1399,N_29883,N_29874);
and UO_1400 (O_1400,N_29803,N_29983);
or UO_1401 (O_1401,N_29909,N_29844);
nor UO_1402 (O_1402,N_29943,N_29844);
xor UO_1403 (O_1403,N_29838,N_29991);
nand UO_1404 (O_1404,N_29977,N_29865);
and UO_1405 (O_1405,N_29951,N_29900);
and UO_1406 (O_1406,N_29881,N_29916);
nand UO_1407 (O_1407,N_29961,N_29919);
nor UO_1408 (O_1408,N_29876,N_29963);
and UO_1409 (O_1409,N_29949,N_29998);
or UO_1410 (O_1410,N_29821,N_29903);
nand UO_1411 (O_1411,N_29932,N_29966);
nor UO_1412 (O_1412,N_29963,N_29816);
xnor UO_1413 (O_1413,N_29914,N_29940);
nand UO_1414 (O_1414,N_29831,N_29867);
nor UO_1415 (O_1415,N_29911,N_29938);
nor UO_1416 (O_1416,N_29894,N_29918);
nand UO_1417 (O_1417,N_29965,N_29805);
or UO_1418 (O_1418,N_29927,N_29978);
nand UO_1419 (O_1419,N_29946,N_29903);
and UO_1420 (O_1420,N_29844,N_29963);
nand UO_1421 (O_1421,N_29904,N_29879);
and UO_1422 (O_1422,N_29847,N_29874);
or UO_1423 (O_1423,N_29914,N_29855);
nor UO_1424 (O_1424,N_29863,N_29840);
nor UO_1425 (O_1425,N_29898,N_29952);
nand UO_1426 (O_1426,N_29800,N_29956);
xnor UO_1427 (O_1427,N_29866,N_29994);
and UO_1428 (O_1428,N_29842,N_29811);
and UO_1429 (O_1429,N_29824,N_29864);
xor UO_1430 (O_1430,N_29837,N_29887);
nand UO_1431 (O_1431,N_29868,N_29872);
or UO_1432 (O_1432,N_29954,N_29948);
or UO_1433 (O_1433,N_29986,N_29802);
or UO_1434 (O_1434,N_29864,N_29886);
xor UO_1435 (O_1435,N_29871,N_29937);
nand UO_1436 (O_1436,N_29969,N_29968);
nand UO_1437 (O_1437,N_29908,N_29846);
nor UO_1438 (O_1438,N_29924,N_29833);
or UO_1439 (O_1439,N_29947,N_29864);
nor UO_1440 (O_1440,N_29963,N_29968);
xnor UO_1441 (O_1441,N_29873,N_29890);
nor UO_1442 (O_1442,N_29951,N_29854);
nand UO_1443 (O_1443,N_29820,N_29810);
nand UO_1444 (O_1444,N_29854,N_29872);
and UO_1445 (O_1445,N_29811,N_29876);
nor UO_1446 (O_1446,N_29976,N_29980);
nor UO_1447 (O_1447,N_29885,N_29867);
or UO_1448 (O_1448,N_29858,N_29848);
or UO_1449 (O_1449,N_29913,N_29855);
and UO_1450 (O_1450,N_29901,N_29814);
nor UO_1451 (O_1451,N_29963,N_29944);
nand UO_1452 (O_1452,N_29920,N_29839);
nor UO_1453 (O_1453,N_29955,N_29914);
and UO_1454 (O_1454,N_29827,N_29954);
nor UO_1455 (O_1455,N_29888,N_29879);
xnor UO_1456 (O_1456,N_29980,N_29954);
or UO_1457 (O_1457,N_29880,N_29884);
or UO_1458 (O_1458,N_29976,N_29895);
and UO_1459 (O_1459,N_29808,N_29867);
xor UO_1460 (O_1460,N_29964,N_29941);
nand UO_1461 (O_1461,N_29973,N_29976);
and UO_1462 (O_1462,N_29811,N_29875);
and UO_1463 (O_1463,N_29912,N_29964);
or UO_1464 (O_1464,N_29952,N_29985);
and UO_1465 (O_1465,N_29858,N_29999);
and UO_1466 (O_1466,N_29933,N_29945);
and UO_1467 (O_1467,N_29946,N_29945);
xnor UO_1468 (O_1468,N_29856,N_29825);
nor UO_1469 (O_1469,N_29898,N_29925);
nand UO_1470 (O_1470,N_29913,N_29878);
or UO_1471 (O_1471,N_29820,N_29878);
xor UO_1472 (O_1472,N_29872,N_29866);
or UO_1473 (O_1473,N_29868,N_29867);
and UO_1474 (O_1474,N_29825,N_29957);
xnor UO_1475 (O_1475,N_29860,N_29841);
nor UO_1476 (O_1476,N_29898,N_29897);
xor UO_1477 (O_1477,N_29965,N_29860);
or UO_1478 (O_1478,N_29938,N_29891);
nand UO_1479 (O_1479,N_29839,N_29808);
nor UO_1480 (O_1480,N_29827,N_29982);
xnor UO_1481 (O_1481,N_29947,N_29900);
nor UO_1482 (O_1482,N_29803,N_29988);
nand UO_1483 (O_1483,N_29974,N_29823);
nor UO_1484 (O_1484,N_29960,N_29903);
or UO_1485 (O_1485,N_29850,N_29971);
or UO_1486 (O_1486,N_29878,N_29811);
nand UO_1487 (O_1487,N_29842,N_29981);
nand UO_1488 (O_1488,N_29814,N_29838);
nor UO_1489 (O_1489,N_29815,N_29938);
nand UO_1490 (O_1490,N_29971,N_29961);
nand UO_1491 (O_1491,N_29948,N_29836);
or UO_1492 (O_1492,N_29905,N_29961);
and UO_1493 (O_1493,N_29946,N_29802);
and UO_1494 (O_1494,N_29836,N_29833);
xor UO_1495 (O_1495,N_29940,N_29874);
and UO_1496 (O_1496,N_29958,N_29865);
nand UO_1497 (O_1497,N_29802,N_29879);
or UO_1498 (O_1498,N_29831,N_29926);
nor UO_1499 (O_1499,N_29971,N_29890);
or UO_1500 (O_1500,N_29981,N_29883);
or UO_1501 (O_1501,N_29815,N_29824);
nor UO_1502 (O_1502,N_29977,N_29891);
nand UO_1503 (O_1503,N_29919,N_29979);
or UO_1504 (O_1504,N_29826,N_29925);
or UO_1505 (O_1505,N_29862,N_29838);
or UO_1506 (O_1506,N_29859,N_29986);
nor UO_1507 (O_1507,N_29855,N_29809);
and UO_1508 (O_1508,N_29881,N_29950);
or UO_1509 (O_1509,N_29922,N_29971);
xor UO_1510 (O_1510,N_29881,N_29800);
nand UO_1511 (O_1511,N_29838,N_29994);
nand UO_1512 (O_1512,N_29858,N_29938);
nand UO_1513 (O_1513,N_29881,N_29892);
or UO_1514 (O_1514,N_29949,N_29842);
or UO_1515 (O_1515,N_29931,N_29846);
or UO_1516 (O_1516,N_29976,N_29951);
or UO_1517 (O_1517,N_29968,N_29890);
nand UO_1518 (O_1518,N_29919,N_29977);
or UO_1519 (O_1519,N_29812,N_29943);
and UO_1520 (O_1520,N_29871,N_29923);
and UO_1521 (O_1521,N_29809,N_29904);
and UO_1522 (O_1522,N_29951,N_29982);
and UO_1523 (O_1523,N_29819,N_29931);
or UO_1524 (O_1524,N_29837,N_29881);
xor UO_1525 (O_1525,N_29810,N_29883);
nor UO_1526 (O_1526,N_29973,N_29906);
and UO_1527 (O_1527,N_29961,N_29921);
or UO_1528 (O_1528,N_29870,N_29971);
nand UO_1529 (O_1529,N_29859,N_29907);
nand UO_1530 (O_1530,N_29904,N_29847);
nor UO_1531 (O_1531,N_29988,N_29846);
and UO_1532 (O_1532,N_29982,N_29800);
nor UO_1533 (O_1533,N_29946,N_29997);
xor UO_1534 (O_1534,N_29899,N_29843);
or UO_1535 (O_1535,N_29824,N_29943);
and UO_1536 (O_1536,N_29932,N_29948);
and UO_1537 (O_1537,N_29809,N_29929);
and UO_1538 (O_1538,N_29980,N_29940);
and UO_1539 (O_1539,N_29930,N_29802);
or UO_1540 (O_1540,N_29821,N_29838);
and UO_1541 (O_1541,N_29993,N_29884);
and UO_1542 (O_1542,N_29908,N_29855);
and UO_1543 (O_1543,N_29903,N_29855);
xnor UO_1544 (O_1544,N_29925,N_29994);
xor UO_1545 (O_1545,N_29813,N_29914);
nand UO_1546 (O_1546,N_29871,N_29965);
nand UO_1547 (O_1547,N_29816,N_29940);
or UO_1548 (O_1548,N_29995,N_29940);
and UO_1549 (O_1549,N_29914,N_29909);
nand UO_1550 (O_1550,N_29914,N_29873);
or UO_1551 (O_1551,N_29904,N_29834);
nand UO_1552 (O_1552,N_29942,N_29859);
nand UO_1553 (O_1553,N_29952,N_29879);
nor UO_1554 (O_1554,N_29954,N_29813);
xor UO_1555 (O_1555,N_29843,N_29943);
and UO_1556 (O_1556,N_29874,N_29917);
nand UO_1557 (O_1557,N_29932,N_29995);
xnor UO_1558 (O_1558,N_29845,N_29841);
xor UO_1559 (O_1559,N_29920,N_29858);
xor UO_1560 (O_1560,N_29977,N_29969);
xor UO_1561 (O_1561,N_29877,N_29974);
and UO_1562 (O_1562,N_29929,N_29993);
xor UO_1563 (O_1563,N_29881,N_29987);
nor UO_1564 (O_1564,N_29823,N_29837);
or UO_1565 (O_1565,N_29978,N_29829);
or UO_1566 (O_1566,N_29945,N_29951);
or UO_1567 (O_1567,N_29863,N_29832);
nand UO_1568 (O_1568,N_29856,N_29896);
or UO_1569 (O_1569,N_29905,N_29962);
and UO_1570 (O_1570,N_29821,N_29861);
or UO_1571 (O_1571,N_29955,N_29896);
xor UO_1572 (O_1572,N_29993,N_29949);
or UO_1573 (O_1573,N_29933,N_29907);
nand UO_1574 (O_1574,N_29808,N_29897);
and UO_1575 (O_1575,N_29958,N_29969);
xnor UO_1576 (O_1576,N_29897,N_29848);
xnor UO_1577 (O_1577,N_29849,N_29977);
or UO_1578 (O_1578,N_29974,N_29879);
xor UO_1579 (O_1579,N_29964,N_29814);
xnor UO_1580 (O_1580,N_29905,N_29980);
nor UO_1581 (O_1581,N_29932,N_29975);
nand UO_1582 (O_1582,N_29912,N_29906);
xor UO_1583 (O_1583,N_29836,N_29806);
nor UO_1584 (O_1584,N_29995,N_29952);
and UO_1585 (O_1585,N_29835,N_29820);
xor UO_1586 (O_1586,N_29853,N_29933);
and UO_1587 (O_1587,N_29906,N_29900);
xor UO_1588 (O_1588,N_29822,N_29903);
nand UO_1589 (O_1589,N_29905,N_29957);
xor UO_1590 (O_1590,N_29863,N_29801);
or UO_1591 (O_1591,N_29862,N_29830);
nor UO_1592 (O_1592,N_29916,N_29853);
and UO_1593 (O_1593,N_29941,N_29938);
and UO_1594 (O_1594,N_29926,N_29823);
or UO_1595 (O_1595,N_29926,N_29830);
and UO_1596 (O_1596,N_29838,N_29940);
or UO_1597 (O_1597,N_29804,N_29860);
xnor UO_1598 (O_1598,N_29937,N_29941);
and UO_1599 (O_1599,N_29980,N_29956);
xor UO_1600 (O_1600,N_29953,N_29919);
xnor UO_1601 (O_1601,N_29972,N_29937);
or UO_1602 (O_1602,N_29943,N_29837);
or UO_1603 (O_1603,N_29927,N_29917);
xor UO_1604 (O_1604,N_29998,N_29807);
xnor UO_1605 (O_1605,N_29847,N_29817);
or UO_1606 (O_1606,N_29843,N_29911);
nor UO_1607 (O_1607,N_29922,N_29986);
and UO_1608 (O_1608,N_29887,N_29844);
or UO_1609 (O_1609,N_29802,N_29876);
or UO_1610 (O_1610,N_29816,N_29855);
nor UO_1611 (O_1611,N_29916,N_29878);
xor UO_1612 (O_1612,N_29931,N_29811);
xor UO_1613 (O_1613,N_29863,N_29898);
xor UO_1614 (O_1614,N_29859,N_29890);
nand UO_1615 (O_1615,N_29942,N_29860);
nand UO_1616 (O_1616,N_29842,N_29961);
and UO_1617 (O_1617,N_29843,N_29825);
and UO_1618 (O_1618,N_29925,N_29953);
nand UO_1619 (O_1619,N_29959,N_29907);
nand UO_1620 (O_1620,N_29856,N_29997);
and UO_1621 (O_1621,N_29978,N_29905);
nor UO_1622 (O_1622,N_29911,N_29917);
xor UO_1623 (O_1623,N_29954,N_29836);
xor UO_1624 (O_1624,N_29938,N_29967);
nor UO_1625 (O_1625,N_29808,N_29930);
nand UO_1626 (O_1626,N_29977,N_29906);
or UO_1627 (O_1627,N_29824,N_29826);
xor UO_1628 (O_1628,N_29841,N_29979);
nand UO_1629 (O_1629,N_29879,N_29812);
or UO_1630 (O_1630,N_29921,N_29818);
and UO_1631 (O_1631,N_29888,N_29904);
nand UO_1632 (O_1632,N_29969,N_29950);
nor UO_1633 (O_1633,N_29943,N_29998);
or UO_1634 (O_1634,N_29973,N_29834);
xnor UO_1635 (O_1635,N_29840,N_29936);
nand UO_1636 (O_1636,N_29974,N_29878);
xor UO_1637 (O_1637,N_29923,N_29949);
nand UO_1638 (O_1638,N_29916,N_29915);
and UO_1639 (O_1639,N_29864,N_29937);
or UO_1640 (O_1640,N_29812,N_29886);
or UO_1641 (O_1641,N_29868,N_29982);
or UO_1642 (O_1642,N_29846,N_29915);
or UO_1643 (O_1643,N_29939,N_29962);
or UO_1644 (O_1644,N_29961,N_29857);
nand UO_1645 (O_1645,N_29844,N_29831);
or UO_1646 (O_1646,N_29978,N_29942);
or UO_1647 (O_1647,N_29936,N_29920);
xor UO_1648 (O_1648,N_29836,N_29912);
nand UO_1649 (O_1649,N_29842,N_29927);
or UO_1650 (O_1650,N_29939,N_29849);
nand UO_1651 (O_1651,N_29824,N_29863);
xor UO_1652 (O_1652,N_29860,N_29829);
and UO_1653 (O_1653,N_29930,N_29984);
nor UO_1654 (O_1654,N_29841,N_29815);
and UO_1655 (O_1655,N_29931,N_29988);
and UO_1656 (O_1656,N_29848,N_29885);
xnor UO_1657 (O_1657,N_29902,N_29986);
or UO_1658 (O_1658,N_29866,N_29995);
nor UO_1659 (O_1659,N_29871,N_29803);
or UO_1660 (O_1660,N_29953,N_29977);
nor UO_1661 (O_1661,N_29988,N_29905);
nor UO_1662 (O_1662,N_29885,N_29969);
and UO_1663 (O_1663,N_29852,N_29901);
or UO_1664 (O_1664,N_29913,N_29992);
and UO_1665 (O_1665,N_29880,N_29954);
or UO_1666 (O_1666,N_29842,N_29926);
nand UO_1667 (O_1667,N_29901,N_29931);
nand UO_1668 (O_1668,N_29925,N_29832);
xnor UO_1669 (O_1669,N_29993,N_29858);
nor UO_1670 (O_1670,N_29875,N_29977);
and UO_1671 (O_1671,N_29822,N_29951);
or UO_1672 (O_1672,N_29997,N_29933);
or UO_1673 (O_1673,N_29994,N_29801);
or UO_1674 (O_1674,N_29909,N_29996);
and UO_1675 (O_1675,N_29831,N_29874);
xor UO_1676 (O_1676,N_29814,N_29875);
xnor UO_1677 (O_1677,N_29902,N_29900);
xnor UO_1678 (O_1678,N_29847,N_29845);
nor UO_1679 (O_1679,N_29927,N_29929);
nand UO_1680 (O_1680,N_29863,N_29938);
and UO_1681 (O_1681,N_29828,N_29999);
and UO_1682 (O_1682,N_29946,N_29858);
nor UO_1683 (O_1683,N_29960,N_29857);
and UO_1684 (O_1684,N_29924,N_29878);
and UO_1685 (O_1685,N_29886,N_29843);
nand UO_1686 (O_1686,N_29869,N_29954);
xor UO_1687 (O_1687,N_29872,N_29915);
xnor UO_1688 (O_1688,N_29899,N_29942);
xor UO_1689 (O_1689,N_29938,N_29880);
xor UO_1690 (O_1690,N_29862,N_29968);
nand UO_1691 (O_1691,N_29898,N_29878);
nand UO_1692 (O_1692,N_29879,N_29819);
nor UO_1693 (O_1693,N_29930,N_29961);
nor UO_1694 (O_1694,N_29911,N_29940);
or UO_1695 (O_1695,N_29907,N_29851);
nor UO_1696 (O_1696,N_29930,N_29956);
nand UO_1697 (O_1697,N_29929,N_29986);
nand UO_1698 (O_1698,N_29852,N_29889);
xnor UO_1699 (O_1699,N_29871,N_29844);
nand UO_1700 (O_1700,N_29868,N_29895);
and UO_1701 (O_1701,N_29822,N_29917);
and UO_1702 (O_1702,N_29865,N_29881);
and UO_1703 (O_1703,N_29810,N_29819);
xnor UO_1704 (O_1704,N_29951,N_29839);
nand UO_1705 (O_1705,N_29981,N_29989);
nand UO_1706 (O_1706,N_29862,N_29988);
or UO_1707 (O_1707,N_29916,N_29864);
xnor UO_1708 (O_1708,N_29840,N_29998);
nor UO_1709 (O_1709,N_29938,N_29960);
nor UO_1710 (O_1710,N_29846,N_29927);
nand UO_1711 (O_1711,N_29924,N_29984);
nor UO_1712 (O_1712,N_29955,N_29950);
nand UO_1713 (O_1713,N_29924,N_29840);
xnor UO_1714 (O_1714,N_29830,N_29909);
or UO_1715 (O_1715,N_29835,N_29830);
and UO_1716 (O_1716,N_29856,N_29888);
xor UO_1717 (O_1717,N_29893,N_29906);
or UO_1718 (O_1718,N_29935,N_29920);
nor UO_1719 (O_1719,N_29829,N_29874);
and UO_1720 (O_1720,N_29971,N_29855);
and UO_1721 (O_1721,N_29967,N_29856);
nor UO_1722 (O_1722,N_29954,N_29912);
and UO_1723 (O_1723,N_29989,N_29888);
nand UO_1724 (O_1724,N_29928,N_29995);
nor UO_1725 (O_1725,N_29876,N_29842);
and UO_1726 (O_1726,N_29975,N_29804);
and UO_1727 (O_1727,N_29901,N_29843);
xor UO_1728 (O_1728,N_29834,N_29948);
or UO_1729 (O_1729,N_29823,N_29818);
and UO_1730 (O_1730,N_29829,N_29812);
nand UO_1731 (O_1731,N_29800,N_29883);
and UO_1732 (O_1732,N_29849,N_29914);
or UO_1733 (O_1733,N_29871,N_29825);
xor UO_1734 (O_1734,N_29921,N_29929);
nor UO_1735 (O_1735,N_29977,N_29852);
and UO_1736 (O_1736,N_29910,N_29884);
nand UO_1737 (O_1737,N_29893,N_29841);
nor UO_1738 (O_1738,N_29883,N_29803);
nand UO_1739 (O_1739,N_29881,N_29896);
nand UO_1740 (O_1740,N_29982,N_29893);
or UO_1741 (O_1741,N_29906,N_29855);
or UO_1742 (O_1742,N_29936,N_29890);
nor UO_1743 (O_1743,N_29931,N_29893);
nor UO_1744 (O_1744,N_29997,N_29829);
nor UO_1745 (O_1745,N_29938,N_29950);
nor UO_1746 (O_1746,N_29969,N_29872);
xor UO_1747 (O_1747,N_29865,N_29930);
and UO_1748 (O_1748,N_29886,N_29975);
or UO_1749 (O_1749,N_29948,N_29965);
nand UO_1750 (O_1750,N_29966,N_29957);
nor UO_1751 (O_1751,N_29945,N_29989);
or UO_1752 (O_1752,N_29986,N_29994);
and UO_1753 (O_1753,N_29968,N_29946);
or UO_1754 (O_1754,N_29933,N_29991);
or UO_1755 (O_1755,N_29840,N_29832);
and UO_1756 (O_1756,N_29875,N_29892);
or UO_1757 (O_1757,N_29989,N_29840);
xor UO_1758 (O_1758,N_29813,N_29826);
or UO_1759 (O_1759,N_29819,N_29955);
and UO_1760 (O_1760,N_29843,N_29945);
nand UO_1761 (O_1761,N_29972,N_29959);
xor UO_1762 (O_1762,N_29905,N_29837);
or UO_1763 (O_1763,N_29869,N_29962);
or UO_1764 (O_1764,N_29962,N_29909);
nand UO_1765 (O_1765,N_29856,N_29988);
nor UO_1766 (O_1766,N_29823,N_29858);
and UO_1767 (O_1767,N_29937,N_29939);
nand UO_1768 (O_1768,N_29969,N_29910);
nand UO_1769 (O_1769,N_29869,N_29882);
xor UO_1770 (O_1770,N_29949,N_29924);
nand UO_1771 (O_1771,N_29916,N_29966);
xnor UO_1772 (O_1772,N_29989,N_29831);
and UO_1773 (O_1773,N_29874,N_29850);
and UO_1774 (O_1774,N_29905,N_29904);
nand UO_1775 (O_1775,N_29946,N_29922);
or UO_1776 (O_1776,N_29917,N_29919);
nor UO_1777 (O_1777,N_29949,N_29958);
and UO_1778 (O_1778,N_29823,N_29907);
or UO_1779 (O_1779,N_29905,N_29940);
nor UO_1780 (O_1780,N_29806,N_29904);
and UO_1781 (O_1781,N_29932,N_29858);
or UO_1782 (O_1782,N_29905,N_29802);
nor UO_1783 (O_1783,N_29902,N_29961);
xnor UO_1784 (O_1784,N_29895,N_29999);
xnor UO_1785 (O_1785,N_29854,N_29823);
nor UO_1786 (O_1786,N_29939,N_29900);
or UO_1787 (O_1787,N_29823,N_29932);
nand UO_1788 (O_1788,N_29927,N_29949);
nor UO_1789 (O_1789,N_29978,N_29894);
nor UO_1790 (O_1790,N_29952,N_29960);
or UO_1791 (O_1791,N_29993,N_29931);
xnor UO_1792 (O_1792,N_29863,N_29983);
or UO_1793 (O_1793,N_29943,N_29950);
and UO_1794 (O_1794,N_29944,N_29885);
nand UO_1795 (O_1795,N_29826,N_29990);
and UO_1796 (O_1796,N_29887,N_29905);
nand UO_1797 (O_1797,N_29809,N_29940);
nand UO_1798 (O_1798,N_29974,N_29824);
xnor UO_1799 (O_1799,N_29911,N_29941);
nor UO_1800 (O_1800,N_29948,N_29896);
nor UO_1801 (O_1801,N_29902,N_29879);
xnor UO_1802 (O_1802,N_29845,N_29831);
nor UO_1803 (O_1803,N_29898,N_29920);
or UO_1804 (O_1804,N_29830,N_29902);
or UO_1805 (O_1805,N_29817,N_29855);
and UO_1806 (O_1806,N_29872,N_29996);
xnor UO_1807 (O_1807,N_29839,N_29851);
or UO_1808 (O_1808,N_29870,N_29953);
or UO_1809 (O_1809,N_29836,N_29855);
nand UO_1810 (O_1810,N_29952,N_29821);
xor UO_1811 (O_1811,N_29845,N_29977);
nand UO_1812 (O_1812,N_29996,N_29821);
xnor UO_1813 (O_1813,N_29988,N_29836);
nand UO_1814 (O_1814,N_29858,N_29842);
xor UO_1815 (O_1815,N_29986,N_29814);
or UO_1816 (O_1816,N_29901,N_29898);
and UO_1817 (O_1817,N_29899,N_29872);
or UO_1818 (O_1818,N_29963,N_29864);
nand UO_1819 (O_1819,N_29997,N_29841);
nor UO_1820 (O_1820,N_29942,N_29878);
or UO_1821 (O_1821,N_29921,N_29807);
or UO_1822 (O_1822,N_29852,N_29929);
nor UO_1823 (O_1823,N_29877,N_29912);
xnor UO_1824 (O_1824,N_29931,N_29859);
or UO_1825 (O_1825,N_29916,N_29805);
nand UO_1826 (O_1826,N_29852,N_29899);
or UO_1827 (O_1827,N_29818,N_29865);
and UO_1828 (O_1828,N_29983,N_29985);
and UO_1829 (O_1829,N_29922,N_29888);
nor UO_1830 (O_1830,N_29995,N_29984);
nand UO_1831 (O_1831,N_29862,N_29828);
or UO_1832 (O_1832,N_29890,N_29951);
nor UO_1833 (O_1833,N_29989,N_29976);
xor UO_1834 (O_1834,N_29867,N_29812);
xor UO_1835 (O_1835,N_29990,N_29805);
nand UO_1836 (O_1836,N_29836,N_29974);
xnor UO_1837 (O_1837,N_29935,N_29916);
nor UO_1838 (O_1838,N_29856,N_29977);
nor UO_1839 (O_1839,N_29916,N_29808);
xor UO_1840 (O_1840,N_29843,N_29936);
and UO_1841 (O_1841,N_29868,N_29805);
and UO_1842 (O_1842,N_29996,N_29921);
nor UO_1843 (O_1843,N_29969,N_29957);
nor UO_1844 (O_1844,N_29899,N_29912);
or UO_1845 (O_1845,N_29931,N_29995);
and UO_1846 (O_1846,N_29867,N_29817);
nand UO_1847 (O_1847,N_29887,N_29879);
and UO_1848 (O_1848,N_29839,N_29854);
and UO_1849 (O_1849,N_29861,N_29837);
nor UO_1850 (O_1850,N_29870,N_29842);
nand UO_1851 (O_1851,N_29882,N_29827);
or UO_1852 (O_1852,N_29986,N_29953);
or UO_1853 (O_1853,N_29842,N_29947);
xor UO_1854 (O_1854,N_29881,N_29982);
and UO_1855 (O_1855,N_29891,N_29814);
nand UO_1856 (O_1856,N_29918,N_29832);
xnor UO_1857 (O_1857,N_29836,N_29888);
nor UO_1858 (O_1858,N_29951,N_29920);
xnor UO_1859 (O_1859,N_29904,N_29916);
nand UO_1860 (O_1860,N_29803,N_29966);
and UO_1861 (O_1861,N_29912,N_29845);
and UO_1862 (O_1862,N_29899,N_29923);
and UO_1863 (O_1863,N_29875,N_29936);
nand UO_1864 (O_1864,N_29967,N_29887);
nor UO_1865 (O_1865,N_29979,N_29969);
or UO_1866 (O_1866,N_29969,N_29857);
xor UO_1867 (O_1867,N_29819,N_29928);
nand UO_1868 (O_1868,N_29892,N_29950);
nand UO_1869 (O_1869,N_29814,N_29904);
nand UO_1870 (O_1870,N_29806,N_29967);
xnor UO_1871 (O_1871,N_29930,N_29906);
nor UO_1872 (O_1872,N_29969,N_29964);
nand UO_1873 (O_1873,N_29906,N_29891);
and UO_1874 (O_1874,N_29998,N_29850);
and UO_1875 (O_1875,N_29820,N_29975);
nor UO_1876 (O_1876,N_29994,N_29875);
nand UO_1877 (O_1877,N_29964,N_29881);
or UO_1878 (O_1878,N_29804,N_29848);
nand UO_1879 (O_1879,N_29968,N_29984);
xnor UO_1880 (O_1880,N_29984,N_29950);
nor UO_1881 (O_1881,N_29954,N_29868);
xnor UO_1882 (O_1882,N_29961,N_29963);
or UO_1883 (O_1883,N_29994,N_29973);
nand UO_1884 (O_1884,N_29826,N_29817);
xor UO_1885 (O_1885,N_29820,N_29983);
xor UO_1886 (O_1886,N_29866,N_29922);
or UO_1887 (O_1887,N_29849,N_29943);
xnor UO_1888 (O_1888,N_29895,N_29880);
nor UO_1889 (O_1889,N_29912,N_29884);
xnor UO_1890 (O_1890,N_29939,N_29802);
nor UO_1891 (O_1891,N_29908,N_29837);
nand UO_1892 (O_1892,N_29909,N_29915);
nand UO_1893 (O_1893,N_29953,N_29948);
xnor UO_1894 (O_1894,N_29800,N_29969);
or UO_1895 (O_1895,N_29952,N_29833);
nand UO_1896 (O_1896,N_29930,N_29977);
xnor UO_1897 (O_1897,N_29818,N_29854);
xor UO_1898 (O_1898,N_29803,N_29874);
nor UO_1899 (O_1899,N_29998,N_29924);
and UO_1900 (O_1900,N_29908,N_29877);
nand UO_1901 (O_1901,N_29812,N_29922);
or UO_1902 (O_1902,N_29929,N_29977);
and UO_1903 (O_1903,N_29896,N_29815);
xnor UO_1904 (O_1904,N_29911,N_29851);
nand UO_1905 (O_1905,N_29938,N_29851);
or UO_1906 (O_1906,N_29803,N_29957);
nor UO_1907 (O_1907,N_29907,N_29914);
nand UO_1908 (O_1908,N_29981,N_29819);
xnor UO_1909 (O_1909,N_29836,N_29838);
nand UO_1910 (O_1910,N_29917,N_29923);
or UO_1911 (O_1911,N_29802,N_29993);
and UO_1912 (O_1912,N_29861,N_29879);
xnor UO_1913 (O_1913,N_29850,N_29825);
and UO_1914 (O_1914,N_29861,N_29967);
nor UO_1915 (O_1915,N_29832,N_29973);
and UO_1916 (O_1916,N_29870,N_29857);
nor UO_1917 (O_1917,N_29839,N_29855);
xnor UO_1918 (O_1918,N_29925,N_29853);
xor UO_1919 (O_1919,N_29979,N_29896);
and UO_1920 (O_1920,N_29953,N_29989);
and UO_1921 (O_1921,N_29820,N_29949);
or UO_1922 (O_1922,N_29895,N_29941);
nor UO_1923 (O_1923,N_29917,N_29837);
nand UO_1924 (O_1924,N_29981,N_29809);
nand UO_1925 (O_1925,N_29819,N_29948);
nand UO_1926 (O_1926,N_29853,N_29995);
or UO_1927 (O_1927,N_29945,N_29864);
nor UO_1928 (O_1928,N_29909,N_29801);
and UO_1929 (O_1929,N_29994,N_29864);
or UO_1930 (O_1930,N_29894,N_29960);
and UO_1931 (O_1931,N_29922,N_29895);
xnor UO_1932 (O_1932,N_29820,N_29978);
nor UO_1933 (O_1933,N_29864,N_29914);
or UO_1934 (O_1934,N_29858,N_29941);
or UO_1935 (O_1935,N_29878,N_29932);
and UO_1936 (O_1936,N_29996,N_29876);
and UO_1937 (O_1937,N_29935,N_29980);
xnor UO_1938 (O_1938,N_29970,N_29827);
xnor UO_1939 (O_1939,N_29918,N_29816);
xnor UO_1940 (O_1940,N_29872,N_29882);
xnor UO_1941 (O_1941,N_29989,N_29869);
or UO_1942 (O_1942,N_29984,N_29857);
or UO_1943 (O_1943,N_29844,N_29937);
nand UO_1944 (O_1944,N_29969,N_29980);
or UO_1945 (O_1945,N_29977,N_29883);
nor UO_1946 (O_1946,N_29810,N_29847);
or UO_1947 (O_1947,N_29858,N_29921);
xnor UO_1948 (O_1948,N_29865,N_29916);
and UO_1949 (O_1949,N_29915,N_29829);
nand UO_1950 (O_1950,N_29897,N_29856);
nor UO_1951 (O_1951,N_29946,N_29970);
and UO_1952 (O_1952,N_29823,N_29862);
xor UO_1953 (O_1953,N_29866,N_29833);
and UO_1954 (O_1954,N_29937,N_29821);
nor UO_1955 (O_1955,N_29997,N_29828);
nand UO_1956 (O_1956,N_29982,N_29961);
nand UO_1957 (O_1957,N_29935,N_29992);
nor UO_1958 (O_1958,N_29926,N_29851);
xnor UO_1959 (O_1959,N_29840,N_29991);
or UO_1960 (O_1960,N_29816,N_29917);
nand UO_1961 (O_1961,N_29898,N_29955);
nand UO_1962 (O_1962,N_29983,N_29847);
nand UO_1963 (O_1963,N_29818,N_29845);
xnor UO_1964 (O_1964,N_29835,N_29974);
nand UO_1965 (O_1965,N_29808,N_29932);
xor UO_1966 (O_1966,N_29963,N_29843);
xnor UO_1967 (O_1967,N_29882,N_29945);
and UO_1968 (O_1968,N_29836,N_29968);
nor UO_1969 (O_1969,N_29997,N_29962);
xnor UO_1970 (O_1970,N_29968,N_29818);
xnor UO_1971 (O_1971,N_29860,N_29805);
nor UO_1972 (O_1972,N_29990,N_29998);
xnor UO_1973 (O_1973,N_29918,N_29956);
xnor UO_1974 (O_1974,N_29879,N_29813);
or UO_1975 (O_1975,N_29928,N_29964);
nand UO_1976 (O_1976,N_29868,N_29901);
and UO_1977 (O_1977,N_29988,N_29875);
nand UO_1978 (O_1978,N_29856,N_29917);
xor UO_1979 (O_1979,N_29952,N_29901);
nand UO_1980 (O_1980,N_29909,N_29871);
and UO_1981 (O_1981,N_29881,N_29851);
xor UO_1982 (O_1982,N_29844,N_29867);
xor UO_1983 (O_1983,N_29978,N_29952);
nor UO_1984 (O_1984,N_29885,N_29978);
or UO_1985 (O_1985,N_29962,N_29974);
nor UO_1986 (O_1986,N_29844,N_29904);
nand UO_1987 (O_1987,N_29932,N_29874);
and UO_1988 (O_1988,N_29846,N_29937);
nor UO_1989 (O_1989,N_29837,N_29845);
or UO_1990 (O_1990,N_29822,N_29904);
or UO_1991 (O_1991,N_29847,N_29851);
and UO_1992 (O_1992,N_29822,N_29841);
nand UO_1993 (O_1993,N_29942,N_29821);
and UO_1994 (O_1994,N_29953,N_29923);
and UO_1995 (O_1995,N_29909,N_29879);
and UO_1996 (O_1996,N_29827,N_29837);
nor UO_1997 (O_1997,N_29945,N_29805);
and UO_1998 (O_1998,N_29818,N_29916);
nor UO_1999 (O_1999,N_29803,N_29884);
or UO_2000 (O_2000,N_29965,N_29955);
nand UO_2001 (O_2001,N_29950,N_29937);
or UO_2002 (O_2002,N_29816,N_29958);
nor UO_2003 (O_2003,N_29837,N_29931);
or UO_2004 (O_2004,N_29817,N_29819);
nor UO_2005 (O_2005,N_29969,N_29987);
nor UO_2006 (O_2006,N_29875,N_29826);
nand UO_2007 (O_2007,N_29942,N_29922);
nand UO_2008 (O_2008,N_29928,N_29838);
or UO_2009 (O_2009,N_29962,N_29864);
or UO_2010 (O_2010,N_29848,N_29834);
nor UO_2011 (O_2011,N_29869,N_29839);
and UO_2012 (O_2012,N_29875,N_29914);
or UO_2013 (O_2013,N_29989,N_29936);
xnor UO_2014 (O_2014,N_29810,N_29897);
or UO_2015 (O_2015,N_29981,N_29983);
nor UO_2016 (O_2016,N_29831,N_29944);
xor UO_2017 (O_2017,N_29805,N_29955);
nand UO_2018 (O_2018,N_29806,N_29968);
xnor UO_2019 (O_2019,N_29921,N_29842);
xnor UO_2020 (O_2020,N_29982,N_29823);
xnor UO_2021 (O_2021,N_29974,N_29925);
or UO_2022 (O_2022,N_29999,N_29857);
nand UO_2023 (O_2023,N_29869,N_29909);
or UO_2024 (O_2024,N_29827,N_29928);
nand UO_2025 (O_2025,N_29805,N_29889);
xor UO_2026 (O_2026,N_29993,N_29904);
or UO_2027 (O_2027,N_29894,N_29998);
or UO_2028 (O_2028,N_29903,N_29976);
nand UO_2029 (O_2029,N_29905,N_29969);
nor UO_2030 (O_2030,N_29907,N_29889);
xor UO_2031 (O_2031,N_29876,N_29945);
or UO_2032 (O_2032,N_29903,N_29974);
nor UO_2033 (O_2033,N_29834,N_29878);
nand UO_2034 (O_2034,N_29967,N_29871);
or UO_2035 (O_2035,N_29891,N_29862);
and UO_2036 (O_2036,N_29889,N_29845);
xor UO_2037 (O_2037,N_29823,N_29979);
or UO_2038 (O_2038,N_29830,N_29916);
and UO_2039 (O_2039,N_29857,N_29925);
or UO_2040 (O_2040,N_29915,N_29934);
nand UO_2041 (O_2041,N_29835,N_29990);
and UO_2042 (O_2042,N_29800,N_29871);
xnor UO_2043 (O_2043,N_29812,N_29848);
xor UO_2044 (O_2044,N_29923,N_29963);
xnor UO_2045 (O_2045,N_29839,N_29882);
and UO_2046 (O_2046,N_29956,N_29863);
xor UO_2047 (O_2047,N_29874,N_29880);
nand UO_2048 (O_2048,N_29941,N_29973);
nor UO_2049 (O_2049,N_29889,N_29939);
nand UO_2050 (O_2050,N_29892,N_29884);
and UO_2051 (O_2051,N_29806,N_29810);
nand UO_2052 (O_2052,N_29825,N_29859);
nand UO_2053 (O_2053,N_29960,N_29974);
nor UO_2054 (O_2054,N_29925,N_29991);
or UO_2055 (O_2055,N_29884,N_29947);
xnor UO_2056 (O_2056,N_29956,N_29921);
nor UO_2057 (O_2057,N_29848,N_29923);
nand UO_2058 (O_2058,N_29885,N_29843);
nand UO_2059 (O_2059,N_29942,N_29828);
or UO_2060 (O_2060,N_29886,N_29973);
or UO_2061 (O_2061,N_29940,N_29983);
nand UO_2062 (O_2062,N_29940,N_29826);
xor UO_2063 (O_2063,N_29890,N_29987);
nor UO_2064 (O_2064,N_29989,N_29863);
nor UO_2065 (O_2065,N_29870,N_29812);
nand UO_2066 (O_2066,N_29932,N_29993);
and UO_2067 (O_2067,N_29901,N_29954);
nor UO_2068 (O_2068,N_29865,N_29842);
nor UO_2069 (O_2069,N_29928,N_29967);
nor UO_2070 (O_2070,N_29988,N_29951);
nand UO_2071 (O_2071,N_29961,N_29956);
xor UO_2072 (O_2072,N_29949,N_29977);
or UO_2073 (O_2073,N_29863,N_29887);
and UO_2074 (O_2074,N_29916,N_29899);
and UO_2075 (O_2075,N_29866,N_29940);
nor UO_2076 (O_2076,N_29984,N_29982);
nor UO_2077 (O_2077,N_29966,N_29842);
and UO_2078 (O_2078,N_29822,N_29958);
and UO_2079 (O_2079,N_29840,N_29946);
nand UO_2080 (O_2080,N_29965,N_29895);
or UO_2081 (O_2081,N_29897,N_29955);
nand UO_2082 (O_2082,N_29815,N_29853);
and UO_2083 (O_2083,N_29842,N_29979);
xnor UO_2084 (O_2084,N_29853,N_29999);
and UO_2085 (O_2085,N_29822,N_29918);
xnor UO_2086 (O_2086,N_29908,N_29857);
nor UO_2087 (O_2087,N_29819,N_29873);
or UO_2088 (O_2088,N_29889,N_29958);
and UO_2089 (O_2089,N_29880,N_29950);
nor UO_2090 (O_2090,N_29870,N_29999);
and UO_2091 (O_2091,N_29942,N_29947);
xor UO_2092 (O_2092,N_29828,N_29844);
xor UO_2093 (O_2093,N_29804,N_29833);
nand UO_2094 (O_2094,N_29944,N_29894);
or UO_2095 (O_2095,N_29992,N_29817);
xor UO_2096 (O_2096,N_29854,N_29835);
nor UO_2097 (O_2097,N_29875,N_29986);
or UO_2098 (O_2098,N_29997,N_29990);
nand UO_2099 (O_2099,N_29990,N_29802);
and UO_2100 (O_2100,N_29832,N_29943);
xor UO_2101 (O_2101,N_29802,N_29942);
and UO_2102 (O_2102,N_29951,N_29972);
nor UO_2103 (O_2103,N_29895,N_29894);
and UO_2104 (O_2104,N_29961,N_29959);
xor UO_2105 (O_2105,N_29873,N_29840);
and UO_2106 (O_2106,N_29887,N_29816);
nor UO_2107 (O_2107,N_29910,N_29824);
xor UO_2108 (O_2108,N_29829,N_29937);
nor UO_2109 (O_2109,N_29936,N_29946);
xnor UO_2110 (O_2110,N_29835,N_29857);
nor UO_2111 (O_2111,N_29985,N_29808);
nand UO_2112 (O_2112,N_29814,N_29869);
nor UO_2113 (O_2113,N_29988,N_29868);
or UO_2114 (O_2114,N_29908,N_29861);
nand UO_2115 (O_2115,N_29897,N_29811);
nand UO_2116 (O_2116,N_29855,N_29876);
or UO_2117 (O_2117,N_29936,N_29919);
nand UO_2118 (O_2118,N_29860,N_29927);
nor UO_2119 (O_2119,N_29940,N_29888);
or UO_2120 (O_2120,N_29985,N_29936);
nor UO_2121 (O_2121,N_29882,N_29876);
nand UO_2122 (O_2122,N_29864,N_29882);
nor UO_2123 (O_2123,N_29830,N_29858);
nand UO_2124 (O_2124,N_29860,N_29991);
xor UO_2125 (O_2125,N_29887,N_29956);
xor UO_2126 (O_2126,N_29854,N_29974);
xor UO_2127 (O_2127,N_29928,N_29888);
nor UO_2128 (O_2128,N_29954,N_29898);
nand UO_2129 (O_2129,N_29856,N_29942);
or UO_2130 (O_2130,N_29943,N_29846);
or UO_2131 (O_2131,N_29905,N_29889);
xor UO_2132 (O_2132,N_29865,N_29845);
and UO_2133 (O_2133,N_29999,N_29808);
nand UO_2134 (O_2134,N_29848,N_29837);
nor UO_2135 (O_2135,N_29987,N_29937);
and UO_2136 (O_2136,N_29958,N_29946);
nor UO_2137 (O_2137,N_29855,N_29990);
and UO_2138 (O_2138,N_29850,N_29877);
or UO_2139 (O_2139,N_29818,N_29811);
nand UO_2140 (O_2140,N_29952,N_29849);
or UO_2141 (O_2141,N_29892,N_29806);
nand UO_2142 (O_2142,N_29935,N_29861);
nor UO_2143 (O_2143,N_29835,N_29839);
nand UO_2144 (O_2144,N_29996,N_29899);
nand UO_2145 (O_2145,N_29843,N_29976);
xnor UO_2146 (O_2146,N_29931,N_29966);
or UO_2147 (O_2147,N_29933,N_29815);
or UO_2148 (O_2148,N_29902,N_29923);
and UO_2149 (O_2149,N_29966,N_29975);
and UO_2150 (O_2150,N_29882,N_29934);
nor UO_2151 (O_2151,N_29866,N_29823);
xnor UO_2152 (O_2152,N_29976,N_29884);
xor UO_2153 (O_2153,N_29905,N_29958);
and UO_2154 (O_2154,N_29810,N_29874);
or UO_2155 (O_2155,N_29881,N_29998);
nor UO_2156 (O_2156,N_29914,N_29825);
xnor UO_2157 (O_2157,N_29885,N_29907);
nor UO_2158 (O_2158,N_29885,N_29862);
nor UO_2159 (O_2159,N_29926,N_29915);
nand UO_2160 (O_2160,N_29989,N_29927);
nor UO_2161 (O_2161,N_29873,N_29895);
nand UO_2162 (O_2162,N_29827,N_29994);
or UO_2163 (O_2163,N_29998,N_29868);
nand UO_2164 (O_2164,N_29849,N_29897);
nand UO_2165 (O_2165,N_29806,N_29837);
or UO_2166 (O_2166,N_29962,N_29898);
and UO_2167 (O_2167,N_29914,N_29856);
or UO_2168 (O_2168,N_29896,N_29890);
or UO_2169 (O_2169,N_29998,N_29889);
and UO_2170 (O_2170,N_29875,N_29964);
xnor UO_2171 (O_2171,N_29816,N_29839);
nor UO_2172 (O_2172,N_29860,N_29931);
or UO_2173 (O_2173,N_29868,N_29959);
nand UO_2174 (O_2174,N_29899,N_29883);
or UO_2175 (O_2175,N_29823,N_29857);
and UO_2176 (O_2176,N_29965,N_29909);
nor UO_2177 (O_2177,N_29888,N_29957);
nor UO_2178 (O_2178,N_29998,N_29829);
or UO_2179 (O_2179,N_29944,N_29887);
and UO_2180 (O_2180,N_29838,N_29910);
or UO_2181 (O_2181,N_29931,N_29996);
xor UO_2182 (O_2182,N_29961,N_29800);
or UO_2183 (O_2183,N_29924,N_29936);
nand UO_2184 (O_2184,N_29839,N_29814);
or UO_2185 (O_2185,N_29806,N_29961);
and UO_2186 (O_2186,N_29821,N_29827);
and UO_2187 (O_2187,N_29878,N_29884);
and UO_2188 (O_2188,N_29905,N_29979);
or UO_2189 (O_2189,N_29962,N_29917);
nor UO_2190 (O_2190,N_29976,N_29961);
nand UO_2191 (O_2191,N_29900,N_29926);
nand UO_2192 (O_2192,N_29849,N_29846);
or UO_2193 (O_2193,N_29899,N_29913);
nor UO_2194 (O_2194,N_29817,N_29934);
xnor UO_2195 (O_2195,N_29880,N_29930);
and UO_2196 (O_2196,N_29947,N_29901);
or UO_2197 (O_2197,N_29924,N_29863);
or UO_2198 (O_2198,N_29882,N_29900);
and UO_2199 (O_2199,N_29948,N_29854);
or UO_2200 (O_2200,N_29855,N_29983);
xor UO_2201 (O_2201,N_29811,N_29895);
xnor UO_2202 (O_2202,N_29913,N_29969);
xnor UO_2203 (O_2203,N_29962,N_29889);
and UO_2204 (O_2204,N_29849,N_29938);
nor UO_2205 (O_2205,N_29826,N_29911);
nand UO_2206 (O_2206,N_29966,N_29862);
nor UO_2207 (O_2207,N_29893,N_29855);
xor UO_2208 (O_2208,N_29971,N_29869);
nor UO_2209 (O_2209,N_29870,N_29912);
or UO_2210 (O_2210,N_29937,N_29820);
or UO_2211 (O_2211,N_29997,N_29925);
nor UO_2212 (O_2212,N_29907,N_29861);
nand UO_2213 (O_2213,N_29978,N_29887);
or UO_2214 (O_2214,N_29833,N_29995);
nand UO_2215 (O_2215,N_29833,N_29873);
xor UO_2216 (O_2216,N_29947,N_29906);
and UO_2217 (O_2217,N_29999,N_29872);
xor UO_2218 (O_2218,N_29953,N_29855);
or UO_2219 (O_2219,N_29980,N_29896);
nor UO_2220 (O_2220,N_29807,N_29822);
and UO_2221 (O_2221,N_29979,N_29857);
or UO_2222 (O_2222,N_29958,N_29830);
nand UO_2223 (O_2223,N_29985,N_29944);
nor UO_2224 (O_2224,N_29890,N_29885);
or UO_2225 (O_2225,N_29899,N_29944);
nand UO_2226 (O_2226,N_29933,N_29981);
and UO_2227 (O_2227,N_29853,N_29855);
nand UO_2228 (O_2228,N_29898,N_29895);
xnor UO_2229 (O_2229,N_29957,N_29804);
xnor UO_2230 (O_2230,N_29916,N_29997);
nor UO_2231 (O_2231,N_29828,N_29897);
or UO_2232 (O_2232,N_29846,N_29814);
and UO_2233 (O_2233,N_29864,N_29912);
nand UO_2234 (O_2234,N_29925,N_29880);
nand UO_2235 (O_2235,N_29815,N_29954);
nor UO_2236 (O_2236,N_29899,N_29851);
and UO_2237 (O_2237,N_29877,N_29953);
or UO_2238 (O_2238,N_29848,N_29948);
and UO_2239 (O_2239,N_29878,N_29991);
nor UO_2240 (O_2240,N_29948,N_29949);
and UO_2241 (O_2241,N_29934,N_29834);
nor UO_2242 (O_2242,N_29926,N_29994);
xnor UO_2243 (O_2243,N_29992,N_29945);
nor UO_2244 (O_2244,N_29853,N_29837);
and UO_2245 (O_2245,N_29895,N_29916);
nor UO_2246 (O_2246,N_29963,N_29912);
and UO_2247 (O_2247,N_29932,N_29922);
and UO_2248 (O_2248,N_29802,N_29880);
nand UO_2249 (O_2249,N_29808,N_29952);
or UO_2250 (O_2250,N_29961,N_29861);
xor UO_2251 (O_2251,N_29887,N_29861);
or UO_2252 (O_2252,N_29902,N_29870);
xor UO_2253 (O_2253,N_29903,N_29829);
and UO_2254 (O_2254,N_29942,N_29923);
nand UO_2255 (O_2255,N_29951,N_29868);
nor UO_2256 (O_2256,N_29813,N_29885);
xor UO_2257 (O_2257,N_29882,N_29807);
xor UO_2258 (O_2258,N_29887,N_29819);
xor UO_2259 (O_2259,N_29999,N_29952);
or UO_2260 (O_2260,N_29800,N_29801);
xor UO_2261 (O_2261,N_29811,N_29865);
and UO_2262 (O_2262,N_29903,N_29867);
xor UO_2263 (O_2263,N_29886,N_29905);
or UO_2264 (O_2264,N_29968,N_29838);
nand UO_2265 (O_2265,N_29827,N_29885);
or UO_2266 (O_2266,N_29854,N_29957);
xor UO_2267 (O_2267,N_29901,N_29834);
or UO_2268 (O_2268,N_29995,N_29868);
nand UO_2269 (O_2269,N_29875,N_29828);
or UO_2270 (O_2270,N_29905,N_29833);
and UO_2271 (O_2271,N_29989,N_29944);
or UO_2272 (O_2272,N_29835,N_29817);
and UO_2273 (O_2273,N_29945,N_29836);
or UO_2274 (O_2274,N_29988,N_29912);
and UO_2275 (O_2275,N_29819,N_29896);
and UO_2276 (O_2276,N_29858,N_29962);
and UO_2277 (O_2277,N_29891,N_29959);
or UO_2278 (O_2278,N_29805,N_29877);
and UO_2279 (O_2279,N_29859,N_29913);
nand UO_2280 (O_2280,N_29836,N_29827);
xnor UO_2281 (O_2281,N_29967,N_29899);
nand UO_2282 (O_2282,N_29970,N_29908);
or UO_2283 (O_2283,N_29803,N_29849);
nand UO_2284 (O_2284,N_29861,N_29998);
nor UO_2285 (O_2285,N_29904,N_29838);
or UO_2286 (O_2286,N_29867,N_29877);
nand UO_2287 (O_2287,N_29844,N_29969);
and UO_2288 (O_2288,N_29835,N_29885);
or UO_2289 (O_2289,N_29818,N_29873);
xnor UO_2290 (O_2290,N_29947,N_29891);
or UO_2291 (O_2291,N_29839,N_29933);
nand UO_2292 (O_2292,N_29814,N_29842);
and UO_2293 (O_2293,N_29986,N_29893);
xnor UO_2294 (O_2294,N_29976,N_29890);
xnor UO_2295 (O_2295,N_29898,N_29883);
nand UO_2296 (O_2296,N_29906,N_29857);
xnor UO_2297 (O_2297,N_29935,N_29872);
nor UO_2298 (O_2298,N_29872,N_29954);
nand UO_2299 (O_2299,N_29972,N_29900);
nor UO_2300 (O_2300,N_29870,N_29834);
nand UO_2301 (O_2301,N_29805,N_29803);
or UO_2302 (O_2302,N_29806,N_29963);
xnor UO_2303 (O_2303,N_29899,N_29805);
or UO_2304 (O_2304,N_29879,N_29899);
nor UO_2305 (O_2305,N_29914,N_29831);
xnor UO_2306 (O_2306,N_29847,N_29979);
nor UO_2307 (O_2307,N_29846,N_29815);
xor UO_2308 (O_2308,N_29860,N_29883);
xnor UO_2309 (O_2309,N_29855,N_29845);
or UO_2310 (O_2310,N_29958,N_29841);
or UO_2311 (O_2311,N_29986,N_29883);
or UO_2312 (O_2312,N_29949,N_29871);
and UO_2313 (O_2313,N_29950,N_29847);
nand UO_2314 (O_2314,N_29872,N_29863);
or UO_2315 (O_2315,N_29996,N_29965);
nand UO_2316 (O_2316,N_29891,N_29813);
nor UO_2317 (O_2317,N_29822,N_29882);
and UO_2318 (O_2318,N_29960,N_29999);
xnor UO_2319 (O_2319,N_29922,N_29925);
nand UO_2320 (O_2320,N_29982,N_29915);
nand UO_2321 (O_2321,N_29808,N_29992);
xor UO_2322 (O_2322,N_29821,N_29855);
and UO_2323 (O_2323,N_29800,N_29959);
and UO_2324 (O_2324,N_29919,N_29907);
or UO_2325 (O_2325,N_29885,N_29923);
nand UO_2326 (O_2326,N_29904,N_29995);
or UO_2327 (O_2327,N_29893,N_29809);
nand UO_2328 (O_2328,N_29889,N_29908);
and UO_2329 (O_2329,N_29957,N_29983);
xor UO_2330 (O_2330,N_29809,N_29806);
and UO_2331 (O_2331,N_29993,N_29863);
xnor UO_2332 (O_2332,N_29903,N_29837);
xor UO_2333 (O_2333,N_29971,N_29902);
nand UO_2334 (O_2334,N_29881,N_29957);
nand UO_2335 (O_2335,N_29891,N_29986);
and UO_2336 (O_2336,N_29869,N_29975);
or UO_2337 (O_2337,N_29980,N_29930);
or UO_2338 (O_2338,N_29827,N_29873);
and UO_2339 (O_2339,N_29899,N_29853);
nand UO_2340 (O_2340,N_29805,N_29931);
and UO_2341 (O_2341,N_29812,N_29842);
xnor UO_2342 (O_2342,N_29988,N_29806);
and UO_2343 (O_2343,N_29862,N_29938);
nor UO_2344 (O_2344,N_29984,N_29879);
and UO_2345 (O_2345,N_29900,N_29887);
xor UO_2346 (O_2346,N_29924,N_29881);
nor UO_2347 (O_2347,N_29890,N_29997);
and UO_2348 (O_2348,N_29852,N_29825);
or UO_2349 (O_2349,N_29815,N_29923);
xnor UO_2350 (O_2350,N_29815,N_29948);
xor UO_2351 (O_2351,N_29802,N_29956);
nor UO_2352 (O_2352,N_29944,N_29814);
nor UO_2353 (O_2353,N_29903,N_29998);
xnor UO_2354 (O_2354,N_29881,N_29969);
nor UO_2355 (O_2355,N_29881,N_29826);
nor UO_2356 (O_2356,N_29959,N_29980);
and UO_2357 (O_2357,N_29898,N_29942);
and UO_2358 (O_2358,N_29872,N_29916);
nand UO_2359 (O_2359,N_29989,N_29855);
or UO_2360 (O_2360,N_29807,N_29877);
and UO_2361 (O_2361,N_29857,N_29918);
xor UO_2362 (O_2362,N_29930,N_29846);
nor UO_2363 (O_2363,N_29880,N_29828);
nand UO_2364 (O_2364,N_29801,N_29870);
xnor UO_2365 (O_2365,N_29835,N_29887);
nor UO_2366 (O_2366,N_29851,N_29966);
nand UO_2367 (O_2367,N_29911,N_29832);
xor UO_2368 (O_2368,N_29914,N_29861);
and UO_2369 (O_2369,N_29889,N_29979);
or UO_2370 (O_2370,N_29893,N_29947);
nand UO_2371 (O_2371,N_29846,N_29840);
nand UO_2372 (O_2372,N_29889,N_29966);
and UO_2373 (O_2373,N_29882,N_29878);
nor UO_2374 (O_2374,N_29947,N_29885);
nand UO_2375 (O_2375,N_29889,N_29869);
or UO_2376 (O_2376,N_29834,N_29914);
xnor UO_2377 (O_2377,N_29919,N_29960);
and UO_2378 (O_2378,N_29907,N_29968);
or UO_2379 (O_2379,N_29932,N_29996);
nand UO_2380 (O_2380,N_29834,N_29817);
nor UO_2381 (O_2381,N_29951,N_29891);
and UO_2382 (O_2382,N_29917,N_29938);
nand UO_2383 (O_2383,N_29868,N_29808);
or UO_2384 (O_2384,N_29958,N_29930);
or UO_2385 (O_2385,N_29830,N_29896);
and UO_2386 (O_2386,N_29887,N_29950);
xor UO_2387 (O_2387,N_29891,N_29838);
and UO_2388 (O_2388,N_29937,N_29931);
nand UO_2389 (O_2389,N_29969,N_29840);
or UO_2390 (O_2390,N_29917,N_29914);
or UO_2391 (O_2391,N_29979,N_29806);
nor UO_2392 (O_2392,N_29858,N_29954);
nand UO_2393 (O_2393,N_29920,N_29851);
nand UO_2394 (O_2394,N_29897,N_29991);
or UO_2395 (O_2395,N_29897,N_29952);
nor UO_2396 (O_2396,N_29917,N_29873);
nor UO_2397 (O_2397,N_29857,N_29815);
xor UO_2398 (O_2398,N_29832,N_29854);
nor UO_2399 (O_2399,N_29924,N_29990);
and UO_2400 (O_2400,N_29966,N_29976);
nand UO_2401 (O_2401,N_29910,N_29923);
nor UO_2402 (O_2402,N_29850,N_29911);
nor UO_2403 (O_2403,N_29931,N_29868);
or UO_2404 (O_2404,N_29977,N_29973);
or UO_2405 (O_2405,N_29977,N_29846);
and UO_2406 (O_2406,N_29989,N_29949);
nor UO_2407 (O_2407,N_29852,N_29965);
xor UO_2408 (O_2408,N_29985,N_29938);
nor UO_2409 (O_2409,N_29929,N_29847);
xnor UO_2410 (O_2410,N_29852,N_29918);
and UO_2411 (O_2411,N_29912,N_29853);
nor UO_2412 (O_2412,N_29980,N_29865);
and UO_2413 (O_2413,N_29921,N_29877);
and UO_2414 (O_2414,N_29888,N_29820);
nor UO_2415 (O_2415,N_29953,N_29835);
nor UO_2416 (O_2416,N_29966,N_29877);
nor UO_2417 (O_2417,N_29993,N_29908);
or UO_2418 (O_2418,N_29948,N_29927);
xnor UO_2419 (O_2419,N_29823,N_29812);
nand UO_2420 (O_2420,N_29931,N_29838);
nand UO_2421 (O_2421,N_29880,N_29865);
and UO_2422 (O_2422,N_29829,N_29853);
and UO_2423 (O_2423,N_29908,N_29968);
and UO_2424 (O_2424,N_29830,N_29842);
nand UO_2425 (O_2425,N_29812,N_29989);
or UO_2426 (O_2426,N_29947,N_29952);
nand UO_2427 (O_2427,N_29867,N_29813);
or UO_2428 (O_2428,N_29856,N_29972);
and UO_2429 (O_2429,N_29915,N_29963);
nor UO_2430 (O_2430,N_29851,N_29986);
or UO_2431 (O_2431,N_29869,N_29943);
or UO_2432 (O_2432,N_29978,N_29886);
and UO_2433 (O_2433,N_29999,N_29924);
nor UO_2434 (O_2434,N_29987,N_29983);
or UO_2435 (O_2435,N_29979,N_29965);
nand UO_2436 (O_2436,N_29974,N_29985);
nand UO_2437 (O_2437,N_29904,N_29945);
nor UO_2438 (O_2438,N_29831,N_29895);
and UO_2439 (O_2439,N_29870,N_29951);
nand UO_2440 (O_2440,N_29848,N_29905);
nand UO_2441 (O_2441,N_29987,N_29887);
and UO_2442 (O_2442,N_29801,N_29996);
xnor UO_2443 (O_2443,N_29825,N_29966);
and UO_2444 (O_2444,N_29830,N_29913);
xor UO_2445 (O_2445,N_29878,N_29806);
or UO_2446 (O_2446,N_29838,N_29895);
and UO_2447 (O_2447,N_29959,N_29950);
nor UO_2448 (O_2448,N_29850,N_29816);
and UO_2449 (O_2449,N_29915,N_29875);
nor UO_2450 (O_2450,N_29888,N_29860);
nand UO_2451 (O_2451,N_29840,N_29824);
nor UO_2452 (O_2452,N_29934,N_29819);
or UO_2453 (O_2453,N_29824,N_29922);
and UO_2454 (O_2454,N_29885,N_29884);
and UO_2455 (O_2455,N_29941,N_29826);
and UO_2456 (O_2456,N_29982,N_29816);
nand UO_2457 (O_2457,N_29848,N_29872);
nor UO_2458 (O_2458,N_29952,N_29805);
or UO_2459 (O_2459,N_29888,N_29819);
or UO_2460 (O_2460,N_29994,N_29900);
nand UO_2461 (O_2461,N_29860,N_29955);
nand UO_2462 (O_2462,N_29986,N_29957);
nand UO_2463 (O_2463,N_29909,N_29808);
nand UO_2464 (O_2464,N_29934,N_29807);
xor UO_2465 (O_2465,N_29873,N_29931);
or UO_2466 (O_2466,N_29891,N_29888);
xnor UO_2467 (O_2467,N_29967,N_29972);
nand UO_2468 (O_2468,N_29835,N_29954);
xor UO_2469 (O_2469,N_29967,N_29805);
or UO_2470 (O_2470,N_29829,N_29994);
nand UO_2471 (O_2471,N_29895,N_29915);
and UO_2472 (O_2472,N_29956,N_29907);
nand UO_2473 (O_2473,N_29826,N_29803);
and UO_2474 (O_2474,N_29939,N_29931);
xnor UO_2475 (O_2475,N_29991,N_29881);
nand UO_2476 (O_2476,N_29948,N_29936);
xor UO_2477 (O_2477,N_29999,N_29985);
or UO_2478 (O_2478,N_29899,N_29817);
nand UO_2479 (O_2479,N_29826,N_29923);
nor UO_2480 (O_2480,N_29875,N_29968);
nor UO_2481 (O_2481,N_29961,N_29924);
nand UO_2482 (O_2482,N_29849,N_29985);
nand UO_2483 (O_2483,N_29957,N_29813);
nand UO_2484 (O_2484,N_29800,N_29850);
nor UO_2485 (O_2485,N_29831,N_29866);
nor UO_2486 (O_2486,N_29891,N_29971);
xor UO_2487 (O_2487,N_29854,N_29849);
nand UO_2488 (O_2488,N_29887,N_29966);
nor UO_2489 (O_2489,N_29973,N_29875);
and UO_2490 (O_2490,N_29821,N_29869);
and UO_2491 (O_2491,N_29895,N_29981);
nand UO_2492 (O_2492,N_29890,N_29847);
or UO_2493 (O_2493,N_29916,N_29882);
or UO_2494 (O_2494,N_29858,N_29961);
or UO_2495 (O_2495,N_29941,N_29991);
or UO_2496 (O_2496,N_29882,N_29952);
nor UO_2497 (O_2497,N_29814,N_29864);
nand UO_2498 (O_2498,N_29903,N_29982);
and UO_2499 (O_2499,N_29840,N_29890);
nor UO_2500 (O_2500,N_29869,N_29879);
nor UO_2501 (O_2501,N_29930,N_29897);
or UO_2502 (O_2502,N_29836,N_29922);
nand UO_2503 (O_2503,N_29863,N_29874);
and UO_2504 (O_2504,N_29952,N_29841);
and UO_2505 (O_2505,N_29917,N_29833);
nor UO_2506 (O_2506,N_29998,N_29837);
or UO_2507 (O_2507,N_29921,N_29838);
nor UO_2508 (O_2508,N_29922,N_29841);
or UO_2509 (O_2509,N_29955,N_29869);
xor UO_2510 (O_2510,N_29909,N_29878);
and UO_2511 (O_2511,N_29822,N_29849);
nand UO_2512 (O_2512,N_29987,N_29873);
xnor UO_2513 (O_2513,N_29898,N_29807);
and UO_2514 (O_2514,N_29966,N_29853);
and UO_2515 (O_2515,N_29881,N_29893);
nand UO_2516 (O_2516,N_29840,N_29902);
and UO_2517 (O_2517,N_29926,N_29841);
or UO_2518 (O_2518,N_29900,N_29820);
or UO_2519 (O_2519,N_29932,N_29934);
and UO_2520 (O_2520,N_29935,N_29885);
nand UO_2521 (O_2521,N_29904,N_29853);
xnor UO_2522 (O_2522,N_29827,N_29890);
or UO_2523 (O_2523,N_29864,N_29953);
and UO_2524 (O_2524,N_29956,N_29804);
nor UO_2525 (O_2525,N_29809,N_29976);
nor UO_2526 (O_2526,N_29948,N_29933);
nor UO_2527 (O_2527,N_29972,N_29862);
nor UO_2528 (O_2528,N_29802,N_29944);
nor UO_2529 (O_2529,N_29804,N_29960);
or UO_2530 (O_2530,N_29971,N_29857);
nand UO_2531 (O_2531,N_29974,N_29826);
and UO_2532 (O_2532,N_29992,N_29846);
or UO_2533 (O_2533,N_29861,N_29878);
nand UO_2534 (O_2534,N_29823,N_29875);
and UO_2535 (O_2535,N_29987,N_29855);
or UO_2536 (O_2536,N_29995,N_29888);
nand UO_2537 (O_2537,N_29929,N_29837);
nor UO_2538 (O_2538,N_29960,N_29850);
xor UO_2539 (O_2539,N_29878,N_29929);
nand UO_2540 (O_2540,N_29871,N_29981);
or UO_2541 (O_2541,N_29894,N_29901);
and UO_2542 (O_2542,N_29938,N_29901);
or UO_2543 (O_2543,N_29802,N_29937);
xnor UO_2544 (O_2544,N_29877,N_29868);
xor UO_2545 (O_2545,N_29873,N_29928);
nand UO_2546 (O_2546,N_29874,N_29861);
or UO_2547 (O_2547,N_29960,N_29830);
nand UO_2548 (O_2548,N_29961,N_29834);
nand UO_2549 (O_2549,N_29917,N_29886);
and UO_2550 (O_2550,N_29998,N_29865);
nor UO_2551 (O_2551,N_29944,N_29858);
and UO_2552 (O_2552,N_29808,N_29977);
xor UO_2553 (O_2553,N_29952,N_29908);
xor UO_2554 (O_2554,N_29859,N_29839);
xor UO_2555 (O_2555,N_29889,N_29860);
xnor UO_2556 (O_2556,N_29901,N_29908);
and UO_2557 (O_2557,N_29998,N_29917);
xor UO_2558 (O_2558,N_29960,N_29962);
or UO_2559 (O_2559,N_29938,N_29986);
nand UO_2560 (O_2560,N_29934,N_29865);
nor UO_2561 (O_2561,N_29920,N_29959);
nor UO_2562 (O_2562,N_29839,N_29824);
and UO_2563 (O_2563,N_29934,N_29908);
nand UO_2564 (O_2564,N_29996,N_29889);
xor UO_2565 (O_2565,N_29896,N_29858);
or UO_2566 (O_2566,N_29824,N_29884);
nand UO_2567 (O_2567,N_29936,N_29901);
or UO_2568 (O_2568,N_29971,N_29954);
or UO_2569 (O_2569,N_29841,N_29866);
or UO_2570 (O_2570,N_29940,N_29923);
or UO_2571 (O_2571,N_29868,N_29989);
nor UO_2572 (O_2572,N_29864,N_29976);
xor UO_2573 (O_2573,N_29866,N_29920);
nand UO_2574 (O_2574,N_29935,N_29880);
nand UO_2575 (O_2575,N_29996,N_29883);
nor UO_2576 (O_2576,N_29910,N_29937);
nor UO_2577 (O_2577,N_29999,N_29821);
nor UO_2578 (O_2578,N_29921,N_29915);
xor UO_2579 (O_2579,N_29874,N_29839);
and UO_2580 (O_2580,N_29919,N_29923);
or UO_2581 (O_2581,N_29958,N_29965);
nor UO_2582 (O_2582,N_29830,N_29998);
xnor UO_2583 (O_2583,N_29826,N_29975);
and UO_2584 (O_2584,N_29914,N_29986);
xor UO_2585 (O_2585,N_29994,N_29944);
nor UO_2586 (O_2586,N_29830,N_29895);
xor UO_2587 (O_2587,N_29853,N_29905);
nand UO_2588 (O_2588,N_29900,N_29829);
nand UO_2589 (O_2589,N_29892,N_29966);
and UO_2590 (O_2590,N_29865,N_29968);
and UO_2591 (O_2591,N_29845,N_29893);
nand UO_2592 (O_2592,N_29918,N_29901);
xor UO_2593 (O_2593,N_29942,N_29815);
and UO_2594 (O_2594,N_29894,N_29861);
nand UO_2595 (O_2595,N_29806,N_29818);
nor UO_2596 (O_2596,N_29924,N_29843);
and UO_2597 (O_2597,N_29925,N_29834);
or UO_2598 (O_2598,N_29940,N_29947);
xor UO_2599 (O_2599,N_29870,N_29940);
nor UO_2600 (O_2600,N_29935,N_29977);
nand UO_2601 (O_2601,N_29818,N_29824);
and UO_2602 (O_2602,N_29901,N_29893);
xnor UO_2603 (O_2603,N_29843,N_29814);
and UO_2604 (O_2604,N_29817,N_29913);
nand UO_2605 (O_2605,N_29874,N_29832);
and UO_2606 (O_2606,N_29824,N_29965);
nand UO_2607 (O_2607,N_29938,N_29906);
nor UO_2608 (O_2608,N_29811,N_29944);
nand UO_2609 (O_2609,N_29915,N_29930);
nor UO_2610 (O_2610,N_29926,N_29821);
or UO_2611 (O_2611,N_29935,N_29874);
nor UO_2612 (O_2612,N_29998,N_29822);
xor UO_2613 (O_2613,N_29994,N_29840);
or UO_2614 (O_2614,N_29965,N_29914);
nand UO_2615 (O_2615,N_29826,N_29926);
nand UO_2616 (O_2616,N_29900,N_29973);
nor UO_2617 (O_2617,N_29854,N_29820);
nand UO_2618 (O_2618,N_29909,N_29953);
or UO_2619 (O_2619,N_29824,N_29955);
or UO_2620 (O_2620,N_29977,N_29824);
xnor UO_2621 (O_2621,N_29806,N_29965);
nor UO_2622 (O_2622,N_29931,N_29983);
nand UO_2623 (O_2623,N_29902,N_29991);
nand UO_2624 (O_2624,N_29892,N_29986);
xor UO_2625 (O_2625,N_29910,N_29951);
xnor UO_2626 (O_2626,N_29808,N_29883);
nor UO_2627 (O_2627,N_29900,N_29883);
xnor UO_2628 (O_2628,N_29973,N_29921);
nor UO_2629 (O_2629,N_29820,N_29944);
nor UO_2630 (O_2630,N_29968,N_29937);
and UO_2631 (O_2631,N_29897,N_29816);
xor UO_2632 (O_2632,N_29881,N_29994);
or UO_2633 (O_2633,N_29818,N_29874);
or UO_2634 (O_2634,N_29969,N_29899);
and UO_2635 (O_2635,N_29817,N_29887);
nor UO_2636 (O_2636,N_29961,N_29822);
nand UO_2637 (O_2637,N_29958,N_29847);
nor UO_2638 (O_2638,N_29979,N_29918);
nor UO_2639 (O_2639,N_29866,N_29802);
or UO_2640 (O_2640,N_29802,N_29868);
and UO_2641 (O_2641,N_29938,N_29934);
or UO_2642 (O_2642,N_29892,N_29985);
xor UO_2643 (O_2643,N_29915,N_29917);
and UO_2644 (O_2644,N_29832,N_29845);
nand UO_2645 (O_2645,N_29952,N_29975);
nor UO_2646 (O_2646,N_29825,N_29963);
and UO_2647 (O_2647,N_29943,N_29928);
nand UO_2648 (O_2648,N_29829,N_29877);
or UO_2649 (O_2649,N_29846,N_29972);
and UO_2650 (O_2650,N_29955,N_29806);
and UO_2651 (O_2651,N_29867,N_29911);
nand UO_2652 (O_2652,N_29852,N_29905);
nor UO_2653 (O_2653,N_29884,N_29997);
xor UO_2654 (O_2654,N_29809,N_29955);
nand UO_2655 (O_2655,N_29948,N_29980);
nand UO_2656 (O_2656,N_29953,N_29890);
nor UO_2657 (O_2657,N_29840,N_29966);
xor UO_2658 (O_2658,N_29803,N_29934);
and UO_2659 (O_2659,N_29975,N_29946);
or UO_2660 (O_2660,N_29929,N_29959);
nand UO_2661 (O_2661,N_29872,N_29964);
xnor UO_2662 (O_2662,N_29840,N_29860);
or UO_2663 (O_2663,N_29912,N_29886);
and UO_2664 (O_2664,N_29958,N_29912);
xor UO_2665 (O_2665,N_29908,N_29977);
and UO_2666 (O_2666,N_29808,N_29967);
nand UO_2667 (O_2667,N_29974,N_29981);
or UO_2668 (O_2668,N_29890,N_29980);
or UO_2669 (O_2669,N_29982,N_29968);
nor UO_2670 (O_2670,N_29855,N_29803);
or UO_2671 (O_2671,N_29925,N_29827);
and UO_2672 (O_2672,N_29935,N_29805);
nand UO_2673 (O_2673,N_29908,N_29886);
or UO_2674 (O_2674,N_29995,N_29979);
nor UO_2675 (O_2675,N_29959,N_29846);
or UO_2676 (O_2676,N_29917,N_29960);
xnor UO_2677 (O_2677,N_29826,N_29994);
and UO_2678 (O_2678,N_29978,N_29874);
nor UO_2679 (O_2679,N_29829,N_29918);
nor UO_2680 (O_2680,N_29902,N_29953);
or UO_2681 (O_2681,N_29965,N_29859);
xnor UO_2682 (O_2682,N_29983,N_29819);
or UO_2683 (O_2683,N_29949,N_29872);
or UO_2684 (O_2684,N_29807,N_29843);
nor UO_2685 (O_2685,N_29891,N_29809);
or UO_2686 (O_2686,N_29894,N_29939);
nor UO_2687 (O_2687,N_29872,N_29901);
and UO_2688 (O_2688,N_29869,N_29922);
nand UO_2689 (O_2689,N_29975,N_29916);
or UO_2690 (O_2690,N_29971,N_29965);
nand UO_2691 (O_2691,N_29878,N_29972);
xor UO_2692 (O_2692,N_29945,N_29856);
nor UO_2693 (O_2693,N_29985,N_29990);
nor UO_2694 (O_2694,N_29976,N_29917);
nor UO_2695 (O_2695,N_29861,N_29965);
or UO_2696 (O_2696,N_29962,N_29961);
or UO_2697 (O_2697,N_29928,N_29931);
and UO_2698 (O_2698,N_29952,N_29949);
nor UO_2699 (O_2699,N_29826,N_29945);
xnor UO_2700 (O_2700,N_29984,N_29977);
nor UO_2701 (O_2701,N_29920,N_29961);
nor UO_2702 (O_2702,N_29946,N_29919);
xnor UO_2703 (O_2703,N_29947,N_29800);
xnor UO_2704 (O_2704,N_29892,N_29944);
xor UO_2705 (O_2705,N_29870,N_29956);
or UO_2706 (O_2706,N_29933,N_29903);
nand UO_2707 (O_2707,N_29812,N_29921);
xnor UO_2708 (O_2708,N_29871,N_29968);
nor UO_2709 (O_2709,N_29982,N_29956);
nand UO_2710 (O_2710,N_29967,N_29873);
xor UO_2711 (O_2711,N_29887,N_29857);
nand UO_2712 (O_2712,N_29963,N_29895);
and UO_2713 (O_2713,N_29949,N_29979);
nor UO_2714 (O_2714,N_29822,N_29972);
xor UO_2715 (O_2715,N_29897,N_29818);
nor UO_2716 (O_2716,N_29803,N_29973);
and UO_2717 (O_2717,N_29811,N_29870);
nand UO_2718 (O_2718,N_29849,N_29986);
nor UO_2719 (O_2719,N_29877,N_29948);
or UO_2720 (O_2720,N_29952,N_29871);
nor UO_2721 (O_2721,N_29920,N_29832);
or UO_2722 (O_2722,N_29810,N_29942);
nor UO_2723 (O_2723,N_29959,N_29884);
or UO_2724 (O_2724,N_29853,N_29890);
xnor UO_2725 (O_2725,N_29997,N_29977);
nor UO_2726 (O_2726,N_29945,N_29937);
and UO_2727 (O_2727,N_29946,N_29981);
nor UO_2728 (O_2728,N_29993,N_29917);
or UO_2729 (O_2729,N_29956,N_29923);
and UO_2730 (O_2730,N_29801,N_29985);
xor UO_2731 (O_2731,N_29963,N_29976);
and UO_2732 (O_2732,N_29843,N_29969);
or UO_2733 (O_2733,N_29893,N_29944);
xnor UO_2734 (O_2734,N_29913,N_29959);
nor UO_2735 (O_2735,N_29865,N_29970);
nor UO_2736 (O_2736,N_29826,N_29804);
nand UO_2737 (O_2737,N_29987,N_29927);
nor UO_2738 (O_2738,N_29962,N_29952);
and UO_2739 (O_2739,N_29892,N_29953);
xor UO_2740 (O_2740,N_29814,N_29888);
or UO_2741 (O_2741,N_29947,N_29807);
nor UO_2742 (O_2742,N_29988,N_29823);
and UO_2743 (O_2743,N_29919,N_29903);
nor UO_2744 (O_2744,N_29826,N_29836);
and UO_2745 (O_2745,N_29848,N_29939);
nor UO_2746 (O_2746,N_29967,N_29888);
or UO_2747 (O_2747,N_29948,N_29844);
nand UO_2748 (O_2748,N_29895,N_29849);
and UO_2749 (O_2749,N_29907,N_29819);
nor UO_2750 (O_2750,N_29969,N_29876);
xor UO_2751 (O_2751,N_29937,N_29810);
and UO_2752 (O_2752,N_29993,N_29820);
nor UO_2753 (O_2753,N_29900,N_29976);
or UO_2754 (O_2754,N_29985,N_29981);
and UO_2755 (O_2755,N_29823,N_29966);
and UO_2756 (O_2756,N_29986,N_29867);
xnor UO_2757 (O_2757,N_29942,N_29907);
or UO_2758 (O_2758,N_29947,N_29937);
nor UO_2759 (O_2759,N_29890,N_29964);
nor UO_2760 (O_2760,N_29806,N_29848);
nand UO_2761 (O_2761,N_29972,N_29984);
and UO_2762 (O_2762,N_29804,N_29814);
xor UO_2763 (O_2763,N_29885,N_29902);
xnor UO_2764 (O_2764,N_29925,N_29988);
xnor UO_2765 (O_2765,N_29890,N_29848);
or UO_2766 (O_2766,N_29820,N_29802);
nand UO_2767 (O_2767,N_29942,N_29883);
nand UO_2768 (O_2768,N_29985,N_29925);
nor UO_2769 (O_2769,N_29971,N_29948);
or UO_2770 (O_2770,N_29933,N_29893);
nand UO_2771 (O_2771,N_29842,N_29849);
and UO_2772 (O_2772,N_29874,N_29990);
nor UO_2773 (O_2773,N_29963,N_29838);
and UO_2774 (O_2774,N_29975,N_29956);
nand UO_2775 (O_2775,N_29837,N_29996);
and UO_2776 (O_2776,N_29829,N_29968);
nor UO_2777 (O_2777,N_29879,N_29980);
nor UO_2778 (O_2778,N_29916,N_29850);
nand UO_2779 (O_2779,N_29880,N_29929);
and UO_2780 (O_2780,N_29803,N_29877);
nor UO_2781 (O_2781,N_29892,N_29825);
nor UO_2782 (O_2782,N_29840,N_29903);
xor UO_2783 (O_2783,N_29963,N_29802);
xor UO_2784 (O_2784,N_29827,N_29907);
nand UO_2785 (O_2785,N_29954,N_29983);
and UO_2786 (O_2786,N_29812,N_29868);
xor UO_2787 (O_2787,N_29928,N_29923);
nor UO_2788 (O_2788,N_29876,N_29830);
xor UO_2789 (O_2789,N_29878,N_29948);
or UO_2790 (O_2790,N_29998,N_29985);
xnor UO_2791 (O_2791,N_29989,N_29985);
nor UO_2792 (O_2792,N_29909,N_29836);
xnor UO_2793 (O_2793,N_29992,N_29910);
nand UO_2794 (O_2794,N_29960,N_29808);
or UO_2795 (O_2795,N_29812,N_29852);
and UO_2796 (O_2796,N_29906,N_29934);
xnor UO_2797 (O_2797,N_29900,N_29988);
xnor UO_2798 (O_2798,N_29817,N_29902);
and UO_2799 (O_2799,N_29909,N_29802);
nor UO_2800 (O_2800,N_29844,N_29982);
and UO_2801 (O_2801,N_29995,N_29877);
and UO_2802 (O_2802,N_29838,N_29874);
nand UO_2803 (O_2803,N_29826,N_29950);
and UO_2804 (O_2804,N_29965,N_29919);
or UO_2805 (O_2805,N_29967,N_29816);
nor UO_2806 (O_2806,N_29883,N_29940);
or UO_2807 (O_2807,N_29961,N_29922);
or UO_2808 (O_2808,N_29889,N_29888);
or UO_2809 (O_2809,N_29914,N_29805);
xor UO_2810 (O_2810,N_29959,N_29960);
nor UO_2811 (O_2811,N_29906,N_29884);
or UO_2812 (O_2812,N_29916,N_29999);
or UO_2813 (O_2813,N_29819,N_29959);
and UO_2814 (O_2814,N_29947,N_29902);
nand UO_2815 (O_2815,N_29901,N_29960);
and UO_2816 (O_2816,N_29904,N_29998);
and UO_2817 (O_2817,N_29858,N_29862);
nor UO_2818 (O_2818,N_29896,N_29861);
xor UO_2819 (O_2819,N_29950,N_29864);
and UO_2820 (O_2820,N_29927,N_29871);
nand UO_2821 (O_2821,N_29895,N_29832);
and UO_2822 (O_2822,N_29950,N_29867);
nand UO_2823 (O_2823,N_29823,N_29815);
and UO_2824 (O_2824,N_29827,N_29939);
or UO_2825 (O_2825,N_29914,N_29963);
xor UO_2826 (O_2826,N_29916,N_29837);
or UO_2827 (O_2827,N_29844,N_29921);
nor UO_2828 (O_2828,N_29912,N_29997);
xnor UO_2829 (O_2829,N_29907,N_29910);
nand UO_2830 (O_2830,N_29985,N_29862);
nand UO_2831 (O_2831,N_29909,N_29823);
nand UO_2832 (O_2832,N_29997,N_29978);
and UO_2833 (O_2833,N_29823,N_29873);
xor UO_2834 (O_2834,N_29891,N_29849);
nor UO_2835 (O_2835,N_29849,N_29994);
nand UO_2836 (O_2836,N_29806,N_29983);
xnor UO_2837 (O_2837,N_29918,N_29917);
nand UO_2838 (O_2838,N_29800,N_29867);
nor UO_2839 (O_2839,N_29823,N_29808);
and UO_2840 (O_2840,N_29826,N_29913);
or UO_2841 (O_2841,N_29832,N_29873);
and UO_2842 (O_2842,N_29813,N_29849);
or UO_2843 (O_2843,N_29883,N_29905);
xnor UO_2844 (O_2844,N_29973,N_29993);
and UO_2845 (O_2845,N_29821,N_29950);
and UO_2846 (O_2846,N_29843,N_29890);
or UO_2847 (O_2847,N_29998,N_29925);
or UO_2848 (O_2848,N_29852,N_29938);
nor UO_2849 (O_2849,N_29847,N_29855);
xnor UO_2850 (O_2850,N_29835,N_29926);
xor UO_2851 (O_2851,N_29903,N_29979);
xor UO_2852 (O_2852,N_29812,N_29960);
nand UO_2853 (O_2853,N_29908,N_29918);
and UO_2854 (O_2854,N_29905,N_29954);
and UO_2855 (O_2855,N_29911,N_29915);
nor UO_2856 (O_2856,N_29805,N_29814);
nor UO_2857 (O_2857,N_29967,N_29988);
nand UO_2858 (O_2858,N_29875,N_29998);
or UO_2859 (O_2859,N_29995,N_29832);
xor UO_2860 (O_2860,N_29811,N_29920);
nor UO_2861 (O_2861,N_29895,N_29952);
xnor UO_2862 (O_2862,N_29874,N_29902);
or UO_2863 (O_2863,N_29834,N_29815);
nor UO_2864 (O_2864,N_29991,N_29995);
nand UO_2865 (O_2865,N_29850,N_29985);
nand UO_2866 (O_2866,N_29834,N_29867);
nand UO_2867 (O_2867,N_29895,N_29968);
or UO_2868 (O_2868,N_29994,N_29899);
or UO_2869 (O_2869,N_29924,N_29849);
nand UO_2870 (O_2870,N_29838,N_29903);
and UO_2871 (O_2871,N_29946,N_29873);
or UO_2872 (O_2872,N_29984,N_29906);
nor UO_2873 (O_2873,N_29997,N_29848);
nor UO_2874 (O_2874,N_29887,N_29852);
xnor UO_2875 (O_2875,N_29874,N_29942);
and UO_2876 (O_2876,N_29926,N_29982);
nand UO_2877 (O_2877,N_29931,N_29943);
nand UO_2878 (O_2878,N_29912,N_29849);
nand UO_2879 (O_2879,N_29861,N_29834);
and UO_2880 (O_2880,N_29917,N_29889);
xor UO_2881 (O_2881,N_29936,N_29828);
or UO_2882 (O_2882,N_29830,N_29961);
xor UO_2883 (O_2883,N_29950,N_29803);
or UO_2884 (O_2884,N_29838,N_29984);
or UO_2885 (O_2885,N_29810,N_29925);
and UO_2886 (O_2886,N_29899,N_29991);
nor UO_2887 (O_2887,N_29834,N_29998);
xnor UO_2888 (O_2888,N_29892,N_29883);
and UO_2889 (O_2889,N_29918,N_29948);
nand UO_2890 (O_2890,N_29981,N_29920);
nand UO_2891 (O_2891,N_29906,N_29921);
and UO_2892 (O_2892,N_29827,N_29800);
nand UO_2893 (O_2893,N_29929,N_29981);
and UO_2894 (O_2894,N_29813,N_29904);
xnor UO_2895 (O_2895,N_29840,N_29942);
and UO_2896 (O_2896,N_29954,N_29959);
nor UO_2897 (O_2897,N_29844,N_29839);
or UO_2898 (O_2898,N_29869,N_29808);
xnor UO_2899 (O_2899,N_29960,N_29825);
and UO_2900 (O_2900,N_29889,N_29912);
xnor UO_2901 (O_2901,N_29868,N_29865);
nand UO_2902 (O_2902,N_29993,N_29860);
nand UO_2903 (O_2903,N_29936,N_29986);
and UO_2904 (O_2904,N_29885,N_29854);
nand UO_2905 (O_2905,N_29951,N_29837);
or UO_2906 (O_2906,N_29921,N_29876);
nand UO_2907 (O_2907,N_29890,N_29831);
xor UO_2908 (O_2908,N_29921,N_29813);
or UO_2909 (O_2909,N_29811,N_29927);
or UO_2910 (O_2910,N_29989,N_29956);
and UO_2911 (O_2911,N_29803,N_29921);
nand UO_2912 (O_2912,N_29902,N_29988);
nor UO_2913 (O_2913,N_29840,N_29856);
nor UO_2914 (O_2914,N_29851,N_29885);
nor UO_2915 (O_2915,N_29921,N_29824);
xnor UO_2916 (O_2916,N_29831,N_29822);
and UO_2917 (O_2917,N_29974,N_29838);
nor UO_2918 (O_2918,N_29839,N_29810);
or UO_2919 (O_2919,N_29937,N_29979);
or UO_2920 (O_2920,N_29916,N_29972);
xor UO_2921 (O_2921,N_29957,N_29848);
xnor UO_2922 (O_2922,N_29971,N_29966);
or UO_2923 (O_2923,N_29941,N_29877);
nor UO_2924 (O_2924,N_29927,N_29998);
nand UO_2925 (O_2925,N_29999,N_29805);
and UO_2926 (O_2926,N_29958,N_29813);
or UO_2927 (O_2927,N_29809,N_29852);
xnor UO_2928 (O_2928,N_29891,N_29993);
or UO_2929 (O_2929,N_29876,N_29901);
nand UO_2930 (O_2930,N_29822,N_29858);
nor UO_2931 (O_2931,N_29966,N_29829);
nor UO_2932 (O_2932,N_29819,N_29805);
nor UO_2933 (O_2933,N_29844,N_29970);
or UO_2934 (O_2934,N_29998,N_29993);
xor UO_2935 (O_2935,N_29923,N_29820);
nor UO_2936 (O_2936,N_29835,N_29942);
nor UO_2937 (O_2937,N_29982,N_29906);
nand UO_2938 (O_2938,N_29928,N_29880);
or UO_2939 (O_2939,N_29931,N_29892);
or UO_2940 (O_2940,N_29856,N_29971);
nand UO_2941 (O_2941,N_29945,N_29898);
nor UO_2942 (O_2942,N_29857,N_29992);
xnor UO_2943 (O_2943,N_29969,N_29992);
xor UO_2944 (O_2944,N_29850,N_29842);
or UO_2945 (O_2945,N_29929,N_29801);
nor UO_2946 (O_2946,N_29966,N_29801);
or UO_2947 (O_2947,N_29938,N_29820);
or UO_2948 (O_2948,N_29814,N_29817);
nand UO_2949 (O_2949,N_29886,N_29913);
xnor UO_2950 (O_2950,N_29899,N_29844);
nor UO_2951 (O_2951,N_29925,N_29848);
xor UO_2952 (O_2952,N_29978,N_29857);
xor UO_2953 (O_2953,N_29941,N_29919);
xor UO_2954 (O_2954,N_29919,N_29845);
xor UO_2955 (O_2955,N_29960,N_29837);
and UO_2956 (O_2956,N_29820,N_29915);
xor UO_2957 (O_2957,N_29998,N_29890);
nor UO_2958 (O_2958,N_29915,N_29981);
and UO_2959 (O_2959,N_29917,N_29949);
nand UO_2960 (O_2960,N_29979,N_29935);
nand UO_2961 (O_2961,N_29901,N_29804);
nand UO_2962 (O_2962,N_29927,N_29937);
xnor UO_2963 (O_2963,N_29803,N_29866);
or UO_2964 (O_2964,N_29812,N_29843);
and UO_2965 (O_2965,N_29835,N_29889);
or UO_2966 (O_2966,N_29921,N_29841);
nand UO_2967 (O_2967,N_29893,N_29971);
nor UO_2968 (O_2968,N_29803,N_29915);
nand UO_2969 (O_2969,N_29865,N_29936);
nand UO_2970 (O_2970,N_29961,N_29978);
nand UO_2971 (O_2971,N_29842,N_29998);
nor UO_2972 (O_2972,N_29938,N_29961);
and UO_2973 (O_2973,N_29856,N_29818);
xnor UO_2974 (O_2974,N_29970,N_29939);
xor UO_2975 (O_2975,N_29977,N_29989);
nand UO_2976 (O_2976,N_29863,N_29927);
nor UO_2977 (O_2977,N_29911,N_29853);
or UO_2978 (O_2978,N_29854,N_29898);
or UO_2979 (O_2979,N_29951,N_29965);
nand UO_2980 (O_2980,N_29875,N_29876);
nor UO_2981 (O_2981,N_29900,N_29935);
or UO_2982 (O_2982,N_29934,N_29844);
and UO_2983 (O_2983,N_29889,N_29885);
and UO_2984 (O_2984,N_29993,N_29985);
and UO_2985 (O_2985,N_29993,N_29959);
xor UO_2986 (O_2986,N_29942,N_29877);
and UO_2987 (O_2987,N_29822,N_29910);
nor UO_2988 (O_2988,N_29808,N_29827);
nand UO_2989 (O_2989,N_29917,N_29984);
nand UO_2990 (O_2990,N_29888,N_29897);
nor UO_2991 (O_2991,N_29956,N_29942);
xor UO_2992 (O_2992,N_29912,N_29905);
nor UO_2993 (O_2993,N_29908,N_29919);
or UO_2994 (O_2994,N_29840,N_29959);
nor UO_2995 (O_2995,N_29846,N_29811);
or UO_2996 (O_2996,N_29903,N_29858);
and UO_2997 (O_2997,N_29948,N_29882);
or UO_2998 (O_2998,N_29909,N_29907);
nor UO_2999 (O_2999,N_29889,N_29964);
nor UO_3000 (O_3000,N_29871,N_29970);
nand UO_3001 (O_3001,N_29981,N_29947);
nor UO_3002 (O_3002,N_29944,N_29839);
xnor UO_3003 (O_3003,N_29972,N_29823);
or UO_3004 (O_3004,N_29982,N_29990);
or UO_3005 (O_3005,N_29878,N_29883);
nor UO_3006 (O_3006,N_29802,N_29839);
xor UO_3007 (O_3007,N_29836,N_29944);
nand UO_3008 (O_3008,N_29858,N_29884);
or UO_3009 (O_3009,N_29968,N_29966);
xnor UO_3010 (O_3010,N_29980,N_29869);
and UO_3011 (O_3011,N_29954,N_29879);
xor UO_3012 (O_3012,N_29870,N_29838);
nor UO_3013 (O_3013,N_29998,N_29898);
xor UO_3014 (O_3014,N_29842,N_29997);
or UO_3015 (O_3015,N_29948,N_29820);
and UO_3016 (O_3016,N_29860,N_29849);
nand UO_3017 (O_3017,N_29873,N_29883);
nand UO_3018 (O_3018,N_29886,N_29906);
and UO_3019 (O_3019,N_29830,N_29911);
nor UO_3020 (O_3020,N_29868,N_29938);
or UO_3021 (O_3021,N_29981,N_29918);
nor UO_3022 (O_3022,N_29963,N_29977);
nor UO_3023 (O_3023,N_29847,N_29808);
or UO_3024 (O_3024,N_29969,N_29837);
and UO_3025 (O_3025,N_29953,N_29920);
nor UO_3026 (O_3026,N_29947,N_29849);
nand UO_3027 (O_3027,N_29904,N_29850);
nand UO_3028 (O_3028,N_29926,N_29850);
xnor UO_3029 (O_3029,N_29927,N_29902);
nand UO_3030 (O_3030,N_29868,N_29823);
xor UO_3031 (O_3031,N_29933,N_29873);
and UO_3032 (O_3032,N_29906,N_29981);
xnor UO_3033 (O_3033,N_29954,N_29923);
and UO_3034 (O_3034,N_29992,N_29947);
and UO_3035 (O_3035,N_29848,N_29981);
xnor UO_3036 (O_3036,N_29896,N_29913);
xor UO_3037 (O_3037,N_29964,N_29820);
or UO_3038 (O_3038,N_29983,N_29828);
or UO_3039 (O_3039,N_29874,N_29912);
or UO_3040 (O_3040,N_29883,N_29814);
xor UO_3041 (O_3041,N_29805,N_29807);
or UO_3042 (O_3042,N_29817,N_29803);
and UO_3043 (O_3043,N_29904,N_29987);
and UO_3044 (O_3044,N_29975,N_29879);
nand UO_3045 (O_3045,N_29807,N_29951);
and UO_3046 (O_3046,N_29946,N_29819);
nand UO_3047 (O_3047,N_29825,N_29928);
nor UO_3048 (O_3048,N_29823,N_29963);
nand UO_3049 (O_3049,N_29921,N_29903);
xor UO_3050 (O_3050,N_29805,N_29842);
nor UO_3051 (O_3051,N_29832,N_29855);
xor UO_3052 (O_3052,N_29875,N_29807);
nand UO_3053 (O_3053,N_29914,N_29888);
and UO_3054 (O_3054,N_29802,N_29999);
nand UO_3055 (O_3055,N_29813,N_29902);
nand UO_3056 (O_3056,N_29942,N_29998);
xnor UO_3057 (O_3057,N_29831,N_29875);
nand UO_3058 (O_3058,N_29827,N_29987);
nand UO_3059 (O_3059,N_29951,N_29869);
nand UO_3060 (O_3060,N_29860,N_29821);
or UO_3061 (O_3061,N_29977,N_29934);
or UO_3062 (O_3062,N_29904,N_29973);
xnor UO_3063 (O_3063,N_29880,N_29970);
or UO_3064 (O_3064,N_29897,N_29961);
and UO_3065 (O_3065,N_29949,N_29884);
and UO_3066 (O_3066,N_29829,N_29984);
nand UO_3067 (O_3067,N_29816,N_29995);
or UO_3068 (O_3068,N_29989,N_29995);
or UO_3069 (O_3069,N_29988,N_29801);
and UO_3070 (O_3070,N_29970,N_29809);
or UO_3071 (O_3071,N_29940,N_29851);
nand UO_3072 (O_3072,N_29936,N_29812);
xor UO_3073 (O_3073,N_29988,N_29995);
xnor UO_3074 (O_3074,N_29939,N_29854);
nand UO_3075 (O_3075,N_29830,N_29954);
and UO_3076 (O_3076,N_29901,N_29827);
nor UO_3077 (O_3077,N_29974,N_29864);
nor UO_3078 (O_3078,N_29830,N_29838);
nand UO_3079 (O_3079,N_29887,N_29921);
nor UO_3080 (O_3080,N_29933,N_29858);
or UO_3081 (O_3081,N_29972,N_29886);
xor UO_3082 (O_3082,N_29858,N_29978);
or UO_3083 (O_3083,N_29913,N_29958);
and UO_3084 (O_3084,N_29848,N_29877);
and UO_3085 (O_3085,N_29988,N_29919);
nand UO_3086 (O_3086,N_29836,N_29977);
nor UO_3087 (O_3087,N_29848,N_29978);
or UO_3088 (O_3088,N_29986,N_29989);
nand UO_3089 (O_3089,N_29862,N_29806);
nand UO_3090 (O_3090,N_29900,N_29864);
or UO_3091 (O_3091,N_29904,N_29936);
and UO_3092 (O_3092,N_29865,N_29843);
nor UO_3093 (O_3093,N_29956,N_29841);
xor UO_3094 (O_3094,N_29874,N_29906);
or UO_3095 (O_3095,N_29994,N_29880);
or UO_3096 (O_3096,N_29892,N_29836);
or UO_3097 (O_3097,N_29956,N_29931);
nand UO_3098 (O_3098,N_29913,N_29818);
nand UO_3099 (O_3099,N_29998,N_29811);
and UO_3100 (O_3100,N_29940,N_29884);
nand UO_3101 (O_3101,N_29936,N_29816);
nand UO_3102 (O_3102,N_29959,N_29971);
and UO_3103 (O_3103,N_29912,N_29842);
and UO_3104 (O_3104,N_29948,N_29891);
or UO_3105 (O_3105,N_29977,N_29932);
or UO_3106 (O_3106,N_29930,N_29815);
or UO_3107 (O_3107,N_29834,N_29976);
xor UO_3108 (O_3108,N_29912,N_29800);
xnor UO_3109 (O_3109,N_29822,N_29826);
or UO_3110 (O_3110,N_29809,N_29931);
nor UO_3111 (O_3111,N_29884,N_29956);
and UO_3112 (O_3112,N_29932,N_29877);
or UO_3113 (O_3113,N_29964,N_29925);
xnor UO_3114 (O_3114,N_29834,N_29960);
nand UO_3115 (O_3115,N_29889,N_29887);
or UO_3116 (O_3116,N_29892,N_29869);
xnor UO_3117 (O_3117,N_29802,N_29809);
or UO_3118 (O_3118,N_29996,N_29838);
and UO_3119 (O_3119,N_29984,N_29940);
and UO_3120 (O_3120,N_29953,N_29987);
nand UO_3121 (O_3121,N_29973,N_29901);
or UO_3122 (O_3122,N_29972,N_29885);
nand UO_3123 (O_3123,N_29958,N_29896);
or UO_3124 (O_3124,N_29829,N_29961);
and UO_3125 (O_3125,N_29825,N_29945);
xor UO_3126 (O_3126,N_29894,N_29997);
or UO_3127 (O_3127,N_29907,N_29896);
nor UO_3128 (O_3128,N_29936,N_29866);
or UO_3129 (O_3129,N_29884,N_29865);
nand UO_3130 (O_3130,N_29859,N_29877);
or UO_3131 (O_3131,N_29861,N_29934);
and UO_3132 (O_3132,N_29938,N_29823);
and UO_3133 (O_3133,N_29931,N_29968);
or UO_3134 (O_3134,N_29973,N_29945);
xor UO_3135 (O_3135,N_29836,N_29841);
nand UO_3136 (O_3136,N_29811,N_29917);
xor UO_3137 (O_3137,N_29904,N_29816);
nand UO_3138 (O_3138,N_29958,N_29955);
nor UO_3139 (O_3139,N_29981,N_29861);
nand UO_3140 (O_3140,N_29814,N_29933);
nand UO_3141 (O_3141,N_29933,N_29909);
nor UO_3142 (O_3142,N_29965,N_29947);
nand UO_3143 (O_3143,N_29910,N_29829);
or UO_3144 (O_3144,N_29946,N_29825);
or UO_3145 (O_3145,N_29804,N_29930);
nor UO_3146 (O_3146,N_29978,N_29850);
nor UO_3147 (O_3147,N_29940,N_29886);
and UO_3148 (O_3148,N_29860,N_29900);
nor UO_3149 (O_3149,N_29807,N_29897);
or UO_3150 (O_3150,N_29915,N_29958);
nand UO_3151 (O_3151,N_29803,N_29845);
xor UO_3152 (O_3152,N_29967,N_29876);
xnor UO_3153 (O_3153,N_29993,N_29971);
xor UO_3154 (O_3154,N_29828,N_29934);
nor UO_3155 (O_3155,N_29806,N_29833);
nor UO_3156 (O_3156,N_29948,N_29976);
nor UO_3157 (O_3157,N_29959,N_29905);
or UO_3158 (O_3158,N_29896,N_29865);
or UO_3159 (O_3159,N_29893,N_29873);
or UO_3160 (O_3160,N_29982,N_29803);
xor UO_3161 (O_3161,N_29916,N_29828);
xnor UO_3162 (O_3162,N_29929,N_29969);
nand UO_3163 (O_3163,N_29971,N_29884);
nor UO_3164 (O_3164,N_29866,N_29955);
or UO_3165 (O_3165,N_29902,N_29958);
nand UO_3166 (O_3166,N_29858,N_29977);
nand UO_3167 (O_3167,N_29904,N_29804);
nand UO_3168 (O_3168,N_29881,N_29931);
or UO_3169 (O_3169,N_29894,N_29888);
or UO_3170 (O_3170,N_29989,N_29886);
nor UO_3171 (O_3171,N_29876,N_29883);
or UO_3172 (O_3172,N_29878,N_29900);
nor UO_3173 (O_3173,N_29903,N_29827);
and UO_3174 (O_3174,N_29929,N_29861);
or UO_3175 (O_3175,N_29815,N_29802);
xnor UO_3176 (O_3176,N_29985,N_29813);
nand UO_3177 (O_3177,N_29838,N_29985);
and UO_3178 (O_3178,N_29963,N_29809);
nor UO_3179 (O_3179,N_29935,N_29804);
xor UO_3180 (O_3180,N_29871,N_29892);
nor UO_3181 (O_3181,N_29985,N_29800);
xor UO_3182 (O_3182,N_29839,N_29881);
or UO_3183 (O_3183,N_29954,N_29887);
nor UO_3184 (O_3184,N_29865,N_29921);
nor UO_3185 (O_3185,N_29970,N_29831);
nor UO_3186 (O_3186,N_29918,N_29913);
nand UO_3187 (O_3187,N_29934,N_29866);
or UO_3188 (O_3188,N_29906,N_29972);
or UO_3189 (O_3189,N_29902,N_29920);
and UO_3190 (O_3190,N_29866,N_29843);
nand UO_3191 (O_3191,N_29912,N_29867);
nor UO_3192 (O_3192,N_29854,N_29943);
nand UO_3193 (O_3193,N_29837,N_29899);
or UO_3194 (O_3194,N_29933,N_29833);
xor UO_3195 (O_3195,N_29973,N_29936);
and UO_3196 (O_3196,N_29925,N_29977);
and UO_3197 (O_3197,N_29857,N_29983);
xor UO_3198 (O_3198,N_29955,N_29902);
nand UO_3199 (O_3199,N_29931,N_29815);
nand UO_3200 (O_3200,N_29863,N_29869);
and UO_3201 (O_3201,N_29873,N_29969);
nor UO_3202 (O_3202,N_29872,N_29906);
nand UO_3203 (O_3203,N_29941,N_29818);
nor UO_3204 (O_3204,N_29944,N_29995);
nor UO_3205 (O_3205,N_29955,N_29971);
xor UO_3206 (O_3206,N_29869,N_29898);
or UO_3207 (O_3207,N_29940,N_29855);
or UO_3208 (O_3208,N_29969,N_29842);
and UO_3209 (O_3209,N_29801,N_29897);
nand UO_3210 (O_3210,N_29844,N_29866);
or UO_3211 (O_3211,N_29847,N_29850);
and UO_3212 (O_3212,N_29868,N_29800);
and UO_3213 (O_3213,N_29848,N_29965);
xnor UO_3214 (O_3214,N_29889,N_29813);
xor UO_3215 (O_3215,N_29993,N_29814);
nand UO_3216 (O_3216,N_29883,N_29836);
nand UO_3217 (O_3217,N_29963,N_29933);
nor UO_3218 (O_3218,N_29883,N_29911);
xor UO_3219 (O_3219,N_29874,N_29826);
and UO_3220 (O_3220,N_29814,N_29896);
nor UO_3221 (O_3221,N_29836,N_29979);
nand UO_3222 (O_3222,N_29944,N_29910);
xnor UO_3223 (O_3223,N_29900,N_29936);
and UO_3224 (O_3224,N_29834,N_29881);
xnor UO_3225 (O_3225,N_29820,N_29897);
nand UO_3226 (O_3226,N_29937,N_29854);
xnor UO_3227 (O_3227,N_29959,N_29886);
and UO_3228 (O_3228,N_29861,N_29913);
nand UO_3229 (O_3229,N_29931,N_29912);
and UO_3230 (O_3230,N_29823,N_29864);
xor UO_3231 (O_3231,N_29841,N_29859);
nor UO_3232 (O_3232,N_29880,N_29901);
nand UO_3233 (O_3233,N_29984,N_29871);
or UO_3234 (O_3234,N_29866,N_29800);
and UO_3235 (O_3235,N_29984,N_29980);
xor UO_3236 (O_3236,N_29890,N_29978);
nand UO_3237 (O_3237,N_29975,N_29953);
nor UO_3238 (O_3238,N_29967,N_29833);
nand UO_3239 (O_3239,N_29865,N_29997);
xnor UO_3240 (O_3240,N_29859,N_29809);
or UO_3241 (O_3241,N_29926,N_29800);
or UO_3242 (O_3242,N_29967,N_29891);
xnor UO_3243 (O_3243,N_29821,N_29938);
or UO_3244 (O_3244,N_29920,N_29932);
nand UO_3245 (O_3245,N_29908,N_29856);
nand UO_3246 (O_3246,N_29935,N_29961);
nor UO_3247 (O_3247,N_29814,N_29909);
or UO_3248 (O_3248,N_29954,N_29918);
xnor UO_3249 (O_3249,N_29858,N_29814);
and UO_3250 (O_3250,N_29871,N_29889);
nor UO_3251 (O_3251,N_29949,N_29843);
nand UO_3252 (O_3252,N_29927,N_29851);
nand UO_3253 (O_3253,N_29910,N_29857);
nand UO_3254 (O_3254,N_29966,N_29845);
or UO_3255 (O_3255,N_29985,N_29939);
or UO_3256 (O_3256,N_29975,N_29834);
xor UO_3257 (O_3257,N_29923,N_29880);
nand UO_3258 (O_3258,N_29863,N_29946);
xnor UO_3259 (O_3259,N_29922,N_29816);
nand UO_3260 (O_3260,N_29856,N_29915);
nand UO_3261 (O_3261,N_29827,N_29853);
nor UO_3262 (O_3262,N_29910,N_29990);
or UO_3263 (O_3263,N_29839,N_29899);
nor UO_3264 (O_3264,N_29884,N_29877);
and UO_3265 (O_3265,N_29824,N_29872);
nand UO_3266 (O_3266,N_29836,N_29935);
and UO_3267 (O_3267,N_29889,N_29890);
or UO_3268 (O_3268,N_29859,N_29928);
nor UO_3269 (O_3269,N_29963,N_29986);
xnor UO_3270 (O_3270,N_29899,N_29815);
nor UO_3271 (O_3271,N_29951,N_29830);
nor UO_3272 (O_3272,N_29862,N_29969);
nor UO_3273 (O_3273,N_29860,N_29963);
or UO_3274 (O_3274,N_29864,N_29821);
xnor UO_3275 (O_3275,N_29999,N_29801);
xor UO_3276 (O_3276,N_29859,N_29995);
xnor UO_3277 (O_3277,N_29813,N_29913);
and UO_3278 (O_3278,N_29863,N_29802);
and UO_3279 (O_3279,N_29917,N_29916);
nor UO_3280 (O_3280,N_29850,N_29962);
nand UO_3281 (O_3281,N_29943,N_29870);
nor UO_3282 (O_3282,N_29805,N_29989);
nand UO_3283 (O_3283,N_29845,N_29848);
and UO_3284 (O_3284,N_29822,N_29993);
nand UO_3285 (O_3285,N_29863,N_29805);
nand UO_3286 (O_3286,N_29903,N_29870);
and UO_3287 (O_3287,N_29811,N_29834);
nor UO_3288 (O_3288,N_29969,N_29988);
or UO_3289 (O_3289,N_29987,N_29805);
nor UO_3290 (O_3290,N_29924,N_29897);
nor UO_3291 (O_3291,N_29997,N_29994);
and UO_3292 (O_3292,N_29801,N_29844);
xor UO_3293 (O_3293,N_29876,N_29833);
nand UO_3294 (O_3294,N_29800,N_29903);
nand UO_3295 (O_3295,N_29929,N_29908);
and UO_3296 (O_3296,N_29880,N_29967);
nand UO_3297 (O_3297,N_29894,N_29831);
or UO_3298 (O_3298,N_29879,N_29916);
nand UO_3299 (O_3299,N_29900,N_29968);
nand UO_3300 (O_3300,N_29971,N_29974);
nor UO_3301 (O_3301,N_29918,N_29856);
nand UO_3302 (O_3302,N_29903,N_29883);
xor UO_3303 (O_3303,N_29886,N_29839);
or UO_3304 (O_3304,N_29972,N_29978);
xnor UO_3305 (O_3305,N_29976,N_29832);
or UO_3306 (O_3306,N_29846,N_29981);
xnor UO_3307 (O_3307,N_29878,N_29877);
or UO_3308 (O_3308,N_29921,N_29855);
xor UO_3309 (O_3309,N_29906,N_29869);
and UO_3310 (O_3310,N_29854,N_29875);
and UO_3311 (O_3311,N_29806,N_29966);
nor UO_3312 (O_3312,N_29918,N_29953);
xor UO_3313 (O_3313,N_29826,N_29847);
nor UO_3314 (O_3314,N_29945,N_29801);
and UO_3315 (O_3315,N_29898,N_29805);
and UO_3316 (O_3316,N_29958,N_29898);
xor UO_3317 (O_3317,N_29999,N_29882);
nand UO_3318 (O_3318,N_29847,N_29836);
nand UO_3319 (O_3319,N_29980,N_29854);
and UO_3320 (O_3320,N_29845,N_29873);
nand UO_3321 (O_3321,N_29885,N_29957);
xor UO_3322 (O_3322,N_29836,N_29942);
and UO_3323 (O_3323,N_29924,N_29809);
xor UO_3324 (O_3324,N_29943,N_29970);
and UO_3325 (O_3325,N_29981,N_29921);
xor UO_3326 (O_3326,N_29919,N_29888);
and UO_3327 (O_3327,N_29926,N_29857);
or UO_3328 (O_3328,N_29989,N_29833);
xor UO_3329 (O_3329,N_29947,N_29987);
nor UO_3330 (O_3330,N_29905,N_29916);
nand UO_3331 (O_3331,N_29960,N_29927);
and UO_3332 (O_3332,N_29854,N_29978);
nor UO_3333 (O_3333,N_29923,N_29889);
or UO_3334 (O_3334,N_29921,N_29972);
nand UO_3335 (O_3335,N_29816,N_29927);
or UO_3336 (O_3336,N_29874,N_29816);
xor UO_3337 (O_3337,N_29917,N_29953);
nand UO_3338 (O_3338,N_29834,N_29833);
or UO_3339 (O_3339,N_29991,N_29803);
and UO_3340 (O_3340,N_29998,N_29883);
xnor UO_3341 (O_3341,N_29973,N_29880);
or UO_3342 (O_3342,N_29825,N_29854);
nand UO_3343 (O_3343,N_29918,N_29903);
and UO_3344 (O_3344,N_29873,N_29821);
or UO_3345 (O_3345,N_29938,N_29916);
nand UO_3346 (O_3346,N_29972,N_29825);
xnor UO_3347 (O_3347,N_29909,N_29942);
xnor UO_3348 (O_3348,N_29949,N_29852);
xnor UO_3349 (O_3349,N_29856,N_29823);
nor UO_3350 (O_3350,N_29901,N_29820);
xor UO_3351 (O_3351,N_29957,N_29846);
or UO_3352 (O_3352,N_29904,N_29874);
nor UO_3353 (O_3353,N_29899,N_29990);
nand UO_3354 (O_3354,N_29828,N_29872);
nand UO_3355 (O_3355,N_29829,N_29908);
xor UO_3356 (O_3356,N_29836,N_29986);
nand UO_3357 (O_3357,N_29927,N_29840);
and UO_3358 (O_3358,N_29808,N_29857);
xor UO_3359 (O_3359,N_29989,N_29917);
and UO_3360 (O_3360,N_29977,N_29890);
and UO_3361 (O_3361,N_29939,N_29877);
nor UO_3362 (O_3362,N_29825,N_29967);
nand UO_3363 (O_3363,N_29836,N_29859);
nand UO_3364 (O_3364,N_29818,N_29863);
nor UO_3365 (O_3365,N_29994,N_29960);
nor UO_3366 (O_3366,N_29868,N_29979);
nor UO_3367 (O_3367,N_29863,N_29944);
nand UO_3368 (O_3368,N_29833,N_29867);
and UO_3369 (O_3369,N_29982,N_29865);
xnor UO_3370 (O_3370,N_29968,N_29909);
xor UO_3371 (O_3371,N_29978,N_29903);
xor UO_3372 (O_3372,N_29901,N_29972);
nand UO_3373 (O_3373,N_29877,N_29830);
nor UO_3374 (O_3374,N_29935,N_29899);
and UO_3375 (O_3375,N_29922,N_29960);
nand UO_3376 (O_3376,N_29985,N_29802);
or UO_3377 (O_3377,N_29907,N_29892);
nor UO_3378 (O_3378,N_29993,N_29928);
nor UO_3379 (O_3379,N_29838,N_29884);
nand UO_3380 (O_3380,N_29832,N_29950);
nand UO_3381 (O_3381,N_29826,N_29862);
nand UO_3382 (O_3382,N_29994,N_29834);
xor UO_3383 (O_3383,N_29941,N_29914);
nand UO_3384 (O_3384,N_29891,N_29802);
nand UO_3385 (O_3385,N_29913,N_29961);
xnor UO_3386 (O_3386,N_29993,N_29958);
xor UO_3387 (O_3387,N_29982,N_29821);
nand UO_3388 (O_3388,N_29933,N_29868);
or UO_3389 (O_3389,N_29807,N_29842);
or UO_3390 (O_3390,N_29806,N_29981);
xor UO_3391 (O_3391,N_29923,N_29936);
nand UO_3392 (O_3392,N_29957,N_29909);
nand UO_3393 (O_3393,N_29858,N_29981);
or UO_3394 (O_3394,N_29823,N_29937);
xor UO_3395 (O_3395,N_29924,N_29806);
xnor UO_3396 (O_3396,N_29985,N_29965);
nand UO_3397 (O_3397,N_29981,N_29804);
nor UO_3398 (O_3398,N_29823,N_29949);
nor UO_3399 (O_3399,N_29811,N_29947);
or UO_3400 (O_3400,N_29876,N_29924);
xnor UO_3401 (O_3401,N_29802,N_29959);
xnor UO_3402 (O_3402,N_29988,N_29882);
nand UO_3403 (O_3403,N_29919,N_29817);
or UO_3404 (O_3404,N_29867,N_29889);
xnor UO_3405 (O_3405,N_29889,N_29893);
nand UO_3406 (O_3406,N_29900,N_29981);
nand UO_3407 (O_3407,N_29802,N_29960);
nand UO_3408 (O_3408,N_29803,N_29989);
and UO_3409 (O_3409,N_29899,N_29958);
or UO_3410 (O_3410,N_29851,N_29813);
xor UO_3411 (O_3411,N_29982,N_29848);
nor UO_3412 (O_3412,N_29931,N_29844);
or UO_3413 (O_3413,N_29872,N_29957);
nand UO_3414 (O_3414,N_29822,N_29966);
xnor UO_3415 (O_3415,N_29824,N_29913);
nor UO_3416 (O_3416,N_29947,N_29894);
nor UO_3417 (O_3417,N_29871,N_29832);
nor UO_3418 (O_3418,N_29957,N_29913);
nand UO_3419 (O_3419,N_29809,N_29985);
nand UO_3420 (O_3420,N_29950,N_29963);
nand UO_3421 (O_3421,N_29893,N_29870);
nor UO_3422 (O_3422,N_29915,N_29996);
xor UO_3423 (O_3423,N_29907,N_29941);
xor UO_3424 (O_3424,N_29834,N_29933);
nor UO_3425 (O_3425,N_29980,N_29835);
and UO_3426 (O_3426,N_29918,N_29993);
and UO_3427 (O_3427,N_29851,N_29952);
nor UO_3428 (O_3428,N_29963,N_29818);
nand UO_3429 (O_3429,N_29888,N_29822);
nor UO_3430 (O_3430,N_29883,N_29846);
xnor UO_3431 (O_3431,N_29817,N_29904);
nor UO_3432 (O_3432,N_29878,N_29848);
xor UO_3433 (O_3433,N_29895,N_29905);
and UO_3434 (O_3434,N_29979,N_29990);
nor UO_3435 (O_3435,N_29892,N_29929);
and UO_3436 (O_3436,N_29855,N_29898);
nor UO_3437 (O_3437,N_29910,N_29954);
nand UO_3438 (O_3438,N_29941,N_29808);
nor UO_3439 (O_3439,N_29999,N_29987);
or UO_3440 (O_3440,N_29969,N_29933);
nor UO_3441 (O_3441,N_29935,N_29971);
xnor UO_3442 (O_3442,N_29834,N_29814);
nand UO_3443 (O_3443,N_29871,N_29922);
and UO_3444 (O_3444,N_29968,N_29897);
and UO_3445 (O_3445,N_29911,N_29910);
and UO_3446 (O_3446,N_29868,N_29857);
nand UO_3447 (O_3447,N_29855,N_29897);
or UO_3448 (O_3448,N_29883,N_29907);
xnor UO_3449 (O_3449,N_29827,N_29819);
or UO_3450 (O_3450,N_29963,N_29910);
or UO_3451 (O_3451,N_29969,N_29981);
nor UO_3452 (O_3452,N_29933,N_29996);
and UO_3453 (O_3453,N_29833,N_29962);
or UO_3454 (O_3454,N_29981,N_29924);
or UO_3455 (O_3455,N_29911,N_29907);
nor UO_3456 (O_3456,N_29989,N_29851);
xnor UO_3457 (O_3457,N_29953,N_29891);
xnor UO_3458 (O_3458,N_29800,N_29872);
nand UO_3459 (O_3459,N_29991,N_29849);
xor UO_3460 (O_3460,N_29895,N_29923);
nand UO_3461 (O_3461,N_29810,N_29833);
nor UO_3462 (O_3462,N_29835,N_29838);
xnor UO_3463 (O_3463,N_29981,N_29930);
nor UO_3464 (O_3464,N_29849,N_29840);
nand UO_3465 (O_3465,N_29995,N_29846);
or UO_3466 (O_3466,N_29989,N_29887);
and UO_3467 (O_3467,N_29902,N_29965);
nand UO_3468 (O_3468,N_29908,N_29960);
and UO_3469 (O_3469,N_29889,N_29865);
nand UO_3470 (O_3470,N_29808,N_29900);
or UO_3471 (O_3471,N_29970,N_29863);
or UO_3472 (O_3472,N_29877,N_29808);
nand UO_3473 (O_3473,N_29846,N_29844);
and UO_3474 (O_3474,N_29911,N_29823);
nand UO_3475 (O_3475,N_29868,N_29880);
and UO_3476 (O_3476,N_29923,N_29904);
and UO_3477 (O_3477,N_29996,N_29840);
nor UO_3478 (O_3478,N_29834,N_29959);
or UO_3479 (O_3479,N_29947,N_29932);
nor UO_3480 (O_3480,N_29853,N_29872);
nand UO_3481 (O_3481,N_29834,N_29847);
xnor UO_3482 (O_3482,N_29849,N_29861);
nand UO_3483 (O_3483,N_29884,N_29905);
or UO_3484 (O_3484,N_29863,N_29888);
or UO_3485 (O_3485,N_29844,N_29865);
xor UO_3486 (O_3486,N_29888,N_29946);
and UO_3487 (O_3487,N_29923,N_29829);
or UO_3488 (O_3488,N_29804,N_29810);
and UO_3489 (O_3489,N_29947,N_29923);
or UO_3490 (O_3490,N_29917,N_29853);
or UO_3491 (O_3491,N_29976,N_29883);
and UO_3492 (O_3492,N_29810,N_29898);
xor UO_3493 (O_3493,N_29915,N_29942);
nand UO_3494 (O_3494,N_29823,N_29924);
xor UO_3495 (O_3495,N_29826,N_29947);
nor UO_3496 (O_3496,N_29888,N_29982);
xor UO_3497 (O_3497,N_29841,N_29906);
xor UO_3498 (O_3498,N_29913,N_29962);
or UO_3499 (O_3499,N_29834,N_29909);
endmodule