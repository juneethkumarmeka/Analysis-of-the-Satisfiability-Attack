module basic_500_3000_500_30_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_140,In_332);
and U1 (N_1,In_478,In_107);
or U2 (N_2,In_263,In_292);
nand U3 (N_3,In_458,In_313);
or U4 (N_4,In_368,In_380);
nor U5 (N_5,In_8,In_320);
nand U6 (N_6,In_479,In_35);
or U7 (N_7,In_208,In_199);
or U8 (N_8,In_346,In_497);
nor U9 (N_9,In_23,In_220);
nor U10 (N_10,In_94,In_11);
nand U11 (N_11,In_46,In_463);
nor U12 (N_12,In_282,In_172);
and U13 (N_13,In_64,In_311);
nand U14 (N_14,In_137,In_59);
or U15 (N_15,In_367,In_249);
nand U16 (N_16,In_81,In_278);
nor U17 (N_17,In_6,In_37);
nor U18 (N_18,In_285,In_103);
nor U19 (N_19,In_41,In_129);
or U20 (N_20,In_425,In_102);
nor U21 (N_21,In_235,In_109);
nand U22 (N_22,In_483,In_353);
or U23 (N_23,In_262,In_275);
xor U24 (N_24,In_99,In_69);
nor U25 (N_25,In_335,In_469);
and U26 (N_26,In_490,In_417);
nor U27 (N_27,In_439,In_218);
nand U28 (N_28,In_92,In_374);
xor U29 (N_29,In_122,In_85);
nor U30 (N_30,In_135,In_47);
nand U31 (N_31,In_229,In_195);
nor U32 (N_32,In_33,In_485);
and U33 (N_33,In_391,In_461);
nor U34 (N_34,In_462,In_434);
nor U35 (N_35,In_392,In_342);
nor U36 (N_36,In_178,In_395);
and U37 (N_37,In_325,In_440);
nor U38 (N_38,In_212,In_101);
nand U39 (N_39,In_71,In_409);
or U40 (N_40,In_192,In_202);
or U41 (N_41,In_309,In_340);
nand U42 (N_42,In_54,In_454);
and U43 (N_43,In_182,In_166);
nor U44 (N_44,In_242,In_393);
nand U45 (N_45,In_245,In_493);
or U46 (N_46,In_260,In_169);
nand U47 (N_47,In_441,In_130);
or U48 (N_48,In_350,In_310);
nand U49 (N_49,In_227,In_293);
and U50 (N_50,In_494,In_489);
and U51 (N_51,In_222,In_327);
or U52 (N_52,In_447,In_82);
nor U53 (N_53,In_34,In_431);
nand U54 (N_54,In_279,In_297);
or U55 (N_55,In_211,In_30);
nand U56 (N_56,In_151,In_432);
nor U57 (N_57,In_487,In_200);
and U58 (N_58,In_345,In_167);
nand U59 (N_59,In_158,In_17);
or U60 (N_60,In_44,In_153);
nand U61 (N_61,In_290,In_257);
or U62 (N_62,In_443,In_196);
and U63 (N_63,In_18,In_55);
and U64 (N_64,In_224,In_465);
nand U65 (N_65,In_435,In_445);
and U66 (N_66,In_201,In_24);
nor U67 (N_67,In_187,In_88);
nor U68 (N_68,In_266,In_217);
nand U69 (N_69,In_337,In_136);
or U70 (N_70,In_170,In_0);
nand U71 (N_71,In_185,In_306);
nand U72 (N_72,In_365,In_300);
and U73 (N_73,In_456,In_22);
and U74 (N_74,In_453,In_119);
nand U75 (N_75,In_142,In_147);
nor U76 (N_76,In_265,In_499);
or U77 (N_77,In_414,In_186);
nand U78 (N_78,In_398,In_57);
and U79 (N_79,In_173,In_160);
nand U80 (N_80,In_312,In_68);
and U81 (N_81,In_205,In_464);
and U82 (N_82,In_386,In_48);
or U83 (N_83,In_385,In_498);
nor U84 (N_84,In_394,In_91);
nand U85 (N_85,In_132,In_214);
nand U86 (N_86,In_271,In_28);
nand U87 (N_87,In_438,In_225);
or U88 (N_88,In_351,In_344);
and U89 (N_89,In_451,In_246);
nand U90 (N_90,In_210,In_481);
nand U91 (N_91,In_449,In_238);
nor U92 (N_92,In_427,In_404);
and U93 (N_93,In_470,In_475);
and U94 (N_94,In_194,In_437);
nor U95 (N_95,In_360,In_89);
nand U96 (N_96,In_250,In_97);
and U97 (N_97,In_412,In_423);
or U98 (N_98,In_161,In_406);
nand U99 (N_99,In_100,In_255);
nand U100 (N_100,In_189,N_91);
nand U101 (N_101,In_356,In_112);
or U102 (N_102,In_256,In_492);
or U103 (N_103,In_314,In_274);
or U104 (N_104,In_86,In_125);
and U105 (N_105,N_11,In_284);
and U106 (N_106,In_116,N_64);
and U107 (N_107,In_93,In_16);
or U108 (N_108,N_63,In_73);
nor U109 (N_109,N_99,In_232);
nand U110 (N_110,In_39,N_96);
nand U111 (N_111,In_436,In_316);
nand U112 (N_112,In_450,N_17);
or U113 (N_113,In_323,In_303);
and U114 (N_114,In_387,N_42);
nor U115 (N_115,In_341,In_78);
and U116 (N_116,In_399,In_5);
nand U117 (N_117,In_400,N_13);
nor U118 (N_118,In_190,In_388);
and U119 (N_119,N_30,N_25);
nand U120 (N_120,In_175,In_236);
xor U121 (N_121,N_72,N_83);
nand U122 (N_122,In_496,N_69);
and U123 (N_123,In_408,In_14);
nand U124 (N_124,In_104,In_413);
and U125 (N_125,In_396,In_482);
nor U126 (N_126,In_298,In_113);
or U127 (N_127,N_53,In_110);
or U128 (N_128,In_241,In_133);
nand U129 (N_129,N_45,In_294);
or U130 (N_130,In_369,In_375);
or U131 (N_131,In_355,In_53);
or U132 (N_132,In_76,In_203);
xnor U133 (N_133,In_253,N_59);
nand U134 (N_134,In_74,N_61);
nor U135 (N_135,In_430,In_145);
or U136 (N_136,N_81,In_467);
or U137 (N_137,In_468,N_1);
or U138 (N_138,In_302,N_35);
nor U139 (N_139,N_37,N_41);
and U140 (N_140,In_19,In_331);
and U141 (N_141,In_382,In_111);
or U142 (N_142,In_179,In_228);
and U143 (N_143,In_273,In_429);
nor U144 (N_144,N_4,N_79);
nand U145 (N_145,In_183,N_0);
nor U146 (N_146,N_48,N_15);
nand U147 (N_147,In_138,In_426);
and U148 (N_148,N_56,In_381);
nand U149 (N_149,In_181,In_163);
or U150 (N_150,N_29,In_491);
xor U151 (N_151,In_370,In_70);
or U152 (N_152,In_308,N_80);
nand U153 (N_153,In_75,In_304);
or U154 (N_154,In_1,In_150);
and U155 (N_155,N_49,In_379);
or U156 (N_156,In_231,In_154);
or U157 (N_157,In_25,N_24);
nand U158 (N_158,In_123,In_319);
nor U159 (N_159,In_358,N_65);
or U160 (N_160,In_288,N_19);
and U161 (N_161,N_84,N_32);
nand U162 (N_162,In_26,In_79);
or U163 (N_163,N_57,In_277);
nand U164 (N_164,In_424,In_317);
nand U165 (N_165,In_329,N_36);
or U166 (N_166,In_108,N_62);
nand U167 (N_167,In_281,In_84);
and U168 (N_168,In_403,In_330);
nand U169 (N_169,In_315,In_239);
xnor U170 (N_170,In_280,In_289);
nand U171 (N_171,In_244,N_74);
and U172 (N_172,In_66,In_171);
or U173 (N_173,In_149,In_444);
or U174 (N_174,In_13,N_50);
nor U175 (N_175,In_197,In_259);
nor U176 (N_176,N_67,N_23);
xor U177 (N_177,In_60,N_7);
nand U178 (N_178,In_383,In_174);
nand U179 (N_179,N_6,In_162);
or U180 (N_180,N_87,In_177);
nor U181 (N_181,In_333,In_49);
nor U182 (N_182,In_452,In_389);
nor U183 (N_183,N_88,In_318);
or U184 (N_184,In_326,N_95);
and U185 (N_185,In_20,In_418);
nor U186 (N_186,In_126,In_143);
nand U187 (N_187,In_204,In_377);
and U188 (N_188,In_419,In_420);
or U189 (N_189,In_480,In_362);
or U190 (N_190,N_39,In_40);
and U191 (N_191,In_219,In_287);
and U192 (N_192,In_267,In_405);
nand U193 (N_193,N_85,In_95);
nor U194 (N_194,In_401,In_428);
and U195 (N_195,In_139,In_234);
and U196 (N_196,In_141,In_477);
or U197 (N_197,In_72,In_361);
nand U198 (N_198,N_66,In_233);
or U199 (N_199,N_9,In_4);
and U200 (N_200,N_5,In_474);
or U201 (N_201,N_107,N_187);
or U202 (N_202,In_105,In_473);
or U203 (N_203,In_216,In_283);
nor U204 (N_204,N_149,In_176);
nand U205 (N_205,N_140,In_61);
nor U206 (N_206,N_147,In_127);
and U207 (N_207,In_29,In_251);
nor U208 (N_208,N_183,N_169);
and U209 (N_209,In_77,N_157);
nor U210 (N_210,In_416,N_136);
and U211 (N_211,In_215,N_128);
or U212 (N_212,N_163,N_162);
and U213 (N_213,In_50,In_359);
nand U214 (N_214,In_45,N_27);
and U215 (N_215,In_305,In_397);
nand U216 (N_216,In_248,In_366);
nand U217 (N_217,In_378,In_193);
nand U218 (N_218,In_357,In_258);
nand U219 (N_219,In_364,In_188);
nor U220 (N_220,In_272,In_270);
or U221 (N_221,N_152,N_137);
nor U222 (N_222,N_191,N_174);
nand U223 (N_223,N_43,In_486);
or U224 (N_224,In_184,In_421);
or U225 (N_225,In_198,In_495);
and U226 (N_226,In_191,N_77);
nand U227 (N_227,In_371,In_12);
nand U228 (N_228,N_180,N_94);
nand U229 (N_229,N_73,N_98);
nor U230 (N_230,In_264,N_143);
nor U231 (N_231,N_44,N_106);
and U232 (N_232,In_252,N_188);
nand U233 (N_233,In_209,In_43);
nor U234 (N_234,N_76,In_124);
nor U235 (N_235,In_21,N_159);
nand U236 (N_236,N_197,In_455);
or U237 (N_237,N_103,In_7);
or U238 (N_238,N_92,In_338);
and U239 (N_239,N_170,N_51);
nor U240 (N_240,In_321,N_199);
and U241 (N_241,N_124,N_114);
or U242 (N_242,N_178,In_295);
or U243 (N_243,In_347,In_269);
and U244 (N_244,In_384,N_139);
nand U245 (N_245,N_26,N_150);
or U246 (N_246,In_422,In_106);
and U247 (N_247,N_161,In_299);
or U248 (N_248,In_373,N_172);
nor U249 (N_249,N_127,N_82);
nand U250 (N_250,N_193,N_198);
nand U251 (N_251,In_51,In_62);
nor U252 (N_252,N_108,N_105);
and U253 (N_253,In_339,In_324);
nor U254 (N_254,N_125,N_86);
nor U255 (N_255,N_184,In_410);
and U256 (N_256,N_129,In_322);
nand U257 (N_257,N_33,In_115);
nor U258 (N_258,N_158,N_22);
nor U259 (N_259,N_177,N_190);
nor U260 (N_260,N_167,N_52);
xnor U261 (N_261,In_80,In_343);
nor U262 (N_262,N_185,In_31);
nor U263 (N_263,In_276,In_448);
nor U264 (N_264,In_472,In_243);
nor U265 (N_265,In_32,N_31);
or U266 (N_266,In_96,In_180);
or U267 (N_267,In_157,N_186);
nand U268 (N_268,N_141,N_134);
or U269 (N_269,In_237,In_471);
and U270 (N_270,N_58,N_132);
and U271 (N_271,N_109,N_138);
and U272 (N_272,N_100,In_328);
nor U273 (N_273,N_34,N_90);
nand U274 (N_274,In_407,N_196);
nand U275 (N_275,In_120,N_126);
and U276 (N_276,In_307,N_121);
nand U277 (N_277,N_112,In_9);
nor U278 (N_278,N_55,In_296);
and U279 (N_279,In_148,In_261);
nor U280 (N_280,In_221,N_168);
or U281 (N_281,In_168,In_488);
nand U282 (N_282,In_376,In_146);
and U283 (N_283,In_98,In_457);
or U284 (N_284,N_21,N_113);
and U285 (N_285,In_15,In_165);
nand U286 (N_286,In_56,N_164);
or U287 (N_287,In_223,N_8);
and U288 (N_288,N_171,N_71);
and U289 (N_289,N_54,N_165);
or U290 (N_290,In_156,N_2);
or U291 (N_291,N_154,In_411);
or U292 (N_292,N_97,N_75);
nand U293 (N_293,In_402,N_194);
nand U294 (N_294,N_116,N_40);
nor U295 (N_295,In_164,N_145);
nor U296 (N_296,N_70,In_446);
and U297 (N_297,In_42,N_111);
nor U298 (N_298,N_146,N_123);
nand U299 (N_299,In_83,In_128);
and U300 (N_300,N_133,In_155);
nand U301 (N_301,N_227,N_297);
nand U302 (N_302,N_144,N_218);
xnor U303 (N_303,N_287,N_166);
nand U304 (N_304,N_160,In_476);
and U305 (N_305,N_195,N_229);
xor U306 (N_306,In_90,N_28);
and U307 (N_307,N_230,N_148);
or U308 (N_308,N_250,N_119);
and U309 (N_309,In_301,N_12);
nor U310 (N_310,In_52,N_243);
and U311 (N_311,N_38,N_155);
and U312 (N_312,In_372,In_254);
nor U313 (N_313,N_68,N_236);
and U314 (N_314,N_276,N_291);
nor U315 (N_315,N_288,N_220);
or U316 (N_316,N_216,N_281);
or U317 (N_317,N_181,N_265);
or U318 (N_318,N_299,N_264);
or U319 (N_319,N_89,In_67);
and U320 (N_320,N_192,In_27);
or U321 (N_321,In_121,N_295);
and U322 (N_322,In_159,In_415);
nand U323 (N_323,In_63,N_239);
or U324 (N_324,In_363,In_117);
or U325 (N_325,N_18,N_237);
nand U326 (N_326,N_251,N_110);
nor U327 (N_327,In_352,N_104);
nand U328 (N_328,N_261,In_336);
nand U329 (N_329,In_36,N_189);
nor U330 (N_330,N_130,N_115);
nand U331 (N_331,N_240,N_258);
and U332 (N_332,N_102,In_334);
nand U333 (N_333,N_200,N_175);
or U334 (N_334,N_10,N_286);
xor U335 (N_335,N_271,N_248);
nand U336 (N_336,N_205,N_173);
and U337 (N_337,N_262,In_58);
or U338 (N_338,In_144,N_274);
or U339 (N_339,N_233,N_293);
and U340 (N_340,N_255,N_231);
or U341 (N_341,In_207,N_228);
nor U342 (N_342,N_254,N_256);
or U343 (N_343,N_93,N_267);
and U344 (N_344,N_266,N_210);
nand U345 (N_345,N_142,N_47);
nand U346 (N_346,N_292,N_280);
and U347 (N_347,In_390,N_277);
and U348 (N_348,N_289,N_269);
or U349 (N_349,N_223,In_230);
or U350 (N_350,In_152,N_16);
or U351 (N_351,N_179,N_122);
and U352 (N_352,In_349,N_238);
nand U353 (N_353,N_232,N_241);
xor U354 (N_354,N_14,N_215);
nor U355 (N_355,N_283,N_290);
nand U356 (N_356,N_212,N_135);
and U357 (N_357,N_245,N_219);
and U358 (N_358,In_466,N_120);
or U359 (N_359,In_65,N_272);
nor U360 (N_360,In_118,N_176);
nand U361 (N_361,N_259,N_285);
nor U362 (N_362,N_46,In_213);
and U363 (N_363,N_214,N_207);
nand U364 (N_364,N_268,N_101);
or U365 (N_365,N_204,N_242);
or U366 (N_366,N_260,N_202);
nor U367 (N_367,In_226,In_354);
xnor U368 (N_368,N_294,N_118);
or U369 (N_369,In_460,In_87);
nand U370 (N_370,N_247,N_201);
nand U371 (N_371,In_206,N_244);
nor U372 (N_372,N_209,N_273);
and U373 (N_373,In_286,N_206);
nor U374 (N_374,N_151,In_131);
or U375 (N_375,N_296,N_235);
nand U376 (N_376,N_203,N_257);
and U377 (N_377,In_38,N_117);
or U378 (N_378,N_156,N_234);
or U379 (N_379,N_263,In_2);
xor U380 (N_380,N_3,N_224);
nor U381 (N_381,In_268,In_484);
nand U382 (N_382,N_20,N_249);
nor U383 (N_383,N_217,N_211);
and U384 (N_384,N_282,In_114);
and U385 (N_385,N_131,In_247);
and U386 (N_386,N_298,In_240);
xor U387 (N_387,In_291,In_3);
and U388 (N_388,N_246,N_284);
or U389 (N_389,N_60,N_182);
and U390 (N_390,N_278,N_222);
and U391 (N_391,N_208,In_348);
and U392 (N_392,N_252,N_253);
nand U393 (N_393,N_270,In_442);
or U394 (N_394,N_225,N_226);
and U395 (N_395,In_134,N_275);
and U396 (N_396,N_78,N_153);
or U397 (N_397,N_279,N_221);
nor U398 (N_398,In_10,N_213);
nand U399 (N_399,In_459,In_433);
or U400 (N_400,N_335,N_365);
nand U401 (N_401,N_329,N_399);
or U402 (N_402,N_342,N_367);
and U403 (N_403,N_318,N_345);
and U404 (N_404,N_389,N_300);
or U405 (N_405,N_387,N_395);
nor U406 (N_406,N_343,N_326);
nor U407 (N_407,N_353,N_306);
and U408 (N_408,N_396,N_327);
nor U409 (N_409,N_358,N_323);
nor U410 (N_410,N_336,N_320);
nand U411 (N_411,N_311,N_317);
and U412 (N_412,N_307,N_360);
and U413 (N_413,N_388,N_355);
xnor U414 (N_414,N_337,N_357);
and U415 (N_415,N_316,N_331);
or U416 (N_416,N_303,N_349);
and U417 (N_417,N_341,N_322);
nand U418 (N_418,N_370,N_375);
nand U419 (N_419,N_369,N_347);
and U420 (N_420,N_305,N_330);
nand U421 (N_421,N_364,N_302);
nor U422 (N_422,N_304,N_379);
or U423 (N_423,N_383,N_366);
nand U424 (N_424,N_376,N_313);
or U425 (N_425,N_324,N_377);
and U426 (N_426,N_392,N_344);
xnor U427 (N_427,N_372,N_381);
nand U428 (N_428,N_378,N_362);
nor U429 (N_429,N_374,N_338);
xnor U430 (N_430,N_354,N_373);
or U431 (N_431,N_328,N_384);
or U432 (N_432,N_359,N_363);
nand U433 (N_433,N_333,N_352);
nor U434 (N_434,N_356,N_346);
nor U435 (N_435,N_348,N_325);
nand U436 (N_436,N_334,N_351);
or U437 (N_437,N_308,N_368);
and U438 (N_438,N_314,N_398);
nor U439 (N_439,N_310,N_332);
or U440 (N_440,N_340,N_380);
or U441 (N_441,N_386,N_371);
and U442 (N_442,N_321,N_382);
nor U443 (N_443,N_309,N_312);
or U444 (N_444,N_319,N_391);
xor U445 (N_445,N_394,N_393);
nor U446 (N_446,N_301,N_397);
and U447 (N_447,N_361,N_339);
nor U448 (N_448,N_315,N_385);
and U449 (N_449,N_350,N_390);
or U450 (N_450,N_340,N_333);
nor U451 (N_451,N_341,N_352);
xor U452 (N_452,N_365,N_371);
and U453 (N_453,N_316,N_395);
and U454 (N_454,N_369,N_325);
nor U455 (N_455,N_324,N_305);
or U456 (N_456,N_322,N_314);
nand U457 (N_457,N_314,N_385);
nand U458 (N_458,N_328,N_392);
nand U459 (N_459,N_348,N_337);
nand U460 (N_460,N_326,N_345);
nor U461 (N_461,N_314,N_368);
nor U462 (N_462,N_353,N_399);
nor U463 (N_463,N_360,N_398);
nand U464 (N_464,N_343,N_354);
nor U465 (N_465,N_364,N_392);
nor U466 (N_466,N_396,N_336);
nand U467 (N_467,N_376,N_356);
or U468 (N_468,N_370,N_311);
and U469 (N_469,N_339,N_304);
nor U470 (N_470,N_372,N_376);
nor U471 (N_471,N_366,N_310);
nand U472 (N_472,N_345,N_351);
xnor U473 (N_473,N_359,N_349);
nand U474 (N_474,N_303,N_370);
nand U475 (N_475,N_338,N_397);
nor U476 (N_476,N_381,N_399);
nor U477 (N_477,N_319,N_389);
nor U478 (N_478,N_361,N_320);
nand U479 (N_479,N_386,N_357);
or U480 (N_480,N_362,N_375);
or U481 (N_481,N_362,N_306);
and U482 (N_482,N_328,N_343);
xnor U483 (N_483,N_366,N_319);
nand U484 (N_484,N_364,N_314);
or U485 (N_485,N_340,N_382);
or U486 (N_486,N_369,N_330);
and U487 (N_487,N_318,N_313);
nand U488 (N_488,N_347,N_368);
and U489 (N_489,N_303,N_314);
or U490 (N_490,N_376,N_329);
or U491 (N_491,N_377,N_359);
nor U492 (N_492,N_364,N_313);
and U493 (N_493,N_304,N_358);
nor U494 (N_494,N_389,N_346);
nand U495 (N_495,N_307,N_383);
or U496 (N_496,N_388,N_393);
and U497 (N_497,N_314,N_330);
and U498 (N_498,N_337,N_360);
and U499 (N_499,N_370,N_352);
and U500 (N_500,N_461,N_448);
nand U501 (N_501,N_409,N_436);
and U502 (N_502,N_497,N_414);
or U503 (N_503,N_485,N_452);
and U504 (N_504,N_421,N_442);
or U505 (N_505,N_403,N_455);
or U506 (N_506,N_410,N_457);
and U507 (N_507,N_454,N_467);
nand U508 (N_508,N_469,N_489);
or U509 (N_509,N_449,N_470);
nand U510 (N_510,N_416,N_496);
and U511 (N_511,N_431,N_479);
and U512 (N_512,N_427,N_456);
nand U513 (N_513,N_451,N_490);
and U514 (N_514,N_458,N_417);
and U515 (N_515,N_411,N_475);
nor U516 (N_516,N_493,N_419);
nor U517 (N_517,N_425,N_499);
nand U518 (N_518,N_400,N_459);
nor U519 (N_519,N_437,N_494);
nand U520 (N_520,N_412,N_420);
and U521 (N_521,N_418,N_404);
nand U522 (N_522,N_428,N_464);
and U523 (N_523,N_447,N_498);
and U524 (N_524,N_434,N_484);
and U525 (N_525,N_483,N_435);
and U526 (N_526,N_480,N_450);
and U527 (N_527,N_487,N_439);
or U528 (N_528,N_477,N_426);
and U529 (N_529,N_438,N_408);
nor U530 (N_530,N_413,N_402);
nand U531 (N_531,N_476,N_460);
and U532 (N_532,N_429,N_432);
nand U533 (N_533,N_422,N_401);
nor U534 (N_534,N_462,N_486);
and U535 (N_535,N_495,N_445);
nor U536 (N_536,N_406,N_430);
or U537 (N_537,N_463,N_405);
or U538 (N_538,N_465,N_471);
and U539 (N_539,N_443,N_488);
and U540 (N_540,N_433,N_407);
nand U541 (N_541,N_481,N_453);
nand U542 (N_542,N_482,N_491);
and U543 (N_543,N_423,N_466);
and U544 (N_544,N_492,N_446);
or U545 (N_545,N_474,N_441);
nand U546 (N_546,N_478,N_444);
nor U547 (N_547,N_424,N_472);
nor U548 (N_548,N_440,N_415);
or U549 (N_549,N_468,N_473);
xor U550 (N_550,N_405,N_434);
and U551 (N_551,N_476,N_483);
nor U552 (N_552,N_467,N_446);
and U553 (N_553,N_419,N_485);
nand U554 (N_554,N_482,N_463);
or U555 (N_555,N_496,N_499);
or U556 (N_556,N_430,N_498);
or U557 (N_557,N_456,N_422);
and U558 (N_558,N_462,N_490);
or U559 (N_559,N_456,N_479);
or U560 (N_560,N_438,N_468);
and U561 (N_561,N_438,N_420);
nand U562 (N_562,N_423,N_495);
nor U563 (N_563,N_417,N_474);
nor U564 (N_564,N_454,N_465);
and U565 (N_565,N_471,N_448);
or U566 (N_566,N_423,N_431);
nand U567 (N_567,N_417,N_407);
xnor U568 (N_568,N_410,N_406);
or U569 (N_569,N_444,N_477);
and U570 (N_570,N_428,N_495);
nor U571 (N_571,N_491,N_436);
nand U572 (N_572,N_438,N_444);
and U573 (N_573,N_448,N_407);
or U574 (N_574,N_458,N_474);
or U575 (N_575,N_488,N_466);
nor U576 (N_576,N_416,N_470);
nand U577 (N_577,N_415,N_444);
and U578 (N_578,N_443,N_434);
and U579 (N_579,N_404,N_406);
and U580 (N_580,N_463,N_498);
or U581 (N_581,N_495,N_435);
and U582 (N_582,N_415,N_408);
or U583 (N_583,N_408,N_492);
nand U584 (N_584,N_403,N_452);
and U585 (N_585,N_415,N_475);
or U586 (N_586,N_493,N_487);
or U587 (N_587,N_477,N_445);
nor U588 (N_588,N_443,N_486);
nor U589 (N_589,N_463,N_452);
nand U590 (N_590,N_444,N_483);
nand U591 (N_591,N_406,N_475);
nor U592 (N_592,N_495,N_464);
nand U593 (N_593,N_440,N_418);
nor U594 (N_594,N_474,N_462);
nand U595 (N_595,N_448,N_493);
nand U596 (N_596,N_479,N_441);
nor U597 (N_597,N_450,N_417);
nand U598 (N_598,N_458,N_407);
nand U599 (N_599,N_408,N_469);
nor U600 (N_600,N_542,N_591);
nand U601 (N_601,N_548,N_563);
nor U602 (N_602,N_567,N_571);
nand U603 (N_603,N_550,N_522);
and U604 (N_604,N_547,N_536);
or U605 (N_605,N_526,N_582);
nand U606 (N_606,N_553,N_579);
nand U607 (N_607,N_588,N_599);
or U608 (N_608,N_574,N_556);
or U609 (N_609,N_557,N_519);
nand U610 (N_610,N_512,N_590);
or U611 (N_611,N_524,N_555);
or U612 (N_612,N_545,N_534);
nand U613 (N_613,N_509,N_538);
nor U614 (N_614,N_592,N_544);
nand U615 (N_615,N_541,N_598);
nand U616 (N_616,N_559,N_546);
nand U617 (N_617,N_510,N_566);
nor U618 (N_618,N_537,N_569);
nand U619 (N_619,N_531,N_511);
nand U620 (N_620,N_551,N_530);
or U621 (N_621,N_507,N_597);
or U622 (N_622,N_521,N_596);
nor U623 (N_623,N_561,N_568);
nor U624 (N_624,N_540,N_580);
nand U625 (N_625,N_527,N_595);
or U626 (N_626,N_528,N_535);
xor U627 (N_627,N_532,N_523);
or U628 (N_628,N_520,N_572);
or U629 (N_629,N_560,N_500);
and U630 (N_630,N_533,N_583);
nand U631 (N_631,N_501,N_552);
and U632 (N_632,N_581,N_584);
nand U633 (N_633,N_593,N_586);
nor U634 (N_634,N_587,N_515);
nor U635 (N_635,N_578,N_589);
and U636 (N_636,N_506,N_539);
and U637 (N_637,N_575,N_517);
nor U638 (N_638,N_549,N_576);
nand U639 (N_639,N_529,N_558);
or U640 (N_640,N_577,N_504);
and U641 (N_641,N_513,N_503);
and U642 (N_642,N_516,N_514);
or U643 (N_643,N_585,N_518);
and U644 (N_644,N_508,N_594);
nand U645 (N_645,N_525,N_564);
or U646 (N_646,N_543,N_565);
nand U647 (N_647,N_570,N_573);
or U648 (N_648,N_562,N_554);
nand U649 (N_649,N_502,N_505);
xnor U650 (N_650,N_540,N_578);
nand U651 (N_651,N_539,N_550);
nand U652 (N_652,N_500,N_591);
and U653 (N_653,N_519,N_596);
and U654 (N_654,N_538,N_535);
nand U655 (N_655,N_564,N_501);
and U656 (N_656,N_599,N_511);
nor U657 (N_657,N_579,N_535);
and U658 (N_658,N_524,N_566);
nand U659 (N_659,N_530,N_584);
nand U660 (N_660,N_590,N_574);
nand U661 (N_661,N_539,N_525);
nand U662 (N_662,N_556,N_568);
and U663 (N_663,N_556,N_592);
or U664 (N_664,N_521,N_558);
nor U665 (N_665,N_580,N_583);
or U666 (N_666,N_593,N_529);
nand U667 (N_667,N_599,N_557);
nor U668 (N_668,N_556,N_545);
and U669 (N_669,N_524,N_571);
nand U670 (N_670,N_587,N_538);
and U671 (N_671,N_577,N_509);
or U672 (N_672,N_501,N_526);
nand U673 (N_673,N_581,N_525);
nand U674 (N_674,N_504,N_500);
nor U675 (N_675,N_529,N_515);
and U676 (N_676,N_523,N_553);
and U677 (N_677,N_586,N_568);
or U678 (N_678,N_592,N_576);
nor U679 (N_679,N_599,N_587);
nor U680 (N_680,N_518,N_510);
nor U681 (N_681,N_508,N_502);
and U682 (N_682,N_518,N_530);
nand U683 (N_683,N_581,N_557);
and U684 (N_684,N_508,N_569);
nor U685 (N_685,N_564,N_589);
or U686 (N_686,N_534,N_573);
nand U687 (N_687,N_546,N_553);
and U688 (N_688,N_549,N_541);
and U689 (N_689,N_579,N_572);
nand U690 (N_690,N_577,N_594);
or U691 (N_691,N_533,N_513);
nand U692 (N_692,N_549,N_546);
nor U693 (N_693,N_542,N_521);
nor U694 (N_694,N_564,N_575);
or U695 (N_695,N_511,N_539);
nand U696 (N_696,N_546,N_570);
or U697 (N_697,N_574,N_572);
and U698 (N_698,N_565,N_544);
nand U699 (N_699,N_564,N_569);
or U700 (N_700,N_681,N_642);
nor U701 (N_701,N_688,N_663);
or U702 (N_702,N_616,N_651);
or U703 (N_703,N_601,N_652);
or U704 (N_704,N_628,N_678);
or U705 (N_705,N_600,N_613);
and U706 (N_706,N_683,N_632);
nor U707 (N_707,N_626,N_636);
or U708 (N_708,N_672,N_620);
nand U709 (N_709,N_694,N_605);
nand U710 (N_710,N_639,N_697);
nor U711 (N_711,N_607,N_604);
nor U712 (N_712,N_679,N_675);
or U713 (N_713,N_647,N_662);
and U714 (N_714,N_656,N_657);
and U715 (N_715,N_624,N_646);
and U716 (N_716,N_634,N_643);
and U717 (N_717,N_669,N_638);
nor U718 (N_718,N_664,N_680);
xor U719 (N_719,N_644,N_625);
nand U720 (N_720,N_650,N_674);
nor U721 (N_721,N_606,N_655);
nor U722 (N_722,N_686,N_692);
or U723 (N_723,N_685,N_677);
nor U724 (N_724,N_693,N_635);
nor U725 (N_725,N_690,N_619);
nor U726 (N_726,N_673,N_684);
and U727 (N_727,N_614,N_610);
or U728 (N_728,N_676,N_691);
and U729 (N_729,N_641,N_666);
nor U730 (N_730,N_687,N_622);
nand U731 (N_731,N_671,N_670);
or U732 (N_732,N_637,N_627);
nor U733 (N_733,N_615,N_609);
or U734 (N_734,N_682,N_695);
or U735 (N_735,N_665,N_698);
nand U736 (N_736,N_630,N_611);
and U737 (N_737,N_653,N_602);
and U738 (N_738,N_648,N_659);
xor U739 (N_739,N_658,N_645);
nor U740 (N_740,N_640,N_623);
nand U741 (N_741,N_612,N_603);
nand U742 (N_742,N_696,N_668);
and U743 (N_743,N_649,N_689);
nand U744 (N_744,N_608,N_667);
and U745 (N_745,N_699,N_661);
nand U746 (N_746,N_629,N_617);
nor U747 (N_747,N_633,N_654);
or U748 (N_748,N_660,N_631);
and U749 (N_749,N_621,N_618);
and U750 (N_750,N_615,N_672);
nor U751 (N_751,N_654,N_653);
nor U752 (N_752,N_670,N_647);
or U753 (N_753,N_674,N_683);
and U754 (N_754,N_621,N_608);
or U755 (N_755,N_676,N_639);
nand U756 (N_756,N_695,N_635);
and U757 (N_757,N_654,N_601);
nand U758 (N_758,N_647,N_677);
nor U759 (N_759,N_607,N_679);
and U760 (N_760,N_626,N_666);
or U761 (N_761,N_620,N_643);
nand U762 (N_762,N_649,N_669);
or U763 (N_763,N_683,N_613);
xor U764 (N_764,N_680,N_628);
nand U765 (N_765,N_660,N_632);
or U766 (N_766,N_640,N_653);
and U767 (N_767,N_608,N_671);
nand U768 (N_768,N_685,N_663);
and U769 (N_769,N_625,N_667);
and U770 (N_770,N_662,N_653);
nor U771 (N_771,N_639,N_698);
nor U772 (N_772,N_618,N_660);
or U773 (N_773,N_621,N_693);
and U774 (N_774,N_603,N_622);
xnor U775 (N_775,N_614,N_601);
nor U776 (N_776,N_667,N_683);
nor U777 (N_777,N_666,N_683);
and U778 (N_778,N_657,N_648);
and U779 (N_779,N_627,N_626);
and U780 (N_780,N_629,N_672);
or U781 (N_781,N_655,N_699);
and U782 (N_782,N_644,N_634);
and U783 (N_783,N_670,N_664);
and U784 (N_784,N_666,N_638);
nor U785 (N_785,N_672,N_655);
and U786 (N_786,N_676,N_677);
nor U787 (N_787,N_633,N_616);
and U788 (N_788,N_608,N_676);
or U789 (N_789,N_678,N_659);
nor U790 (N_790,N_649,N_608);
nor U791 (N_791,N_633,N_634);
or U792 (N_792,N_649,N_625);
or U793 (N_793,N_699,N_652);
nand U794 (N_794,N_633,N_662);
and U795 (N_795,N_639,N_692);
nand U796 (N_796,N_620,N_609);
nand U797 (N_797,N_616,N_626);
nand U798 (N_798,N_670,N_681);
and U799 (N_799,N_662,N_686);
nor U800 (N_800,N_725,N_706);
nor U801 (N_801,N_780,N_718);
and U802 (N_802,N_733,N_737);
and U803 (N_803,N_772,N_766);
nor U804 (N_804,N_715,N_752);
nor U805 (N_805,N_764,N_713);
nand U806 (N_806,N_778,N_787);
nor U807 (N_807,N_756,N_746);
nand U808 (N_808,N_717,N_769);
xnor U809 (N_809,N_760,N_730);
nor U810 (N_810,N_736,N_792);
or U811 (N_811,N_793,N_757);
and U812 (N_812,N_726,N_739);
and U813 (N_813,N_732,N_724);
and U814 (N_814,N_765,N_742);
and U815 (N_815,N_731,N_729);
or U816 (N_816,N_723,N_781);
nand U817 (N_817,N_788,N_782);
nand U818 (N_818,N_721,N_776);
and U819 (N_819,N_709,N_702);
and U820 (N_820,N_738,N_791);
and U821 (N_821,N_798,N_763);
and U822 (N_822,N_704,N_700);
or U823 (N_823,N_761,N_748);
or U824 (N_824,N_777,N_707);
and U825 (N_825,N_749,N_786);
nand U826 (N_826,N_753,N_796);
and U827 (N_827,N_779,N_743);
or U828 (N_828,N_774,N_705);
and U829 (N_829,N_744,N_703);
nand U830 (N_830,N_741,N_799);
or U831 (N_831,N_727,N_783);
nor U832 (N_832,N_735,N_762);
or U833 (N_833,N_775,N_789);
or U834 (N_834,N_745,N_790);
and U835 (N_835,N_747,N_784);
and U836 (N_836,N_755,N_714);
or U837 (N_837,N_768,N_750);
nor U838 (N_838,N_728,N_710);
nand U839 (N_839,N_785,N_719);
and U840 (N_840,N_770,N_734);
nand U841 (N_841,N_711,N_722);
nand U842 (N_842,N_795,N_754);
nor U843 (N_843,N_773,N_759);
nor U844 (N_844,N_716,N_797);
or U845 (N_845,N_751,N_712);
nand U846 (N_846,N_794,N_767);
and U847 (N_847,N_740,N_758);
nor U848 (N_848,N_708,N_720);
or U849 (N_849,N_771,N_701);
nand U850 (N_850,N_797,N_770);
nand U851 (N_851,N_732,N_744);
or U852 (N_852,N_717,N_729);
and U853 (N_853,N_706,N_790);
or U854 (N_854,N_730,N_768);
nor U855 (N_855,N_716,N_763);
nand U856 (N_856,N_797,N_725);
nor U857 (N_857,N_739,N_781);
or U858 (N_858,N_707,N_734);
nand U859 (N_859,N_717,N_735);
nor U860 (N_860,N_760,N_731);
nand U861 (N_861,N_790,N_723);
nor U862 (N_862,N_710,N_737);
or U863 (N_863,N_798,N_742);
or U864 (N_864,N_748,N_728);
nor U865 (N_865,N_712,N_703);
and U866 (N_866,N_782,N_745);
or U867 (N_867,N_789,N_704);
nor U868 (N_868,N_770,N_715);
nand U869 (N_869,N_773,N_799);
and U870 (N_870,N_705,N_740);
nor U871 (N_871,N_751,N_738);
nor U872 (N_872,N_790,N_716);
or U873 (N_873,N_709,N_711);
nor U874 (N_874,N_715,N_780);
or U875 (N_875,N_771,N_765);
nand U876 (N_876,N_796,N_771);
or U877 (N_877,N_750,N_735);
nand U878 (N_878,N_787,N_791);
or U879 (N_879,N_701,N_785);
or U880 (N_880,N_701,N_772);
nand U881 (N_881,N_745,N_713);
nor U882 (N_882,N_713,N_784);
and U883 (N_883,N_781,N_780);
nor U884 (N_884,N_772,N_717);
nor U885 (N_885,N_794,N_749);
nand U886 (N_886,N_737,N_757);
nand U887 (N_887,N_720,N_709);
or U888 (N_888,N_783,N_769);
nor U889 (N_889,N_765,N_719);
xor U890 (N_890,N_748,N_799);
or U891 (N_891,N_712,N_783);
or U892 (N_892,N_709,N_748);
or U893 (N_893,N_775,N_724);
nor U894 (N_894,N_796,N_797);
nand U895 (N_895,N_759,N_723);
and U896 (N_896,N_721,N_713);
or U897 (N_897,N_736,N_720);
and U898 (N_898,N_749,N_743);
or U899 (N_899,N_736,N_719);
nand U900 (N_900,N_879,N_842);
and U901 (N_901,N_850,N_802);
or U902 (N_902,N_826,N_852);
and U903 (N_903,N_815,N_804);
nor U904 (N_904,N_840,N_808);
xnor U905 (N_905,N_849,N_800);
nor U906 (N_906,N_891,N_874);
or U907 (N_907,N_817,N_878);
or U908 (N_908,N_807,N_816);
or U909 (N_909,N_871,N_832);
and U910 (N_910,N_863,N_846);
and U911 (N_911,N_867,N_823);
nor U912 (N_912,N_845,N_833);
xnor U913 (N_913,N_885,N_895);
nand U914 (N_914,N_828,N_890);
nor U915 (N_915,N_825,N_824);
or U916 (N_916,N_892,N_834);
nand U917 (N_917,N_810,N_898);
and U918 (N_918,N_883,N_887);
nor U919 (N_919,N_855,N_866);
and U920 (N_920,N_827,N_872);
and U921 (N_921,N_813,N_812);
and U922 (N_922,N_856,N_820);
or U923 (N_923,N_847,N_844);
xor U924 (N_924,N_830,N_839);
nand U925 (N_925,N_899,N_848);
and U926 (N_926,N_809,N_884);
xor U927 (N_927,N_819,N_875);
nand U928 (N_928,N_893,N_853);
or U929 (N_929,N_805,N_857);
nor U930 (N_930,N_861,N_886);
and U931 (N_931,N_851,N_801);
nand U932 (N_932,N_831,N_889);
and U933 (N_933,N_859,N_860);
nor U934 (N_934,N_803,N_869);
and U935 (N_935,N_877,N_837);
or U936 (N_936,N_868,N_864);
nor U937 (N_937,N_836,N_881);
and U938 (N_938,N_876,N_888);
nand U939 (N_939,N_897,N_838);
nand U940 (N_940,N_896,N_829);
nand U941 (N_941,N_862,N_858);
nor U942 (N_942,N_870,N_854);
and U943 (N_943,N_818,N_880);
nor U944 (N_944,N_894,N_811);
nor U945 (N_945,N_822,N_873);
nor U946 (N_946,N_821,N_865);
or U947 (N_947,N_806,N_835);
nor U948 (N_948,N_841,N_843);
or U949 (N_949,N_814,N_882);
and U950 (N_950,N_830,N_858);
nor U951 (N_951,N_880,N_848);
or U952 (N_952,N_803,N_847);
and U953 (N_953,N_884,N_868);
nor U954 (N_954,N_801,N_874);
or U955 (N_955,N_845,N_884);
nand U956 (N_956,N_826,N_877);
nor U957 (N_957,N_826,N_897);
xor U958 (N_958,N_800,N_844);
nand U959 (N_959,N_812,N_832);
nor U960 (N_960,N_824,N_885);
nor U961 (N_961,N_896,N_849);
and U962 (N_962,N_866,N_891);
xor U963 (N_963,N_820,N_873);
nand U964 (N_964,N_894,N_899);
or U965 (N_965,N_846,N_820);
nand U966 (N_966,N_889,N_886);
or U967 (N_967,N_880,N_866);
and U968 (N_968,N_869,N_852);
or U969 (N_969,N_814,N_869);
nand U970 (N_970,N_806,N_898);
nand U971 (N_971,N_874,N_803);
xnor U972 (N_972,N_898,N_841);
nand U973 (N_973,N_841,N_873);
and U974 (N_974,N_856,N_808);
nand U975 (N_975,N_852,N_838);
nor U976 (N_976,N_823,N_808);
nand U977 (N_977,N_817,N_898);
nand U978 (N_978,N_847,N_831);
nor U979 (N_979,N_801,N_867);
or U980 (N_980,N_863,N_878);
nand U981 (N_981,N_867,N_870);
and U982 (N_982,N_813,N_887);
nor U983 (N_983,N_820,N_810);
nand U984 (N_984,N_867,N_875);
nor U985 (N_985,N_892,N_843);
and U986 (N_986,N_812,N_873);
and U987 (N_987,N_840,N_885);
nor U988 (N_988,N_817,N_859);
nor U989 (N_989,N_808,N_866);
and U990 (N_990,N_875,N_847);
nor U991 (N_991,N_853,N_870);
or U992 (N_992,N_810,N_811);
or U993 (N_993,N_837,N_832);
or U994 (N_994,N_887,N_803);
nand U995 (N_995,N_831,N_804);
and U996 (N_996,N_822,N_831);
and U997 (N_997,N_876,N_869);
nand U998 (N_998,N_803,N_864);
nand U999 (N_999,N_858,N_809);
or U1000 (N_1000,N_909,N_922);
or U1001 (N_1001,N_972,N_937);
nor U1002 (N_1002,N_991,N_994);
nor U1003 (N_1003,N_916,N_911);
nand U1004 (N_1004,N_958,N_927);
or U1005 (N_1005,N_944,N_970);
nor U1006 (N_1006,N_966,N_988);
and U1007 (N_1007,N_912,N_957);
nand U1008 (N_1008,N_982,N_981);
and U1009 (N_1009,N_949,N_997);
and U1010 (N_1010,N_998,N_955);
and U1011 (N_1011,N_904,N_952);
nand U1012 (N_1012,N_920,N_928);
nand U1013 (N_1013,N_942,N_987);
nor U1014 (N_1014,N_975,N_978);
nor U1015 (N_1015,N_940,N_954);
or U1016 (N_1016,N_933,N_961);
nor U1017 (N_1017,N_973,N_980);
or U1018 (N_1018,N_946,N_924);
nand U1019 (N_1019,N_979,N_930);
nor U1020 (N_1020,N_907,N_974);
nand U1021 (N_1021,N_932,N_929);
and U1022 (N_1022,N_931,N_919);
nand U1023 (N_1023,N_965,N_914);
and U1024 (N_1024,N_934,N_905);
or U1025 (N_1025,N_938,N_976);
or U1026 (N_1026,N_915,N_971);
nor U1027 (N_1027,N_983,N_951);
and U1028 (N_1028,N_967,N_950);
and U1029 (N_1029,N_996,N_993);
nand U1030 (N_1030,N_941,N_902);
or U1031 (N_1031,N_908,N_985);
xnor U1032 (N_1032,N_953,N_918);
or U1033 (N_1033,N_963,N_984);
or U1034 (N_1034,N_901,N_968);
nand U1035 (N_1035,N_921,N_917);
nand U1036 (N_1036,N_989,N_962);
xnor U1037 (N_1037,N_969,N_960);
and U1038 (N_1038,N_913,N_935);
nand U1039 (N_1039,N_925,N_939);
nand U1040 (N_1040,N_926,N_936);
nor U1041 (N_1041,N_977,N_945);
and U1042 (N_1042,N_964,N_992);
nor U1043 (N_1043,N_947,N_990);
nand U1044 (N_1044,N_995,N_999);
nand U1045 (N_1045,N_900,N_910);
or U1046 (N_1046,N_923,N_943);
or U1047 (N_1047,N_986,N_948);
and U1048 (N_1048,N_959,N_906);
and U1049 (N_1049,N_903,N_956);
nor U1050 (N_1050,N_981,N_977);
or U1051 (N_1051,N_967,N_995);
nor U1052 (N_1052,N_927,N_921);
and U1053 (N_1053,N_930,N_969);
and U1054 (N_1054,N_999,N_905);
and U1055 (N_1055,N_979,N_919);
xnor U1056 (N_1056,N_973,N_922);
nor U1057 (N_1057,N_939,N_949);
or U1058 (N_1058,N_962,N_903);
and U1059 (N_1059,N_983,N_995);
and U1060 (N_1060,N_930,N_947);
nor U1061 (N_1061,N_938,N_932);
nor U1062 (N_1062,N_924,N_966);
or U1063 (N_1063,N_938,N_946);
and U1064 (N_1064,N_933,N_996);
or U1065 (N_1065,N_950,N_959);
and U1066 (N_1066,N_954,N_992);
nand U1067 (N_1067,N_915,N_933);
nand U1068 (N_1068,N_932,N_925);
nand U1069 (N_1069,N_944,N_901);
nor U1070 (N_1070,N_983,N_972);
nand U1071 (N_1071,N_967,N_949);
nor U1072 (N_1072,N_952,N_958);
and U1073 (N_1073,N_982,N_965);
xor U1074 (N_1074,N_960,N_911);
and U1075 (N_1075,N_953,N_938);
xnor U1076 (N_1076,N_982,N_992);
nand U1077 (N_1077,N_994,N_955);
nand U1078 (N_1078,N_975,N_927);
nor U1079 (N_1079,N_953,N_926);
nand U1080 (N_1080,N_947,N_901);
or U1081 (N_1081,N_937,N_905);
nand U1082 (N_1082,N_908,N_913);
nor U1083 (N_1083,N_967,N_997);
or U1084 (N_1084,N_935,N_941);
and U1085 (N_1085,N_912,N_950);
xnor U1086 (N_1086,N_900,N_939);
nand U1087 (N_1087,N_934,N_912);
or U1088 (N_1088,N_930,N_992);
or U1089 (N_1089,N_922,N_977);
or U1090 (N_1090,N_908,N_945);
and U1091 (N_1091,N_903,N_973);
nor U1092 (N_1092,N_923,N_914);
or U1093 (N_1093,N_995,N_943);
xnor U1094 (N_1094,N_925,N_923);
or U1095 (N_1095,N_989,N_916);
or U1096 (N_1096,N_955,N_932);
or U1097 (N_1097,N_983,N_942);
or U1098 (N_1098,N_959,N_952);
nor U1099 (N_1099,N_979,N_947);
nand U1100 (N_1100,N_1083,N_1038);
nor U1101 (N_1101,N_1000,N_1001);
or U1102 (N_1102,N_1020,N_1042);
or U1103 (N_1103,N_1035,N_1071);
nor U1104 (N_1104,N_1014,N_1079);
and U1105 (N_1105,N_1072,N_1027);
nor U1106 (N_1106,N_1056,N_1043);
nor U1107 (N_1107,N_1099,N_1007);
nand U1108 (N_1108,N_1077,N_1095);
nor U1109 (N_1109,N_1082,N_1004);
nand U1110 (N_1110,N_1045,N_1049);
and U1111 (N_1111,N_1025,N_1070);
nand U1112 (N_1112,N_1006,N_1030);
nor U1113 (N_1113,N_1063,N_1033);
xnor U1114 (N_1114,N_1075,N_1058);
and U1115 (N_1115,N_1005,N_1066);
nor U1116 (N_1116,N_1003,N_1022);
or U1117 (N_1117,N_1009,N_1029);
and U1118 (N_1118,N_1039,N_1054);
nor U1119 (N_1119,N_1073,N_1018);
and U1120 (N_1120,N_1037,N_1047);
nand U1121 (N_1121,N_1080,N_1060);
nand U1122 (N_1122,N_1008,N_1028);
or U1123 (N_1123,N_1044,N_1097);
and U1124 (N_1124,N_1088,N_1057);
or U1125 (N_1125,N_1062,N_1064);
nor U1126 (N_1126,N_1052,N_1051);
xnor U1127 (N_1127,N_1032,N_1016);
nand U1128 (N_1128,N_1026,N_1085);
nand U1129 (N_1129,N_1041,N_1086);
xor U1130 (N_1130,N_1096,N_1050);
and U1131 (N_1131,N_1040,N_1021);
nor U1132 (N_1132,N_1011,N_1087);
or U1133 (N_1133,N_1048,N_1076);
nand U1134 (N_1134,N_1031,N_1002);
and U1135 (N_1135,N_1092,N_1068);
and U1136 (N_1136,N_1067,N_1091);
nand U1137 (N_1137,N_1017,N_1089);
and U1138 (N_1138,N_1053,N_1046);
nor U1139 (N_1139,N_1036,N_1013);
and U1140 (N_1140,N_1012,N_1069);
and U1141 (N_1141,N_1015,N_1090);
nand U1142 (N_1142,N_1061,N_1024);
nor U1143 (N_1143,N_1059,N_1098);
or U1144 (N_1144,N_1093,N_1019);
or U1145 (N_1145,N_1074,N_1065);
nand U1146 (N_1146,N_1010,N_1055);
nor U1147 (N_1147,N_1094,N_1034);
xor U1148 (N_1148,N_1081,N_1023);
nand U1149 (N_1149,N_1078,N_1084);
and U1150 (N_1150,N_1043,N_1061);
xor U1151 (N_1151,N_1014,N_1088);
nor U1152 (N_1152,N_1069,N_1076);
nand U1153 (N_1153,N_1050,N_1043);
nand U1154 (N_1154,N_1005,N_1072);
nand U1155 (N_1155,N_1076,N_1068);
and U1156 (N_1156,N_1042,N_1047);
xnor U1157 (N_1157,N_1073,N_1017);
and U1158 (N_1158,N_1036,N_1062);
or U1159 (N_1159,N_1085,N_1064);
nor U1160 (N_1160,N_1073,N_1050);
and U1161 (N_1161,N_1081,N_1094);
or U1162 (N_1162,N_1022,N_1048);
nand U1163 (N_1163,N_1070,N_1069);
and U1164 (N_1164,N_1075,N_1004);
and U1165 (N_1165,N_1001,N_1073);
and U1166 (N_1166,N_1003,N_1051);
or U1167 (N_1167,N_1014,N_1043);
and U1168 (N_1168,N_1023,N_1024);
nor U1169 (N_1169,N_1000,N_1098);
or U1170 (N_1170,N_1046,N_1026);
or U1171 (N_1171,N_1021,N_1025);
nand U1172 (N_1172,N_1096,N_1061);
nand U1173 (N_1173,N_1009,N_1005);
xnor U1174 (N_1174,N_1050,N_1005);
or U1175 (N_1175,N_1086,N_1030);
and U1176 (N_1176,N_1083,N_1003);
nand U1177 (N_1177,N_1098,N_1067);
nor U1178 (N_1178,N_1007,N_1066);
nand U1179 (N_1179,N_1049,N_1029);
and U1180 (N_1180,N_1045,N_1028);
nor U1181 (N_1181,N_1047,N_1090);
or U1182 (N_1182,N_1088,N_1076);
nor U1183 (N_1183,N_1060,N_1042);
and U1184 (N_1184,N_1063,N_1047);
and U1185 (N_1185,N_1088,N_1098);
or U1186 (N_1186,N_1020,N_1003);
nor U1187 (N_1187,N_1098,N_1090);
or U1188 (N_1188,N_1060,N_1004);
and U1189 (N_1189,N_1074,N_1070);
or U1190 (N_1190,N_1049,N_1096);
nand U1191 (N_1191,N_1034,N_1033);
nand U1192 (N_1192,N_1081,N_1056);
and U1193 (N_1193,N_1099,N_1084);
and U1194 (N_1194,N_1070,N_1057);
and U1195 (N_1195,N_1052,N_1067);
or U1196 (N_1196,N_1036,N_1015);
nand U1197 (N_1197,N_1074,N_1034);
and U1198 (N_1198,N_1017,N_1000);
or U1199 (N_1199,N_1045,N_1054);
and U1200 (N_1200,N_1130,N_1148);
nand U1201 (N_1201,N_1110,N_1112);
nand U1202 (N_1202,N_1188,N_1151);
nand U1203 (N_1203,N_1144,N_1194);
and U1204 (N_1204,N_1101,N_1184);
nor U1205 (N_1205,N_1199,N_1172);
or U1206 (N_1206,N_1161,N_1193);
xnor U1207 (N_1207,N_1155,N_1189);
or U1208 (N_1208,N_1134,N_1106);
or U1209 (N_1209,N_1179,N_1137);
nor U1210 (N_1210,N_1141,N_1177);
nor U1211 (N_1211,N_1173,N_1181);
nand U1212 (N_1212,N_1187,N_1128);
nand U1213 (N_1213,N_1158,N_1191);
nor U1214 (N_1214,N_1147,N_1162);
or U1215 (N_1215,N_1104,N_1183);
or U1216 (N_1216,N_1135,N_1160);
and U1217 (N_1217,N_1157,N_1127);
or U1218 (N_1218,N_1165,N_1136);
or U1219 (N_1219,N_1195,N_1196);
nor U1220 (N_1220,N_1175,N_1111);
and U1221 (N_1221,N_1107,N_1114);
nor U1222 (N_1222,N_1124,N_1109);
or U1223 (N_1223,N_1108,N_1156);
or U1224 (N_1224,N_1198,N_1145);
or U1225 (N_1225,N_1117,N_1190);
nand U1226 (N_1226,N_1143,N_1105);
nor U1227 (N_1227,N_1166,N_1153);
nor U1228 (N_1228,N_1182,N_1164);
and U1229 (N_1229,N_1100,N_1131);
nor U1230 (N_1230,N_1150,N_1192);
nand U1231 (N_1231,N_1170,N_1154);
nand U1232 (N_1232,N_1103,N_1120);
nand U1233 (N_1233,N_1163,N_1123);
or U1234 (N_1234,N_1159,N_1149);
nor U1235 (N_1235,N_1139,N_1176);
or U1236 (N_1236,N_1180,N_1186);
nand U1237 (N_1237,N_1174,N_1132);
nand U1238 (N_1238,N_1113,N_1133);
nand U1239 (N_1239,N_1152,N_1169);
and U1240 (N_1240,N_1142,N_1140);
or U1241 (N_1241,N_1129,N_1197);
and U1242 (N_1242,N_1102,N_1126);
or U1243 (N_1243,N_1115,N_1121);
or U1244 (N_1244,N_1138,N_1168);
nor U1245 (N_1245,N_1116,N_1171);
xor U1246 (N_1246,N_1185,N_1119);
nor U1247 (N_1247,N_1146,N_1178);
and U1248 (N_1248,N_1118,N_1122);
xnor U1249 (N_1249,N_1167,N_1125);
or U1250 (N_1250,N_1155,N_1191);
and U1251 (N_1251,N_1109,N_1105);
or U1252 (N_1252,N_1138,N_1157);
and U1253 (N_1253,N_1118,N_1194);
nor U1254 (N_1254,N_1117,N_1149);
or U1255 (N_1255,N_1110,N_1103);
or U1256 (N_1256,N_1192,N_1129);
or U1257 (N_1257,N_1138,N_1137);
nand U1258 (N_1258,N_1130,N_1179);
nand U1259 (N_1259,N_1165,N_1161);
and U1260 (N_1260,N_1150,N_1100);
or U1261 (N_1261,N_1188,N_1153);
and U1262 (N_1262,N_1162,N_1175);
nor U1263 (N_1263,N_1107,N_1189);
or U1264 (N_1264,N_1153,N_1105);
xnor U1265 (N_1265,N_1176,N_1124);
and U1266 (N_1266,N_1158,N_1153);
nor U1267 (N_1267,N_1120,N_1123);
or U1268 (N_1268,N_1106,N_1168);
or U1269 (N_1269,N_1181,N_1143);
nor U1270 (N_1270,N_1139,N_1179);
nand U1271 (N_1271,N_1145,N_1195);
nand U1272 (N_1272,N_1145,N_1178);
or U1273 (N_1273,N_1157,N_1133);
nor U1274 (N_1274,N_1150,N_1102);
and U1275 (N_1275,N_1163,N_1118);
or U1276 (N_1276,N_1185,N_1165);
and U1277 (N_1277,N_1184,N_1148);
nor U1278 (N_1278,N_1114,N_1173);
or U1279 (N_1279,N_1191,N_1123);
nor U1280 (N_1280,N_1182,N_1124);
nor U1281 (N_1281,N_1163,N_1139);
nand U1282 (N_1282,N_1180,N_1136);
nor U1283 (N_1283,N_1156,N_1136);
nor U1284 (N_1284,N_1100,N_1130);
nand U1285 (N_1285,N_1119,N_1173);
or U1286 (N_1286,N_1141,N_1122);
and U1287 (N_1287,N_1180,N_1179);
or U1288 (N_1288,N_1105,N_1166);
or U1289 (N_1289,N_1118,N_1127);
nand U1290 (N_1290,N_1121,N_1144);
and U1291 (N_1291,N_1114,N_1106);
or U1292 (N_1292,N_1187,N_1195);
and U1293 (N_1293,N_1106,N_1115);
or U1294 (N_1294,N_1193,N_1192);
nand U1295 (N_1295,N_1102,N_1136);
or U1296 (N_1296,N_1177,N_1175);
and U1297 (N_1297,N_1128,N_1116);
or U1298 (N_1298,N_1159,N_1179);
nand U1299 (N_1299,N_1122,N_1110);
or U1300 (N_1300,N_1213,N_1202);
nand U1301 (N_1301,N_1249,N_1283);
nand U1302 (N_1302,N_1244,N_1203);
and U1303 (N_1303,N_1254,N_1210);
or U1304 (N_1304,N_1239,N_1257);
or U1305 (N_1305,N_1215,N_1299);
or U1306 (N_1306,N_1242,N_1209);
nor U1307 (N_1307,N_1258,N_1245);
nand U1308 (N_1308,N_1201,N_1216);
or U1309 (N_1309,N_1217,N_1279);
nand U1310 (N_1310,N_1265,N_1241);
and U1311 (N_1311,N_1273,N_1234);
nor U1312 (N_1312,N_1207,N_1218);
or U1313 (N_1313,N_1205,N_1272);
or U1314 (N_1314,N_1286,N_1208);
nor U1315 (N_1315,N_1219,N_1206);
nor U1316 (N_1316,N_1295,N_1292);
or U1317 (N_1317,N_1296,N_1264);
or U1318 (N_1318,N_1277,N_1280);
nand U1319 (N_1319,N_1268,N_1220);
nor U1320 (N_1320,N_1289,N_1236);
and U1321 (N_1321,N_1260,N_1246);
xnor U1322 (N_1322,N_1243,N_1224);
nor U1323 (N_1323,N_1255,N_1287);
nand U1324 (N_1324,N_1297,N_1285);
nor U1325 (N_1325,N_1212,N_1253);
nor U1326 (N_1326,N_1270,N_1291);
nand U1327 (N_1327,N_1235,N_1238);
and U1328 (N_1328,N_1269,N_1223);
and U1329 (N_1329,N_1227,N_1267);
nor U1330 (N_1330,N_1232,N_1230);
nand U1331 (N_1331,N_1261,N_1233);
nand U1332 (N_1332,N_1250,N_1262);
or U1333 (N_1333,N_1252,N_1211);
or U1334 (N_1334,N_1259,N_1274);
nand U1335 (N_1335,N_1221,N_1293);
nand U1336 (N_1336,N_1251,N_1226);
nand U1337 (N_1337,N_1298,N_1256);
nor U1338 (N_1338,N_1284,N_1266);
or U1339 (N_1339,N_1214,N_1228);
nand U1340 (N_1340,N_1200,N_1204);
or U1341 (N_1341,N_1222,N_1247);
nand U1342 (N_1342,N_1263,N_1225);
or U1343 (N_1343,N_1294,N_1278);
and U1344 (N_1344,N_1229,N_1231);
and U1345 (N_1345,N_1276,N_1281);
nand U1346 (N_1346,N_1248,N_1240);
or U1347 (N_1347,N_1271,N_1290);
nor U1348 (N_1348,N_1237,N_1275);
nand U1349 (N_1349,N_1282,N_1288);
nand U1350 (N_1350,N_1256,N_1254);
nor U1351 (N_1351,N_1262,N_1233);
nand U1352 (N_1352,N_1217,N_1207);
or U1353 (N_1353,N_1250,N_1297);
nand U1354 (N_1354,N_1258,N_1211);
and U1355 (N_1355,N_1255,N_1209);
or U1356 (N_1356,N_1292,N_1248);
nor U1357 (N_1357,N_1269,N_1245);
nor U1358 (N_1358,N_1236,N_1203);
and U1359 (N_1359,N_1265,N_1266);
nand U1360 (N_1360,N_1217,N_1222);
nor U1361 (N_1361,N_1258,N_1200);
or U1362 (N_1362,N_1298,N_1231);
or U1363 (N_1363,N_1263,N_1215);
nor U1364 (N_1364,N_1201,N_1262);
nor U1365 (N_1365,N_1221,N_1251);
or U1366 (N_1366,N_1297,N_1233);
nand U1367 (N_1367,N_1222,N_1227);
and U1368 (N_1368,N_1294,N_1279);
or U1369 (N_1369,N_1271,N_1237);
and U1370 (N_1370,N_1290,N_1224);
nand U1371 (N_1371,N_1263,N_1201);
nor U1372 (N_1372,N_1250,N_1205);
nor U1373 (N_1373,N_1283,N_1228);
nor U1374 (N_1374,N_1272,N_1212);
or U1375 (N_1375,N_1271,N_1239);
nand U1376 (N_1376,N_1255,N_1200);
xnor U1377 (N_1377,N_1285,N_1269);
and U1378 (N_1378,N_1209,N_1285);
nand U1379 (N_1379,N_1227,N_1289);
nand U1380 (N_1380,N_1240,N_1252);
nand U1381 (N_1381,N_1225,N_1208);
nor U1382 (N_1382,N_1211,N_1269);
nor U1383 (N_1383,N_1247,N_1287);
and U1384 (N_1384,N_1294,N_1209);
or U1385 (N_1385,N_1292,N_1209);
or U1386 (N_1386,N_1212,N_1215);
and U1387 (N_1387,N_1230,N_1277);
and U1388 (N_1388,N_1237,N_1260);
and U1389 (N_1389,N_1250,N_1254);
nor U1390 (N_1390,N_1246,N_1207);
and U1391 (N_1391,N_1234,N_1250);
xor U1392 (N_1392,N_1261,N_1218);
and U1393 (N_1393,N_1209,N_1261);
or U1394 (N_1394,N_1277,N_1214);
or U1395 (N_1395,N_1225,N_1298);
or U1396 (N_1396,N_1230,N_1262);
or U1397 (N_1397,N_1232,N_1220);
nor U1398 (N_1398,N_1283,N_1280);
or U1399 (N_1399,N_1210,N_1232);
nor U1400 (N_1400,N_1320,N_1334);
nor U1401 (N_1401,N_1373,N_1367);
nor U1402 (N_1402,N_1384,N_1363);
and U1403 (N_1403,N_1398,N_1396);
and U1404 (N_1404,N_1343,N_1355);
xor U1405 (N_1405,N_1309,N_1395);
nor U1406 (N_1406,N_1324,N_1341);
nand U1407 (N_1407,N_1399,N_1357);
nor U1408 (N_1408,N_1331,N_1305);
nor U1409 (N_1409,N_1323,N_1347);
nand U1410 (N_1410,N_1374,N_1372);
and U1411 (N_1411,N_1319,N_1386);
or U1412 (N_1412,N_1371,N_1356);
or U1413 (N_1413,N_1389,N_1311);
nand U1414 (N_1414,N_1333,N_1313);
and U1415 (N_1415,N_1383,N_1344);
or U1416 (N_1416,N_1361,N_1364);
nor U1417 (N_1417,N_1397,N_1329);
nor U1418 (N_1418,N_1304,N_1394);
and U1419 (N_1419,N_1376,N_1314);
nor U1420 (N_1420,N_1349,N_1327);
or U1421 (N_1421,N_1370,N_1351);
nand U1422 (N_1422,N_1317,N_1303);
or U1423 (N_1423,N_1316,N_1381);
nand U1424 (N_1424,N_1391,N_1359);
nand U1425 (N_1425,N_1346,N_1382);
nor U1426 (N_1426,N_1368,N_1328);
nor U1427 (N_1427,N_1369,N_1390);
or U1428 (N_1428,N_1360,N_1393);
nand U1429 (N_1429,N_1307,N_1308);
nand U1430 (N_1430,N_1350,N_1337);
and U1431 (N_1431,N_1339,N_1322);
nand U1432 (N_1432,N_1300,N_1326);
or U1433 (N_1433,N_1336,N_1378);
nand U1434 (N_1434,N_1358,N_1353);
or U1435 (N_1435,N_1377,N_1354);
or U1436 (N_1436,N_1338,N_1345);
nor U1437 (N_1437,N_1301,N_1302);
nand U1438 (N_1438,N_1387,N_1330);
nor U1439 (N_1439,N_1366,N_1312);
or U1440 (N_1440,N_1348,N_1385);
nand U1441 (N_1441,N_1325,N_1340);
and U1442 (N_1442,N_1392,N_1332);
nor U1443 (N_1443,N_1306,N_1388);
nand U1444 (N_1444,N_1335,N_1318);
or U1445 (N_1445,N_1352,N_1380);
nand U1446 (N_1446,N_1321,N_1362);
or U1447 (N_1447,N_1365,N_1310);
nand U1448 (N_1448,N_1315,N_1375);
nor U1449 (N_1449,N_1342,N_1379);
nand U1450 (N_1450,N_1377,N_1388);
and U1451 (N_1451,N_1326,N_1373);
and U1452 (N_1452,N_1387,N_1353);
and U1453 (N_1453,N_1313,N_1305);
and U1454 (N_1454,N_1381,N_1317);
and U1455 (N_1455,N_1383,N_1327);
nand U1456 (N_1456,N_1362,N_1315);
nor U1457 (N_1457,N_1339,N_1382);
nand U1458 (N_1458,N_1311,N_1388);
nor U1459 (N_1459,N_1313,N_1369);
and U1460 (N_1460,N_1371,N_1342);
nor U1461 (N_1461,N_1336,N_1362);
nor U1462 (N_1462,N_1346,N_1361);
and U1463 (N_1463,N_1368,N_1355);
or U1464 (N_1464,N_1361,N_1340);
or U1465 (N_1465,N_1312,N_1369);
or U1466 (N_1466,N_1388,N_1359);
nor U1467 (N_1467,N_1377,N_1386);
nand U1468 (N_1468,N_1394,N_1305);
nor U1469 (N_1469,N_1319,N_1379);
nand U1470 (N_1470,N_1336,N_1347);
and U1471 (N_1471,N_1373,N_1376);
nand U1472 (N_1472,N_1305,N_1397);
nor U1473 (N_1473,N_1373,N_1344);
or U1474 (N_1474,N_1320,N_1307);
or U1475 (N_1475,N_1394,N_1316);
xnor U1476 (N_1476,N_1323,N_1322);
nor U1477 (N_1477,N_1334,N_1374);
nor U1478 (N_1478,N_1326,N_1398);
or U1479 (N_1479,N_1339,N_1385);
or U1480 (N_1480,N_1373,N_1337);
and U1481 (N_1481,N_1345,N_1371);
nor U1482 (N_1482,N_1381,N_1327);
or U1483 (N_1483,N_1398,N_1337);
nor U1484 (N_1484,N_1397,N_1339);
nand U1485 (N_1485,N_1300,N_1366);
nand U1486 (N_1486,N_1388,N_1345);
and U1487 (N_1487,N_1336,N_1368);
nor U1488 (N_1488,N_1312,N_1361);
or U1489 (N_1489,N_1311,N_1349);
nand U1490 (N_1490,N_1315,N_1331);
nand U1491 (N_1491,N_1347,N_1358);
or U1492 (N_1492,N_1360,N_1357);
or U1493 (N_1493,N_1322,N_1387);
nand U1494 (N_1494,N_1334,N_1369);
nor U1495 (N_1495,N_1300,N_1327);
nand U1496 (N_1496,N_1376,N_1355);
or U1497 (N_1497,N_1315,N_1368);
nor U1498 (N_1498,N_1383,N_1345);
or U1499 (N_1499,N_1339,N_1374);
nand U1500 (N_1500,N_1470,N_1414);
or U1501 (N_1501,N_1449,N_1443);
and U1502 (N_1502,N_1413,N_1483);
or U1503 (N_1503,N_1447,N_1405);
or U1504 (N_1504,N_1490,N_1478);
or U1505 (N_1505,N_1431,N_1499);
or U1506 (N_1506,N_1426,N_1428);
nand U1507 (N_1507,N_1464,N_1412);
nor U1508 (N_1508,N_1438,N_1466);
or U1509 (N_1509,N_1458,N_1404);
nand U1510 (N_1510,N_1430,N_1422);
or U1511 (N_1511,N_1460,N_1463);
and U1512 (N_1512,N_1493,N_1435);
nor U1513 (N_1513,N_1419,N_1467);
and U1514 (N_1514,N_1473,N_1498);
nor U1515 (N_1515,N_1417,N_1420);
and U1516 (N_1516,N_1400,N_1471);
nand U1517 (N_1517,N_1454,N_1481);
nand U1518 (N_1518,N_1432,N_1456);
or U1519 (N_1519,N_1444,N_1486);
and U1520 (N_1520,N_1459,N_1427);
nor U1521 (N_1521,N_1415,N_1429);
and U1522 (N_1522,N_1479,N_1434);
and U1523 (N_1523,N_1461,N_1406);
nor U1524 (N_1524,N_1453,N_1497);
or U1525 (N_1525,N_1475,N_1441);
or U1526 (N_1526,N_1424,N_1448);
or U1527 (N_1527,N_1446,N_1425);
and U1528 (N_1528,N_1480,N_1442);
nand U1529 (N_1529,N_1439,N_1418);
nor U1530 (N_1530,N_1437,N_1484);
nand U1531 (N_1531,N_1474,N_1410);
or U1532 (N_1532,N_1476,N_1465);
nand U1533 (N_1533,N_1407,N_1495);
or U1534 (N_1534,N_1403,N_1482);
or U1535 (N_1535,N_1457,N_1416);
and U1536 (N_1536,N_1402,N_1487);
nand U1537 (N_1537,N_1409,N_1452);
nand U1538 (N_1538,N_1492,N_1451);
and U1539 (N_1539,N_1445,N_1401);
and U1540 (N_1540,N_1491,N_1440);
and U1541 (N_1541,N_1455,N_1411);
nand U1542 (N_1542,N_1472,N_1433);
or U1543 (N_1543,N_1477,N_1496);
nor U1544 (N_1544,N_1468,N_1436);
or U1545 (N_1545,N_1450,N_1489);
or U1546 (N_1546,N_1421,N_1494);
and U1547 (N_1547,N_1485,N_1488);
or U1548 (N_1548,N_1469,N_1423);
or U1549 (N_1549,N_1462,N_1408);
or U1550 (N_1550,N_1412,N_1462);
nor U1551 (N_1551,N_1499,N_1450);
nor U1552 (N_1552,N_1476,N_1405);
nand U1553 (N_1553,N_1487,N_1431);
and U1554 (N_1554,N_1488,N_1487);
or U1555 (N_1555,N_1400,N_1488);
nand U1556 (N_1556,N_1417,N_1469);
or U1557 (N_1557,N_1438,N_1482);
and U1558 (N_1558,N_1481,N_1483);
nand U1559 (N_1559,N_1487,N_1435);
nand U1560 (N_1560,N_1406,N_1469);
and U1561 (N_1561,N_1496,N_1497);
or U1562 (N_1562,N_1468,N_1483);
or U1563 (N_1563,N_1459,N_1433);
and U1564 (N_1564,N_1449,N_1439);
and U1565 (N_1565,N_1441,N_1420);
and U1566 (N_1566,N_1494,N_1483);
nand U1567 (N_1567,N_1470,N_1493);
nand U1568 (N_1568,N_1494,N_1423);
or U1569 (N_1569,N_1432,N_1406);
nor U1570 (N_1570,N_1439,N_1424);
xor U1571 (N_1571,N_1416,N_1434);
nand U1572 (N_1572,N_1431,N_1439);
nand U1573 (N_1573,N_1407,N_1481);
and U1574 (N_1574,N_1478,N_1461);
or U1575 (N_1575,N_1413,N_1489);
nor U1576 (N_1576,N_1483,N_1491);
nand U1577 (N_1577,N_1424,N_1489);
and U1578 (N_1578,N_1429,N_1436);
and U1579 (N_1579,N_1438,N_1420);
or U1580 (N_1580,N_1414,N_1406);
xnor U1581 (N_1581,N_1432,N_1476);
xor U1582 (N_1582,N_1494,N_1410);
and U1583 (N_1583,N_1490,N_1439);
or U1584 (N_1584,N_1483,N_1403);
and U1585 (N_1585,N_1494,N_1471);
nand U1586 (N_1586,N_1431,N_1428);
nand U1587 (N_1587,N_1403,N_1477);
nand U1588 (N_1588,N_1430,N_1467);
nor U1589 (N_1589,N_1440,N_1411);
or U1590 (N_1590,N_1465,N_1449);
nor U1591 (N_1591,N_1468,N_1424);
and U1592 (N_1592,N_1423,N_1409);
or U1593 (N_1593,N_1434,N_1493);
nand U1594 (N_1594,N_1429,N_1492);
and U1595 (N_1595,N_1416,N_1486);
nand U1596 (N_1596,N_1461,N_1442);
or U1597 (N_1597,N_1447,N_1457);
nand U1598 (N_1598,N_1430,N_1400);
nand U1599 (N_1599,N_1401,N_1436);
nand U1600 (N_1600,N_1573,N_1565);
and U1601 (N_1601,N_1572,N_1590);
or U1602 (N_1602,N_1562,N_1555);
or U1603 (N_1603,N_1557,N_1540);
or U1604 (N_1604,N_1541,N_1570);
or U1605 (N_1605,N_1509,N_1505);
or U1606 (N_1606,N_1546,N_1550);
and U1607 (N_1607,N_1584,N_1560);
or U1608 (N_1608,N_1585,N_1551);
or U1609 (N_1609,N_1574,N_1580);
and U1610 (N_1610,N_1535,N_1524);
nand U1611 (N_1611,N_1503,N_1598);
or U1612 (N_1612,N_1587,N_1523);
and U1613 (N_1613,N_1538,N_1553);
and U1614 (N_1614,N_1531,N_1508);
or U1615 (N_1615,N_1589,N_1593);
and U1616 (N_1616,N_1561,N_1504);
nand U1617 (N_1617,N_1594,N_1571);
nand U1618 (N_1618,N_1554,N_1542);
nand U1619 (N_1619,N_1596,N_1525);
nor U1620 (N_1620,N_1543,N_1513);
nor U1621 (N_1621,N_1521,N_1556);
and U1622 (N_1622,N_1586,N_1578);
or U1623 (N_1623,N_1592,N_1519);
or U1624 (N_1624,N_1597,N_1518);
and U1625 (N_1625,N_1510,N_1577);
and U1626 (N_1626,N_1545,N_1549);
nand U1627 (N_1627,N_1563,N_1530);
nand U1628 (N_1628,N_1502,N_1595);
and U1629 (N_1629,N_1537,N_1599);
nand U1630 (N_1630,N_1569,N_1564);
nand U1631 (N_1631,N_1516,N_1501);
nor U1632 (N_1632,N_1576,N_1512);
xnor U1633 (N_1633,N_1514,N_1506);
nand U1634 (N_1634,N_1533,N_1575);
or U1635 (N_1635,N_1520,N_1588);
nor U1636 (N_1636,N_1500,N_1529);
or U1637 (N_1637,N_1527,N_1526);
nor U1638 (N_1638,N_1511,N_1591);
and U1639 (N_1639,N_1522,N_1539);
nor U1640 (N_1640,N_1544,N_1579);
nor U1641 (N_1641,N_1552,N_1507);
nor U1642 (N_1642,N_1581,N_1547);
nor U1643 (N_1643,N_1582,N_1558);
and U1644 (N_1644,N_1548,N_1559);
nor U1645 (N_1645,N_1515,N_1534);
or U1646 (N_1646,N_1567,N_1536);
nor U1647 (N_1647,N_1583,N_1528);
xnor U1648 (N_1648,N_1566,N_1517);
and U1649 (N_1649,N_1568,N_1532);
nor U1650 (N_1650,N_1591,N_1563);
or U1651 (N_1651,N_1582,N_1568);
and U1652 (N_1652,N_1501,N_1592);
and U1653 (N_1653,N_1599,N_1516);
and U1654 (N_1654,N_1567,N_1532);
nand U1655 (N_1655,N_1514,N_1569);
nor U1656 (N_1656,N_1549,N_1566);
or U1657 (N_1657,N_1501,N_1574);
nand U1658 (N_1658,N_1506,N_1565);
or U1659 (N_1659,N_1564,N_1592);
nand U1660 (N_1660,N_1575,N_1528);
and U1661 (N_1661,N_1526,N_1517);
nand U1662 (N_1662,N_1541,N_1574);
nand U1663 (N_1663,N_1542,N_1514);
nor U1664 (N_1664,N_1510,N_1558);
and U1665 (N_1665,N_1517,N_1535);
and U1666 (N_1666,N_1517,N_1524);
or U1667 (N_1667,N_1554,N_1540);
and U1668 (N_1668,N_1584,N_1577);
or U1669 (N_1669,N_1587,N_1508);
nand U1670 (N_1670,N_1510,N_1596);
xor U1671 (N_1671,N_1507,N_1570);
nand U1672 (N_1672,N_1545,N_1524);
or U1673 (N_1673,N_1587,N_1532);
and U1674 (N_1674,N_1530,N_1574);
and U1675 (N_1675,N_1581,N_1531);
nand U1676 (N_1676,N_1526,N_1586);
and U1677 (N_1677,N_1503,N_1595);
nor U1678 (N_1678,N_1557,N_1538);
nand U1679 (N_1679,N_1599,N_1520);
or U1680 (N_1680,N_1575,N_1518);
and U1681 (N_1681,N_1526,N_1522);
nand U1682 (N_1682,N_1556,N_1577);
and U1683 (N_1683,N_1504,N_1551);
nand U1684 (N_1684,N_1525,N_1566);
and U1685 (N_1685,N_1552,N_1549);
and U1686 (N_1686,N_1530,N_1550);
nand U1687 (N_1687,N_1564,N_1554);
nand U1688 (N_1688,N_1554,N_1534);
and U1689 (N_1689,N_1540,N_1590);
or U1690 (N_1690,N_1514,N_1556);
nor U1691 (N_1691,N_1522,N_1529);
and U1692 (N_1692,N_1513,N_1588);
and U1693 (N_1693,N_1590,N_1522);
or U1694 (N_1694,N_1514,N_1591);
nand U1695 (N_1695,N_1582,N_1564);
and U1696 (N_1696,N_1542,N_1503);
and U1697 (N_1697,N_1593,N_1521);
and U1698 (N_1698,N_1579,N_1574);
nor U1699 (N_1699,N_1504,N_1533);
nor U1700 (N_1700,N_1605,N_1638);
nor U1701 (N_1701,N_1662,N_1698);
nor U1702 (N_1702,N_1684,N_1602);
or U1703 (N_1703,N_1601,N_1603);
xnor U1704 (N_1704,N_1647,N_1641);
and U1705 (N_1705,N_1658,N_1681);
and U1706 (N_1706,N_1648,N_1651);
or U1707 (N_1707,N_1674,N_1610);
and U1708 (N_1708,N_1693,N_1654);
or U1709 (N_1709,N_1615,N_1628);
and U1710 (N_1710,N_1606,N_1653);
nor U1711 (N_1711,N_1696,N_1614);
nand U1712 (N_1712,N_1600,N_1652);
nand U1713 (N_1713,N_1666,N_1687);
nor U1714 (N_1714,N_1669,N_1676);
or U1715 (N_1715,N_1612,N_1631);
nor U1716 (N_1716,N_1619,N_1649);
and U1717 (N_1717,N_1624,N_1673);
and U1718 (N_1718,N_1639,N_1692);
nor U1719 (N_1719,N_1630,N_1618);
nor U1720 (N_1720,N_1689,N_1663);
nor U1721 (N_1721,N_1626,N_1617);
and U1722 (N_1722,N_1661,N_1691);
or U1723 (N_1723,N_1613,N_1625);
nor U1724 (N_1724,N_1622,N_1620);
and U1725 (N_1725,N_1694,N_1607);
and U1726 (N_1726,N_1643,N_1670);
and U1727 (N_1727,N_1677,N_1688);
or U1728 (N_1728,N_1645,N_1675);
xor U1729 (N_1729,N_1636,N_1635);
or U1730 (N_1730,N_1629,N_1634);
nand U1731 (N_1731,N_1627,N_1637);
nor U1732 (N_1732,N_1611,N_1621);
nand U1733 (N_1733,N_1604,N_1667);
nand U1734 (N_1734,N_1665,N_1679);
and U1735 (N_1735,N_1672,N_1686);
nor U1736 (N_1736,N_1608,N_1680);
xor U1737 (N_1737,N_1633,N_1632);
and U1738 (N_1738,N_1642,N_1678);
nand U1739 (N_1739,N_1609,N_1656);
nor U1740 (N_1740,N_1668,N_1660);
or U1741 (N_1741,N_1697,N_1671);
or U1742 (N_1742,N_1699,N_1659);
nor U1743 (N_1743,N_1640,N_1664);
nand U1744 (N_1744,N_1623,N_1690);
or U1745 (N_1745,N_1616,N_1650);
and U1746 (N_1746,N_1646,N_1695);
nor U1747 (N_1747,N_1685,N_1655);
and U1748 (N_1748,N_1644,N_1657);
nor U1749 (N_1749,N_1683,N_1682);
nand U1750 (N_1750,N_1630,N_1668);
or U1751 (N_1751,N_1661,N_1620);
or U1752 (N_1752,N_1653,N_1621);
nand U1753 (N_1753,N_1677,N_1694);
nor U1754 (N_1754,N_1639,N_1686);
xor U1755 (N_1755,N_1685,N_1634);
and U1756 (N_1756,N_1649,N_1609);
nor U1757 (N_1757,N_1612,N_1698);
and U1758 (N_1758,N_1644,N_1672);
and U1759 (N_1759,N_1635,N_1687);
or U1760 (N_1760,N_1691,N_1689);
or U1761 (N_1761,N_1662,N_1627);
nor U1762 (N_1762,N_1689,N_1693);
nor U1763 (N_1763,N_1698,N_1658);
nand U1764 (N_1764,N_1620,N_1680);
nor U1765 (N_1765,N_1625,N_1684);
and U1766 (N_1766,N_1609,N_1660);
or U1767 (N_1767,N_1664,N_1645);
and U1768 (N_1768,N_1663,N_1622);
nor U1769 (N_1769,N_1688,N_1699);
nor U1770 (N_1770,N_1659,N_1651);
and U1771 (N_1771,N_1603,N_1694);
and U1772 (N_1772,N_1658,N_1618);
and U1773 (N_1773,N_1653,N_1602);
nand U1774 (N_1774,N_1667,N_1658);
nor U1775 (N_1775,N_1683,N_1656);
nand U1776 (N_1776,N_1620,N_1668);
nand U1777 (N_1777,N_1608,N_1600);
or U1778 (N_1778,N_1646,N_1692);
and U1779 (N_1779,N_1614,N_1638);
or U1780 (N_1780,N_1687,N_1625);
nor U1781 (N_1781,N_1645,N_1635);
or U1782 (N_1782,N_1631,N_1665);
or U1783 (N_1783,N_1641,N_1638);
nor U1784 (N_1784,N_1687,N_1643);
and U1785 (N_1785,N_1631,N_1684);
nand U1786 (N_1786,N_1664,N_1661);
or U1787 (N_1787,N_1634,N_1619);
nor U1788 (N_1788,N_1634,N_1674);
or U1789 (N_1789,N_1665,N_1638);
or U1790 (N_1790,N_1656,N_1662);
nor U1791 (N_1791,N_1695,N_1669);
and U1792 (N_1792,N_1612,N_1613);
nand U1793 (N_1793,N_1689,N_1670);
xnor U1794 (N_1794,N_1639,N_1683);
or U1795 (N_1795,N_1631,N_1639);
nor U1796 (N_1796,N_1670,N_1671);
nand U1797 (N_1797,N_1620,N_1674);
or U1798 (N_1798,N_1677,N_1643);
nand U1799 (N_1799,N_1660,N_1617);
nor U1800 (N_1800,N_1759,N_1739);
and U1801 (N_1801,N_1729,N_1754);
xor U1802 (N_1802,N_1774,N_1716);
nand U1803 (N_1803,N_1728,N_1736);
or U1804 (N_1804,N_1789,N_1795);
and U1805 (N_1805,N_1794,N_1737);
or U1806 (N_1806,N_1787,N_1743);
nand U1807 (N_1807,N_1749,N_1724);
or U1808 (N_1808,N_1735,N_1700);
and U1809 (N_1809,N_1767,N_1725);
and U1810 (N_1810,N_1793,N_1712);
or U1811 (N_1811,N_1753,N_1779);
nand U1812 (N_1812,N_1764,N_1792);
nand U1813 (N_1813,N_1780,N_1721);
nor U1814 (N_1814,N_1732,N_1741);
nand U1815 (N_1815,N_1709,N_1762);
or U1816 (N_1816,N_1751,N_1782);
nor U1817 (N_1817,N_1788,N_1771);
or U1818 (N_1818,N_1748,N_1718);
xnor U1819 (N_1819,N_1702,N_1778);
or U1820 (N_1820,N_1776,N_1710);
nand U1821 (N_1821,N_1786,N_1744);
nand U1822 (N_1822,N_1731,N_1797);
and U1823 (N_1823,N_1756,N_1703);
nand U1824 (N_1824,N_1770,N_1706);
xnor U1825 (N_1825,N_1761,N_1752);
nand U1826 (N_1826,N_1798,N_1757);
nand U1827 (N_1827,N_1747,N_1708);
and U1828 (N_1828,N_1773,N_1701);
nand U1829 (N_1829,N_1730,N_1772);
and U1830 (N_1830,N_1766,N_1723);
nor U1831 (N_1831,N_1717,N_1765);
or U1832 (N_1832,N_1742,N_1745);
xnor U1833 (N_1833,N_1799,N_1705);
nand U1834 (N_1834,N_1740,N_1785);
nand U1835 (N_1835,N_1790,N_1768);
nand U1836 (N_1836,N_1760,N_1733);
and U1837 (N_1837,N_1715,N_1704);
nor U1838 (N_1838,N_1726,N_1727);
or U1839 (N_1839,N_1755,N_1738);
or U1840 (N_1840,N_1720,N_1783);
nand U1841 (N_1841,N_1746,N_1714);
nor U1842 (N_1842,N_1713,N_1784);
nand U1843 (N_1843,N_1796,N_1711);
nor U1844 (N_1844,N_1769,N_1734);
and U1845 (N_1845,N_1758,N_1707);
nand U1846 (N_1846,N_1781,N_1750);
nand U1847 (N_1847,N_1777,N_1719);
or U1848 (N_1848,N_1763,N_1722);
nor U1849 (N_1849,N_1775,N_1791);
nor U1850 (N_1850,N_1738,N_1734);
nor U1851 (N_1851,N_1754,N_1760);
or U1852 (N_1852,N_1755,N_1734);
or U1853 (N_1853,N_1788,N_1703);
nor U1854 (N_1854,N_1711,N_1786);
nor U1855 (N_1855,N_1747,N_1748);
or U1856 (N_1856,N_1760,N_1771);
nand U1857 (N_1857,N_1753,N_1740);
and U1858 (N_1858,N_1779,N_1792);
nand U1859 (N_1859,N_1748,N_1717);
nand U1860 (N_1860,N_1789,N_1796);
nor U1861 (N_1861,N_1747,N_1735);
nand U1862 (N_1862,N_1706,N_1746);
or U1863 (N_1863,N_1709,N_1720);
and U1864 (N_1864,N_1771,N_1747);
or U1865 (N_1865,N_1784,N_1775);
and U1866 (N_1866,N_1711,N_1751);
and U1867 (N_1867,N_1729,N_1719);
and U1868 (N_1868,N_1783,N_1794);
nand U1869 (N_1869,N_1767,N_1746);
nand U1870 (N_1870,N_1748,N_1783);
and U1871 (N_1871,N_1779,N_1749);
or U1872 (N_1872,N_1799,N_1731);
and U1873 (N_1873,N_1706,N_1785);
and U1874 (N_1874,N_1758,N_1751);
or U1875 (N_1875,N_1743,N_1709);
or U1876 (N_1876,N_1748,N_1792);
nor U1877 (N_1877,N_1714,N_1739);
and U1878 (N_1878,N_1700,N_1724);
nor U1879 (N_1879,N_1702,N_1706);
nand U1880 (N_1880,N_1715,N_1719);
nor U1881 (N_1881,N_1797,N_1767);
nor U1882 (N_1882,N_1715,N_1741);
nor U1883 (N_1883,N_1764,N_1785);
or U1884 (N_1884,N_1742,N_1757);
xnor U1885 (N_1885,N_1703,N_1708);
nand U1886 (N_1886,N_1748,N_1710);
or U1887 (N_1887,N_1705,N_1741);
and U1888 (N_1888,N_1708,N_1767);
and U1889 (N_1889,N_1754,N_1714);
or U1890 (N_1890,N_1760,N_1763);
nor U1891 (N_1891,N_1760,N_1716);
nand U1892 (N_1892,N_1795,N_1746);
or U1893 (N_1893,N_1796,N_1764);
and U1894 (N_1894,N_1730,N_1714);
nor U1895 (N_1895,N_1738,N_1767);
or U1896 (N_1896,N_1700,N_1758);
or U1897 (N_1897,N_1754,N_1704);
nand U1898 (N_1898,N_1778,N_1707);
or U1899 (N_1899,N_1792,N_1780);
and U1900 (N_1900,N_1808,N_1857);
nor U1901 (N_1901,N_1805,N_1844);
or U1902 (N_1902,N_1806,N_1887);
nor U1903 (N_1903,N_1847,N_1876);
nand U1904 (N_1904,N_1855,N_1836);
or U1905 (N_1905,N_1897,N_1851);
nand U1906 (N_1906,N_1818,N_1868);
nand U1907 (N_1907,N_1810,N_1819);
and U1908 (N_1908,N_1875,N_1895);
nor U1909 (N_1909,N_1801,N_1879);
or U1910 (N_1910,N_1811,N_1830);
nand U1911 (N_1911,N_1852,N_1842);
nor U1912 (N_1912,N_1816,N_1812);
or U1913 (N_1913,N_1892,N_1854);
and U1914 (N_1914,N_1845,N_1821);
nand U1915 (N_1915,N_1846,N_1856);
or U1916 (N_1916,N_1886,N_1804);
or U1917 (N_1917,N_1849,N_1825);
or U1918 (N_1918,N_1809,N_1807);
or U1919 (N_1919,N_1848,N_1888);
nor U1920 (N_1920,N_1822,N_1863);
nor U1921 (N_1921,N_1874,N_1889);
and U1922 (N_1922,N_1861,N_1814);
or U1923 (N_1923,N_1866,N_1803);
nor U1924 (N_1924,N_1834,N_1867);
nor U1925 (N_1925,N_1817,N_1864);
and U1926 (N_1926,N_1841,N_1877);
or U1927 (N_1927,N_1835,N_1898);
nand U1928 (N_1928,N_1865,N_1813);
nand U1929 (N_1929,N_1823,N_1832);
nand U1930 (N_1930,N_1884,N_1839);
or U1931 (N_1931,N_1827,N_1893);
or U1932 (N_1932,N_1891,N_1838);
and U1933 (N_1933,N_1890,N_1831);
or U1934 (N_1934,N_1862,N_1815);
nor U1935 (N_1935,N_1885,N_1882);
nand U1936 (N_1936,N_1881,N_1870);
nand U1937 (N_1937,N_1883,N_1802);
nand U1938 (N_1938,N_1833,N_1824);
or U1939 (N_1939,N_1828,N_1829);
nand U1940 (N_1940,N_1894,N_1820);
and U1941 (N_1941,N_1899,N_1878);
or U1942 (N_1942,N_1826,N_1880);
nor U1943 (N_1943,N_1800,N_1837);
or U1944 (N_1944,N_1869,N_1859);
nor U1945 (N_1945,N_1860,N_1872);
and U1946 (N_1946,N_1853,N_1858);
or U1947 (N_1947,N_1843,N_1896);
or U1948 (N_1948,N_1871,N_1850);
or U1949 (N_1949,N_1840,N_1873);
nand U1950 (N_1950,N_1872,N_1887);
and U1951 (N_1951,N_1815,N_1847);
nor U1952 (N_1952,N_1856,N_1805);
and U1953 (N_1953,N_1894,N_1828);
or U1954 (N_1954,N_1873,N_1821);
and U1955 (N_1955,N_1870,N_1821);
or U1956 (N_1956,N_1898,N_1863);
or U1957 (N_1957,N_1875,N_1811);
nor U1958 (N_1958,N_1828,N_1898);
nand U1959 (N_1959,N_1880,N_1800);
or U1960 (N_1960,N_1885,N_1806);
nor U1961 (N_1961,N_1811,N_1822);
and U1962 (N_1962,N_1871,N_1812);
and U1963 (N_1963,N_1862,N_1836);
or U1964 (N_1964,N_1889,N_1803);
or U1965 (N_1965,N_1813,N_1863);
or U1966 (N_1966,N_1895,N_1814);
or U1967 (N_1967,N_1897,N_1885);
and U1968 (N_1968,N_1890,N_1835);
xnor U1969 (N_1969,N_1880,N_1809);
nor U1970 (N_1970,N_1839,N_1883);
and U1971 (N_1971,N_1861,N_1848);
and U1972 (N_1972,N_1876,N_1857);
and U1973 (N_1973,N_1890,N_1876);
nor U1974 (N_1974,N_1822,N_1852);
or U1975 (N_1975,N_1816,N_1809);
nand U1976 (N_1976,N_1842,N_1894);
nand U1977 (N_1977,N_1843,N_1816);
or U1978 (N_1978,N_1803,N_1838);
or U1979 (N_1979,N_1886,N_1821);
or U1980 (N_1980,N_1801,N_1834);
nand U1981 (N_1981,N_1896,N_1827);
nor U1982 (N_1982,N_1893,N_1846);
and U1983 (N_1983,N_1853,N_1814);
nor U1984 (N_1984,N_1879,N_1804);
or U1985 (N_1985,N_1825,N_1842);
and U1986 (N_1986,N_1821,N_1832);
nand U1987 (N_1987,N_1831,N_1853);
or U1988 (N_1988,N_1800,N_1824);
nor U1989 (N_1989,N_1890,N_1880);
xor U1990 (N_1990,N_1809,N_1817);
and U1991 (N_1991,N_1823,N_1813);
nor U1992 (N_1992,N_1877,N_1830);
nor U1993 (N_1993,N_1872,N_1878);
nor U1994 (N_1994,N_1822,N_1854);
nor U1995 (N_1995,N_1802,N_1864);
nand U1996 (N_1996,N_1822,N_1877);
or U1997 (N_1997,N_1887,N_1839);
nor U1998 (N_1998,N_1875,N_1808);
or U1999 (N_1999,N_1883,N_1805);
nand U2000 (N_2000,N_1934,N_1988);
and U2001 (N_2001,N_1930,N_1979);
and U2002 (N_2002,N_1976,N_1998);
nor U2003 (N_2003,N_1995,N_1902);
nand U2004 (N_2004,N_1993,N_1955);
nor U2005 (N_2005,N_1969,N_1954);
nor U2006 (N_2006,N_1926,N_1981);
xor U2007 (N_2007,N_1933,N_1911);
or U2008 (N_2008,N_1980,N_1903);
nand U2009 (N_2009,N_1962,N_1935);
nor U2010 (N_2010,N_1917,N_1967);
or U2011 (N_2011,N_1974,N_1984);
nand U2012 (N_2012,N_1941,N_1948);
nand U2013 (N_2013,N_1959,N_1982);
and U2014 (N_2014,N_1960,N_1924);
or U2015 (N_2015,N_1910,N_1907);
nand U2016 (N_2016,N_1921,N_1949);
nand U2017 (N_2017,N_1920,N_1925);
nand U2018 (N_2018,N_1991,N_1950);
and U2019 (N_2019,N_1973,N_1970);
or U2020 (N_2020,N_1928,N_1940);
or U2021 (N_2021,N_1985,N_1947);
nand U2022 (N_2022,N_1905,N_1972);
nand U2023 (N_2023,N_1983,N_1963);
nor U2024 (N_2024,N_1964,N_1989);
and U2025 (N_2025,N_1965,N_1992);
nor U2026 (N_2026,N_1906,N_1929);
or U2027 (N_2027,N_1938,N_1999);
nand U2028 (N_2028,N_1997,N_1939);
nor U2029 (N_2029,N_1958,N_1919);
and U2030 (N_2030,N_1943,N_1957);
or U2031 (N_2031,N_1942,N_1912);
xor U2032 (N_2032,N_1901,N_1986);
nand U2033 (N_2033,N_1990,N_1944);
nor U2034 (N_2034,N_1968,N_1918);
nor U2035 (N_2035,N_1971,N_1946);
nor U2036 (N_2036,N_1916,N_1923);
nor U2037 (N_2037,N_1953,N_1951);
nor U2038 (N_2038,N_1961,N_1913);
nor U2039 (N_2039,N_1909,N_1996);
and U2040 (N_2040,N_1915,N_1977);
nand U2041 (N_2041,N_1956,N_1994);
nor U2042 (N_2042,N_1945,N_1978);
nand U2043 (N_2043,N_1900,N_1908);
and U2044 (N_2044,N_1931,N_1932);
or U2045 (N_2045,N_1936,N_1927);
nor U2046 (N_2046,N_1975,N_1937);
and U2047 (N_2047,N_1904,N_1987);
nor U2048 (N_2048,N_1966,N_1952);
nand U2049 (N_2049,N_1922,N_1914);
nor U2050 (N_2050,N_1954,N_1909);
and U2051 (N_2051,N_1919,N_1921);
nand U2052 (N_2052,N_1987,N_1984);
or U2053 (N_2053,N_1950,N_1973);
nor U2054 (N_2054,N_1946,N_1969);
and U2055 (N_2055,N_1923,N_1984);
or U2056 (N_2056,N_1989,N_1906);
nor U2057 (N_2057,N_1990,N_1993);
nor U2058 (N_2058,N_1922,N_1978);
nor U2059 (N_2059,N_1973,N_1938);
nand U2060 (N_2060,N_1970,N_1965);
and U2061 (N_2061,N_1946,N_1920);
and U2062 (N_2062,N_1984,N_1996);
or U2063 (N_2063,N_1957,N_1970);
nor U2064 (N_2064,N_1913,N_1978);
and U2065 (N_2065,N_1985,N_1990);
nor U2066 (N_2066,N_1936,N_1924);
xnor U2067 (N_2067,N_1951,N_1993);
or U2068 (N_2068,N_1926,N_1920);
or U2069 (N_2069,N_1972,N_1924);
and U2070 (N_2070,N_1952,N_1907);
and U2071 (N_2071,N_1945,N_1975);
or U2072 (N_2072,N_1980,N_1942);
nor U2073 (N_2073,N_1966,N_1920);
and U2074 (N_2074,N_1927,N_1965);
or U2075 (N_2075,N_1990,N_1901);
and U2076 (N_2076,N_1994,N_1925);
or U2077 (N_2077,N_1970,N_1966);
nand U2078 (N_2078,N_1907,N_1925);
nand U2079 (N_2079,N_1964,N_1978);
nand U2080 (N_2080,N_1958,N_1901);
or U2081 (N_2081,N_1983,N_1977);
nand U2082 (N_2082,N_1995,N_1900);
nor U2083 (N_2083,N_1912,N_1965);
nor U2084 (N_2084,N_1910,N_1936);
or U2085 (N_2085,N_1917,N_1971);
nor U2086 (N_2086,N_1956,N_1993);
and U2087 (N_2087,N_1968,N_1947);
and U2088 (N_2088,N_1934,N_1936);
and U2089 (N_2089,N_1956,N_1974);
nor U2090 (N_2090,N_1931,N_1915);
and U2091 (N_2091,N_1905,N_1929);
nor U2092 (N_2092,N_1939,N_1932);
or U2093 (N_2093,N_1933,N_1945);
nand U2094 (N_2094,N_1934,N_1924);
or U2095 (N_2095,N_1912,N_1918);
or U2096 (N_2096,N_1990,N_1946);
nand U2097 (N_2097,N_1927,N_1962);
and U2098 (N_2098,N_1950,N_1949);
nand U2099 (N_2099,N_1971,N_1975);
or U2100 (N_2100,N_2014,N_2025);
and U2101 (N_2101,N_2079,N_2055);
nand U2102 (N_2102,N_2081,N_2040);
nor U2103 (N_2103,N_2058,N_2007);
nand U2104 (N_2104,N_2041,N_2053);
nand U2105 (N_2105,N_2090,N_2066);
and U2106 (N_2106,N_2091,N_2011);
xnor U2107 (N_2107,N_2031,N_2000);
and U2108 (N_2108,N_2047,N_2003);
nor U2109 (N_2109,N_2051,N_2042);
or U2110 (N_2110,N_2088,N_2065);
or U2111 (N_2111,N_2052,N_2092);
and U2112 (N_2112,N_2071,N_2077);
or U2113 (N_2113,N_2069,N_2016);
nor U2114 (N_2114,N_2029,N_2057);
or U2115 (N_2115,N_2074,N_2084);
or U2116 (N_2116,N_2082,N_2044);
nand U2117 (N_2117,N_2061,N_2012);
nor U2118 (N_2118,N_2089,N_2018);
and U2119 (N_2119,N_2002,N_2085);
xor U2120 (N_2120,N_2070,N_2067);
or U2121 (N_2121,N_2022,N_2097);
or U2122 (N_2122,N_2036,N_2098);
or U2123 (N_2123,N_2063,N_2035);
or U2124 (N_2124,N_2075,N_2095);
or U2125 (N_2125,N_2083,N_2060);
and U2126 (N_2126,N_2059,N_2076);
nand U2127 (N_2127,N_2005,N_2064);
or U2128 (N_2128,N_2078,N_2050);
and U2129 (N_2129,N_2015,N_2054);
or U2130 (N_2130,N_2045,N_2038);
and U2131 (N_2131,N_2039,N_2032);
or U2132 (N_2132,N_2010,N_2046);
nor U2133 (N_2133,N_2087,N_2004);
nor U2134 (N_2134,N_2026,N_2006);
and U2135 (N_2135,N_2033,N_2030);
or U2136 (N_2136,N_2056,N_2001);
or U2137 (N_2137,N_2072,N_2099);
and U2138 (N_2138,N_2062,N_2093);
nand U2139 (N_2139,N_2023,N_2049);
nand U2140 (N_2140,N_2034,N_2027);
or U2141 (N_2141,N_2009,N_2024);
nor U2142 (N_2142,N_2021,N_2094);
and U2143 (N_2143,N_2028,N_2017);
nor U2144 (N_2144,N_2008,N_2096);
or U2145 (N_2145,N_2043,N_2080);
and U2146 (N_2146,N_2086,N_2020);
nand U2147 (N_2147,N_2037,N_2019);
or U2148 (N_2148,N_2048,N_2073);
or U2149 (N_2149,N_2013,N_2068);
or U2150 (N_2150,N_2095,N_2056);
and U2151 (N_2151,N_2021,N_2060);
nand U2152 (N_2152,N_2097,N_2020);
nor U2153 (N_2153,N_2058,N_2022);
nand U2154 (N_2154,N_2076,N_2034);
or U2155 (N_2155,N_2076,N_2040);
or U2156 (N_2156,N_2097,N_2007);
nand U2157 (N_2157,N_2030,N_2099);
and U2158 (N_2158,N_2055,N_2088);
and U2159 (N_2159,N_2059,N_2024);
or U2160 (N_2160,N_2016,N_2018);
and U2161 (N_2161,N_2000,N_2049);
or U2162 (N_2162,N_2050,N_2095);
nor U2163 (N_2163,N_2071,N_2058);
or U2164 (N_2164,N_2029,N_2021);
or U2165 (N_2165,N_2051,N_2065);
and U2166 (N_2166,N_2002,N_2054);
nor U2167 (N_2167,N_2011,N_2099);
nor U2168 (N_2168,N_2016,N_2097);
and U2169 (N_2169,N_2077,N_2021);
or U2170 (N_2170,N_2043,N_2002);
and U2171 (N_2171,N_2004,N_2073);
and U2172 (N_2172,N_2017,N_2057);
and U2173 (N_2173,N_2086,N_2058);
or U2174 (N_2174,N_2041,N_2001);
nor U2175 (N_2175,N_2099,N_2067);
nor U2176 (N_2176,N_2084,N_2067);
nor U2177 (N_2177,N_2059,N_2023);
nand U2178 (N_2178,N_2089,N_2038);
nor U2179 (N_2179,N_2097,N_2025);
and U2180 (N_2180,N_2059,N_2025);
and U2181 (N_2181,N_2084,N_2095);
nor U2182 (N_2182,N_2032,N_2070);
and U2183 (N_2183,N_2018,N_2081);
nor U2184 (N_2184,N_2050,N_2068);
nand U2185 (N_2185,N_2046,N_2054);
and U2186 (N_2186,N_2051,N_2059);
and U2187 (N_2187,N_2060,N_2032);
and U2188 (N_2188,N_2024,N_2001);
nand U2189 (N_2189,N_2016,N_2054);
nand U2190 (N_2190,N_2014,N_2076);
nand U2191 (N_2191,N_2002,N_2051);
and U2192 (N_2192,N_2084,N_2048);
and U2193 (N_2193,N_2056,N_2018);
nand U2194 (N_2194,N_2075,N_2070);
nor U2195 (N_2195,N_2020,N_2008);
and U2196 (N_2196,N_2089,N_2011);
nor U2197 (N_2197,N_2020,N_2048);
nor U2198 (N_2198,N_2061,N_2048);
and U2199 (N_2199,N_2069,N_2083);
nand U2200 (N_2200,N_2174,N_2180);
nand U2201 (N_2201,N_2149,N_2166);
nor U2202 (N_2202,N_2109,N_2185);
and U2203 (N_2203,N_2115,N_2116);
nor U2204 (N_2204,N_2191,N_2194);
nor U2205 (N_2205,N_2163,N_2175);
and U2206 (N_2206,N_2140,N_2179);
nand U2207 (N_2207,N_2154,N_2146);
or U2208 (N_2208,N_2165,N_2128);
nor U2209 (N_2209,N_2152,N_2170);
xor U2210 (N_2210,N_2169,N_2150);
and U2211 (N_2211,N_2196,N_2189);
nand U2212 (N_2212,N_2104,N_2178);
nand U2213 (N_2213,N_2122,N_2105);
or U2214 (N_2214,N_2133,N_2101);
nor U2215 (N_2215,N_2124,N_2148);
nand U2216 (N_2216,N_2142,N_2119);
and U2217 (N_2217,N_2144,N_2182);
nor U2218 (N_2218,N_2141,N_2187);
or U2219 (N_2219,N_2177,N_2172);
and U2220 (N_2220,N_2156,N_2193);
nand U2221 (N_2221,N_2186,N_2147);
and U2222 (N_2222,N_2120,N_2138);
nand U2223 (N_2223,N_2197,N_2168);
or U2224 (N_2224,N_2112,N_2143);
nor U2225 (N_2225,N_2151,N_2162);
and U2226 (N_2226,N_2167,N_2192);
nor U2227 (N_2227,N_2126,N_2130);
or U2228 (N_2228,N_2114,N_2164);
nor U2229 (N_2229,N_2155,N_2123);
nand U2230 (N_2230,N_2113,N_2139);
nor U2231 (N_2231,N_2190,N_2184);
nor U2232 (N_2232,N_2183,N_2136);
and U2233 (N_2233,N_2117,N_2102);
nand U2234 (N_2234,N_2176,N_2106);
nor U2235 (N_2235,N_2118,N_2131);
nor U2236 (N_2236,N_2129,N_2137);
nor U2237 (N_2237,N_2111,N_2121);
nand U2238 (N_2238,N_2160,N_2100);
nor U2239 (N_2239,N_2103,N_2199);
xnor U2240 (N_2240,N_2135,N_2159);
or U2241 (N_2241,N_2173,N_2158);
and U2242 (N_2242,N_2145,N_2157);
nand U2243 (N_2243,N_2195,N_2132);
nor U2244 (N_2244,N_2110,N_2127);
xnor U2245 (N_2245,N_2161,N_2198);
nor U2246 (N_2246,N_2125,N_2188);
nand U2247 (N_2247,N_2107,N_2108);
or U2248 (N_2248,N_2153,N_2171);
nand U2249 (N_2249,N_2134,N_2181);
nand U2250 (N_2250,N_2105,N_2189);
and U2251 (N_2251,N_2198,N_2191);
nor U2252 (N_2252,N_2172,N_2186);
and U2253 (N_2253,N_2175,N_2147);
or U2254 (N_2254,N_2198,N_2181);
nor U2255 (N_2255,N_2185,N_2194);
nand U2256 (N_2256,N_2151,N_2138);
nor U2257 (N_2257,N_2148,N_2168);
xnor U2258 (N_2258,N_2140,N_2198);
or U2259 (N_2259,N_2167,N_2121);
and U2260 (N_2260,N_2194,N_2108);
or U2261 (N_2261,N_2154,N_2161);
nor U2262 (N_2262,N_2190,N_2171);
and U2263 (N_2263,N_2155,N_2198);
nor U2264 (N_2264,N_2161,N_2132);
or U2265 (N_2265,N_2171,N_2130);
nand U2266 (N_2266,N_2185,N_2156);
or U2267 (N_2267,N_2160,N_2115);
and U2268 (N_2268,N_2152,N_2124);
nand U2269 (N_2269,N_2138,N_2110);
and U2270 (N_2270,N_2177,N_2113);
or U2271 (N_2271,N_2119,N_2143);
or U2272 (N_2272,N_2169,N_2107);
and U2273 (N_2273,N_2122,N_2126);
nor U2274 (N_2274,N_2145,N_2198);
nand U2275 (N_2275,N_2122,N_2112);
nor U2276 (N_2276,N_2109,N_2186);
nor U2277 (N_2277,N_2102,N_2119);
and U2278 (N_2278,N_2194,N_2142);
or U2279 (N_2279,N_2125,N_2150);
nor U2280 (N_2280,N_2120,N_2168);
nor U2281 (N_2281,N_2118,N_2146);
nand U2282 (N_2282,N_2101,N_2116);
nor U2283 (N_2283,N_2133,N_2102);
or U2284 (N_2284,N_2162,N_2172);
and U2285 (N_2285,N_2130,N_2198);
and U2286 (N_2286,N_2172,N_2102);
xnor U2287 (N_2287,N_2100,N_2112);
xnor U2288 (N_2288,N_2112,N_2117);
or U2289 (N_2289,N_2136,N_2194);
nor U2290 (N_2290,N_2115,N_2114);
or U2291 (N_2291,N_2178,N_2194);
nor U2292 (N_2292,N_2157,N_2183);
and U2293 (N_2293,N_2148,N_2190);
nor U2294 (N_2294,N_2152,N_2189);
and U2295 (N_2295,N_2150,N_2121);
and U2296 (N_2296,N_2162,N_2180);
nor U2297 (N_2297,N_2129,N_2127);
and U2298 (N_2298,N_2191,N_2193);
and U2299 (N_2299,N_2183,N_2147);
or U2300 (N_2300,N_2217,N_2245);
nor U2301 (N_2301,N_2284,N_2283);
or U2302 (N_2302,N_2263,N_2273);
and U2303 (N_2303,N_2293,N_2244);
or U2304 (N_2304,N_2221,N_2226);
nor U2305 (N_2305,N_2270,N_2216);
and U2306 (N_2306,N_2276,N_2213);
and U2307 (N_2307,N_2246,N_2242);
nor U2308 (N_2308,N_2297,N_2210);
and U2309 (N_2309,N_2208,N_2206);
and U2310 (N_2310,N_2259,N_2275);
or U2311 (N_2311,N_2218,N_2209);
nand U2312 (N_2312,N_2233,N_2268);
nand U2313 (N_2313,N_2261,N_2249);
nor U2314 (N_2314,N_2205,N_2203);
xnor U2315 (N_2315,N_2241,N_2232);
and U2316 (N_2316,N_2267,N_2282);
and U2317 (N_2317,N_2288,N_2201);
nor U2318 (N_2318,N_2262,N_2214);
nor U2319 (N_2319,N_2274,N_2234);
nand U2320 (N_2320,N_2231,N_2212);
and U2321 (N_2321,N_2230,N_2298);
nand U2322 (N_2322,N_2222,N_2252);
and U2323 (N_2323,N_2204,N_2223);
nand U2324 (N_2324,N_2251,N_2265);
and U2325 (N_2325,N_2280,N_2299);
or U2326 (N_2326,N_2240,N_2294);
or U2327 (N_2327,N_2224,N_2235);
xnor U2328 (N_2328,N_2290,N_2292);
nand U2329 (N_2329,N_2256,N_2287);
and U2330 (N_2330,N_2227,N_2281);
or U2331 (N_2331,N_2220,N_2207);
nand U2332 (N_2332,N_2247,N_2264);
nand U2333 (N_2333,N_2257,N_2271);
or U2334 (N_2334,N_2295,N_2200);
nor U2335 (N_2335,N_2279,N_2272);
and U2336 (N_2336,N_2266,N_2258);
nand U2337 (N_2337,N_2236,N_2243);
nor U2338 (N_2338,N_2229,N_2286);
nand U2339 (N_2339,N_2238,N_2219);
nor U2340 (N_2340,N_2250,N_2296);
nor U2341 (N_2341,N_2248,N_2291);
and U2342 (N_2342,N_2255,N_2225);
and U2343 (N_2343,N_2285,N_2278);
and U2344 (N_2344,N_2253,N_2237);
xor U2345 (N_2345,N_2289,N_2260);
nand U2346 (N_2346,N_2277,N_2215);
nor U2347 (N_2347,N_2239,N_2269);
and U2348 (N_2348,N_2228,N_2211);
nor U2349 (N_2349,N_2202,N_2254);
nor U2350 (N_2350,N_2270,N_2257);
and U2351 (N_2351,N_2261,N_2272);
nand U2352 (N_2352,N_2274,N_2230);
or U2353 (N_2353,N_2285,N_2290);
nor U2354 (N_2354,N_2295,N_2266);
nand U2355 (N_2355,N_2258,N_2298);
nand U2356 (N_2356,N_2267,N_2240);
nor U2357 (N_2357,N_2225,N_2264);
and U2358 (N_2358,N_2259,N_2217);
nand U2359 (N_2359,N_2243,N_2260);
nand U2360 (N_2360,N_2262,N_2296);
nand U2361 (N_2361,N_2224,N_2269);
nor U2362 (N_2362,N_2259,N_2204);
and U2363 (N_2363,N_2283,N_2201);
and U2364 (N_2364,N_2284,N_2233);
and U2365 (N_2365,N_2243,N_2253);
xor U2366 (N_2366,N_2289,N_2218);
xnor U2367 (N_2367,N_2231,N_2298);
and U2368 (N_2368,N_2279,N_2216);
nor U2369 (N_2369,N_2219,N_2204);
and U2370 (N_2370,N_2280,N_2233);
or U2371 (N_2371,N_2214,N_2203);
nand U2372 (N_2372,N_2227,N_2206);
nand U2373 (N_2373,N_2227,N_2298);
nand U2374 (N_2374,N_2208,N_2255);
and U2375 (N_2375,N_2211,N_2281);
or U2376 (N_2376,N_2283,N_2263);
and U2377 (N_2377,N_2276,N_2226);
nand U2378 (N_2378,N_2252,N_2277);
or U2379 (N_2379,N_2284,N_2216);
or U2380 (N_2380,N_2262,N_2291);
or U2381 (N_2381,N_2256,N_2297);
nor U2382 (N_2382,N_2216,N_2212);
nor U2383 (N_2383,N_2253,N_2263);
xor U2384 (N_2384,N_2256,N_2226);
xnor U2385 (N_2385,N_2262,N_2230);
nand U2386 (N_2386,N_2270,N_2252);
and U2387 (N_2387,N_2240,N_2247);
and U2388 (N_2388,N_2263,N_2203);
and U2389 (N_2389,N_2273,N_2201);
and U2390 (N_2390,N_2228,N_2249);
or U2391 (N_2391,N_2232,N_2264);
and U2392 (N_2392,N_2245,N_2253);
and U2393 (N_2393,N_2238,N_2277);
and U2394 (N_2394,N_2241,N_2278);
nand U2395 (N_2395,N_2220,N_2212);
xnor U2396 (N_2396,N_2231,N_2299);
nand U2397 (N_2397,N_2223,N_2253);
nor U2398 (N_2398,N_2215,N_2251);
xor U2399 (N_2399,N_2276,N_2271);
nand U2400 (N_2400,N_2308,N_2369);
or U2401 (N_2401,N_2338,N_2346);
nor U2402 (N_2402,N_2341,N_2335);
nand U2403 (N_2403,N_2358,N_2371);
nor U2404 (N_2404,N_2325,N_2359);
and U2405 (N_2405,N_2333,N_2382);
nor U2406 (N_2406,N_2378,N_2389);
or U2407 (N_2407,N_2303,N_2367);
nor U2408 (N_2408,N_2376,N_2336);
xnor U2409 (N_2409,N_2394,N_2344);
or U2410 (N_2410,N_2320,N_2321);
nor U2411 (N_2411,N_2391,N_2319);
or U2412 (N_2412,N_2315,N_2395);
nor U2413 (N_2413,N_2350,N_2360);
and U2414 (N_2414,N_2398,N_2313);
or U2415 (N_2415,N_2329,N_2381);
or U2416 (N_2416,N_2301,N_2396);
nor U2417 (N_2417,N_2397,N_2343);
nand U2418 (N_2418,N_2372,N_2383);
nor U2419 (N_2419,N_2388,N_2379);
or U2420 (N_2420,N_2323,N_2355);
nor U2421 (N_2421,N_2345,N_2361);
nor U2422 (N_2422,N_2331,N_2328);
nor U2423 (N_2423,N_2309,N_2370);
nand U2424 (N_2424,N_2374,N_2368);
and U2425 (N_2425,N_2304,N_2364);
and U2426 (N_2426,N_2332,N_2324);
nor U2427 (N_2427,N_2316,N_2390);
and U2428 (N_2428,N_2349,N_2392);
and U2429 (N_2429,N_2363,N_2305);
and U2430 (N_2430,N_2353,N_2330);
and U2431 (N_2431,N_2334,N_2311);
or U2432 (N_2432,N_2393,N_2377);
or U2433 (N_2433,N_2399,N_2386);
and U2434 (N_2434,N_2302,N_2342);
and U2435 (N_2435,N_2322,N_2375);
or U2436 (N_2436,N_2318,N_2380);
and U2437 (N_2437,N_2307,N_2312);
nor U2438 (N_2438,N_2366,N_2347);
and U2439 (N_2439,N_2365,N_2357);
nand U2440 (N_2440,N_2362,N_2351);
or U2441 (N_2441,N_2314,N_2300);
and U2442 (N_2442,N_2356,N_2354);
nand U2443 (N_2443,N_2337,N_2348);
nand U2444 (N_2444,N_2339,N_2310);
nand U2445 (N_2445,N_2326,N_2340);
or U2446 (N_2446,N_2384,N_2327);
nand U2447 (N_2447,N_2317,N_2385);
or U2448 (N_2448,N_2352,N_2306);
or U2449 (N_2449,N_2387,N_2373);
xor U2450 (N_2450,N_2340,N_2351);
nand U2451 (N_2451,N_2388,N_2342);
nand U2452 (N_2452,N_2394,N_2339);
nor U2453 (N_2453,N_2329,N_2378);
or U2454 (N_2454,N_2399,N_2327);
and U2455 (N_2455,N_2374,N_2359);
xor U2456 (N_2456,N_2319,N_2384);
or U2457 (N_2457,N_2357,N_2393);
nor U2458 (N_2458,N_2354,N_2304);
and U2459 (N_2459,N_2338,N_2370);
or U2460 (N_2460,N_2363,N_2378);
or U2461 (N_2461,N_2308,N_2306);
xnor U2462 (N_2462,N_2300,N_2353);
nor U2463 (N_2463,N_2331,N_2316);
nand U2464 (N_2464,N_2373,N_2300);
and U2465 (N_2465,N_2375,N_2341);
nor U2466 (N_2466,N_2371,N_2369);
and U2467 (N_2467,N_2303,N_2398);
nor U2468 (N_2468,N_2380,N_2377);
and U2469 (N_2469,N_2318,N_2345);
nor U2470 (N_2470,N_2370,N_2328);
nand U2471 (N_2471,N_2329,N_2312);
or U2472 (N_2472,N_2397,N_2312);
or U2473 (N_2473,N_2330,N_2377);
nor U2474 (N_2474,N_2373,N_2363);
nor U2475 (N_2475,N_2329,N_2314);
nand U2476 (N_2476,N_2358,N_2319);
nand U2477 (N_2477,N_2398,N_2385);
and U2478 (N_2478,N_2351,N_2390);
and U2479 (N_2479,N_2391,N_2367);
or U2480 (N_2480,N_2314,N_2390);
nand U2481 (N_2481,N_2311,N_2373);
or U2482 (N_2482,N_2388,N_2380);
nand U2483 (N_2483,N_2397,N_2395);
nor U2484 (N_2484,N_2366,N_2314);
nand U2485 (N_2485,N_2308,N_2398);
nor U2486 (N_2486,N_2329,N_2313);
nand U2487 (N_2487,N_2359,N_2321);
or U2488 (N_2488,N_2380,N_2363);
nor U2489 (N_2489,N_2387,N_2377);
or U2490 (N_2490,N_2304,N_2395);
nand U2491 (N_2491,N_2320,N_2356);
nor U2492 (N_2492,N_2392,N_2348);
nor U2493 (N_2493,N_2358,N_2309);
nand U2494 (N_2494,N_2387,N_2365);
nor U2495 (N_2495,N_2308,N_2395);
or U2496 (N_2496,N_2394,N_2333);
xor U2497 (N_2497,N_2395,N_2353);
nor U2498 (N_2498,N_2305,N_2349);
nor U2499 (N_2499,N_2366,N_2342);
nor U2500 (N_2500,N_2411,N_2499);
or U2501 (N_2501,N_2412,N_2492);
or U2502 (N_2502,N_2400,N_2402);
and U2503 (N_2503,N_2447,N_2488);
and U2504 (N_2504,N_2477,N_2448);
nor U2505 (N_2505,N_2493,N_2433);
or U2506 (N_2506,N_2443,N_2476);
and U2507 (N_2507,N_2482,N_2490);
nor U2508 (N_2508,N_2416,N_2481);
or U2509 (N_2509,N_2422,N_2409);
or U2510 (N_2510,N_2486,N_2419);
or U2511 (N_2511,N_2489,N_2496);
and U2512 (N_2512,N_2446,N_2436);
nor U2513 (N_2513,N_2473,N_2435);
nor U2514 (N_2514,N_2420,N_2410);
nand U2515 (N_2515,N_2415,N_2495);
nand U2516 (N_2516,N_2479,N_2406);
or U2517 (N_2517,N_2467,N_2472);
nand U2518 (N_2518,N_2439,N_2461);
or U2519 (N_2519,N_2465,N_2426);
nand U2520 (N_2520,N_2414,N_2483);
nor U2521 (N_2521,N_2418,N_2445);
nor U2522 (N_2522,N_2438,N_2404);
nand U2523 (N_2523,N_2442,N_2454);
nand U2524 (N_2524,N_2452,N_2408);
or U2525 (N_2525,N_2437,N_2475);
or U2526 (N_2526,N_2421,N_2471);
and U2527 (N_2527,N_2485,N_2462);
nand U2528 (N_2528,N_2413,N_2458);
and U2529 (N_2529,N_2453,N_2487);
nand U2530 (N_2530,N_2430,N_2460);
nor U2531 (N_2531,N_2450,N_2405);
or U2532 (N_2532,N_2470,N_2457);
or U2533 (N_2533,N_2449,N_2464);
nor U2534 (N_2534,N_2425,N_2440);
nor U2535 (N_2535,N_2459,N_2401);
nor U2536 (N_2536,N_2403,N_2494);
nand U2537 (N_2537,N_2456,N_2427);
nand U2538 (N_2538,N_2474,N_2431);
and U2539 (N_2539,N_2444,N_2480);
and U2540 (N_2540,N_2455,N_2424);
nand U2541 (N_2541,N_2469,N_2451);
nand U2542 (N_2542,N_2498,N_2429);
or U2543 (N_2543,N_2468,N_2466);
and U2544 (N_2544,N_2428,N_2463);
nand U2545 (N_2545,N_2407,N_2478);
xnor U2546 (N_2546,N_2491,N_2423);
nand U2547 (N_2547,N_2441,N_2484);
and U2548 (N_2548,N_2432,N_2417);
nand U2549 (N_2549,N_2434,N_2497);
xor U2550 (N_2550,N_2460,N_2467);
nor U2551 (N_2551,N_2469,N_2466);
nand U2552 (N_2552,N_2415,N_2434);
or U2553 (N_2553,N_2429,N_2424);
nor U2554 (N_2554,N_2401,N_2434);
nand U2555 (N_2555,N_2423,N_2426);
nor U2556 (N_2556,N_2435,N_2457);
or U2557 (N_2557,N_2439,N_2442);
xor U2558 (N_2558,N_2456,N_2463);
and U2559 (N_2559,N_2498,N_2408);
nor U2560 (N_2560,N_2410,N_2478);
nand U2561 (N_2561,N_2443,N_2440);
or U2562 (N_2562,N_2424,N_2467);
or U2563 (N_2563,N_2455,N_2493);
nor U2564 (N_2564,N_2465,N_2492);
nor U2565 (N_2565,N_2445,N_2433);
nor U2566 (N_2566,N_2418,N_2400);
nand U2567 (N_2567,N_2473,N_2474);
and U2568 (N_2568,N_2442,N_2452);
nor U2569 (N_2569,N_2441,N_2491);
nor U2570 (N_2570,N_2450,N_2415);
nand U2571 (N_2571,N_2455,N_2457);
or U2572 (N_2572,N_2414,N_2404);
nand U2573 (N_2573,N_2437,N_2482);
nor U2574 (N_2574,N_2423,N_2499);
nand U2575 (N_2575,N_2447,N_2413);
nand U2576 (N_2576,N_2486,N_2457);
nand U2577 (N_2577,N_2483,N_2487);
and U2578 (N_2578,N_2447,N_2486);
or U2579 (N_2579,N_2425,N_2415);
nand U2580 (N_2580,N_2410,N_2487);
nand U2581 (N_2581,N_2492,N_2424);
and U2582 (N_2582,N_2493,N_2445);
nor U2583 (N_2583,N_2498,N_2497);
nand U2584 (N_2584,N_2400,N_2472);
nor U2585 (N_2585,N_2439,N_2469);
nand U2586 (N_2586,N_2403,N_2419);
nor U2587 (N_2587,N_2469,N_2438);
and U2588 (N_2588,N_2442,N_2437);
nand U2589 (N_2589,N_2476,N_2419);
and U2590 (N_2590,N_2403,N_2410);
or U2591 (N_2591,N_2408,N_2434);
or U2592 (N_2592,N_2456,N_2458);
nor U2593 (N_2593,N_2459,N_2478);
nor U2594 (N_2594,N_2479,N_2442);
nor U2595 (N_2595,N_2461,N_2420);
or U2596 (N_2596,N_2480,N_2414);
or U2597 (N_2597,N_2429,N_2439);
and U2598 (N_2598,N_2498,N_2492);
and U2599 (N_2599,N_2464,N_2433);
and U2600 (N_2600,N_2549,N_2592);
and U2601 (N_2601,N_2551,N_2535);
xor U2602 (N_2602,N_2539,N_2519);
nand U2603 (N_2603,N_2580,N_2589);
or U2604 (N_2604,N_2513,N_2544);
nor U2605 (N_2605,N_2560,N_2538);
or U2606 (N_2606,N_2502,N_2555);
nand U2607 (N_2607,N_2565,N_2591);
and U2608 (N_2608,N_2588,N_2501);
and U2609 (N_2609,N_2561,N_2599);
or U2610 (N_2610,N_2563,N_2533);
and U2611 (N_2611,N_2597,N_2567);
and U2612 (N_2612,N_2527,N_2569);
or U2613 (N_2613,N_2552,N_2584);
or U2614 (N_2614,N_2521,N_2506);
nor U2615 (N_2615,N_2548,N_2558);
nand U2616 (N_2616,N_2523,N_2574);
and U2617 (N_2617,N_2570,N_2520);
and U2618 (N_2618,N_2590,N_2526);
nand U2619 (N_2619,N_2524,N_2556);
xor U2620 (N_2620,N_2509,N_2528);
nand U2621 (N_2621,N_2529,N_2582);
nand U2622 (N_2622,N_2553,N_2571);
nor U2623 (N_2623,N_2579,N_2568);
and U2624 (N_2624,N_2546,N_2508);
and U2625 (N_2625,N_2505,N_2596);
nand U2626 (N_2626,N_2598,N_2543);
nand U2627 (N_2627,N_2542,N_2550);
nand U2628 (N_2628,N_2566,N_2578);
nor U2629 (N_2629,N_2525,N_2587);
or U2630 (N_2630,N_2516,N_2573);
nand U2631 (N_2631,N_2500,N_2547);
nand U2632 (N_2632,N_2504,N_2557);
or U2633 (N_2633,N_2576,N_2522);
and U2634 (N_2634,N_2594,N_2536);
and U2635 (N_2635,N_2595,N_2559);
or U2636 (N_2636,N_2562,N_2583);
nand U2637 (N_2637,N_2537,N_2530);
and U2638 (N_2638,N_2503,N_2577);
or U2639 (N_2639,N_2515,N_2581);
and U2640 (N_2640,N_2531,N_2586);
and U2641 (N_2641,N_2545,N_2554);
or U2642 (N_2642,N_2517,N_2534);
nor U2643 (N_2643,N_2532,N_2512);
and U2644 (N_2644,N_2510,N_2564);
and U2645 (N_2645,N_2585,N_2572);
or U2646 (N_2646,N_2541,N_2511);
and U2647 (N_2647,N_2514,N_2518);
nor U2648 (N_2648,N_2593,N_2575);
nor U2649 (N_2649,N_2507,N_2540);
nor U2650 (N_2650,N_2575,N_2506);
nor U2651 (N_2651,N_2575,N_2567);
nand U2652 (N_2652,N_2528,N_2531);
nor U2653 (N_2653,N_2577,N_2545);
nand U2654 (N_2654,N_2507,N_2598);
xor U2655 (N_2655,N_2534,N_2591);
nor U2656 (N_2656,N_2502,N_2519);
xor U2657 (N_2657,N_2531,N_2502);
nand U2658 (N_2658,N_2569,N_2570);
nand U2659 (N_2659,N_2529,N_2508);
nor U2660 (N_2660,N_2523,N_2586);
nand U2661 (N_2661,N_2505,N_2511);
nand U2662 (N_2662,N_2549,N_2555);
nand U2663 (N_2663,N_2538,N_2508);
nand U2664 (N_2664,N_2591,N_2517);
nand U2665 (N_2665,N_2581,N_2571);
and U2666 (N_2666,N_2513,N_2591);
nand U2667 (N_2667,N_2513,N_2507);
nand U2668 (N_2668,N_2590,N_2539);
and U2669 (N_2669,N_2586,N_2597);
or U2670 (N_2670,N_2585,N_2554);
or U2671 (N_2671,N_2558,N_2581);
and U2672 (N_2672,N_2568,N_2500);
or U2673 (N_2673,N_2574,N_2569);
nor U2674 (N_2674,N_2506,N_2510);
and U2675 (N_2675,N_2523,N_2562);
xnor U2676 (N_2676,N_2541,N_2544);
or U2677 (N_2677,N_2556,N_2530);
nor U2678 (N_2678,N_2571,N_2519);
nor U2679 (N_2679,N_2535,N_2525);
and U2680 (N_2680,N_2533,N_2579);
nor U2681 (N_2681,N_2556,N_2550);
and U2682 (N_2682,N_2585,N_2573);
and U2683 (N_2683,N_2580,N_2552);
nor U2684 (N_2684,N_2546,N_2505);
and U2685 (N_2685,N_2562,N_2524);
nor U2686 (N_2686,N_2571,N_2580);
nand U2687 (N_2687,N_2519,N_2596);
xor U2688 (N_2688,N_2550,N_2575);
and U2689 (N_2689,N_2596,N_2567);
nand U2690 (N_2690,N_2548,N_2505);
and U2691 (N_2691,N_2552,N_2533);
or U2692 (N_2692,N_2515,N_2599);
and U2693 (N_2693,N_2587,N_2507);
or U2694 (N_2694,N_2569,N_2545);
and U2695 (N_2695,N_2537,N_2533);
and U2696 (N_2696,N_2500,N_2574);
nand U2697 (N_2697,N_2503,N_2562);
and U2698 (N_2698,N_2502,N_2529);
or U2699 (N_2699,N_2547,N_2506);
nand U2700 (N_2700,N_2678,N_2658);
nor U2701 (N_2701,N_2670,N_2676);
nor U2702 (N_2702,N_2677,N_2692);
nor U2703 (N_2703,N_2665,N_2602);
nor U2704 (N_2704,N_2610,N_2654);
or U2705 (N_2705,N_2668,N_2627);
and U2706 (N_2706,N_2637,N_2675);
and U2707 (N_2707,N_2685,N_2659);
xnor U2708 (N_2708,N_2674,N_2657);
nor U2709 (N_2709,N_2624,N_2672);
nand U2710 (N_2710,N_2614,N_2619);
and U2711 (N_2711,N_2691,N_2636);
or U2712 (N_2712,N_2641,N_2605);
nor U2713 (N_2713,N_2651,N_2673);
nand U2714 (N_2714,N_2604,N_2699);
or U2715 (N_2715,N_2679,N_2638);
and U2716 (N_2716,N_2615,N_2655);
and U2717 (N_2717,N_2649,N_2629);
and U2718 (N_2718,N_2687,N_2646);
or U2719 (N_2719,N_2648,N_2669);
nor U2720 (N_2720,N_2639,N_2623);
nand U2721 (N_2721,N_2695,N_2616);
or U2722 (N_2722,N_2671,N_2686);
nor U2723 (N_2723,N_2612,N_2681);
nand U2724 (N_2724,N_2644,N_2663);
nand U2725 (N_2725,N_2631,N_2664);
and U2726 (N_2726,N_2613,N_2633);
nand U2727 (N_2727,N_2652,N_2643);
xnor U2728 (N_2728,N_2688,N_2625);
or U2729 (N_2729,N_2683,N_2606);
nand U2730 (N_2730,N_2667,N_2660);
nor U2731 (N_2731,N_2608,N_2656);
nand U2732 (N_2732,N_2621,N_2642);
or U2733 (N_2733,N_2680,N_2647);
and U2734 (N_2734,N_2662,N_2607);
nor U2735 (N_2735,N_2626,N_2618);
nor U2736 (N_2736,N_2690,N_2611);
nand U2737 (N_2737,N_2696,N_2600);
nor U2738 (N_2738,N_2620,N_2628);
and U2739 (N_2739,N_2661,N_2697);
or U2740 (N_2740,N_2666,N_2694);
and U2741 (N_2741,N_2645,N_2653);
nand U2742 (N_2742,N_2622,N_2650);
nor U2743 (N_2743,N_2617,N_2630);
or U2744 (N_2744,N_2682,N_2640);
nand U2745 (N_2745,N_2689,N_2693);
and U2746 (N_2746,N_2609,N_2698);
and U2747 (N_2747,N_2603,N_2601);
nand U2748 (N_2748,N_2635,N_2632);
nand U2749 (N_2749,N_2634,N_2684);
nand U2750 (N_2750,N_2675,N_2606);
or U2751 (N_2751,N_2667,N_2676);
nor U2752 (N_2752,N_2699,N_2641);
or U2753 (N_2753,N_2637,N_2678);
or U2754 (N_2754,N_2650,N_2691);
or U2755 (N_2755,N_2610,N_2625);
and U2756 (N_2756,N_2641,N_2630);
and U2757 (N_2757,N_2681,N_2663);
nand U2758 (N_2758,N_2631,N_2673);
nand U2759 (N_2759,N_2607,N_2630);
or U2760 (N_2760,N_2617,N_2625);
and U2761 (N_2761,N_2622,N_2689);
nand U2762 (N_2762,N_2672,N_2627);
or U2763 (N_2763,N_2650,N_2633);
nor U2764 (N_2764,N_2682,N_2692);
and U2765 (N_2765,N_2677,N_2633);
nor U2766 (N_2766,N_2622,N_2696);
xor U2767 (N_2767,N_2637,N_2605);
and U2768 (N_2768,N_2662,N_2600);
nor U2769 (N_2769,N_2666,N_2685);
nor U2770 (N_2770,N_2647,N_2642);
xor U2771 (N_2771,N_2696,N_2676);
xor U2772 (N_2772,N_2605,N_2667);
nand U2773 (N_2773,N_2625,N_2619);
or U2774 (N_2774,N_2685,N_2665);
xor U2775 (N_2775,N_2663,N_2620);
and U2776 (N_2776,N_2650,N_2675);
nor U2777 (N_2777,N_2600,N_2684);
and U2778 (N_2778,N_2693,N_2641);
nand U2779 (N_2779,N_2603,N_2664);
or U2780 (N_2780,N_2679,N_2624);
or U2781 (N_2781,N_2620,N_2667);
nor U2782 (N_2782,N_2611,N_2677);
and U2783 (N_2783,N_2621,N_2618);
or U2784 (N_2784,N_2657,N_2660);
nor U2785 (N_2785,N_2657,N_2690);
nand U2786 (N_2786,N_2643,N_2626);
and U2787 (N_2787,N_2668,N_2684);
nand U2788 (N_2788,N_2659,N_2606);
or U2789 (N_2789,N_2608,N_2601);
nand U2790 (N_2790,N_2605,N_2674);
and U2791 (N_2791,N_2616,N_2625);
nand U2792 (N_2792,N_2635,N_2620);
nor U2793 (N_2793,N_2685,N_2660);
nand U2794 (N_2794,N_2625,N_2656);
nor U2795 (N_2795,N_2635,N_2690);
xnor U2796 (N_2796,N_2606,N_2667);
or U2797 (N_2797,N_2627,N_2638);
and U2798 (N_2798,N_2637,N_2600);
nand U2799 (N_2799,N_2611,N_2649);
and U2800 (N_2800,N_2745,N_2756);
or U2801 (N_2801,N_2719,N_2792);
nor U2802 (N_2802,N_2738,N_2771);
and U2803 (N_2803,N_2734,N_2723);
or U2804 (N_2804,N_2711,N_2799);
nor U2805 (N_2805,N_2741,N_2717);
or U2806 (N_2806,N_2758,N_2729);
nand U2807 (N_2807,N_2700,N_2753);
nand U2808 (N_2808,N_2733,N_2772);
or U2809 (N_2809,N_2722,N_2790);
and U2810 (N_2810,N_2794,N_2735);
nor U2811 (N_2811,N_2774,N_2730);
nand U2812 (N_2812,N_2778,N_2702);
nand U2813 (N_2813,N_2761,N_2750);
or U2814 (N_2814,N_2786,N_2707);
or U2815 (N_2815,N_2769,N_2773);
and U2816 (N_2816,N_2710,N_2787);
or U2817 (N_2817,N_2767,N_2713);
and U2818 (N_2818,N_2764,N_2725);
and U2819 (N_2819,N_2740,N_2744);
nor U2820 (N_2820,N_2765,N_2793);
nor U2821 (N_2821,N_2749,N_2739);
nand U2822 (N_2822,N_2766,N_2776);
and U2823 (N_2823,N_2720,N_2703);
nand U2824 (N_2824,N_2781,N_2770);
nand U2825 (N_2825,N_2726,N_2754);
and U2826 (N_2826,N_2718,N_2760);
and U2827 (N_2827,N_2712,N_2706);
nand U2828 (N_2828,N_2746,N_2732);
nor U2829 (N_2829,N_2791,N_2788);
nor U2830 (N_2830,N_2731,N_2796);
or U2831 (N_2831,N_2751,N_2709);
nor U2832 (N_2832,N_2701,N_2742);
or U2833 (N_2833,N_2779,N_2798);
nor U2834 (N_2834,N_2752,N_2763);
or U2835 (N_2835,N_2705,N_2789);
nand U2836 (N_2836,N_2775,N_2716);
or U2837 (N_2837,N_2708,N_2728);
or U2838 (N_2838,N_2777,N_2755);
nand U2839 (N_2839,N_2737,N_2736);
and U2840 (N_2840,N_2780,N_2768);
nor U2841 (N_2841,N_2762,N_2748);
and U2842 (N_2842,N_2724,N_2782);
and U2843 (N_2843,N_2721,N_2759);
nand U2844 (N_2844,N_2784,N_2785);
xor U2845 (N_2845,N_2795,N_2743);
nand U2846 (N_2846,N_2704,N_2783);
or U2847 (N_2847,N_2715,N_2747);
nand U2848 (N_2848,N_2714,N_2797);
or U2849 (N_2849,N_2727,N_2757);
nand U2850 (N_2850,N_2711,N_2742);
nand U2851 (N_2851,N_2717,N_2784);
or U2852 (N_2852,N_2786,N_2794);
nand U2853 (N_2853,N_2788,N_2771);
nor U2854 (N_2854,N_2719,N_2720);
nand U2855 (N_2855,N_2744,N_2783);
and U2856 (N_2856,N_2724,N_2757);
or U2857 (N_2857,N_2783,N_2721);
and U2858 (N_2858,N_2715,N_2780);
and U2859 (N_2859,N_2797,N_2743);
or U2860 (N_2860,N_2703,N_2796);
nand U2861 (N_2861,N_2751,N_2786);
xnor U2862 (N_2862,N_2713,N_2712);
nand U2863 (N_2863,N_2722,N_2739);
and U2864 (N_2864,N_2774,N_2734);
nand U2865 (N_2865,N_2797,N_2780);
nand U2866 (N_2866,N_2750,N_2713);
nand U2867 (N_2867,N_2730,N_2766);
and U2868 (N_2868,N_2712,N_2700);
nand U2869 (N_2869,N_2797,N_2769);
and U2870 (N_2870,N_2727,N_2717);
nand U2871 (N_2871,N_2758,N_2772);
nor U2872 (N_2872,N_2715,N_2756);
xor U2873 (N_2873,N_2705,N_2708);
or U2874 (N_2874,N_2709,N_2785);
and U2875 (N_2875,N_2773,N_2702);
nand U2876 (N_2876,N_2784,N_2740);
nand U2877 (N_2877,N_2761,N_2730);
and U2878 (N_2878,N_2782,N_2742);
nand U2879 (N_2879,N_2765,N_2772);
or U2880 (N_2880,N_2717,N_2716);
and U2881 (N_2881,N_2786,N_2746);
nor U2882 (N_2882,N_2774,N_2718);
nand U2883 (N_2883,N_2707,N_2723);
nor U2884 (N_2884,N_2779,N_2751);
nor U2885 (N_2885,N_2732,N_2730);
or U2886 (N_2886,N_2712,N_2755);
xor U2887 (N_2887,N_2722,N_2764);
nor U2888 (N_2888,N_2728,N_2709);
or U2889 (N_2889,N_2725,N_2742);
or U2890 (N_2890,N_2784,N_2739);
and U2891 (N_2891,N_2731,N_2754);
nand U2892 (N_2892,N_2715,N_2788);
or U2893 (N_2893,N_2777,N_2717);
or U2894 (N_2894,N_2766,N_2771);
nand U2895 (N_2895,N_2779,N_2709);
and U2896 (N_2896,N_2759,N_2772);
and U2897 (N_2897,N_2725,N_2755);
or U2898 (N_2898,N_2768,N_2709);
nor U2899 (N_2899,N_2701,N_2728);
or U2900 (N_2900,N_2825,N_2865);
or U2901 (N_2901,N_2886,N_2813);
nand U2902 (N_2902,N_2847,N_2842);
or U2903 (N_2903,N_2863,N_2840);
or U2904 (N_2904,N_2881,N_2826);
and U2905 (N_2905,N_2843,N_2801);
and U2906 (N_2906,N_2874,N_2853);
or U2907 (N_2907,N_2873,N_2832);
nor U2908 (N_2908,N_2878,N_2850);
or U2909 (N_2909,N_2810,N_2804);
nor U2910 (N_2910,N_2855,N_2802);
or U2911 (N_2911,N_2818,N_2864);
nand U2912 (N_2912,N_2882,N_2861);
nor U2913 (N_2913,N_2817,N_2837);
nor U2914 (N_2914,N_2869,N_2806);
nand U2915 (N_2915,N_2833,N_2834);
and U2916 (N_2916,N_2872,N_2859);
nor U2917 (N_2917,N_2815,N_2820);
nor U2918 (N_2918,N_2805,N_2896);
nor U2919 (N_2919,N_2808,N_2895);
and U2920 (N_2920,N_2821,N_2898);
or U2921 (N_2921,N_2862,N_2852);
or U2922 (N_2922,N_2858,N_2851);
or U2923 (N_2923,N_2884,N_2824);
nor U2924 (N_2924,N_2890,N_2835);
and U2925 (N_2925,N_2831,N_2827);
nor U2926 (N_2926,N_2887,N_2845);
and U2927 (N_2927,N_2854,N_2894);
nand U2928 (N_2928,N_2844,N_2899);
nand U2929 (N_2929,N_2841,N_2891);
and U2930 (N_2930,N_2889,N_2814);
or U2931 (N_2931,N_2877,N_2860);
nor U2932 (N_2932,N_2892,N_2867);
or U2933 (N_2933,N_2819,N_2897);
or U2934 (N_2934,N_2839,N_2846);
and U2935 (N_2935,N_2836,N_2811);
and U2936 (N_2936,N_2807,N_2879);
and U2937 (N_2937,N_2856,N_2857);
nor U2938 (N_2938,N_2883,N_2822);
nand U2939 (N_2939,N_2888,N_2800);
and U2940 (N_2940,N_2870,N_2816);
nor U2941 (N_2941,N_2809,N_2830);
nand U2942 (N_2942,N_2871,N_2823);
and U2943 (N_2943,N_2875,N_2803);
nor U2944 (N_2944,N_2849,N_2885);
or U2945 (N_2945,N_2812,N_2828);
or U2946 (N_2946,N_2829,N_2868);
nor U2947 (N_2947,N_2876,N_2866);
nand U2948 (N_2948,N_2880,N_2848);
xnor U2949 (N_2949,N_2838,N_2893);
and U2950 (N_2950,N_2822,N_2897);
nand U2951 (N_2951,N_2848,N_2852);
or U2952 (N_2952,N_2849,N_2895);
nand U2953 (N_2953,N_2819,N_2809);
or U2954 (N_2954,N_2874,N_2877);
or U2955 (N_2955,N_2896,N_2835);
nor U2956 (N_2956,N_2843,N_2810);
or U2957 (N_2957,N_2854,N_2888);
and U2958 (N_2958,N_2845,N_2899);
or U2959 (N_2959,N_2809,N_2812);
nand U2960 (N_2960,N_2894,N_2855);
nand U2961 (N_2961,N_2882,N_2832);
or U2962 (N_2962,N_2880,N_2882);
nor U2963 (N_2963,N_2881,N_2806);
nor U2964 (N_2964,N_2847,N_2811);
nand U2965 (N_2965,N_2822,N_2843);
nand U2966 (N_2966,N_2895,N_2801);
and U2967 (N_2967,N_2863,N_2882);
or U2968 (N_2968,N_2891,N_2826);
and U2969 (N_2969,N_2805,N_2898);
or U2970 (N_2970,N_2834,N_2800);
xor U2971 (N_2971,N_2844,N_2882);
or U2972 (N_2972,N_2838,N_2828);
nand U2973 (N_2973,N_2852,N_2804);
or U2974 (N_2974,N_2852,N_2892);
nand U2975 (N_2975,N_2899,N_2892);
and U2976 (N_2976,N_2866,N_2826);
and U2977 (N_2977,N_2887,N_2839);
and U2978 (N_2978,N_2830,N_2873);
or U2979 (N_2979,N_2851,N_2897);
xor U2980 (N_2980,N_2862,N_2802);
nor U2981 (N_2981,N_2824,N_2858);
and U2982 (N_2982,N_2804,N_2850);
nand U2983 (N_2983,N_2868,N_2846);
nor U2984 (N_2984,N_2892,N_2864);
and U2985 (N_2985,N_2874,N_2833);
nor U2986 (N_2986,N_2823,N_2856);
nor U2987 (N_2987,N_2892,N_2838);
and U2988 (N_2988,N_2839,N_2806);
or U2989 (N_2989,N_2816,N_2846);
or U2990 (N_2990,N_2835,N_2887);
and U2991 (N_2991,N_2807,N_2814);
or U2992 (N_2992,N_2801,N_2893);
nor U2993 (N_2993,N_2815,N_2866);
nor U2994 (N_2994,N_2801,N_2876);
and U2995 (N_2995,N_2804,N_2878);
nor U2996 (N_2996,N_2846,N_2823);
xnor U2997 (N_2997,N_2872,N_2835);
and U2998 (N_2998,N_2898,N_2806);
or U2999 (N_2999,N_2859,N_2860);
or UO_0 (O_0,N_2966,N_2924);
or UO_1 (O_1,N_2931,N_2920);
nor UO_2 (O_2,N_2955,N_2913);
and UO_3 (O_3,N_2927,N_2947);
nand UO_4 (O_4,N_2929,N_2923);
nor UO_5 (O_5,N_2901,N_2951);
nand UO_6 (O_6,N_2902,N_2928);
or UO_7 (O_7,N_2991,N_2919);
nand UO_8 (O_8,N_2941,N_2987);
nand UO_9 (O_9,N_2990,N_2940);
and UO_10 (O_10,N_2982,N_2962);
or UO_11 (O_11,N_2996,N_2969);
and UO_12 (O_12,N_2983,N_2944);
and UO_13 (O_13,N_2912,N_2945);
and UO_14 (O_14,N_2922,N_2998);
nor UO_15 (O_15,N_2921,N_2993);
or UO_16 (O_16,N_2988,N_2992);
or UO_17 (O_17,N_2915,N_2950);
nand UO_18 (O_18,N_2900,N_2925);
nand UO_19 (O_19,N_2999,N_2909);
or UO_20 (O_20,N_2984,N_2981);
nor UO_21 (O_21,N_2961,N_2978);
nor UO_22 (O_22,N_2973,N_2917);
and UO_23 (O_23,N_2953,N_2918);
xor UO_24 (O_24,N_2936,N_2938);
or UO_25 (O_25,N_2904,N_2935);
or UO_26 (O_26,N_2970,N_2934);
nor UO_27 (O_27,N_2952,N_2907);
and UO_28 (O_28,N_2972,N_2989);
and UO_29 (O_29,N_2963,N_2948);
nor UO_30 (O_30,N_2926,N_2905);
and UO_31 (O_31,N_2967,N_2911);
and UO_32 (O_32,N_2914,N_2997);
nor UO_33 (O_33,N_2986,N_2930);
or UO_34 (O_34,N_2943,N_2916);
and UO_35 (O_35,N_2965,N_2995);
and UO_36 (O_36,N_2939,N_2979);
nand UO_37 (O_37,N_2959,N_2949);
nor UO_38 (O_38,N_2977,N_2910);
nor UO_39 (O_39,N_2908,N_2960);
nand UO_40 (O_40,N_2964,N_2974);
and UO_41 (O_41,N_2975,N_2933);
nand UO_42 (O_42,N_2946,N_2932);
and UO_43 (O_43,N_2985,N_2971);
nor UO_44 (O_44,N_2903,N_2942);
or UO_45 (O_45,N_2954,N_2994);
nand UO_46 (O_46,N_2968,N_2957);
and UO_47 (O_47,N_2906,N_2958);
nand UO_48 (O_48,N_2976,N_2937);
nand UO_49 (O_49,N_2956,N_2980);
xor UO_50 (O_50,N_2951,N_2971);
and UO_51 (O_51,N_2926,N_2962);
nor UO_52 (O_52,N_2952,N_2972);
nor UO_53 (O_53,N_2982,N_2947);
nor UO_54 (O_54,N_2944,N_2961);
nor UO_55 (O_55,N_2925,N_2937);
nand UO_56 (O_56,N_2931,N_2953);
nor UO_57 (O_57,N_2947,N_2959);
or UO_58 (O_58,N_2994,N_2976);
and UO_59 (O_59,N_2941,N_2930);
nor UO_60 (O_60,N_2920,N_2983);
nor UO_61 (O_61,N_2963,N_2952);
or UO_62 (O_62,N_2911,N_2987);
nand UO_63 (O_63,N_2928,N_2995);
nor UO_64 (O_64,N_2922,N_2928);
nand UO_65 (O_65,N_2928,N_2934);
nand UO_66 (O_66,N_2981,N_2985);
and UO_67 (O_67,N_2933,N_2993);
nor UO_68 (O_68,N_2954,N_2937);
nand UO_69 (O_69,N_2933,N_2910);
and UO_70 (O_70,N_2948,N_2976);
or UO_71 (O_71,N_2950,N_2918);
nand UO_72 (O_72,N_2922,N_2990);
and UO_73 (O_73,N_2909,N_2926);
and UO_74 (O_74,N_2995,N_2985);
nor UO_75 (O_75,N_2946,N_2967);
and UO_76 (O_76,N_2994,N_2902);
and UO_77 (O_77,N_2943,N_2955);
or UO_78 (O_78,N_2955,N_2946);
and UO_79 (O_79,N_2979,N_2936);
nand UO_80 (O_80,N_2931,N_2924);
nand UO_81 (O_81,N_2924,N_2913);
and UO_82 (O_82,N_2986,N_2987);
nor UO_83 (O_83,N_2925,N_2942);
or UO_84 (O_84,N_2995,N_2975);
or UO_85 (O_85,N_2970,N_2906);
and UO_86 (O_86,N_2984,N_2952);
and UO_87 (O_87,N_2915,N_2946);
nand UO_88 (O_88,N_2913,N_2962);
nand UO_89 (O_89,N_2921,N_2939);
nor UO_90 (O_90,N_2901,N_2926);
or UO_91 (O_91,N_2978,N_2921);
or UO_92 (O_92,N_2932,N_2914);
nor UO_93 (O_93,N_2940,N_2965);
nand UO_94 (O_94,N_2903,N_2995);
and UO_95 (O_95,N_2980,N_2995);
nand UO_96 (O_96,N_2944,N_2933);
or UO_97 (O_97,N_2961,N_2959);
and UO_98 (O_98,N_2988,N_2907);
nor UO_99 (O_99,N_2982,N_2946);
and UO_100 (O_100,N_2994,N_2946);
and UO_101 (O_101,N_2926,N_2933);
nand UO_102 (O_102,N_2982,N_2936);
nor UO_103 (O_103,N_2917,N_2979);
and UO_104 (O_104,N_2957,N_2935);
nor UO_105 (O_105,N_2929,N_2933);
nand UO_106 (O_106,N_2907,N_2996);
or UO_107 (O_107,N_2976,N_2943);
nor UO_108 (O_108,N_2955,N_2981);
nand UO_109 (O_109,N_2939,N_2991);
and UO_110 (O_110,N_2986,N_2950);
nand UO_111 (O_111,N_2939,N_2961);
nor UO_112 (O_112,N_2949,N_2936);
and UO_113 (O_113,N_2999,N_2979);
nor UO_114 (O_114,N_2915,N_2942);
nor UO_115 (O_115,N_2937,N_2981);
and UO_116 (O_116,N_2968,N_2998);
and UO_117 (O_117,N_2932,N_2969);
nand UO_118 (O_118,N_2960,N_2957);
and UO_119 (O_119,N_2901,N_2985);
or UO_120 (O_120,N_2972,N_2980);
or UO_121 (O_121,N_2982,N_2952);
nor UO_122 (O_122,N_2942,N_2967);
nor UO_123 (O_123,N_2934,N_2993);
and UO_124 (O_124,N_2932,N_2905);
nor UO_125 (O_125,N_2910,N_2926);
and UO_126 (O_126,N_2950,N_2995);
nand UO_127 (O_127,N_2936,N_2975);
nor UO_128 (O_128,N_2974,N_2963);
and UO_129 (O_129,N_2943,N_2922);
or UO_130 (O_130,N_2952,N_2921);
and UO_131 (O_131,N_2966,N_2953);
or UO_132 (O_132,N_2930,N_2928);
or UO_133 (O_133,N_2943,N_2995);
nor UO_134 (O_134,N_2954,N_2972);
nor UO_135 (O_135,N_2913,N_2915);
nor UO_136 (O_136,N_2911,N_2936);
and UO_137 (O_137,N_2919,N_2980);
nand UO_138 (O_138,N_2927,N_2968);
and UO_139 (O_139,N_2913,N_2947);
and UO_140 (O_140,N_2961,N_2911);
nor UO_141 (O_141,N_2957,N_2900);
nor UO_142 (O_142,N_2935,N_2975);
nand UO_143 (O_143,N_2935,N_2927);
and UO_144 (O_144,N_2971,N_2994);
or UO_145 (O_145,N_2966,N_2960);
nor UO_146 (O_146,N_2929,N_2954);
and UO_147 (O_147,N_2930,N_2918);
nand UO_148 (O_148,N_2989,N_2932);
and UO_149 (O_149,N_2947,N_2967);
nand UO_150 (O_150,N_2953,N_2906);
nor UO_151 (O_151,N_2944,N_2997);
nand UO_152 (O_152,N_2983,N_2955);
and UO_153 (O_153,N_2992,N_2973);
nand UO_154 (O_154,N_2944,N_2919);
or UO_155 (O_155,N_2915,N_2987);
and UO_156 (O_156,N_2987,N_2960);
nand UO_157 (O_157,N_2959,N_2969);
nand UO_158 (O_158,N_2959,N_2928);
or UO_159 (O_159,N_2901,N_2918);
or UO_160 (O_160,N_2968,N_2993);
and UO_161 (O_161,N_2930,N_2900);
nand UO_162 (O_162,N_2940,N_2902);
or UO_163 (O_163,N_2960,N_2975);
and UO_164 (O_164,N_2937,N_2967);
nor UO_165 (O_165,N_2962,N_2957);
and UO_166 (O_166,N_2937,N_2968);
nor UO_167 (O_167,N_2978,N_2908);
nor UO_168 (O_168,N_2981,N_2966);
nor UO_169 (O_169,N_2961,N_2971);
or UO_170 (O_170,N_2974,N_2931);
or UO_171 (O_171,N_2989,N_2936);
or UO_172 (O_172,N_2997,N_2904);
nand UO_173 (O_173,N_2945,N_2999);
or UO_174 (O_174,N_2922,N_2941);
or UO_175 (O_175,N_2982,N_2920);
nand UO_176 (O_176,N_2913,N_2959);
and UO_177 (O_177,N_2975,N_2942);
xor UO_178 (O_178,N_2927,N_2900);
and UO_179 (O_179,N_2925,N_2927);
nand UO_180 (O_180,N_2927,N_2988);
nand UO_181 (O_181,N_2941,N_2932);
and UO_182 (O_182,N_2975,N_2957);
nand UO_183 (O_183,N_2979,N_2969);
nand UO_184 (O_184,N_2920,N_2995);
nand UO_185 (O_185,N_2993,N_2979);
nor UO_186 (O_186,N_2921,N_2987);
nor UO_187 (O_187,N_2917,N_2926);
nand UO_188 (O_188,N_2917,N_2988);
nand UO_189 (O_189,N_2901,N_2962);
nor UO_190 (O_190,N_2979,N_2992);
or UO_191 (O_191,N_2989,N_2939);
and UO_192 (O_192,N_2908,N_2976);
nand UO_193 (O_193,N_2936,N_2930);
nor UO_194 (O_194,N_2986,N_2988);
and UO_195 (O_195,N_2946,N_2936);
nor UO_196 (O_196,N_2979,N_2964);
and UO_197 (O_197,N_2994,N_2908);
nand UO_198 (O_198,N_2925,N_2938);
and UO_199 (O_199,N_2920,N_2942);
and UO_200 (O_200,N_2987,N_2966);
xnor UO_201 (O_201,N_2913,N_2960);
xnor UO_202 (O_202,N_2949,N_2973);
or UO_203 (O_203,N_2956,N_2920);
or UO_204 (O_204,N_2957,N_2944);
and UO_205 (O_205,N_2941,N_2953);
nand UO_206 (O_206,N_2918,N_2928);
nand UO_207 (O_207,N_2947,N_2938);
or UO_208 (O_208,N_2951,N_2946);
and UO_209 (O_209,N_2957,N_2961);
and UO_210 (O_210,N_2970,N_2904);
or UO_211 (O_211,N_2953,N_2920);
or UO_212 (O_212,N_2991,N_2926);
nand UO_213 (O_213,N_2941,N_2934);
and UO_214 (O_214,N_2990,N_2912);
and UO_215 (O_215,N_2915,N_2997);
or UO_216 (O_216,N_2941,N_2904);
nand UO_217 (O_217,N_2985,N_2912);
or UO_218 (O_218,N_2925,N_2926);
and UO_219 (O_219,N_2926,N_2936);
nor UO_220 (O_220,N_2981,N_2995);
and UO_221 (O_221,N_2957,N_2954);
or UO_222 (O_222,N_2951,N_2915);
nor UO_223 (O_223,N_2969,N_2918);
nand UO_224 (O_224,N_2972,N_2924);
xnor UO_225 (O_225,N_2903,N_2994);
nand UO_226 (O_226,N_2945,N_2985);
xnor UO_227 (O_227,N_2937,N_2972);
nor UO_228 (O_228,N_2950,N_2943);
nor UO_229 (O_229,N_2987,N_2919);
or UO_230 (O_230,N_2926,N_2996);
or UO_231 (O_231,N_2999,N_2946);
and UO_232 (O_232,N_2911,N_2998);
or UO_233 (O_233,N_2970,N_2930);
nor UO_234 (O_234,N_2974,N_2918);
nor UO_235 (O_235,N_2973,N_2953);
nor UO_236 (O_236,N_2978,N_2958);
or UO_237 (O_237,N_2949,N_2929);
nand UO_238 (O_238,N_2973,N_2920);
and UO_239 (O_239,N_2940,N_2995);
xnor UO_240 (O_240,N_2922,N_2999);
or UO_241 (O_241,N_2968,N_2942);
nor UO_242 (O_242,N_2913,N_2977);
or UO_243 (O_243,N_2923,N_2986);
nand UO_244 (O_244,N_2941,N_2935);
and UO_245 (O_245,N_2904,N_2931);
and UO_246 (O_246,N_2954,N_2906);
or UO_247 (O_247,N_2975,N_2977);
or UO_248 (O_248,N_2904,N_2974);
and UO_249 (O_249,N_2947,N_2908);
and UO_250 (O_250,N_2915,N_2995);
and UO_251 (O_251,N_2967,N_2972);
nand UO_252 (O_252,N_2985,N_2942);
and UO_253 (O_253,N_2957,N_2985);
nand UO_254 (O_254,N_2980,N_2952);
or UO_255 (O_255,N_2991,N_2920);
nor UO_256 (O_256,N_2949,N_2989);
nor UO_257 (O_257,N_2941,N_2916);
nand UO_258 (O_258,N_2944,N_2980);
nand UO_259 (O_259,N_2962,N_2977);
nand UO_260 (O_260,N_2907,N_2906);
nand UO_261 (O_261,N_2934,N_2931);
nand UO_262 (O_262,N_2988,N_2946);
or UO_263 (O_263,N_2969,N_2968);
or UO_264 (O_264,N_2964,N_2973);
nand UO_265 (O_265,N_2996,N_2956);
or UO_266 (O_266,N_2963,N_2904);
nor UO_267 (O_267,N_2996,N_2977);
nor UO_268 (O_268,N_2941,N_2919);
nor UO_269 (O_269,N_2973,N_2956);
and UO_270 (O_270,N_2934,N_2992);
nand UO_271 (O_271,N_2941,N_2997);
nor UO_272 (O_272,N_2938,N_2903);
nor UO_273 (O_273,N_2907,N_2962);
and UO_274 (O_274,N_2945,N_2964);
or UO_275 (O_275,N_2976,N_2987);
and UO_276 (O_276,N_2997,N_2948);
or UO_277 (O_277,N_2928,N_2941);
nor UO_278 (O_278,N_2925,N_2967);
nand UO_279 (O_279,N_2995,N_2929);
or UO_280 (O_280,N_2945,N_2996);
nor UO_281 (O_281,N_2909,N_2931);
nand UO_282 (O_282,N_2909,N_2919);
and UO_283 (O_283,N_2933,N_2997);
and UO_284 (O_284,N_2993,N_2998);
xnor UO_285 (O_285,N_2983,N_2963);
nand UO_286 (O_286,N_2933,N_2912);
nand UO_287 (O_287,N_2961,N_2942);
and UO_288 (O_288,N_2991,N_2990);
and UO_289 (O_289,N_2903,N_2973);
and UO_290 (O_290,N_2936,N_2992);
and UO_291 (O_291,N_2941,N_2983);
nor UO_292 (O_292,N_2965,N_2902);
nand UO_293 (O_293,N_2990,N_2913);
or UO_294 (O_294,N_2902,N_2947);
or UO_295 (O_295,N_2902,N_2910);
nor UO_296 (O_296,N_2985,N_2960);
nor UO_297 (O_297,N_2964,N_2972);
nor UO_298 (O_298,N_2967,N_2994);
and UO_299 (O_299,N_2957,N_2977);
or UO_300 (O_300,N_2998,N_2981);
nor UO_301 (O_301,N_2918,N_2959);
nand UO_302 (O_302,N_2989,N_2970);
or UO_303 (O_303,N_2913,N_2909);
nand UO_304 (O_304,N_2998,N_2990);
nand UO_305 (O_305,N_2910,N_2989);
and UO_306 (O_306,N_2953,N_2911);
nand UO_307 (O_307,N_2964,N_2932);
nand UO_308 (O_308,N_2969,N_2955);
or UO_309 (O_309,N_2944,N_2949);
xor UO_310 (O_310,N_2943,N_2992);
or UO_311 (O_311,N_2941,N_2931);
nand UO_312 (O_312,N_2905,N_2948);
or UO_313 (O_313,N_2942,N_2940);
nor UO_314 (O_314,N_2988,N_2976);
nand UO_315 (O_315,N_2927,N_2946);
or UO_316 (O_316,N_2992,N_2980);
nor UO_317 (O_317,N_2937,N_2987);
and UO_318 (O_318,N_2968,N_2994);
nor UO_319 (O_319,N_2957,N_2995);
or UO_320 (O_320,N_2990,N_2902);
or UO_321 (O_321,N_2981,N_2987);
or UO_322 (O_322,N_2976,N_2941);
and UO_323 (O_323,N_2952,N_2919);
and UO_324 (O_324,N_2933,N_2963);
nor UO_325 (O_325,N_2906,N_2979);
and UO_326 (O_326,N_2963,N_2999);
nor UO_327 (O_327,N_2906,N_2985);
and UO_328 (O_328,N_2989,N_2958);
and UO_329 (O_329,N_2933,N_2990);
or UO_330 (O_330,N_2969,N_2951);
or UO_331 (O_331,N_2961,N_2968);
or UO_332 (O_332,N_2954,N_2913);
xnor UO_333 (O_333,N_2904,N_2948);
or UO_334 (O_334,N_2935,N_2986);
and UO_335 (O_335,N_2995,N_2951);
nand UO_336 (O_336,N_2965,N_2963);
and UO_337 (O_337,N_2968,N_2956);
nor UO_338 (O_338,N_2921,N_2930);
nor UO_339 (O_339,N_2904,N_2933);
nor UO_340 (O_340,N_2964,N_2998);
nor UO_341 (O_341,N_2911,N_2994);
and UO_342 (O_342,N_2902,N_2971);
nand UO_343 (O_343,N_2946,N_2909);
nor UO_344 (O_344,N_2997,N_2928);
nor UO_345 (O_345,N_2952,N_2974);
nor UO_346 (O_346,N_2941,N_2967);
nor UO_347 (O_347,N_2990,N_2999);
and UO_348 (O_348,N_2951,N_2949);
and UO_349 (O_349,N_2972,N_2944);
nor UO_350 (O_350,N_2911,N_2973);
nor UO_351 (O_351,N_2958,N_2917);
and UO_352 (O_352,N_2955,N_2954);
or UO_353 (O_353,N_2968,N_2967);
and UO_354 (O_354,N_2925,N_2951);
or UO_355 (O_355,N_2923,N_2954);
or UO_356 (O_356,N_2914,N_2938);
nor UO_357 (O_357,N_2938,N_2916);
and UO_358 (O_358,N_2925,N_2963);
or UO_359 (O_359,N_2931,N_2959);
and UO_360 (O_360,N_2945,N_2965);
xnor UO_361 (O_361,N_2948,N_2973);
nand UO_362 (O_362,N_2984,N_2925);
xor UO_363 (O_363,N_2993,N_2996);
and UO_364 (O_364,N_2995,N_2926);
nand UO_365 (O_365,N_2905,N_2911);
nor UO_366 (O_366,N_2916,N_2978);
or UO_367 (O_367,N_2942,N_2929);
or UO_368 (O_368,N_2937,N_2906);
or UO_369 (O_369,N_2902,N_2942);
nand UO_370 (O_370,N_2914,N_2949);
or UO_371 (O_371,N_2947,N_2926);
nand UO_372 (O_372,N_2948,N_2969);
nand UO_373 (O_373,N_2983,N_2901);
and UO_374 (O_374,N_2925,N_2931);
nor UO_375 (O_375,N_2900,N_2993);
nand UO_376 (O_376,N_2988,N_2970);
nor UO_377 (O_377,N_2945,N_2933);
nand UO_378 (O_378,N_2961,N_2929);
and UO_379 (O_379,N_2934,N_2996);
and UO_380 (O_380,N_2954,N_2991);
nand UO_381 (O_381,N_2923,N_2906);
and UO_382 (O_382,N_2999,N_2912);
and UO_383 (O_383,N_2992,N_2993);
and UO_384 (O_384,N_2999,N_2917);
and UO_385 (O_385,N_2975,N_2925);
nand UO_386 (O_386,N_2933,N_2949);
or UO_387 (O_387,N_2969,N_2990);
and UO_388 (O_388,N_2942,N_2927);
or UO_389 (O_389,N_2938,N_2905);
nor UO_390 (O_390,N_2994,N_2900);
and UO_391 (O_391,N_2954,N_2918);
nor UO_392 (O_392,N_2912,N_2987);
nand UO_393 (O_393,N_2998,N_2924);
nor UO_394 (O_394,N_2996,N_2952);
or UO_395 (O_395,N_2978,N_2980);
nand UO_396 (O_396,N_2938,N_2962);
and UO_397 (O_397,N_2945,N_2917);
nor UO_398 (O_398,N_2966,N_2963);
nand UO_399 (O_399,N_2989,N_2971);
or UO_400 (O_400,N_2903,N_2960);
nor UO_401 (O_401,N_2928,N_2908);
and UO_402 (O_402,N_2980,N_2935);
nor UO_403 (O_403,N_2906,N_2999);
and UO_404 (O_404,N_2942,N_2979);
nor UO_405 (O_405,N_2949,N_2980);
nor UO_406 (O_406,N_2937,N_2910);
nor UO_407 (O_407,N_2997,N_2996);
or UO_408 (O_408,N_2948,N_2919);
or UO_409 (O_409,N_2945,N_2943);
nor UO_410 (O_410,N_2980,N_2959);
and UO_411 (O_411,N_2951,N_2937);
nor UO_412 (O_412,N_2938,N_2964);
nor UO_413 (O_413,N_2982,N_2979);
nor UO_414 (O_414,N_2946,N_2981);
and UO_415 (O_415,N_2938,N_2998);
nand UO_416 (O_416,N_2968,N_2933);
nand UO_417 (O_417,N_2914,N_2951);
nor UO_418 (O_418,N_2979,N_2911);
nor UO_419 (O_419,N_2983,N_2961);
or UO_420 (O_420,N_2928,N_2932);
nor UO_421 (O_421,N_2943,N_2989);
or UO_422 (O_422,N_2988,N_2996);
nand UO_423 (O_423,N_2957,N_2973);
nor UO_424 (O_424,N_2941,N_2956);
and UO_425 (O_425,N_2999,N_2934);
xnor UO_426 (O_426,N_2906,N_2911);
nand UO_427 (O_427,N_2904,N_2914);
nand UO_428 (O_428,N_2909,N_2952);
and UO_429 (O_429,N_2907,N_2961);
xnor UO_430 (O_430,N_2977,N_2955);
nand UO_431 (O_431,N_2934,N_2969);
nand UO_432 (O_432,N_2963,N_2926);
nand UO_433 (O_433,N_2949,N_2939);
nand UO_434 (O_434,N_2903,N_2975);
nand UO_435 (O_435,N_2928,N_2989);
nor UO_436 (O_436,N_2944,N_2992);
and UO_437 (O_437,N_2939,N_2988);
or UO_438 (O_438,N_2950,N_2971);
nand UO_439 (O_439,N_2909,N_2975);
nor UO_440 (O_440,N_2910,N_2982);
nor UO_441 (O_441,N_2909,N_2956);
nor UO_442 (O_442,N_2994,N_2934);
nand UO_443 (O_443,N_2970,N_2951);
nor UO_444 (O_444,N_2906,N_2996);
and UO_445 (O_445,N_2903,N_2962);
nand UO_446 (O_446,N_2925,N_2997);
and UO_447 (O_447,N_2989,N_2996);
and UO_448 (O_448,N_2999,N_2902);
nor UO_449 (O_449,N_2935,N_2996);
nor UO_450 (O_450,N_2952,N_2990);
and UO_451 (O_451,N_2975,N_2906);
and UO_452 (O_452,N_2984,N_2948);
or UO_453 (O_453,N_2958,N_2903);
nor UO_454 (O_454,N_2982,N_2992);
or UO_455 (O_455,N_2970,N_2944);
or UO_456 (O_456,N_2940,N_2906);
nor UO_457 (O_457,N_2995,N_2937);
nand UO_458 (O_458,N_2989,N_2911);
and UO_459 (O_459,N_2962,N_2908);
nand UO_460 (O_460,N_2989,N_2948);
or UO_461 (O_461,N_2926,N_2916);
or UO_462 (O_462,N_2933,N_2936);
nor UO_463 (O_463,N_2948,N_2910);
nand UO_464 (O_464,N_2912,N_2930);
and UO_465 (O_465,N_2982,N_2900);
or UO_466 (O_466,N_2959,N_2993);
nand UO_467 (O_467,N_2982,N_2934);
or UO_468 (O_468,N_2931,N_2975);
and UO_469 (O_469,N_2938,N_2966);
xnor UO_470 (O_470,N_2988,N_2960);
and UO_471 (O_471,N_2908,N_2970);
and UO_472 (O_472,N_2998,N_2991);
and UO_473 (O_473,N_2980,N_2991);
nor UO_474 (O_474,N_2949,N_2998);
nand UO_475 (O_475,N_2978,N_2914);
or UO_476 (O_476,N_2903,N_2935);
or UO_477 (O_477,N_2998,N_2941);
and UO_478 (O_478,N_2972,N_2966);
or UO_479 (O_479,N_2924,N_2938);
or UO_480 (O_480,N_2943,N_2981);
and UO_481 (O_481,N_2971,N_2953);
xnor UO_482 (O_482,N_2985,N_2910);
nand UO_483 (O_483,N_2968,N_2902);
nor UO_484 (O_484,N_2994,N_2925);
nand UO_485 (O_485,N_2993,N_2925);
and UO_486 (O_486,N_2918,N_2975);
and UO_487 (O_487,N_2914,N_2976);
nand UO_488 (O_488,N_2903,N_2909);
or UO_489 (O_489,N_2984,N_2999);
xnor UO_490 (O_490,N_2992,N_2955);
and UO_491 (O_491,N_2975,N_2989);
nand UO_492 (O_492,N_2976,N_2963);
nor UO_493 (O_493,N_2945,N_2991);
xor UO_494 (O_494,N_2945,N_2972);
nand UO_495 (O_495,N_2976,N_2906);
nand UO_496 (O_496,N_2946,N_2943);
nand UO_497 (O_497,N_2954,N_2921);
nor UO_498 (O_498,N_2943,N_2991);
nand UO_499 (O_499,N_2997,N_2985);
endmodule