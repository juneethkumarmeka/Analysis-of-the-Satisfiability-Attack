module basic_1000_10000_1500_5_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_74,In_496);
or U1 (N_1,In_517,In_82);
xor U2 (N_2,In_850,In_615);
and U3 (N_3,In_765,In_640);
nor U4 (N_4,In_446,In_706);
and U5 (N_5,In_494,In_536);
or U6 (N_6,In_318,In_397);
or U7 (N_7,In_844,In_443);
nand U8 (N_8,In_588,In_973);
nor U9 (N_9,In_945,In_981);
and U10 (N_10,In_840,In_559);
nor U11 (N_11,In_628,In_569);
nand U12 (N_12,In_238,In_266);
nor U13 (N_13,In_191,In_552);
and U14 (N_14,In_324,In_198);
and U15 (N_15,In_599,In_880);
nand U16 (N_16,In_763,In_235);
nor U17 (N_17,In_886,In_783);
nor U18 (N_18,In_375,In_951);
and U19 (N_19,In_79,In_121);
nor U20 (N_20,In_584,In_190);
or U21 (N_21,In_719,In_51);
or U22 (N_22,In_729,In_126);
or U23 (N_23,In_222,In_711);
nor U24 (N_24,In_727,In_777);
nor U25 (N_25,In_811,In_693);
nor U26 (N_26,In_644,In_671);
nor U27 (N_27,In_463,In_650);
and U28 (N_28,In_660,In_932);
and U29 (N_29,In_974,In_534);
and U30 (N_30,In_741,In_259);
or U31 (N_31,In_39,In_393);
nand U32 (N_32,In_349,In_515);
and U33 (N_33,In_771,In_999);
and U34 (N_34,In_456,In_164);
nand U35 (N_35,In_337,In_381);
nor U36 (N_36,In_824,In_89);
and U37 (N_37,In_917,In_80);
and U38 (N_38,In_27,In_817);
nor U39 (N_39,In_251,In_66);
nor U40 (N_40,In_41,In_600);
or U41 (N_41,In_208,In_395);
or U42 (N_42,In_949,In_321);
nor U43 (N_43,In_407,In_968);
and U44 (N_44,In_519,In_952);
or U45 (N_45,In_231,In_891);
nor U46 (N_46,In_866,In_295);
and U47 (N_47,In_62,In_530);
nand U48 (N_48,In_377,In_832);
or U49 (N_49,In_421,In_218);
nor U50 (N_50,In_331,In_400);
nand U51 (N_51,In_94,In_829);
nor U52 (N_52,In_963,In_885);
nand U53 (N_53,In_123,In_914);
nor U54 (N_54,In_948,In_790);
or U55 (N_55,In_367,In_453);
nor U56 (N_56,In_928,In_326);
and U57 (N_57,In_839,In_184);
and U58 (N_58,In_204,In_301);
nor U59 (N_59,In_735,In_428);
nand U60 (N_60,In_927,In_987);
or U61 (N_61,In_631,In_835);
xor U62 (N_62,In_618,In_846);
and U63 (N_63,In_293,In_21);
and U64 (N_64,In_842,In_937);
and U65 (N_65,In_838,In_700);
or U66 (N_66,In_214,In_554);
nand U67 (N_67,In_713,In_680);
or U68 (N_68,In_168,In_721);
nor U69 (N_69,In_853,In_95);
and U70 (N_70,In_77,In_905);
and U71 (N_71,In_84,In_360);
nor U72 (N_72,In_101,In_724);
or U73 (N_73,In_356,In_148);
nand U74 (N_74,In_57,In_419);
nand U75 (N_75,In_75,In_977);
nand U76 (N_76,In_647,In_431);
nand U77 (N_77,In_2,In_207);
or U78 (N_78,In_612,In_466);
or U79 (N_79,In_223,In_504);
and U80 (N_80,In_328,In_372);
and U81 (N_81,In_820,In_49);
or U82 (N_82,In_776,In_830);
nor U83 (N_83,In_117,In_452);
and U84 (N_84,In_394,In_998);
or U85 (N_85,In_209,In_910);
nor U86 (N_86,In_547,In_578);
and U87 (N_87,In_734,In_666);
or U88 (N_88,In_169,In_882);
nor U89 (N_89,In_594,In_151);
xnor U90 (N_90,In_247,In_900);
nand U91 (N_91,In_980,In_934);
nand U92 (N_92,In_874,In_961);
and U93 (N_93,In_658,In_971);
and U94 (N_94,In_8,In_71);
or U95 (N_95,In_587,In_665);
or U96 (N_96,In_877,In_156);
nand U97 (N_97,In_787,In_480);
and U98 (N_98,In_916,In_100);
or U99 (N_99,In_386,In_500);
nand U100 (N_100,In_43,In_864);
and U101 (N_101,In_33,In_601);
and U102 (N_102,In_709,In_592);
nor U103 (N_103,In_149,In_779);
and U104 (N_104,In_186,In_183);
nand U105 (N_105,In_956,In_361);
nand U106 (N_106,In_250,In_76);
or U107 (N_107,In_826,In_298);
and U108 (N_108,In_226,In_253);
or U109 (N_109,In_683,In_83);
nand U110 (N_110,In_457,In_307);
nor U111 (N_111,In_472,In_962);
nor U112 (N_112,In_580,In_823);
nand U113 (N_113,In_303,In_335);
or U114 (N_114,In_553,In_933);
or U115 (N_115,In_718,In_378);
or U116 (N_116,In_809,In_436);
or U117 (N_117,In_475,In_343);
or U118 (N_118,In_451,In_345);
nand U119 (N_119,In_525,In_764);
or U120 (N_120,In_920,In_55);
and U121 (N_121,In_696,In_740);
nand U122 (N_122,In_884,In_358);
nor U123 (N_123,In_330,In_205);
and U124 (N_124,In_791,In_966);
xor U125 (N_125,In_810,In_73);
or U126 (N_126,In_264,In_234);
or U127 (N_127,In_166,In_284);
nand U128 (N_128,In_701,In_54);
nand U129 (N_129,In_953,In_622);
nand U130 (N_130,In_571,In_526);
nor U131 (N_131,In_538,In_371);
nand U132 (N_132,In_181,In_221);
and U133 (N_133,In_570,In_36);
nand U134 (N_134,In_742,In_909);
nand U135 (N_135,In_300,In_179);
or U136 (N_136,In_678,In_363);
nand U137 (N_137,In_297,In_566);
xnor U138 (N_138,In_674,In_340);
or U139 (N_139,In_528,In_10);
and U140 (N_140,In_894,In_362);
nand U141 (N_141,In_629,In_778);
nand U142 (N_142,In_261,In_286);
nor U143 (N_143,In_40,In_522);
and U144 (N_144,In_178,In_61);
nand U145 (N_145,In_746,In_269);
and U146 (N_146,In_964,In_643);
nor U147 (N_147,In_762,In_210);
and U148 (N_148,In_280,In_401);
nand U149 (N_149,In_785,In_497);
nand U150 (N_150,In_403,In_883);
or U151 (N_151,In_415,In_505);
nor U152 (N_152,In_144,In_263);
nand U153 (N_153,In_37,In_573);
nand U154 (N_154,In_710,In_511);
and U155 (N_155,In_26,In_461);
and U156 (N_156,In_348,In_873);
nand U157 (N_157,In_69,In_754);
or U158 (N_158,In_814,In_414);
or U159 (N_159,In_444,In_723);
xnor U160 (N_160,In_143,In_512);
xnor U161 (N_161,In_901,In_849);
nand U162 (N_162,In_477,In_299);
nand U163 (N_163,In_613,In_341);
nor U164 (N_164,In_581,In_260);
xor U165 (N_165,In_589,In_115);
and U166 (N_166,In_922,In_568);
and U167 (N_167,In_879,In_120);
nand U168 (N_168,In_462,In_501);
xor U169 (N_169,In_564,In_675);
or U170 (N_170,In_116,In_273);
and U171 (N_171,In_926,In_244);
nand U172 (N_172,In_216,In_805);
or U173 (N_173,In_486,In_543);
nor U174 (N_174,In_138,In_249);
nor U175 (N_175,In_203,In_441);
or U176 (N_176,In_549,In_426);
nor U177 (N_177,In_510,In_382);
nand U178 (N_178,In_540,In_858);
nand U179 (N_179,In_969,In_294);
and U180 (N_180,In_45,In_482);
or U181 (N_181,In_656,In_445);
nor U182 (N_182,In_760,In_550);
nor U183 (N_183,In_11,In_370);
or U184 (N_184,In_459,In_781);
nand U185 (N_185,In_878,In_392);
or U186 (N_186,In_344,In_730);
and U187 (N_187,In_887,In_376);
or U188 (N_188,In_274,In_602);
nand U189 (N_189,In_744,In_911);
nor U190 (N_190,In_815,In_336);
xnor U191 (N_191,In_489,In_774);
or U192 (N_192,In_270,In_984);
nand U193 (N_193,In_645,In_87);
nand U194 (N_194,In_346,In_338);
or U195 (N_195,In_994,In_308);
nor U196 (N_196,In_197,In_989);
and U197 (N_197,In_368,In_576);
nand U198 (N_198,In_31,In_978);
and U199 (N_199,In_503,In_470);
and U200 (N_200,In_843,In_305);
nand U201 (N_201,In_315,In_256);
nand U202 (N_202,In_872,In_942);
and U203 (N_203,In_556,In_567);
nor U204 (N_204,In_857,In_114);
nor U205 (N_205,In_617,In_819);
or U206 (N_206,In_131,In_146);
nand U207 (N_207,In_365,In_689);
and U208 (N_208,In_159,In_703);
xnor U209 (N_209,In_194,In_185);
or U210 (N_210,In_474,In_807);
and U211 (N_211,In_786,In_309);
and U212 (N_212,In_670,In_232);
nor U213 (N_213,In_416,In_586);
or U214 (N_214,In_485,In_772);
nand U215 (N_215,In_769,In_35);
and U216 (N_216,In_246,In_107);
nand U217 (N_217,In_768,In_306);
or U218 (N_218,In_320,In_739);
nand U219 (N_219,In_682,In_919);
and U220 (N_220,In_423,In_420);
and U221 (N_221,In_852,In_720);
nor U222 (N_222,In_471,In_609);
nor U223 (N_223,In_48,In_292);
nor U224 (N_224,In_545,In_625);
xnor U225 (N_225,In_68,In_333);
nand U226 (N_226,In_875,In_685);
or U227 (N_227,In_982,In_946);
and U228 (N_228,In_304,In_582);
nor U229 (N_229,In_369,In_385);
nor U230 (N_230,In_859,In_947);
nand U231 (N_231,In_141,In_161);
nand U232 (N_232,In_175,In_498);
or U233 (N_233,In_507,In_440);
nor U234 (N_234,In_708,In_491);
nor U235 (N_235,In_354,In_590);
and U236 (N_236,In_533,In_20);
and U237 (N_237,In_229,In_792);
nand U238 (N_238,In_940,In_111);
and U239 (N_239,In_476,In_364);
and U240 (N_240,In_782,In_240);
nand U241 (N_241,In_108,In_521);
nor U242 (N_242,In_193,In_142);
and U243 (N_243,In_469,In_122);
nor U244 (N_244,In_285,In_473);
and U245 (N_245,In_862,In_788);
nand U246 (N_246,In_833,In_467);
nor U247 (N_247,In_103,In_213);
or U248 (N_248,In_755,In_661);
nor U249 (N_249,In_509,In_25);
nand U250 (N_250,In_158,In_139);
nor U251 (N_251,In_383,In_912);
or U252 (N_252,In_225,In_145);
and U253 (N_253,In_702,In_125);
nor U254 (N_254,In_109,In_520);
nor U255 (N_255,In_219,In_13);
nand U256 (N_256,In_483,In_130);
or U257 (N_257,In_325,In_624);
nand U258 (N_258,In_93,In_698);
or U259 (N_259,In_621,In_632);
nand U260 (N_260,In_944,In_47);
nand U261 (N_261,In_557,In_747);
nor U262 (N_262,In_611,In_282);
or U263 (N_263,In_64,In_635);
nand U264 (N_264,In_699,In_366);
and U265 (N_265,In_943,In_954);
and U266 (N_266,In_695,In_634);
or U267 (N_267,In_672,In_34);
nand U268 (N_268,In_268,In_535);
and U269 (N_269,In_63,In_892);
nand U270 (N_270,In_44,In_733);
nand U271 (N_271,In_737,In_265);
and U272 (N_272,In_479,In_639);
nor U273 (N_273,In_707,In_508);
nand U274 (N_274,In_90,In_432);
and U275 (N_275,In_437,In_118);
nand U276 (N_276,In_854,In_748);
or U277 (N_277,In_132,In_743);
nor U278 (N_278,In_384,In_638);
nor U279 (N_279,In_38,In_607);
nor U280 (N_280,In_930,In_716);
nand U281 (N_281,In_342,In_690);
and U282 (N_282,In_499,In_646);
nor U283 (N_283,In_88,In_583);
nand U284 (N_284,In_565,In_195);
nor U285 (N_285,In_58,In_825);
and U286 (N_286,In_429,In_784);
nor U287 (N_287,In_860,In_488);
nand U288 (N_288,In_373,In_279);
or U289 (N_289,In_939,In_449);
and U290 (N_290,In_12,In_187);
and U291 (N_291,In_399,In_626);
nand U292 (N_292,In_201,In_4);
or U293 (N_293,In_271,In_722);
and U294 (N_294,In_861,In_598);
nor U295 (N_295,In_30,In_418);
nor U296 (N_296,In_70,In_359);
nor U297 (N_297,In_59,In_135);
or U298 (N_298,In_527,In_424);
nand U299 (N_299,In_889,In_91);
or U300 (N_300,In_616,In_906);
nor U301 (N_301,In_233,In_697);
or U302 (N_302,In_379,In_561);
and U303 (N_303,In_562,In_996);
or U304 (N_304,In_908,In_97);
nand U305 (N_305,In_633,In_202);
and U306 (N_306,In_291,In_907);
and U307 (N_307,In_78,In_228);
nor U308 (N_308,In_258,In_694);
or U309 (N_309,In_523,In_923);
or U310 (N_310,In_623,In_18);
or U311 (N_311,In_657,In_925);
or U312 (N_312,In_112,In_975);
or U313 (N_313,In_514,In_728);
nor U314 (N_314,In_7,In_606);
nand U315 (N_315,In_837,In_119);
or U316 (N_316,In_649,In_990);
nor U317 (N_317,In_691,In_575);
nor U318 (N_318,In_24,In_319);
nor U319 (N_319,In_967,In_745);
and U320 (N_320,In_795,In_171);
or U321 (N_321,In_230,In_398);
nor U322 (N_322,In_841,In_972);
nand U323 (N_323,In_750,In_402);
nand U324 (N_324,In_808,In_460);
and U325 (N_325,In_705,In_935);
nand U326 (N_326,In_200,In_794);
or U327 (N_327,In_81,In_749);
or U328 (N_328,In_302,In_993);
and U329 (N_329,In_322,In_775);
or U330 (N_330,In_409,In_215);
nor U331 (N_331,In_224,In_995);
or U332 (N_332,In_313,In_127);
nor U333 (N_333,In_537,In_714);
nor U334 (N_334,In_16,In_150);
or U335 (N_335,In_664,In_813);
and U336 (N_336,In_597,In_140);
and U337 (N_337,In_174,In_417);
nor U338 (N_338,In_681,In_98);
and U339 (N_339,In_574,In_277);
and U340 (N_340,In_991,In_992);
xor U341 (N_341,In_405,In_104);
and U342 (N_342,In_532,In_72);
xor U343 (N_343,In_152,In_113);
or U344 (N_344,In_822,In_789);
nor U345 (N_345,In_541,In_668);
or U346 (N_346,In_856,In_248);
nand U347 (N_347,In_896,In_812);
nand U348 (N_348,In_481,In_314);
or U349 (N_349,In_903,In_913);
nor U350 (N_350,In_902,In_206);
or U351 (N_351,In_938,In_888);
and U352 (N_352,In_836,In_726);
nand U353 (N_353,In_281,In_28);
nor U354 (N_354,In_275,In_921);
nand U355 (N_355,In_834,In_351);
and U356 (N_356,In_797,In_220);
nand U357 (N_357,In_867,In_958);
nor U358 (N_358,In_334,In_546);
or U359 (N_359,In_404,In_352);
and U360 (N_360,In_177,In_761);
nor U361 (N_361,In_450,In_110);
nor U362 (N_362,In_237,In_603);
nor U363 (N_363,In_516,In_92);
nor U364 (N_364,In_767,In_374);
or U365 (N_365,In_847,In_757);
nand U366 (N_366,In_798,In_801);
and U367 (N_367,In_236,In_715);
nand U368 (N_368,In_593,In_329);
or U369 (N_369,In_257,In_23);
or U370 (N_370,In_136,In_42);
nor U371 (N_371,In_439,In_890);
or U372 (N_372,In_262,In_14);
and U373 (N_373,In_447,In_756);
or U374 (N_374,In_411,In_673);
or U375 (N_375,In_642,In_86);
and U376 (N_376,In_17,In_65);
nor U377 (N_377,In_732,In_390);
and U378 (N_378,In_278,In_272);
nor U379 (N_379,In_391,In_725);
nand U380 (N_380,In_929,In_15);
nand U381 (N_381,In_555,In_147);
nor U382 (N_382,In_712,In_848);
nor U383 (N_383,In_46,In_563);
or U384 (N_384,In_736,In_827);
and U385 (N_385,In_869,In_153);
or U386 (N_386,In_659,In_134);
or U387 (N_387,In_350,In_170);
and U388 (N_388,In_154,In_608);
or U389 (N_389,In_495,In_9);
nand U390 (N_390,In_851,In_493);
nor U391 (N_391,In_614,In_960);
or U392 (N_392,In_551,In_752);
or U393 (N_393,In_196,In_67);
nor U394 (N_394,In_396,In_806);
nand U395 (N_395,In_430,In_312);
and U396 (N_396,In_679,In_327);
nand U397 (N_397,In_243,In_893);
and U398 (N_398,In_669,In_448);
or U399 (N_399,In_529,In_636);
nor U400 (N_400,In_959,In_988);
and U401 (N_401,In_105,In_96);
nor U402 (N_402,In_317,In_871);
or U403 (N_403,In_753,In_19);
and U404 (N_404,In_408,In_276);
nand U405 (N_405,In_357,In_738);
nor U406 (N_406,In_957,In_759);
nor U407 (N_407,In_663,In_800);
nor U408 (N_408,In_986,In_435);
nand U409 (N_409,In_212,In_818);
and U410 (N_410,In_897,In_267);
or U411 (N_411,In_976,In_610);
nor U412 (N_412,In_189,In_124);
nor U413 (N_413,In_662,In_502);
xor U414 (N_414,In_845,In_455);
nand U415 (N_415,In_780,In_924);
nor U416 (N_416,In_157,In_56);
or U417 (N_417,In_667,In_311);
or U418 (N_418,In_163,In_487);
nand U419 (N_419,In_751,In_442);
nand U420 (N_420,In_137,In_687);
and U421 (N_421,In_283,In_241);
nor U422 (N_422,In_985,In_128);
and U423 (N_423,In_388,In_255);
nor U424 (N_424,In_353,In_686);
or U425 (N_425,In_160,In_637);
and U426 (N_426,In_918,In_60);
and U427 (N_427,In_427,In_355);
nand U428 (N_428,In_245,In_192);
or U429 (N_429,In_99,In_676);
nand U430 (N_430,In_677,In_412);
or U431 (N_431,In_796,In_85);
or U432 (N_432,In_413,In_870);
or U433 (N_433,In_5,In_425);
and U434 (N_434,In_524,In_310);
and U435 (N_435,In_895,In_188);
nand U436 (N_436,In_828,In_288);
nand U437 (N_437,In_692,In_438);
and U438 (N_438,In_865,In_287);
nand U439 (N_439,In_855,In_254);
nand U440 (N_440,In_799,In_955);
nand U441 (N_441,In_0,In_290);
or U442 (N_442,In_106,In_539);
or U443 (N_443,In_478,In_468);
or U444 (N_444,In_605,In_684);
nor U445 (N_445,In_899,In_717);
nand U446 (N_446,In_1,In_558);
nand U447 (N_447,In_931,In_513);
and U448 (N_448,In_387,In_591);
xnor U449 (N_449,In_518,In_465);
or U450 (N_450,In_490,In_560);
or U451 (N_451,In_252,In_688);
nor U452 (N_452,In_389,In_965);
nor U453 (N_453,In_876,In_803);
nand U454 (N_454,In_102,In_641);
nand U455 (N_455,In_332,In_29);
and U456 (N_456,In_804,In_542);
nand U457 (N_457,In_52,In_380);
nand U458 (N_458,In_211,In_410);
nand U459 (N_459,In_406,In_464);
and U460 (N_460,In_793,In_648);
nand U461 (N_461,In_651,In_199);
and U462 (N_462,In_572,In_347);
nand U463 (N_463,In_173,In_133);
nor U464 (N_464,In_619,In_296);
nand U465 (N_465,In_289,In_983);
or U466 (N_466,In_898,In_577);
nand U467 (N_467,In_531,In_458);
nand U468 (N_468,In_758,In_53);
nor U469 (N_469,In_773,In_585);
nor U470 (N_470,In_620,In_997);
nor U471 (N_471,In_596,In_816);
and U472 (N_472,In_323,In_162);
and U473 (N_473,In_492,In_484);
nor U474 (N_474,In_434,In_979);
or U475 (N_475,In_422,In_655);
and U476 (N_476,In_182,In_32);
or U477 (N_477,In_652,In_766);
or U478 (N_478,In_653,In_544);
nor U479 (N_479,In_654,In_604);
nand U480 (N_480,In_704,In_770);
nand U481 (N_481,In_881,In_506);
nand U482 (N_482,In_165,In_50);
or U483 (N_483,In_227,In_217);
or U484 (N_484,In_176,In_950);
and U485 (N_485,In_915,In_595);
and U486 (N_486,In_433,In_630);
nand U487 (N_487,In_941,In_339);
nor U488 (N_488,In_316,In_904);
nand U489 (N_489,In_129,In_802);
nor U490 (N_490,In_548,In_731);
nor U491 (N_491,In_180,In_579);
nor U492 (N_492,In_167,In_22);
and U493 (N_493,In_936,In_242);
nand U494 (N_494,In_863,In_970);
nand U495 (N_495,In_831,In_3);
and U496 (N_496,In_868,In_155);
nor U497 (N_497,In_821,In_239);
nand U498 (N_498,In_172,In_627);
nor U499 (N_499,In_454,In_6);
and U500 (N_500,In_425,In_216);
and U501 (N_501,In_448,In_365);
or U502 (N_502,In_319,In_242);
nand U503 (N_503,In_422,In_788);
nand U504 (N_504,In_239,In_624);
nor U505 (N_505,In_395,In_272);
nand U506 (N_506,In_769,In_841);
or U507 (N_507,In_254,In_629);
nand U508 (N_508,In_578,In_541);
and U509 (N_509,In_764,In_273);
and U510 (N_510,In_38,In_549);
nor U511 (N_511,In_497,In_452);
nor U512 (N_512,In_369,In_658);
nor U513 (N_513,In_435,In_69);
nor U514 (N_514,In_8,In_937);
nor U515 (N_515,In_499,In_630);
or U516 (N_516,In_17,In_275);
or U517 (N_517,In_342,In_200);
or U518 (N_518,In_861,In_755);
and U519 (N_519,In_41,In_834);
and U520 (N_520,In_233,In_525);
and U521 (N_521,In_45,In_189);
nand U522 (N_522,In_62,In_182);
nor U523 (N_523,In_150,In_775);
nor U524 (N_524,In_398,In_759);
or U525 (N_525,In_121,In_208);
nand U526 (N_526,In_940,In_693);
nor U527 (N_527,In_5,In_435);
nand U528 (N_528,In_86,In_628);
nand U529 (N_529,In_604,In_605);
and U530 (N_530,In_283,In_229);
or U531 (N_531,In_291,In_767);
nor U532 (N_532,In_536,In_607);
or U533 (N_533,In_282,In_913);
nand U534 (N_534,In_939,In_750);
or U535 (N_535,In_995,In_158);
or U536 (N_536,In_139,In_998);
nand U537 (N_537,In_329,In_197);
or U538 (N_538,In_652,In_268);
or U539 (N_539,In_831,In_374);
nand U540 (N_540,In_963,In_613);
nor U541 (N_541,In_16,In_564);
nor U542 (N_542,In_183,In_847);
and U543 (N_543,In_802,In_33);
xnor U544 (N_544,In_891,In_441);
and U545 (N_545,In_62,In_186);
nor U546 (N_546,In_146,In_759);
or U547 (N_547,In_972,In_640);
or U548 (N_548,In_801,In_943);
nor U549 (N_549,In_327,In_550);
nor U550 (N_550,In_281,In_662);
or U551 (N_551,In_342,In_499);
and U552 (N_552,In_293,In_149);
and U553 (N_553,In_53,In_870);
and U554 (N_554,In_602,In_1);
and U555 (N_555,In_937,In_553);
and U556 (N_556,In_309,In_622);
nand U557 (N_557,In_615,In_797);
nand U558 (N_558,In_92,In_508);
nand U559 (N_559,In_752,In_540);
nand U560 (N_560,In_329,In_458);
and U561 (N_561,In_991,In_143);
nand U562 (N_562,In_152,In_682);
nand U563 (N_563,In_753,In_875);
nor U564 (N_564,In_171,In_207);
and U565 (N_565,In_924,In_140);
and U566 (N_566,In_731,In_6);
nand U567 (N_567,In_954,In_933);
nor U568 (N_568,In_732,In_539);
and U569 (N_569,In_843,In_662);
or U570 (N_570,In_214,In_849);
nand U571 (N_571,In_211,In_672);
or U572 (N_572,In_104,In_392);
and U573 (N_573,In_907,In_839);
or U574 (N_574,In_813,In_89);
nor U575 (N_575,In_119,In_730);
or U576 (N_576,In_78,In_217);
nand U577 (N_577,In_145,In_318);
nor U578 (N_578,In_659,In_176);
xor U579 (N_579,In_315,In_560);
nand U580 (N_580,In_229,In_851);
nor U581 (N_581,In_442,In_471);
or U582 (N_582,In_446,In_0);
nor U583 (N_583,In_604,In_581);
nor U584 (N_584,In_673,In_62);
nand U585 (N_585,In_520,In_435);
nand U586 (N_586,In_594,In_853);
nor U587 (N_587,In_111,In_927);
nand U588 (N_588,In_484,In_661);
nor U589 (N_589,In_323,In_23);
nor U590 (N_590,In_983,In_213);
or U591 (N_591,In_644,In_264);
or U592 (N_592,In_932,In_28);
or U593 (N_593,In_781,In_397);
nand U594 (N_594,In_125,In_982);
nand U595 (N_595,In_255,In_139);
and U596 (N_596,In_866,In_456);
and U597 (N_597,In_611,In_95);
or U598 (N_598,In_368,In_714);
nor U599 (N_599,In_370,In_884);
and U600 (N_600,In_601,In_584);
nor U601 (N_601,In_104,In_935);
and U602 (N_602,In_830,In_433);
or U603 (N_603,In_734,In_911);
nand U604 (N_604,In_577,In_387);
nand U605 (N_605,In_603,In_309);
xor U606 (N_606,In_866,In_163);
nand U607 (N_607,In_878,In_214);
nor U608 (N_608,In_928,In_912);
nand U609 (N_609,In_286,In_131);
or U610 (N_610,In_471,In_246);
xor U611 (N_611,In_412,In_455);
and U612 (N_612,In_542,In_643);
nand U613 (N_613,In_807,In_145);
or U614 (N_614,In_404,In_177);
and U615 (N_615,In_485,In_208);
or U616 (N_616,In_450,In_91);
nor U617 (N_617,In_959,In_896);
nor U618 (N_618,In_559,In_529);
xnor U619 (N_619,In_646,In_536);
and U620 (N_620,In_537,In_110);
and U621 (N_621,In_212,In_924);
nor U622 (N_622,In_10,In_582);
nor U623 (N_623,In_689,In_967);
or U624 (N_624,In_777,In_130);
or U625 (N_625,In_137,In_717);
nand U626 (N_626,In_626,In_359);
or U627 (N_627,In_95,In_614);
xnor U628 (N_628,In_963,In_865);
nor U629 (N_629,In_798,In_459);
and U630 (N_630,In_719,In_935);
and U631 (N_631,In_327,In_500);
or U632 (N_632,In_312,In_657);
and U633 (N_633,In_953,In_517);
nand U634 (N_634,In_358,In_331);
or U635 (N_635,In_577,In_212);
nand U636 (N_636,In_685,In_498);
nand U637 (N_637,In_939,In_677);
or U638 (N_638,In_683,In_290);
and U639 (N_639,In_550,In_102);
nor U640 (N_640,In_597,In_357);
nand U641 (N_641,In_158,In_377);
and U642 (N_642,In_994,In_444);
and U643 (N_643,In_400,In_763);
or U644 (N_644,In_572,In_485);
nand U645 (N_645,In_635,In_795);
nand U646 (N_646,In_643,In_176);
or U647 (N_647,In_341,In_329);
and U648 (N_648,In_813,In_314);
nand U649 (N_649,In_751,In_622);
and U650 (N_650,In_329,In_821);
or U651 (N_651,In_496,In_170);
nand U652 (N_652,In_225,In_286);
nand U653 (N_653,In_39,In_943);
nand U654 (N_654,In_640,In_635);
or U655 (N_655,In_787,In_641);
or U656 (N_656,In_714,In_160);
and U657 (N_657,In_290,In_734);
nor U658 (N_658,In_4,In_593);
and U659 (N_659,In_871,In_604);
and U660 (N_660,In_168,In_522);
and U661 (N_661,In_291,In_562);
or U662 (N_662,In_846,In_687);
or U663 (N_663,In_87,In_764);
nand U664 (N_664,In_500,In_860);
or U665 (N_665,In_233,In_932);
and U666 (N_666,In_778,In_259);
and U667 (N_667,In_890,In_995);
and U668 (N_668,In_680,In_596);
or U669 (N_669,In_409,In_310);
and U670 (N_670,In_954,In_268);
xnor U671 (N_671,In_448,In_96);
or U672 (N_672,In_60,In_451);
nor U673 (N_673,In_82,In_316);
or U674 (N_674,In_672,In_485);
and U675 (N_675,In_960,In_709);
and U676 (N_676,In_688,In_40);
or U677 (N_677,In_476,In_103);
or U678 (N_678,In_525,In_88);
nand U679 (N_679,In_158,In_709);
nand U680 (N_680,In_800,In_281);
or U681 (N_681,In_444,In_955);
and U682 (N_682,In_226,In_967);
and U683 (N_683,In_649,In_747);
and U684 (N_684,In_985,In_438);
nand U685 (N_685,In_920,In_461);
nor U686 (N_686,In_20,In_112);
or U687 (N_687,In_613,In_87);
or U688 (N_688,In_510,In_871);
and U689 (N_689,In_578,In_953);
nor U690 (N_690,In_260,In_908);
or U691 (N_691,In_266,In_179);
or U692 (N_692,In_518,In_922);
and U693 (N_693,In_712,In_627);
nand U694 (N_694,In_852,In_696);
and U695 (N_695,In_689,In_449);
nand U696 (N_696,In_90,In_122);
and U697 (N_697,In_970,In_746);
nand U698 (N_698,In_940,In_573);
or U699 (N_699,In_217,In_931);
nand U700 (N_700,In_121,In_367);
and U701 (N_701,In_259,In_686);
nand U702 (N_702,In_771,In_973);
or U703 (N_703,In_850,In_739);
or U704 (N_704,In_509,In_894);
or U705 (N_705,In_763,In_857);
or U706 (N_706,In_832,In_141);
and U707 (N_707,In_437,In_244);
nor U708 (N_708,In_139,In_327);
xor U709 (N_709,In_675,In_500);
nor U710 (N_710,In_665,In_733);
and U711 (N_711,In_935,In_594);
or U712 (N_712,In_581,In_15);
or U713 (N_713,In_536,In_630);
and U714 (N_714,In_394,In_902);
or U715 (N_715,In_969,In_765);
nand U716 (N_716,In_621,In_149);
or U717 (N_717,In_608,In_558);
xor U718 (N_718,In_349,In_347);
nor U719 (N_719,In_680,In_436);
or U720 (N_720,In_395,In_270);
nand U721 (N_721,In_375,In_34);
nand U722 (N_722,In_338,In_164);
and U723 (N_723,In_704,In_503);
nor U724 (N_724,In_347,In_113);
nand U725 (N_725,In_952,In_951);
nor U726 (N_726,In_272,In_583);
or U727 (N_727,In_884,In_663);
or U728 (N_728,In_705,In_638);
nor U729 (N_729,In_991,In_190);
and U730 (N_730,In_557,In_52);
nor U731 (N_731,In_872,In_563);
or U732 (N_732,In_691,In_547);
and U733 (N_733,In_671,In_637);
nor U734 (N_734,In_870,In_313);
nand U735 (N_735,In_555,In_493);
and U736 (N_736,In_867,In_158);
or U737 (N_737,In_124,In_426);
or U738 (N_738,In_118,In_982);
and U739 (N_739,In_159,In_186);
nor U740 (N_740,In_979,In_155);
nand U741 (N_741,In_965,In_815);
and U742 (N_742,In_426,In_744);
nor U743 (N_743,In_828,In_204);
or U744 (N_744,In_639,In_0);
and U745 (N_745,In_310,In_707);
nand U746 (N_746,In_535,In_862);
nand U747 (N_747,In_473,In_271);
nand U748 (N_748,In_73,In_281);
nand U749 (N_749,In_452,In_866);
nor U750 (N_750,In_171,In_752);
nand U751 (N_751,In_427,In_610);
or U752 (N_752,In_184,In_408);
and U753 (N_753,In_925,In_280);
and U754 (N_754,In_342,In_91);
or U755 (N_755,In_980,In_336);
xnor U756 (N_756,In_894,In_936);
and U757 (N_757,In_480,In_177);
or U758 (N_758,In_643,In_108);
or U759 (N_759,In_508,In_104);
nor U760 (N_760,In_795,In_608);
nor U761 (N_761,In_154,In_732);
and U762 (N_762,In_593,In_766);
nand U763 (N_763,In_354,In_406);
and U764 (N_764,In_626,In_984);
and U765 (N_765,In_844,In_357);
nor U766 (N_766,In_893,In_450);
nand U767 (N_767,In_549,In_802);
and U768 (N_768,In_216,In_295);
xnor U769 (N_769,In_736,In_338);
and U770 (N_770,In_787,In_487);
nor U771 (N_771,In_89,In_202);
nor U772 (N_772,In_233,In_600);
nand U773 (N_773,In_1,In_887);
or U774 (N_774,In_617,In_893);
or U775 (N_775,In_29,In_168);
and U776 (N_776,In_102,In_904);
nor U777 (N_777,In_736,In_761);
xor U778 (N_778,In_463,In_201);
nand U779 (N_779,In_817,In_299);
or U780 (N_780,In_896,In_427);
nand U781 (N_781,In_686,In_666);
nor U782 (N_782,In_733,In_798);
nor U783 (N_783,In_520,In_157);
nor U784 (N_784,In_654,In_476);
or U785 (N_785,In_923,In_663);
and U786 (N_786,In_411,In_486);
nor U787 (N_787,In_175,In_56);
nor U788 (N_788,In_928,In_643);
nor U789 (N_789,In_645,In_294);
or U790 (N_790,In_629,In_324);
nor U791 (N_791,In_727,In_873);
nor U792 (N_792,In_495,In_284);
nand U793 (N_793,In_112,In_9);
and U794 (N_794,In_576,In_874);
and U795 (N_795,In_231,In_301);
nor U796 (N_796,In_15,In_775);
and U797 (N_797,In_969,In_130);
nand U798 (N_798,In_735,In_147);
nand U799 (N_799,In_886,In_933);
or U800 (N_800,In_254,In_736);
nand U801 (N_801,In_749,In_149);
or U802 (N_802,In_465,In_730);
nand U803 (N_803,In_272,In_27);
or U804 (N_804,In_822,In_508);
or U805 (N_805,In_627,In_722);
nand U806 (N_806,In_962,In_524);
and U807 (N_807,In_687,In_559);
nand U808 (N_808,In_904,In_828);
or U809 (N_809,In_521,In_634);
nand U810 (N_810,In_518,In_707);
or U811 (N_811,In_405,In_253);
or U812 (N_812,In_127,In_573);
and U813 (N_813,In_771,In_640);
nor U814 (N_814,In_850,In_601);
or U815 (N_815,In_40,In_904);
nor U816 (N_816,In_755,In_771);
nand U817 (N_817,In_81,In_382);
nor U818 (N_818,In_446,In_691);
or U819 (N_819,In_33,In_226);
nand U820 (N_820,In_299,In_260);
nand U821 (N_821,In_866,In_25);
or U822 (N_822,In_526,In_593);
xnor U823 (N_823,In_719,In_45);
nor U824 (N_824,In_829,In_726);
nor U825 (N_825,In_489,In_626);
and U826 (N_826,In_614,In_359);
nor U827 (N_827,In_870,In_435);
nand U828 (N_828,In_271,In_664);
nor U829 (N_829,In_786,In_680);
and U830 (N_830,In_172,In_89);
and U831 (N_831,In_752,In_840);
and U832 (N_832,In_859,In_278);
and U833 (N_833,In_29,In_353);
or U834 (N_834,In_773,In_59);
and U835 (N_835,In_828,In_451);
nor U836 (N_836,In_439,In_338);
nor U837 (N_837,In_958,In_966);
nor U838 (N_838,In_464,In_471);
and U839 (N_839,In_928,In_871);
or U840 (N_840,In_106,In_530);
and U841 (N_841,In_465,In_347);
nand U842 (N_842,In_83,In_134);
nor U843 (N_843,In_244,In_931);
and U844 (N_844,In_277,In_200);
nand U845 (N_845,In_444,In_206);
or U846 (N_846,In_941,In_917);
or U847 (N_847,In_945,In_69);
nand U848 (N_848,In_445,In_297);
or U849 (N_849,In_89,In_95);
or U850 (N_850,In_424,In_242);
or U851 (N_851,In_867,In_22);
nand U852 (N_852,In_150,In_474);
and U853 (N_853,In_531,In_252);
or U854 (N_854,In_791,In_279);
nand U855 (N_855,In_874,In_959);
or U856 (N_856,In_127,In_394);
nand U857 (N_857,In_802,In_918);
and U858 (N_858,In_637,In_977);
nor U859 (N_859,In_263,In_265);
nor U860 (N_860,In_234,In_467);
or U861 (N_861,In_291,In_475);
xor U862 (N_862,In_867,In_159);
or U863 (N_863,In_134,In_55);
nand U864 (N_864,In_857,In_276);
or U865 (N_865,In_42,In_966);
nor U866 (N_866,In_631,In_58);
nor U867 (N_867,In_602,In_959);
or U868 (N_868,In_784,In_773);
or U869 (N_869,In_123,In_378);
and U870 (N_870,In_232,In_420);
or U871 (N_871,In_248,In_878);
or U872 (N_872,In_187,In_36);
or U873 (N_873,In_265,In_31);
or U874 (N_874,In_889,In_134);
and U875 (N_875,In_312,In_760);
nand U876 (N_876,In_143,In_767);
or U877 (N_877,In_411,In_843);
and U878 (N_878,In_785,In_608);
xor U879 (N_879,In_457,In_222);
or U880 (N_880,In_293,In_516);
and U881 (N_881,In_840,In_261);
or U882 (N_882,In_587,In_797);
and U883 (N_883,In_944,In_63);
and U884 (N_884,In_612,In_220);
or U885 (N_885,In_180,In_388);
xnor U886 (N_886,In_197,In_190);
or U887 (N_887,In_28,In_637);
or U888 (N_888,In_352,In_851);
nand U889 (N_889,In_161,In_800);
or U890 (N_890,In_447,In_551);
or U891 (N_891,In_456,In_70);
xnor U892 (N_892,In_734,In_769);
and U893 (N_893,In_64,In_359);
nand U894 (N_894,In_545,In_382);
nand U895 (N_895,In_639,In_818);
nor U896 (N_896,In_924,In_696);
xor U897 (N_897,In_610,In_40);
nand U898 (N_898,In_27,In_25);
nor U899 (N_899,In_198,In_415);
nand U900 (N_900,In_948,In_305);
or U901 (N_901,In_383,In_505);
and U902 (N_902,In_783,In_90);
or U903 (N_903,In_250,In_358);
and U904 (N_904,In_910,In_444);
nand U905 (N_905,In_353,In_114);
nor U906 (N_906,In_1,In_515);
nand U907 (N_907,In_361,In_821);
nand U908 (N_908,In_931,In_679);
nand U909 (N_909,In_271,In_819);
nand U910 (N_910,In_399,In_312);
or U911 (N_911,In_850,In_516);
and U912 (N_912,In_318,In_112);
nand U913 (N_913,In_961,In_462);
nand U914 (N_914,In_343,In_518);
and U915 (N_915,In_847,In_288);
or U916 (N_916,In_137,In_133);
or U917 (N_917,In_737,In_994);
nor U918 (N_918,In_445,In_905);
or U919 (N_919,In_97,In_906);
or U920 (N_920,In_885,In_170);
nand U921 (N_921,In_813,In_920);
nand U922 (N_922,In_855,In_53);
and U923 (N_923,In_319,In_610);
or U924 (N_924,In_475,In_879);
nor U925 (N_925,In_491,In_153);
nand U926 (N_926,In_128,In_178);
nor U927 (N_927,In_998,In_153);
and U928 (N_928,In_89,In_833);
nor U929 (N_929,In_654,In_280);
and U930 (N_930,In_628,In_752);
nand U931 (N_931,In_999,In_544);
nor U932 (N_932,In_489,In_289);
and U933 (N_933,In_720,In_331);
and U934 (N_934,In_412,In_448);
nor U935 (N_935,In_54,In_563);
nor U936 (N_936,In_224,In_300);
nand U937 (N_937,In_97,In_739);
nor U938 (N_938,In_663,In_575);
nor U939 (N_939,In_907,In_178);
nor U940 (N_940,In_497,In_291);
nor U941 (N_941,In_442,In_492);
nor U942 (N_942,In_254,In_692);
xnor U943 (N_943,In_171,In_943);
nand U944 (N_944,In_164,In_295);
xnor U945 (N_945,In_224,In_71);
or U946 (N_946,In_114,In_537);
or U947 (N_947,In_467,In_599);
nor U948 (N_948,In_121,In_46);
and U949 (N_949,In_678,In_961);
and U950 (N_950,In_52,In_717);
nor U951 (N_951,In_889,In_629);
or U952 (N_952,In_455,In_723);
and U953 (N_953,In_773,In_673);
nand U954 (N_954,In_381,In_935);
and U955 (N_955,In_40,In_89);
nor U956 (N_956,In_13,In_841);
and U957 (N_957,In_207,In_401);
and U958 (N_958,In_369,In_124);
nor U959 (N_959,In_414,In_453);
nand U960 (N_960,In_669,In_446);
nand U961 (N_961,In_631,In_927);
nand U962 (N_962,In_678,In_258);
xor U963 (N_963,In_682,In_327);
nand U964 (N_964,In_686,In_476);
or U965 (N_965,In_973,In_360);
and U966 (N_966,In_937,In_249);
and U967 (N_967,In_271,In_948);
nor U968 (N_968,In_453,In_978);
nand U969 (N_969,In_876,In_407);
or U970 (N_970,In_25,In_826);
or U971 (N_971,In_434,In_905);
nor U972 (N_972,In_746,In_895);
and U973 (N_973,In_807,In_742);
and U974 (N_974,In_270,In_528);
and U975 (N_975,In_370,In_6);
or U976 (N_976,In_112,In_479);
nand U977 (N_977,In_314,In_216);
xnor U978 (N_978,In_640,In_85);
or U979 (N_979,In_126,In_327);
nor U980 (N_980,In_78,In_463);
or U981 (N_981,In_666,In_629);
nand U982 (N_982,In_497,In_468);
or U983 (N_983,In_785,In_777);
nor U984 (N_984,In_184,In_783);
nor U985 (N_985,In_27,In_503);
or U986 (N_986,In_158,In_337);
nand U987 (N_987,In_976,In_697);
or U988 (N_988,In_300,In_149);
nand U989 (N_989,In_159,In_191);
nor U990 (N_990,In_737,In_315);
or U991 (N_991,In_315,In_980);
nor U992 (N_992,In_513,In_505);
and U993 (N_993,In_791,In_784);
nand U994 (N_994,In_19,In_133);
and U995 (N_995,In_229,In_706);
nor U996 (N_996,In_916,In_323);
and U997 (N_997,In_533,In_957);
nor U998 (N_998,In_735,In_854);
nand U999 (N_999,In_762,In_67);
nor U1000 (N_1000,In_537,In_686);
or U1001 (N_1001,In_739,In_479);
xor U1002 (N_1002,In_65,In_802);
or U1003 (N_1003,In_535,In_964);
nor U1004 (N_1004,In_298,In_332);
or U1005 (N_1005,In_273,In_660);
nand U1006 (N_1006,In_503,In_952);
nor U1007 (N_1007,In_913,In_317);
or U1008 (N_1008,In_710,In_926);
nand U1009 (N_1009,In_627,In_589);
nand U1010 (N_1010,In_277,In_868);
and U1011 (N_1011,In_741,In_157);
nor U1012 (N_1012,In_577,In_923);
nor U1013 (N_1013,In_796,In_606);
and U1014 (N_1014,In_747,In_952);
and U1015 (N_1015,In_28,In_104);
nor U1016 (N_1016,In_554,In_88);
nand U1017 (N_1017,In_430,In_307);
or U1018 (N_1018,In_353,In_781);
and U1019 (N_1019,In_129,In_447);
and U1020 (N_1020,In_556,In_774);
nor U1021 (N_1021,In_304,In_90);
nand U1022 (N_1022,In_106,In_53);
or U1023 (N_1023,In_214,In_511);
or U1024 (N_1024,In_672,In_299);
or U1025 (N_1025,In_341,In_325);
nand U1026 (N_1026,In_640,In_87);
or U1027 (N_1027,In_174,In_651);
and U1028 (N_1028,In_310,In_29);
nand U1029 (N_1029,In_437,In_152);
nand U1030 (N_1030,In_839,In_87);
and U1031 (N_1031,In_958,In_830);
and U1032 (N_1032,In_486,In_669);
and U1033 (N_1033,In_786,In_287);
nor U1034 (N_1034,In_699,In_903);
or U1035 (N_1035,In_748,In_892);
xnor U1036 (N_1036,In_277,In_782);
nand U1037 (N_1037,In_996,In_69);
or U1038 (N_1038,In_530,In_359);
or U1039 (N_1039,In_768,In_244);
nand U1040 (N_1040,In_324,In_975);
nand U1041 (N_1041,In_157,In_29);
nand U1042 (N_1042,In_672,In_709);
and U1043 (N_1043,In_40,In_888);
and U1044 (N_1044,In_259,In_281);
or U1045 (N_1045,In_628,In_287);
or U1046 (N_1046,In_731,In_0);
nor U1047 (N_1047,In_852,In_342);
nor U1048 (N_1048,In_393,In_136);
and U1049 (N_1049,In_622,In_284);
and U1050 (N_1050,In_959,In_660);
or U1051 (N_1051,In_621,In_710);
or U1052 (N_1052,In_682,In_917);
nor U1053 (N_1053,In_282,In_804);
or U1054 (N_1054,In_428,In_438);
or U1055 (N_1055,In_368,In_30);
and U1056 (N_1056,In_115,In_911);
or U1057 (N_1057,In_113,In_643);
nand U1058 (N_1058,In_127,In_150);
and U1059 (N_1059,In_78,In_579);
nor U1060 (N_1060,In_364,In_867);
or U1061 (N_1061,In_877,In_147);
nor U1062 (N_1062,In_289,In_846);
nor U1063 (N_1063,In_90,In_569);
or U1064 (N_1064,In_303,In_339);
or U1065 (N_1065,In_953,In_749);
nor U1066 (N_1066,In_846,In_836);
or U1067 (N_1067,In_773,In_532);
nand U1068 (N_1068,In_112,In_91);
or U1069 (N_1069,In_282,In_344);
nor U1070 (N_1070,In_671,In_189);
and U1071 (N_1071,In_202,In_27);
xnor U1072 (N_1072,In_891,In_1);
and U1073 (N_1073,In_836,In_237);
and U1074 (N_1074,In_312,In_521);
nor U1075 (N_1075,In_321,In_809);
nor U1076 (N_1076,In_98,In_560);
nand U1077 (N_1077,In_555,In_838);
or U1078 (N_1078,In_445,In_9);
or U1079 (N_1079,In_769,In_951);
nand U1080 (N_1080,In_442,In_716);
nand U1081 (N_1081,In_763,In_669);
and U1082 (N_1082,In_410,In_198);
or U1083 (N_1083,In_567,In_592);
and U1084 (N_1084,In_662,In_371);
nor U1085 (N_1085,In_81,In_794);
and U1086 (N_1086,In_939,In_156);
nor U1087 (N_1087,In_881,In_989);
or U1088 (N_1088,In_948,In_312);
and U1089 (N_1089,In_498,In_296);
or U1090 (N_1090,In_909,In_280);
nand U1091 (N_1091,In_770,In_284);
nand U1092 (N_1092,In_917,In_755);
nor U1093 (N_1093,In_477,In_807);
nor U1094 (N_1094,In_459,In_47);
or U1095 (N_1095,In_283,In_676);
or U1096 (N_1096,In_166,In_56);
nand U1097 (N_1097,In_935,In_979);
and U1098 (N_1098,In_869,In_491);
or U1099 (N_1099,In_616,In_940);
nand U1100 (N_1100,In_740,In_692);
nand U1101 (N_1101,In_828,In_55);
xor U1102 (N_1102,In_401,In_287);
and U1103 (N_1103,In_374,In_492);
xor U1104 (N_1104,In_15,In_626);
xor U1105 (N_1105,In_325,In_732);
nand U1106 (N_1106,In_262,In_275);
and U1107 (N_1107,In_207,In_829);
and U1108 (N_1108,In_391,In_564);
nor U1109 (N_1109,In_762,In_626);
or U1110 (N_1110,In_113,In_323);
nand U1111 (N_1111,In_69,In_858);
nor U1112 (N_1112,In_978,In_424);
and U1113 (N_1113,In_477,In_539);
and U1114 (N_1114,In_274,In_515);
or U1115 (N_1115,In_607,In_333);
and U1116 (N_1116,In_480,In_977);
nor U1117 (N_1117,In_967,In_780);
or U1118 (N_1118,In_367,In_137);
nand U1119 (N_1119,In_557,In_752);
nor U1120 (N_1120,In_622,In_536);
and U1121 (N_1121,In_339,In_911);
or U1122 (N_1122,In_804,In_553);
and U1123 (N_1123,In_778,In_411);
or U1124 (N_1124,In_974,In_524);
xor U1125 (N_1125,In_321,In_730);
or U1126 (N_1126,In_800,In_594);
or U1127 (N_1127,In_534,In_592);
nor U1128 (N_1128,In_328,In_58);
nand U1129 (N_1129,In_357,In_533);
nor U1130 (N_1130,In_528,In_462);
nand U1131 (N_1131,In_630,In_893);
nor U1132 (N_1132,In_947,In_612);
nor U1133 (N_1133,In_430,In_184);
nor U1134 (N_1134,In_408,In_16);
and U1135 (N_1135,In_379,In_972);
nor U1136 (N_1136,In_621,In_103);
nor U1137 (N_1137,In_660,In_365);
or U1138 (N_1138,In_282,In_365);
nor U1139 (N_1139,In_713,In_681);
nand U1140 (N_1140,In_161,In_71);
nand U1141 (N_1141,In_302,In_442);
or U1142 (N_1142,In_219,In_294);
nor U1143 (N_1143,In_809,In_68);
nand U1144 (N_1144,In_910,In_321);
nand U1145 (N_1145,In_799,In_447);
nor U1146 (N_1146,In_136,In_760);
nand U1147 (N_1147,In_211,In_735);
nor U1148 (N_1148,In_478,In_959);
nand U1149 (N_1149,In_68,In_742);
or U1150 (N_1150,In_934,In_399);
or U1151 (N_1151,In_634,In_901);
nor U1152 (N_1152,In_416,In_785);
nor U1153 (N_1153,In_935,In_121);
or U1154 (N_1154,In_817,In_693);
nand U1155 (N_1155,In_19,In_891);
nand U1156 (N_1156,In_995,In_775);
and U1157 (N_1157,In_609,In_394);
nand U1158 (N_1158,In_932,In_495);
or U1159 (N_1159,In_751,In_223);
nor U1160 (N_1160,In_250,In_314);
nand U1161 (N_1161,In_959,In_72);
or U1162 (N_1162,In_979,In_563);
nor U1163 (N_1163,In_501,In_372);
nand U1164 (N_1164,In_500,In_598);
nor U1165 (N_1165,In_901,In_109);
nor U1166 (N_1166,In_950,In_89);
and U1167 (N_1167,In_782,In_53);
and U1168 (N_1168,In_581,In_580);
and U1169 (N_1169,In_26,In_457);
or U1170 (N_1170,In_199,In_614);
and U1171 (N_1171,In_78,In_153);
and U1172 (N_1172,In_470,In_851);
and U1173 (N_1173,In_57,In_704);
nand U1174 (N_1174,In_964,In_303);
and U1175 (N_1175,In_97,In_554);
or U1176 (N_1176,In_345,In_820);
and U1177 (N_1177,In_328,In_148);
and U1178 (N_1178,In_636,In_182);
and U1179 (N_1179,In_409,In_206);
and U1180 (N_1180,In_731,In_411);
nor U1181 (N_1181,In_228,In_991);
nand U1182 (N_1182,In_315,In_454);
xor U1183 (N_1183,In_158,In_594);
nor U1184 (N_1184,In_895,In_614);
and U1185 (N_1185,In_85,In_604);
nand U1186 (N_1186,In_192,In_148);
nor U1187 (N_1187,In_183,In_903);
or U1188 (N_1188,In_710,In_144);
and U1189 (N_1189,In_901,In_842);
nand U1190 (N_1190,In_784,In_249);
nand U1191 (N_1191,In_350,In_318);
and U1192 (N_1192,In_322,In_931);
or U1193 (N_1193,In_905,In_918);
nor U1194 (N_1194,In_656,In_505);
nand U1195 (N_1195,In_543,In_430);
or U1196 (N_1196,In_843,In_701);
and U1197 (N_1197,In_774,In_997);
and U1198 (N_1198,In_758,In_583);
nor U1199 (N_1199,In_316,In_400);
and U1200 (N_1200,In_786,In_462);
nand U1201 (N_1201,In_742,In_551);
and U1202 (N_1202,In_732,In_277);
or U1203 (N_1203,In_708,In_813);
nor U1204 (N_1204,In_12,In_689);
or U1205 (N_1205,In_248,In_83);
nand U1206 (N_1206,In_656,In_327);
and U1207 (N_1207,In_558,In_948);
nor U1208 (N_1208,In_962,In_206);
or U1209 (N_1209,In_716,In_360);
nand U1210 (N_1210,In_994,In_670);
and U1211 (N_1211,In_719,In_887);
and U1212 (N_1212,In_18,In_162);
nor U1213 (N_1213,In_989,In_345);
or U1214 (N_1214,In_66,In_177);
and U1215 (N_1215,In_293,In_614);
nand U1216 (N_1216,In_947,In_56);
and U1217 (N_1217,In_78,In_461);
and U1218 (N_1218,In_255,In_445);
xor U1219 (N_1219,In_223,In_606);
nor U1220 (N_1220,In_844,In_304);
xor U1221 (N_1221,In_155,In_515);
and U1222 (N_1222,In_352,In_228);
nand U1223 (N_1223,In_247,In_979);
nand U1224 (N_1224,In_875,In_970);
or U1225 (N_1225,In_732,In_72);
xor U1226 (N_1226,In_565,In_610);
nor U1227 (N_1227,In_926,In_587);
nand U1228 (N_1228,In_643,In_479);
or U1229 (N_1229,In_622,In_345);
nand U1230 (N_1230,In_392,In_856);
and U1231 (N_1231,In_648,In_821);
or U1232 (N_1232,In_764,In_255);
and U1233 (N_1233,In_63,In_795);
and U1234 (N_1234,In_488,In_603);
nor U1235 (N_1235,In_201,In_52);
and U1236 (N_1236,In_218,In_543);
or U1237 (N_1237,In_69,In_242);
xnor U1238 (N_1238,In_247,In_265);
or U1239 (N_1239,In_658,In_680);
and U1240 (N_1240,In_447,In_537);
nand U1241 (N_1241,In_882,In_303);
and U1242 (N_1242,In_917,In_807);
nor U1243 (N_1243,In_642,In_17);
and U1244 (N_1244,In_780,In_91);
and U1245 (N_1245,In_153,In_150);
nand U1246 (N_1246,In_310,In_393);
or U1247 (N_1247,In_108,In_858);
and U1248 (N_1248,In_71,In_229);
or U1249 (N_1249,In_529,In_897);
or U1250 (N_1250,In_255,In_594);
nor U1251 (N_1251,In_556,In_787);
and U1252 (N_1252,In_127,In_139);
and U1253 (N_1253,In_615,In_854);
or U1254 (N_1254,In_162,In_797);
nand U1255 (N_1255,In_726,In_256);
or U1256 (N_1256,In_861,In_225);
nand U1257 (N_1257,In_402,In_901);
nand U1258 (N_1258,In_184,In_392);
nor U1259 (N_1259,In_305,In_115);
xnor U1260 (N_1260,In_899,In_497);
or U1261 (N_1261,In_716,In_31);
nor U1262 (N_1262,In_64,In_369);
or U1263 (N_1263,In_948,In_929);
and U1264 (N_1264,In_377,In_227);
or U1265 (N_1265,In_575,In_973);
nor U1266 (N_1266,In_885,In_945);
or U1267 (N_1267,In_804,In_43);
or U1268 (N_1268,In_863,In_23);
or U1269 (N_1269,In_79,In_534);
or U1270 (N_1270,In_631,In_941);
or U1271 (N_1271,In_257,In_99);
and U1272 (N_1272,In_916,In_420);
and U1273 (N_1273,In_706,In_168);
or U1274 (N_1274,In_251,In_571);
nor U1275 (N_1275,In_652,In_755);
xnor U1276 (N_1276,In_962,In_464);
or U1277 (N_1277,In_637,In_350);
nor U1278 (N_1278,In_473,In_892);
nor U1279 (N_1279,In_435,In_433);
or U1280 (N_1280,In_232,In_35);
and U1281 (N_1281,In_257,In_712);
and U1282 (N_1282,In_247,In_686);
xor U1283 (N_1283,In_999,In_181);
and U1284 (N_1284,In_236,In_431);
or U1285 (N_1285,In_36,In_839);
or U1286 (N_1286,In_777,In_999);
or U1287 (N_1287,In_990,In_451);
or U1288 (N_1288,In_245,In_647);
or U1289 (N_1289,In_340,In_863);
or U1290 (N_1290,In_227,In_849);
and U1291 (N_1291,In_405,In_354);
or U1292 (N_1292,In_640,In_2);
nor U1293 (N_1293,In_247,In_866);
nor U1294 (N_1294,In_667,In_987);
and U1295 (N_1295,In_833,In_269);
nor U1296 (N_1296,In_689,In_92);
or U1297 (N_1297,In_567,In_694);
or U1298 (N_1298,In_664,In_347);
nor U1299 (N_1299,In_395,In_624);
or U1300 (N_1300,In_785,In_346);
nand U1301 (N_1301,In_153,In_486);
nand U1302 (N_1302,In_532,In_329);
nor U1303 (N_1303,In_720,In_639);
nand U1304 (N_1304,In_489,In_119);
or U1305 (N_1305,In_972,In_287);
or U1306 (N_1306,In_625,In_770);
or U1307 (N_1307,In_430,In_817);
nor U1308 (N_1308,In_623,In_273);
nor U1309 (N_1309,In_449,In_657);
or U1310 (N_1310,In_423,In_907);
or U1311 (N_1311,In_108,In_294);
or U1312 (N_1312,In_355,In_234);
and U1313 (N_1313,In_536,In_491);
nor U1314 (N_1314,In_78,In_838);
nor U1315 (N_1315,In_46,In_51);
nor U1316 (N_1316,In_722,In_968);
or U1317 (N_1317,In_564,In_532);
nand U1318 (N_1318,In_600,In_662);
nor U1319 (N_1319,In_215,In_214);
nand U1320 (N_1320,In_672,In_335);
and U1321 (N_1321,In_997,In_655);
xor U1322 (N_1322,In_500,In_110);
or U1323 (N_1323,In_656,In_53);
nand U1324 (N_1324,In_51,In_495);
nor U1325 (N_1325,In_978,In_391);
or U1326 (N_1326,In_465,In_428);
or U1327 (N_1327,In_669,In_464);
and U1328 (N_1328,In_116,In_733);
xor U1329 (N_1329,In_235,In_993);
nand U1330 (N_1330,In_286,In_723);
and U1331 (N_1331,In_837,In_325);
or U1332 (N_1332,In_37,In_359);
xor U1333 (N_1333,In_502,In_435);
nor U1334 (N_1334,In_120,In_825);
nor U1335 (N_1335,In_795,In_302);
nand U1336 (N_1336,In_229,In_86);
or U1337 (N_1337,In_79,In_420);
nand U1338 (N_1338,In_50,In_614);
nand U1339 (N_1339,In_353,In_42);
or U1340 (N_1340,In_704,In_166);
and U1341 (N_1341,In_180,In_443);
or U1342 (N_1342,In_126,In_866);
or U1343 (N_1343,In_407,In_524);
nor U1344 (N_1344,In_741,In_832);
or U1345 (N_1345,In_73,In_118);
and U1346 (N_1346,In_45,In_584);
nand U1347 (N_1347,In_809,In_863);
and U1348 (N_1348,In_209,In_930);
and U1349 (N_1349,In_88,In_732);
nand U1350 (N_1350,In_864,In_697);
nor U1351 (N_1351,In_887,In_726);
xor U1352 (N_1352,In_250,In_560);
nand U1353 (N_1353,In_991,In_218);
nand U1354 (N_1354,In_297,In_958);
or U1355 (N_1355,In_150,In_238);
or U1356 (N_1356,In_962,In_618);
and U1357 (N_1357,In_265,In_255);
and U1358 (N_1358,In_962,In_93);
and U1359 (N_1359,In_815,In_668);
nor U1360 (N_1360,In_259,In_212);
or U1361 (N_1361,In_40,In_723);
and U1362 (N_1362,In_447,In_59);
nand U1363 (N_1363,In_937,In_50);
or U1364 (N_1364,In_497,In_718);
nor U1365 (N_1365,In_941,In_855);
nor U1366 (N_1366,In_826,In_623);
nand U1367 (N_1367,In_782,In_458);
or U1368 (N_1368,In_282,In_758);
or U1369 (N_1369,In_518,In_186);
or U1370 (N_1370,In_216,In_342);
or U1371 (N_1371,In_946,In_236);
nand U1372 (N_1372,In_897,In_740);
nand U1373 (N_1373,In_880,In_818);
nand U1374 (N_1374,In_966,In_620);
nand U1375 (N_1375,In_364,In_249);
nor U1376 (N_1376,In_892,In_678);
and U1377 (N_1377,In_538,In_993);
and U1378 (N_1378,In_332,In_469);
nand U1379 (N_1379,In_653,In_177);
nand U1380 (N_1380,In_425,In_206);
nor U1381 (N_1381,In_937,In_490);
nand U1382 (N_1382,In_901,In_724);
and U1383 (N_1383,In_21,In_475);
nor U1384 (N_1384,In_263,In_919);
or U1385 (N_1385,In_644,In_904);
or U1386 (N_1386,In_857,In_529);
nor U1387 (N_1387,In_945,In_21);
and U1388 (N_1388,In_832,In_86);
and U1389 (N_1389,In_405,In_921);
or U1390 (N_1390,In_211,In_144);
nand U1391 (N_1391,In_769,In_526);
or U1392 (N_1392,In_399,In_842);
nand U1393 (N_1393,In_734,In_814);
or U1394 (N_1394,In_854,In_600);
and U1395 (N_1395,In_240,In_690);
and U1396 (N_1396,In_647,In_403);
and U1397 (N_1397,In_624,In_244);
or U1398 (N_1398,In_538,In_438);
and U1399 (N_1399,In_894,In_597);
nor U1400 (N_1400,In_323,In_492);
and U1401 (N_1401,In_701,In_675);
or U1402 (N_1402,In_991,In_224);
or U1403 (N_1403,In_132,In_100);
and U1404 (N_1404,In_472,In_198);
nor U1405 (N_1405,In_626,In_877);
or U1406 (N_1406,In_915,In_471);
or U1407 (N_1407,In_837,In_78);
nor U1408 (N_1408,In_499,In_322);
nand U1409 (N_1409,In_216,In_331);
and U1410 (N_1410,In_810,In_676);
and U1411 (N_1411,In_169,In_600);
and U1412 (N_1412,In_995,In_497);
nand U1413 (N_1413,In_264,In_455);
and U1414 (N_1414,In_646,In_879);
and U1415 (N_1415,In_817,In_376);
nor U1416 (N_1416,In_62,In_52);
nor U1417 (N_1417,In_714,In_517);
or U1418 (N_1418,In_27,In_395);
nand U1419 (N_1419,In_510,In_478);
or U1420 (N_1420,In_263,In_985);
nand U1421 (N_1421,In_931,In_196);
and U1422 (N_1422,In_809,In_223);
nand U1423 (N_1423,In_468,In_363);
and U1424 (N_1424,In_509,In_306);
nand U1425 (N_1425,In_680,In_617);
and U1426 (N_1426,In_662,In_38);
nand U1427 (N_1427,In_50,In_701);
nand U1428 (N_1428,In_702,In_132);
and U1429 (N_1429,In_432,In_354);
nand U1430 (N_1430,In_421,In_818);
nand U1431 (N_1431,In_6,In_363);
nor U1432 (N_1432,In_848,In_385);
nand U1433 (N_1433,In_280,In_210);
nor U1434 (N_1434,In_888,In_782);
nor U1435 (N_1435,In_302,In_965);
nor U1436 (N_1436,In_386,In_767);
and U1437 (N_1437,In_319,In_335);
nor U1438 (N_1438,In_933,In_635);
nand U1439 (N_1439,In_127,In_584);
nor U1440 (N_1440,In_686,In_613);
xor U1441 (N_1441,In_9,In_930);
or U1442 (N_1442,In_199,In_517);
nand U1443 (N_1443,In_24,In_441);
xnor U1444 (N_1444,In_857,In_262);
nand U1445 (N_1445,In_164,In_475);
nor U1446 (N_1446,In_359,In_394);
nor U1447 (N_1447,In_523,In_495);
nor U1448 (N_1448,In_405,In_199);
and U1449 (N_1449,In_520,In_462);
and U1450 (N_1450,In_285,In_720);
or U1451 (N_1451,In_442,In_146);
nand U1452 (N_1452,In_186,In_248);
or U1453 (N_1453,In_873,In_231);
nand U1454 (N_1454,In_851,In_79);
nand U1455 (N_1455,In_149,In_623);
or U1456 (N_1456,In_336,In_674);
and U1457 (N_1457,In_411,In_45);
and U1458 (N_1458,In_737,In_436);
and U1459 (N_1459,In_459,In_457);
nand U1460 (N_1460,In_850,In_326);
nand U1461 (N_1461,In_748,In_358);
nor U1462 (N_1462,In_437,In_540);
and U1463 (N_1463,In_452,In_539);
nand U1464 (N_1464,In_790,In_58);
or U1465 (N_1465,In_398,In_643);
or U1466 (N_1466,In_611,In_813);
nand U1467 (N_1467,In_431,In_406);
nand U1468 (N_1468,In_343,In_951);
nand U1469 (N_1469,In_766,In_460);
or U1470 (N_1470,In_737,In_221);
nor U1471 (N_1471,In_551,In_460);
and U1472 (N_1472,In_787,In_823);
nand U1473 (N_1473,In_6,In_159);
and U1474 (N_1474,In_396,In_869);
nand U1475 (N_1475,In_707,In_301);
nand U1476 (N_1476,In_713,In_784);
nor U1477 (N_1477,In_59,In_236);
nor U1478 (N_1478,In_262,In_627);
and U1479 (N_1479,In_351,In_888);
nand U1480 (N_1480,In_405,In_723);
nand U1481 (N_1481,In_82,In_151);
nand U1482 (N_1482,In_314,In_385);
or U1483 (N_1483,In_677,In_818);
xnor U1484 (N_1484,In_85,In_774);
or U1485 (N_1485,In_355,In_546);
xnor U1486 (N_1486,In_689,In_405);
and U1487 (N_1487,In_505,In_863);
nand U1488 (N_1488,In_529,In_738);
nor U1489 (N_1489,In_757,In_407);
xnor U1490 (N_1490,In_193,In_758);
nor U1491 (N_1491,In_516,In_172);
or U1492 (N_1492,In_759,In_767);
or U1493 (N_1493,In_975,In_898);
nand U1494 (N_1494,In_291,In_188);
and U1495 (N_1495,In_146,In_170);
or U1496 (N_1496,In_134,In_761);
nor U1497 (N_1497,In_201,In_506);
or U1498 (N_1498,In_966,In_573);
nor U1499 (N_1499,In_200,In_552);
nand U1500 (N_1500,In_623,In_482);
or U1501 (N_1501,In_558,In_435);
nand U1502 (N_1502,In_863,In_228);
nor U1503 (N_1503,In_879,In_567);
nor U1504 (N_1504,In_166,In_532);
nor U1505 (N_1505,In_228,In_423);
nor U1506 (N_1506,In_88,In_31);
nand U1507 (N_1507,In_233,In_616);
nand U1508 (N_1508,In_828,In_882);
and U1509 (N_1509,In_426,In_543);
nor U1510 (N_1510,In_748,In_601);
and U1511 (N_1511,In_638,In_761);
nand U1512 (N_1512,In_49,In_635);
nor U1513 (N_1513,In_649,In_494);
nor U1514 (N_1514,In_834,In_422);
nor U1515 (N_1515,In_125,In_841);
nand U1516 (N_1516,In_222,In_710);
and U1517 (N_1517,In_846,In_492);
xor U1518 (N_1518,In_892,In_101);
and U1519 (N_1519,In_59,In_420);
nand U1520 (N_1520,In_644,In_369);
nand U1521 (N_1521,In_7,In_887);
nor U1522 (N_1522,In_720,In_346);
nand U1523 (N_1523,In_182,In_585);
xor U1524 (N_1524,In_61,In_41);
and U1525 (N_1525,In_42,In_803);
nor U1526 (N_1526,In_960,In_171);
nand U1527 (N_1527,In_100,In_3);
or U1528 (N_1528,In_429,In_638);
or U1529 (N_1529,In_660,In_850);
and U1530 (N_1530,In_303,In_466);
nand U1531 (N_1531,In_722,In_514);
nor U1532 (N_1532,In_610,In_129);
nor U1533 (N_1533,In_35,In_478);
and U1534 (N_1534,In_586,In_350);
nand U1535 (N_1535,In_705,In_604);
nand U1536 (N_1536,In_367,In_447);
or U1537 (N_1537,In_348,In_18);
or U1538 (N_1538,In_851,In_802);
xor U1539 (N_1539,In_401,In_225);
or U1540 (N_1540,In_418,In_882);
and U1541 (N_1541,In_385,In_717);
nand U1542 (N_1542,In_440,In_693);
nor U1543 (N_1543,In_611,In_485);
or U1544 (N_1544,In_199,In_88);
nor U1545 (N_1545,In_948,In_694);
nor U1546 (N_1546,In_361,In_567);
or U1547 (N_1547,In_992,In_503);
or U1548 (N_1548,In_318,In_87);
nand U1549 (N_1549,In_484,In_173);
nor U1550 (N_1550,In_590,In_903);
nand U1551 (N_1551,In_803,In_347);
nor U1552 (N_1552,In_346,In_616);
nor U1553 (N_1553,In_697,In_626);
or U1554 (N_1554,In_248,In_886);
and U1555 (N_1555,In_434,In_538);
nor U1556 (N_1556,In_207,In_447);
and U1557 (N_1557,In_633,In_451);
nor U1558 (N_1558,In_128,In_523);
nor U1559 (N_1559,In_302,In_11);
or U1560 (N_1560,In_34,In_348);
nor U1561 (N_1561,In_996,In_183);
or U1562 (N_1562,In_607,In_267);
nor U1563 (N_1563,In_407,In_71);
nor U1564 (N_1564,In_88,In_178);
and U1565 (N_1565,In_632,In_169);
and U1566 (N_1566,In_654,In_650);
nand U1567 (N_1567,In_145,In_856);
nand U1568 (N_1568,In_744,In_16);
nand U1569 (N_1569,In_146,In_781);
nor U1570 (N_1570,In_511,In_329);
and U1571 (N_1571,In_344,In_381);
nor U1572 (N_1572,In_225,In_782);
nand U1573 (N_1573,In_921,In_49);
and U1574 (N_1574,In_613,In_364);
or U1575 (N_1575,In_663,In_336);
nand U1576 (N_1576,In_993,In_249);
or U1577 (N_1577,In_592,In_566);
nor U1578 (N_1578,In_719,In_279);
or U1579 (N_1579,In_174,In_338);
or U1580 (N_1580,In_788,In_873);
and U1581 (N_1581,In_800,In_672);
nand U1582 (N_1582,In_230,In_292);
or U1583 (N_1583,In_326,In_300);
nor U1584 (N_1584,In_474,In_802);
nor U1585 (N_1585,In_811,In_79);
nand U1586 (N_1586,In_140,In_304);
and U1587 (N_1587,In_843,In_667);
nand U1588 (N_1588,In_607,In_967);
and U1589 (N_1589,In_880,In_277);
nor U1590 (N_1590,In_846,In_845);
or U1591 (N_1591,In_271,In_150);
or U1592 (N_1592,In_747,In_441);
nand U1593 (N_1593,In_268,In_598);
or U1594 (N_1594,In_447,In_264);
or U1595 (N_1595,In_890,In_916);
nand U1596 (N_1596,In_246,In_425);
nand U1597 (N_1597,In_634,In_347);
or U1598 (N_1598,In_959,In_856);
and U1599 (N_1599,In_124,In_107);
nand U1600 (N_1600,In_393,In_553);
or U1601 (N_1601,In_12,In_588);
or U1602 (N_1602,In_479,In_872);
and U1603 (N_1603,In_827,In_702);
nand U1604 (N_1604,In_986,In_87);
and U1605 (N_1605,In_379,In_86);
nor U1606 (N_1606,In_261,In_209);
nand U1607 (N_1607,In_839,In_344);
nor U1608 (N_1608,In_835,In_256);
nor U1609 (N_1609,In_295,In_398);
or U1610 (N_1610,In_641,In_100);
or U1611 (N_1611,In_407,In_261);
nor U1612 (N_1612,In_224,In_513);
and U1613 (N_1613,In_979,In_505);
or U1614 (N_1614,In_534,In_652);
nand U1615 (N_1615,In_672,In_64);
or U1616 (N_1616,In_489,In_75);
nor U1617 (N_1617,In_330,In_728);
or U1618 (N_1618,In_588,In_440);
nand U1619 (N_1619,In_328,In_49);
and U1620 (N_1620,In_816,In_533);
and U1621 (N_1621,In_199,In_346);
nor U1622 (N_1622,In_111,In_480);
nor U1623 (N_1623,In_560,In_184);
and U1624 (N_1624,In_599,In_331);
nand U1625 (N_1625,In_578,In_925);
xor U1626 (N_1626,In_749,In_410);
or U1627 (N_1627,In_610,In_875);
nand U1628 (N_1628,In_324,In_524);
or U1629 (N_1629,In_892,In_623);
and U1630 (N_1630,In_386,In_40);
nor U1631 (N_1631,In_527,In_876);
nand U1632 (N_1632,In_204,In_295);
or U1633 (N_1633,In_934,In_639);
or U1634 (N_1634,In_676,In_734);
and U1635 (N_1635,In_303,In_344);
nand U1636 (N_1636,In_845,In_666);
or U1637 (N_1637,In_883,In_393);
nor U1638 (N_1638,In_960,In_445);
and U1639 (N_1639,In_313,In_164);
nand U1640 (N_1640,In_770,In_298);
nor U1641 (N_1641,In_446,In_284);
or U1642 (N_1642,In_121,In_241);
nand U1643 (N_1643,In_289,In_555);
or U1644 (N_1644,In_598,In_246);
nand U1645 (N_1645,In_435,In_701);
nand U1646 (N_1646,In_607,In_626);
and U1647 (N_1647,In_797,In_941);
nor U1648 (N_1648,In_283,In_375);
nand U1649 (N_1649,In_699,In_287);
or U1650 (N_1650,In_375,In_971);
nor U1651 (N_1651,In_517,In_315);
and U1652 (N_1652,In_130,In_471);
nor U1653 (N_1653,In_33,In_797);
nand U1654 (N_1654,In_601,In_541);
or U1655 (N_1655,In_702,In_754);
nand U1656 (N_1656,In_116,In_985);
and U1657 (N_1657,In_139,In_653);
nor U1658 (N_1658,In_625,In_816);
or U1659 (N_1659,In_980,In_916);
nor U1660 (N_1660,In_855,In_387);
or U1661 (N_1661,In_360,In_465);
or U1662 (N_1662,In_428,In_718);
nand U1663 (N_1663,In_4,In_709);
xor U1664 (N_1664,In_33,In_41);
nor U1665 (N_1665,In_323,In_511);
nand U1666 (N_1666,In_465,In_246);
nand U1667 (N_1667,In_957,In_716);
or U1668 (N_1668,In_783,In_943);
nor U1669 (N_1669,In_407,In_279);
and U1670 (N_1670,In_418,In_48);
nand U1671 (N_1671,In_296,In_721);
nand U1672 (N_1672,In_419,In_622);
or U1673 (N_1673,In_580,In_157);
and U1674 (N_1674,In_763,In_367);
or U1675 (N_1675,In_20,In_125);
or U1676 (N_1676,In_152,In_77);
nand U1677 (N_1677,In_484,In_820);
or U1678 (N_1678,In_651,In_128);
nand U1679 (N_1679,In_719,In_8);
or U1680 (N_1680,In_476,In_504);
and U1681 (N_1681,In_312,In_786);
nor U1682 (N_1682,In_736,In_955);
and U1683 (N_1683,In_607,In_917);
and U1684 (N_1684,In_812,In_106);
or U1685 (N_1685,In_865,In_546);
nand U1686 (N_1686,In_5,In_709);
nand U1687 (N_1687,In_732,In_194);
nand U1688 (N_1688,In_18,In_578);
or U1689 (N_1689,In_687,In_746);
or U1690 (N_1690,In_917,In_18);
and U1691 (N_1691,In_234,In_702);
nand U1692 (N_1692,In_17,In_115);
nand U1693 (N_1693,In_769,In_268);
or U1694 (N_1694,In_965,In_377);
or U1695 (N_1695,In_796,In_177);
nor U1696 (N_1696,In_205,In_23);
or U1697 (N_1697,In_373,In_422);
nor U1698 (N_1698,In_612,In_595);
or U1699 (N_1699,In_652,In_207);
nand U1700 (N_1700,In_592,In_930);
nor U1701 (N_1701,In_849,In_714);
nand U1702 (N_1702,In_879,In_69);
and U1703 (N_1703,In_755,In_600);
or U1704 (N_1704,In_800,In_868);
nor U1705 (N_1705,In_615,In_712);
or U1706 (N_1706,In_239,In_189);
nand U1707 (N_1707,In_940,In_722);
or U1708 (N_1708,In_651,In_307);
and U1709 (N_1709,In_100,In_922);
or U1710 (N_1710,In_936,In_958);
and U1711 (N_1711,In_345,In_552);
or U1712 (N_1712,In_892,In_316);
or U1713 (N_1713,In_695,In_566);
and U1714 (N_1714,In_153,In_921);
and U1715 (N_1715,In_155,In_763);
and U1716 (N_1716,In_770,In_204);
nor U1717 (N_1717,In_767,In_660);
or U1718 (N_1718,In_321,In_675);
nor U1719 (N_1719,In_426,In_853);
and U1720 (N_1720,In_817,In_247);
and U1721 (N_1721,In_209,In_11);
or U1722 (N_1722,In_884,In_705);
nand U1723 (N_1723,In_340,In_912);
or U1724 (N_1724,In_194,In_31);
nand U1725 (N_1725,In_434,In_889);
nand U1726 (N_1726,In_14,In_212);
and U1727 (N_1727,In_759,In_557);
and U1728 (N_1728,In_953,In_321);
or U1729 (N_1729,In_672,In_472);
and U1730 (N_1730,In_282,In_725);
and U1731 (N_1731,In_57,In_45);
nor U1732 (N_1732,In_460,In_260);
nor U1733 (N_1733,In_888,In_100);
nor U1734 (N_1734,In_234,In_258);
nor U1735 (N_1735,In_568,In_25);
nand U1736 (N_1736,In_139,In_674);
or U1737 (N_1737,In_121,In_45);
or U1738 (N_1738,In_41,In_737);
nor U1739 (N_1739,In_636,In_105);
or U1740 (N_1740,In_40,In_441);
nor U1741 (N_1741,In_633,In_81);
nand U1742 (N_1742,In_261,In_584);
or U1743 (N_1743,In_963,In_789);
and U1744 (N_1744,In_57,In_262);
or U1745 (N_1745,In_394,In_2);
nand U1746 (N_1746,In_386,In_183);
or U1747 (N_1747,In_147,In_987);
nor U1748 (N_1748,In_881,In_770);
or U1749 (N_1749,In_549,In_173);
nand U1750 (N_1750,In_1,In_133);
and U1751 (N_1751,In_409,In_763);
nor U1752 (N_1752,In_328,In_120);
and U1753 (N_1753,In_571,In_220);
nor U1754 (N_1754,In_459,In_311);
xnor U1755 (N_1755,In_116,In_566);
xor U1756 (N_1756,In_370,In_835);
nor U1757 (N_1757,In_344,In_877);
nor U1758 (N_1758,In_667,In_357);
or U1759 (N_1759,In_480,In_326);
and U1760 (N_1760,In_954,In_430);
and U1761 (N_1761,In_968,In_452);
nand U1762 (N_1762,In_989,In_648);
and U1763 (N_1763,In_776,In_711);
or U1764 (N_1764,In_983,In_235);
and U1765 (N_1765,In_292,In_914);
nor U1766 (N_1766,In_133,In_427);
nand U1767 (N_1767,In_984,In_344);
xnor U1768 (N_1768,In_18,In_433);
nand U1769 (N_1769,In_807,In_290);
or U1770 (N_1770,In_25,In_697);
nand U1771 (N_1771,In_852,In_266);
nand U1772 (N_1772,In_973,In_835);
nand U1773 (N_1773,In_313,In_336);
nor U1774 (N_1774,In_409,In_145);
and U1775 (N_1775,In_724,In_782);
nand U1776 (N_1776,In_289,In_98);
nor U1777 (N_1777,In_916,In_762);
nor U1778 (N_1778,In_636,In_512);
nor U1779 (N_1779,In_463,In_490);
and U1780 (N_1780,In_380,In_803);
nand U1781 (N_1781,In_137,In_731);
nand U1782 (N_1782,In_434,In_936);
and U1783 (N_1783,In_459,In_616);
and U1784 (N_1784,In_557,In_221);
nor U1785 (N_1785,In_571,In_859);
nor U1786 (N_1786,In_977,In_315);
or U1787 (N_1787,In_150,In_45);
nand U1788 (N_1788,In_388,In_156);
nor U1789 (N_1789,In_257,In_40);
and U1790 (N_1790,In_897,In_310);
and U1791 (N_1791,In_724,In_884);
nand U1792 (N_1792,In_320,In_244);
nand U1793 (N_1793,In_670,In_609);
or U1794 (N_1794,In_397,In_598);
nor U1795 (N_1795,In_512,In_651);
nor U1796 (N_1796,In_737,In_949);
or U1797 (N_1797,In_788,In_727);
and U1798 (N_1798,In_735,In_232);
and U1799 (N_1799,In_7,In_100);
nor U1800 (N_1800,In_226,In_665);
or U1801 (N_1801,In_71,In_1);
nor U1802 (N_1802,In_16,In_942);
or U1803 (N_1803,In_554,In_742);
nand U1804 (N_1804,In_459,In_340);
nor U1805 (N_1805,In_105,In_98);
nand U1806 (N_1806,In_100,In_337);
nor U1807 (N_1807,In_653,In_835);
and U1808 (N_1808,In_944,In_493);
nor U1809 (N_1809,In_78,In_711);
nor U1810 (N_1810,In_205,In_51);
nor U1811 (N_1811,In_821,In_145);
xor U1812 (N_1812,In_902,In_784);
nand U1813 (N_1813,In_861,In_237);
nor U1814 (N_1814,In_436,In_964);
xnor U1815 (N_1815,In_815,In_126);
nand U1816 (N_1816,In_333,In_572);
nand U1817 (N_1817,In_506,In_796);
and U1818 (N_1818,In_12,In_286);
and U1819 (N_1819,In_561,In_773);
and U1820 (N_1820,In_911,In_435);
and U1821 (N_1821,In_446,In_629);
nand U1822 (N_1822,In_23,In_77);
nor U1823 (N_1823,In_362,In_415);
nand U1824 (N_1824,In_723,In_918);
nor U1825 (N_1825,In_872,In_464);
nor U1826 (N_1826,In_836,In_816);
nor U1827 (N_1827,In_598,In_451);
xor U1828 (N_1828,In_351,In_613);
nor U1829 (N_1829,In_652,In_997);
and U1830 (N_1830,In_252,In_476);
nand U1831 (N_1831,In_477,In_652);
and U1832 (N_1832,In_84,In_647);
nor U1833 (N_1833,In_892,In_140);
and U1834 (N_1834,In_312,In_265);
or U1835 (N_1835,In_322,In_975);
or U1836 (N_1836,In_273,In_225);
and U1837 (N_1837,In_895,In_86);
and U1838 (N_1838,In_28,In_105);
or U1839 (N_1839,In_93,In_633);
and U1840 (N_1840,In_275,In_376);
nand U1841 (N_1841,In_388,In_743);
nand U1842 (N_1842,In_509,In_650);
and U1843 (N_1843,In_300,In_419);
or U1844 (N_1844,In_201,In_624);
and U1845 (N_1845,In_943,In_277);
nand U1846 (N_1846,In_787,In_921);
or U1847 (N_1847,In_626,In_979);
nand U1848 (N_1848,In_162,In_987);
xor U1849 (N_1849,In_973,In_792);
nand U1850 (N_1850,In_353,In_692);
and U1851 (N_1851,In_239,In_831);
nand U1852 (N_1852,In_253,In_234);
nand U1853 (N_1853,In_623,In_420);
or U1854 (N_1854,In_811,In_944);
or U1855 (N_1855,In_539,In_189);
nand U1856 (N_1856,In_787,In_809);
or U1857 (N_1857,In_922,In_355);
nor U1858 (N_1858,In_129,In_459);
and U1859 (N_1859,In_518,In_306);
nand U1860 (N_1860,In_226,In_215);
or U1861 (N_1861,In_243,In_41);
nand U1862 (N_1862,In_180,In_831);
or U1863 (N_1863,In_286,In_777);
nor U1864 (N_1864,In_375,In_587);
nand U1865 (N_1865,In_117,In_73);
or U1866 (N_1866,In_50,In_718);
nor U1867 (N_1867,In_231,In_851);
and U1868 (N_1868,In_969,In_775);
nand U1869 (N_1869,In_521,In_243);
or U1870 (N_1870,In_520,In_214);
xnor U1871 (N_1871,In_196,In_93);
nor U1872 (N_1872,In_208,In_598);
and U1873 (N_1873,In_403,In_101);
nor U1874 (N_1874,In_178,In_8);
nor U1875 (N_1875,In_401,In_846);
nor U1876 (N_1876,In_93,In_972);
or U1877 (N_1877,In_105,In_263);
and U1878 (N_1878,In_83,In_874);
nor U1879 (N_1879,In_681,In_309);
or U1880 (N_1880,In_573,In_938);
nor U1881 (N_1881,In_718,In_696);
or U1882 (N_1882,In_229,In_614);
nand U1883 (N_1883,In_850,In_452);
and U1884 (N_1884,In_183,In_772);
and U1885 (N_1885,In_813,In_829);
nand U1886 (N_1886,In_313,In_4);
or U1887 (N_1887,In_789,In_352);
nand U1888 (N_1888,In_716,In_150);
and U1889 (N_1889,In_25,In_508);
nand U1890 (N_1890,In_313,In_631);
xnor U1891 (N_1891,In_508,In_318);
xnor U1892 (N_1892,In_29,In_624);
nand U1893 (N_1893,In_456,In_500);
or U1894 (N_1894,In_98,In_502);
nor U1895 (N_1895,In_423,In_167);
and U1896 (N_1896,In_917,In_964);
and U1897 (N_1897,In_43,In_321);
nand U1898 (N_1898,In_871,In_727);
nor U1899 (N_1899,In_782,In_901);
nand U1900 (N_1900,In_322,In_406);
or U1901 (N_1901,In_35,In_437);
nand U1902 (N_1902,In_91,In_748);
or U1903 (N_1903,In_711,In_58);
nand U1904 (N_1904,In_632,In_789);
nand U1905 (N_1905,In_516,In_175);
nand U1906 (N_1906,In_4,In_80);
nand U1907 (N_1907,In_586,In_895);
nor U1908 (N_1908,In_136,In_523);
and U1909 (N_1909,In_88,In_429);
nor U1910 (N_1910,In_101,In_782);
nor U1911 (N_1911,In_68,In_704);
nand U1912 (N_1912,In_981,In_317);
nand U1913 (N_1913,In_603,In_434);
nor U1914 (N_1914,In_596,In_933);
or U1915 (N_1915,In_368,In_360);
xor U1916 (N_1916,In_422,In_729);
or U1917 (N_1917,In_408,In_535);
nand U1918 (N_1918,In_873,In_862);
or U1919 (N_1919,In_492,In_742);
nor U1920 (N_1920,In_77,In_221);
nor U1921 (N_1921,In_890,In_954);
or U1922 (N_1922,In_191,In_300);
nor U1923 (N_1923,In_402,In_896);
or U1924 (N_1924,In_342,In_791);
and U1925 (N_1925,In_633,In_542);
and U1926 (N_1926,In_22,In_231);
or U1927 (N_1927,In_38,In_162);
or U1928 (N_1928,In_893,In_760);
or U1929 (N_1929,In_522,In_328);
nor U1930 (N_1930,In_331,In_439);
and U1931 (N_1931,In_573,In_665);
nor U1932 (N_1932,In_440,In_757);
nand U1933 (N_1933,In_553,In_564);
and U1934 (N_1934,In_801,In_257);
or U1935 (N_1935,In_832,In_526);
and U1936 (N_1936,In_4,In_514);
or U1937 (N_1937,In_448,In_348);
nor U1938 (N_1938,In_488,In_190);
or U1939 (N_1939,In_233,In_243);
nor U1940 (N_1940,In_390,In_304);
or U1941 (N_1941,In_928,In_275);
nor U1942 (N_1942,In_541,In_176);
nor U1943 (N_1943,In_57,In_47);
nand U1944 (N_1944,In_838,In_857);
and U1945 (N_1945,In_705,In_543);
nand U1946 (N_1946,In_812,In_842);
nor U1947 (N_1947,In_100,In_395);
nor U1948 (N_1948,In_373,In_655);
nor U1949 (N_1949,In_974,In_841);
and U1950 (N_1950,In_283,In_775);
or U1951 (N_1951,In_906,In_417);
nor U1952 (N_1952,In_752,In_920);
nor U1953 (N_1953,In_812,In_389);
nor U1954 (N_1954,In_904,In_903);
or U1955 (N_1955,In_985,In_694);
and U1956 (N_1956,In_525,In_555);
nor U1957 (N_1957,In_375,In_331);
nor U1958 (N_1958,In_845,In_423);
nor U1959 (N_1959,In_142,In_937);
and U1960 (N_1960,In_79,In_528);
nand U1961 (N_1961,In_128,In_763);
and U1962 (N_1962,In_348,In_731);
and U1963 (N_1963,In_98,In_614);
and U1964 (N_1964,In_731,In_857);
nand U1965 (N_1965,In_691,In_277);
nor U1966 (N_1966,In_517,In_349);
nor U1967 (N_1967,In_419,In_220);
or U1968 (N_1968,In_730,In_545);
or U1969 (N_1969,In_935,In_389);
nand U1970 (N_1970,In_169,In_60);
nor U1971 (N_1971,In_59,In_851);
and U1972 (N_1972,In_897,In_775);
and U1973 (N_1973,In_924,In_659);
or U1974 (N_1974,In_944,In_708);
and U1975 (N_1975,In_211,In_723);
and U1976 (N_1976,In_862,In_774);
or U1977 (N_1977,In_713,In_380);
nor U1978 (N_1978,In_312,In_619);
or U1979 (N_1979,In_324,In_659);
and U1980 (N_1980,In_661,In_230);
or U1981 (N_1981,In_624,In_598);
xor U1982 (N_1982,In_157,In_570);
nor U1983 (N_1983,In_762,In_193);
nand U1984 (N_1984,In_967,In_774);
and U1985 (N_1985,In_226,In_817);
nand U1986 (N_1986,In_164,In_359);
nand U1987 (N_1987,In_397,In_349);
and U1988 (N_1988,In_640,In_749);
and U1989 (N_1989,In_504,In_213);
and U1990 (N_1990,In_133,In_690);
nand U1991 (N_1991,In_395,In_425);
nand U1992 (N_1992,In_517,In_254);
or U1993 (N_1993,In_582,In_723);
or U1994 (N_1994,In_713,In_431);
xor U1995 (N_1995,In_151,In_657);
or U1996 (N_1996,In_192,In_69);
nor U1997 (N_1997,In_835,In_878);
nand U1998 (N_1998,In_651,In_954);
nor U1999 (N_1999,In_770,In_138);
or U2000 (N_2000,N_1632,N_1948);
xor U2001 (N_2001,N_1487,N_644);
or U2002 (N_2002,N_1030,N_503);
and U2003 (N_2003,N_1119,N_308);
nor U2004 (N_2004,N_206,N_316);
or U2005 (N_2005,N_596,N_1663);
and U2006 (N_2006,N_1051,N_593);
nand U2007 (N_2007,N_60,N_698);
nand U2008 (N_2008,N_586,N_1822);
or U2009 (N_2009,N_330,N_115);
nand U2010 (N_2010,N_938,N_84);
and U2011 (N_2011,N_315,N_5);
or U2012 (N_2012,N_1209,N_1234);
and U2013 (N_2013,N_673,N_625);
or U2014 (N_2014,N_936,N_656);
or U2015 (N_2015,N_931,N_1521);
nor U2016 (N_2016,N_164,N_255);
xnor U2017 (N_2017,N_1771,N_1984);
nand U2018 (N_2018,N_1802,N_1781);
or U2019 (N_2019,N_1720,N_1257);
or U2020 (N_2020,N_839,N_1329);
xnor U2021 (N_2021,N_1456,N_437);
and U2022 (N_2022,N_1689,N_957);
nor U2023 (N_2023,N_1612,N_1816);
and U2024 (N_2024,N_1215,N_101);
or U2025 (N_2025,N_968,N_710);
nand U2026 (N_2026,N_1007,N_1682);
and U2027 (N_2027,N_1295,N_896);
and U2028 (N_2028,N_1551,N_218);
and U2029 (N_2029,N_554,N_1541);
nor U2030 (N_2030,N_1873,N_1472);
or U2031 (N_2031,N_1388,N_298);
nand U2032 (N_2032,N_264,N_239);
or U2033 (N_2033,N_834,N_857);
or U2034 (N_2034,N_749,N_181);
nand U2035 (N_2035,N_195,N_464);
nand U2036 (N_2036,N_1213,N_555);
nor U2037 (N_2037,N_1005,N_1300);
and U2038 (N_2038,N_138,N_948);
xor U2039 (N_2039,N_974,N_1639);
nand U2040 (N_2040,N_1634,N_1233);
nand U2041 (N_2041,N_1885,N_960);
nand U2042 (N_2042,N_530,N_782);
nor U2043 (N_2043,N_790,N_990);
and U2044 (N_2044,N_478,N_860);
nand U2045 (N_2045,N_1704,N_1597);
nor U2046 (N_2046,N_1672,N_1364);
nor U2047 (N_2047,N_760,N_898);
nor U2048 (N_2048,N_764,N_1272);
nand U2049 (N_2049,N_1509,N_1365);
nor U2050 (N_2050,N_1435,N_301);
or U2051 (N_2051,N_809,N_328);
and U2052 (N_2052,N_525,N_432);
or U2053 (N_2053,N_325,N_279);
and U2054 (N_2054,N_1746,N_191);
nand U2055 (N_2055,N_230,N_311);
or U2056 (N_2056,N_1384,N_462);
or U2057 (N_2057,N_352,N_709);
nand U2058 (N_2058,N_1316,N_1350);
xnor U2059 (N_2059,N_193,N_558);
and U2060 (N_2060,N_28,N_632);
nand U2061 (N_2061,N_306,N_141);
or U2062 (N_2062,N_1359,N_12);
and U2063 (N_2063,N_1477,N_535);
or U2064 (N_2064,N_336,N_1382);
nand U2065 (N_2065,N_47,N_1309);
xnor U2066 (N_2066,N_34,N_1320);
or U2067 (N_2067,N_980,N_1627);
or U2068 (N_2068,N_1910,N_488);
or U2069 (N_2069,N_1953,N_4);
or U2070 (N_2070,N_649,N_1163);
and U2071 (N_2071,N_1537,N_543);
nand U2072 (N_2072,N_946,N_1017);
nor U2073 (N_2073,N_811,N_1305);
nand U2074 (N_2074,N_1648,N_1080);
and U2075 (N_2075,N_1540,N_1990);
or U2076 (N_2076,N_480,N_774);
and U2077 (N_2077,N_914,N_819);
xor U2078 (N_2078,N_1250,N_1795);
nand U2079 (N_2079,N_1614,N_1923);
and U2080 (N_2080,N_1688,N_1633);
nor U2081 (N_2081,N_1308,N_307);
xnor U2082 (N_2082,N_1941,N_147);
and U2083 (N_2083,N_73,N_196);
nand U2084 (N_2084,N_1399,N_995);
and U2085 (N_2085,N_601,N_581);
nand U2086 (N_2086,N_551,N_1480);
nand U2087 (N_2087,N_1160,N_1381);
or U2088 (N_2088,N_272,N_384);
xor U2089 (N_2089,N_1149,N_1865);
or U2090 (N_2090,N_1545,N_1071);
or U2091 (N_2091,N_1932,N_192);
or U2092 (N_2092,N_747,N_637);
or U2093 (N_2093,N_1556,N_1060);
and U2094 (N_2094,N_420,N_1067);
xor U2095 (N_2095,N_1488,N_470);
nor U2096 (N_2096,N_1579,N_456);
nand U2097 (N_2097,N_189,N_728);
and U2098 (N_2098,N_969,N_81);
or U2099 (N_2099,N_1539,N_1425);
nor U2100 (N_2100,N_492,N_1064);
nand U2101 (N_2101,N_234,N_227);
or U2102 (N_2102,N_1286,N_259);
or U2103 (N_2103,N_1889,N_416);
or U2104 (N_2104,N_263,N_63);
and U2105 (N_2105,N_1188,N_1332);
nand U2106 (N_2106,N_734,N_987);
nor U2107 (N_2107,N_1905,N_50);
nor U2108 (N_2108,N_1219,N_814);
nand U2109 (N_2109,N_651,N_286);
nor U2110 (N_2110,N_105,N_215);
nor U2111 (N_2111,N_1061,N_937);
and U2112 (N_2112,N_1036,N_855);
and U2113 (N_2113,N_1445,N_1430);
or U2114 (N_2114,N_1956,N_1117);
nor U2115 (N_2115,N_1709,N_729);
and U2116 (N_2116,N_1723,N_213);
and U2117 (N_2117,N_468,N_1434);
nor U2118 (N_2118,N_1127,N_662);
nor U2119 (N_2119,N_413,N_208);
nor U2120 (N_2120,N_891,N_1992);
or U2121 (N_2121,N_807,N_1996);
nand U2122 (N_2122,N_1534,N_604);
or U2123 (N_2123,N_199,N_1289);
nand U2124 (N_2124,N_587,N_216);
or U2125 (N_2125,N_1745,N_482);
nor U2126 (N_2126,N_1360,N_858);
and U2127 (N_2127,N_403,N_1401);
and U2128 (N_2128,N_1535,N_1713);
or U2129 (N_2129,N_813,N_843);
or U2130 (N_2130,N_930,N_859);
and U2131 (N_2131,N_761,N_675);
or U2132 (N_2132,N_725,N_571);
nand U2133 (N_2133,N_1249,N_1896);
nor U2134 (N_2134,N_1311,N_1392);
or U2135 (N_2135,N_884,N_682);
or U2136 (N_2136,N_477,N_320);
nand U2137 (N_2137,N_514,N_1624);
nor U2138 (N_2138,N_1684,N_1602);
and U2139 (N_2139,N_1362,N_1253);
or U2140 (N_2140,N_917,N_576);
nand U2141 (N_2141,N_1568,N_1070);
or U2142 (N_2142,N_1090,N_1096);
and U2143 (N_2143,N_1210,N_1622);
xor U2144 (N_2144,N_523,N_1776);
or U2145 (N_2145,N_185,N_552);
or U2146 (N_2146,N_1811,N_282);
nand U2147 (N_2147,N_267,N_258);
and U2148 (N_2148,N_635,N_22);
nand U2149 (N_2149,N_1890,N_841);
nand U2150 (N_2150,N_1443,N_1863);
nand U2151 (N_2151,N_619,N_1471);
and U2152 (N_2152,N_408,N_902);
xor U2153 (N_2153,N_1710,N_20);
nor U2154 (N_2154,N_1719,N_1231);
nand U2155 (N_2155,N_1722,N_302);
or U2156 (N_2156,N_1888,N_1928);
and U2157 (N_2157,N_580,N_585);
or U2158 (N_2158,N_1201,N_1742);
nand U2159 (N_2159,N_1094,N_1275);
and U2160 (N_2160,N_487,N_1529);
or U2161 (N_2161,N_54,N_61);
nand U2162 (N_2162,N_64,N_1118);
xnor U2163 (N_2163,N_1176,N_907);
nand U2164 (N_2164,N_612,N_1357);
and U2165 (N_2165,N_1769,N_935);
or U2166 (N_2166,N_693,N_1516);
nand U2167 (N_2167,N_1258,N_963);
or U2168 (N_2168,N_1151,N_1171);
or U2169 (N_2169,N_1240,N_1823);
or U2170 (N_2170,N_1423,N_1157);
nor U2171 (N_2171,N_1661,N_1730);
nor U2172 (N_2172,N_1807,N_1611);
or U2173 (N_2173,N_1121,N_285);
or U2174 (N_2174,N_1904,N_512);
and U2175 (N_2175,N_1462,N_1840);
nor U2176 (N_2176,N_1637,N_1490);
or U2177 (N_2177,N_1892,N_1921);
nor U2178 (N_2178,N_1854,N_1454);
nor U2179 (N_2179,N_1759,N_1660);
or U2180 (N_2180,N_1417,N_1869);
nor U2181 (N_2181,N_549,N_1919);
nor U2182 (N_2182,N_242,N_1803);
or U2183 (N_2183,N_789,N_1830);
nor U2184 (N_2184,N_335,N_1544);
or U2185 (N_2185,N_249,N_1626);
and U2186 (N_2186,N_89,N_1299);
nand U2187 (N_2187,N_850,N_1038);
nor U2188 (N_2188,N_655,N_1666);
nand U2189 (N_2189,N_1824,N_1025);
and U2190 (N_2190,N_1532,N_7);
and U2191 (N_2191,N_844,N_326);
nand U2192 (N_2192,N_1277,N_1778);
nor U2193 (N_2193,N_915,N_1266);
nand U2194 (N_2194,N_846,N_1328);
or U2195 (N_2195,N_357,N_531);
and U2196 (N_2196,N_1492,N_1594);
and U2197 (N_2197,N_36,N_1465);
or U2198 (N_2198,N_117,N_1796);
nor U2199 (N_2199,N_1877,N_735);
nand U2200 (N_2200,N_1139,N_457);
nand U2201 (N_2201,N_703,N_1994);
or U2202 (N_2202,N_1385,N_1741);
or U2203 (N_2203,N_909,N_296);
nand U2204 (N_2204,N_1172,N_1668);
nand U2205 (N_2205,N_1931,N_1676);
nor U2206 (N_2206,N_21,N_1882);
and U2207 (N_2207,N_1954,N_1558);
nand U2208 (N_2208,N_1788,N_69);
xor U2209 (N_2209,N_1271,N_892);
nor U2210 (N_2210,N_928,N_941);
and U2211 (N_2211,N_808,N_180);
and U2212 (N_2212,N_1567,N_1886);
nand U2213 (N_2213,N_1203,N_1174);
nand U2214 (N_2214,N_1031,N_23);
nand U2215 (N_2215,N_680,N_954);
nand U2216 (N_2216,N_704,N_889);
nor U2217 (N_2217,N_1899,N_225);
nor U2218 (N_2218,N_1609,N_1424);
nand U2219 (N_2219,N_1015,N_454);
nand U2220 (N_2220,N_484,N_1331);
nand U2221 (N_2221,N_1217,N_871);
nand U2222 (N_2222,N_1747,N_578);
and U2223 (N_2223,N_1893,N_256);
and U2224 (N_2224,N_284,N_1458);
and U2225 (N_2225,N_1297,N_1256);
nand U2226 (N_2226,N_1377,N_1003);
and U2227 (N_2227,N_1596,N_1555);
xor U2228 (N_2228,N_59,N_469);
nand U2229 (N_2229,N_205,N_607);
xor U2230 (N_2230,N_1026,N_33);
or U2231 (N_2231,N_1798,N_711);
and U2232 (N_2232,N_1683,N_1033);
and U2233 (N_2233,N_186,N_510);
nand U2234 (N_2234,N_1336,N_1756);
and U2235 (N_2235,N_986,N_1570);
nand U2236 (N_2236,N_1323,N_828);
and U2237 (N_2237,N_273,N_519);
and U2238 (N_2238,N_803,N_1418);
nor U2239 (N_2239,N_658,N_545);
nand U2240 (N_2240,N_300,N_622);
and U2241 (N_2241,N_1924,N_661);
nor U2242 (N_2242,N_1693,N_900);
nand U2243 (N_2243,N_110,N_847);
or U2244 (N_2244,N_82,N_1261);
and U2245 (N_2245,N_1585,N_573);
nand U2246 (N_2246,N_1734,N_1623);
nor U2247 (N_2247,N_1664,N_1589);
nor U2248 (N_2248,N_832,N_237);
or U2249 (N_2249,N_1575,N_1608);
nor U2250 (N_2250,N_241,N_1055);
nand U2251 (N_2251,N_627,N_885);
nor U2252 (N_2252,N_495,N_289);
nand U2253 (N_2253,N_348,N_13);
nand U2254 (N_2254,N_1832,N_1048);
nor U2255 (N_2255,N_1503,N_618);
or U2256 (N_2256,N_1346,N_43);
nand U2257 (N_2257,N_985,N_1629);
nor U2258 (N_2258,N_827,N_727);
and U2259 (N_2259,N_1313,N_1922);
nor U2260 (N_2260,N_1238,N_1826);
and U2261 (N_2261,N_598,N_1968);
and U2262 (N_2262,N_1505,N_85);
nand U2263 (N_2263,N_78,N_9);
nand U2264 (N_2264,N_1691,N_1089);
or U2265 (N_2265,N_1744,N_1366);
nor U2266 (N_2266,N_415,N_419);
and U2267 (N_2267,N_610,N_767);
and U2268 (N_2268,N_1519,N_1547);
xor U2269 (N_2269,N_203,N_1194);
nor U2270 (N_2270,N_564,N_904);
nand U2271 (N_2271,N_426,N_982);
nand U2272 (N_2272,N_1501,N_507);
xnor U2273 (N_2273,N_1002,N_380);
and U2274 (N_2274,N_1613,N_68);
and U2275 (N_2275,N_1718,N_1173);
and U2276 (N_2276,N_1461,N_116);
xor U2277 (N_2277,N_1175,N_1894);
nand U2278 (N_2278,N_1592,N_642);
nand U2279 (N_2279,N_467,N_1391);
or U2280 (N_2280,N_1239,N_453);
nor U2281 (N_2281,N_19,N_1694);
and U2282 (N_2282,N_1785,N_1775);
nand U2283 (N_2283,N_162,N_1670);
nand U2284 (N_2284,N_1810,N_1936);
nor U2285 (N_2285,N_765,N_1153);
nand U2286 (N_2286,N_1463,N_643);
nand U2287 (N_2287,N_364,N_833);
nand U2288 (N_2288,N_1967,N_210);
nor U2289 (N_2289,N_1935,N_1337);
nand U2290 (N_2290,N_1779,N_1696);
nor U2291 (N_2291,N_449,N_1053);
nand U2292 (N_2292,N_528,N_310);
nor U2293 (N_2293,N_1436,N_1278);
or U2294 (N_2294,N_1442,N_1034);
nand U2295 (N_2295,N_1560,N_166);
and U2296 (N_2296,N_1232,N_959);
nand U2297 (N_2297,N_243,N_1222);
nor U2298 (N_2298,N_1485,N_795);
or U2299 (N_2299,N_1847,N_1962);
nor U2300 (N_2300,N_992,N_483);
nor U2301 (N_2301,N_390,N_741);
nor U2302 (N_2302,N_971,N_41);
and U2303 (N_2303,N_40,N_471);
nor U2304 (N_2304,N_594,N_1342);
and U2305 (N_2305,N_772,N_1991);
nor U2306 (N_2306,N_951,N_1900);
or U2307 (N_2307,N_908,N_745);
or U2308 (N_2308,N_1557,N_1081);
or U2309 (N_2309,N_424,N_111);
nor U2310 (N_2310,N_1134,N_52);
nor U2311 (N_2311,N_31,N_718);
nand U2312 (N_2312,N_1563,N_1907);
nor U2313 (N_2313,N_169,N_107);
and U2314 (N_2314,N_1884,N_716);
or U2315 (N_2315,N_1791,N_1843);
or U2316 (N_2316,N_967,N_1164);
nor U2317 (N_2317,N_83,N_1000);
nor U2318 (N_2318,N_473,N_24);
and U2319 (N_2319,N_1552,N_1269);
or U2320 (N_2320,N_57,N_1595);
and U2321 (N_2321,N_151,N_1404);
nor U2322 (N_2322,N_821,N_268);
nor U2323 (N_2323,N_1829,N_639);
and U2324 (N_2324,N_1988,N_1444);
and U2325 (N_2325,N_1934,N_421);
and U2326 (N_2326,N_972,N_630);
or U2327 (N_2327,N_1448,N_640);
and U2328 (N_2328,N_438,N_1671);
or U2329 (N_2329,N_723,N_1517);
nor U2330 (N_2330,N_1335,N_125);
or U2331 (N_2331,N_479,N_918);
nand U2332 (N_2332,N_344,N_1695);
and U2333 (N_2333,N_1100,N_67);
nor U2334 (N_2334,N_266,N_906);
nand U2335 (N_2335,N_608,N_1380);
and U2336 (N_2336,N_1603,N_18);
and U2337 (N_2337,N_2,N_290);
nor U2338 (N_2338,N_1878,N_1280);
nand U2339 (N_2339,N_1341,N_1735);
nor U2340 (N_2340,N_161,N_93);
and U2341 (N_2341,N_773,N_1394);
nand U2342 (N_2342,N_897,N_1374);
or U2343 (N_2343,N_1196,N_669);
or U2344 (N_2344,N_739,N_339);
and U2345 (N_2345,N_155,N_647);
and U2346 (N_2346,N_1851,N_231);
nand U2347 (N_2347,N_1993,N_431);
or U2348 (N_2348,N_667,N_781);
or U2349 (N_2349,N_830,N_1506);
and U2350 (N_2350,N_1014,N_1553);
and U2351 (N_2351,N_1729,N_1112);
and U2352 (N_2352,N_1420,N_520);
and U2353 (N_2353,N_1581,N_1766);
nand U2354 (N_2354,N_1918,N_1494);
nand U2355 (N_2355,N_1059,N_371);
and U2356 (N_2356,N_502,N_880);
and U2357 (N_2357,N_204,N_657);
and U2358 (N_2358,N_574,N_572);
nor U2359 (N_2359,N_942,N_688);
nand U2360 (N_2360,N_1835,N_1211);
nand U2361 (N_2361,N_1431,N_1441);
or U2362 (N_2362,N_1065,N_1428);
or U2363 (N_2363,N_1144,N_1113);
or U2364 (N_2364,N_1937,N_776);
or U2365 (N_2365,N_566,N_1757);
nor U2366 (N_2366,N_626,N_1191);
nand U2367 (N_2367,N_428,N_1842);
nand U2368 (N_2368,N_1006,N_753);
nor U2369 (N_2369,N_613,N_804);
nand U2370 (N_2370,N_197,N_695);
nand U2371 (N_2371,N_1912,N_958);
or U2372 (N_2372,N_1214,N_899);
or U2373 (N_2373,N_25,N_317);
nor U2374 (N_2374,N_1680,N_389);
or U2375 (N_2375,N_1022,N_10);
nand U2376 (N_2376,N_236,N_229);
nand U2377 (N_2377,N_1600,N_226);
or U2378 (N_2378,N_1062,N_313);
nor U2379 (N_2379,N_177,N_391);
or U2380 (N_2380,N_383,N_1057);
nor U2381 (N_2381,N_250,N_1643);
nand U2382 (N_2382,N_363,N_1264);
nor U2383 (N_2383,N_1287,N_715);
nor U2384 (N_2384,N_679,N_1288);
nor U2385 (N_2385,N_876,N_337);
nor U2386 (N_2386,N_1049,N_1263);
nand U2387 (N_2387,N_1260,N_1860);
nor U2388 (N_2388,N_1507,N_1774);
nor U2389 (N_2389,N_80,N_1760);
nand U2390 (N_2390,N_1982,N_1977);
or U2391 (N_2391,N_1412,N_783);
and U2392 (N_2392,N_271,N_377);
nor U2393 (N_2393,N_1833,N_1107);
or U2394 (N_2394,N_55,N_748);
nor U2395 (N_2395,N_713,N_374);
nand U2396 (N_2396,N_913,N_1001);
or U2397 (N_2397,N_890,N_198);
nor U2398 (N_2398,N_112,N_1724);
or U2399 (N_2399,N_1284,N_1591);
nor U2400 (N_2400,N_121,N_559);
or U2401 (N_2401,N_402,N_1765);
nor U2402 (N_2402,N_1523,N_623);
nor U2403 (N_2403,N_700,N_706);
nor U2404 (N_2404,N_1702,N_346);
or U2405 (N_2405,N_815,N_1242);
nor U2406 (N_2406,N_497,N_1016);
nor U2407 (N_2407,N_1512,N_1819);
or U2408 (N_2408,N_590,N_35);
nor U2409 (N_2409,N_276,N_1911);
nand U2410 (N_2410,N_966,N_367);
or U2411 (N_2411,N_1920,N_1572);
nor U2412 (N_2412,N_816,N_1812);
nor U2413 (N_2413,N_1123,N_1302);
nand U2414 (N_2414,N_755,N_1244);
nand U2415 (N_2415,N_1616,N_1493);
nand U2416 (N_2416,N_146,N_1453);
nand U2417 (N_2417,N_631,N_1158);
or U2418 (N_2418,N_222,N_1700);
and U2419 (N_2419,N_98,N_1136);
nor U2420 (N_2420,N_1262,N_1584);
nor U2421 (N_2421,N_1971,N_1421);
nand U2422 (N_2422,N_997,N_1981);
nor U2423 (N_2423,N_820,N_1446);
nor U2424 (N_2424,N_1129,N_1915);
nand U2425 (N_2425,N_131,N_163);
and U2426 (N_2426,N_1133,N_746);
and U2427 (N_2427,N_1698,N_1020);
nor U2428 (N_2428,N_94,N_616);
nand U2429 (N_2429,N_397,N_600);
and U2430 (N_2430,N_1849,N_1372);
or U2431 (N_2431,N_1874,N_425);
nand U2432 (N_2432,N_1780,N_947);
nand U2433 (N_2433,N_1768,N_257);
nor U2434 (N_2434,N_584,N_235);
and U2435 (N_2435,N_1043,N_934);
nor U2436 (N_2436,N_702,N_220);
nor U2437 (N_2437,N_304,N_165);
nand U2438 (N_2438,N_851,N_309);
nand U2439 (N_2439,N_565,N_1538);
and U2440 (N_2440,N_1390,N_674);
nand U2441 (N_2441,N_933,N_1793);
or U2442 (N_2442,N_1880,N_866);
and U2443 (N_2443,N_356,N_318);
nor U2444 (N_2444,N_1195,N_1944);
nand U2445 (N_2445,N_1711,N_1598);
nor U2446 (N_2446,N_1571,N_148);
or U2447 (N_2447,N_925,N_534);
xnor U2448 (N_2448,N_614,N_228);
nor U2449 (N_2449,N_677,N_1871);
nor U2450 (N_2450,N_1228,N_1947);
xnor U2451 (N_2451,N_1743,N_1838);
nor U2452 (N_2452,N_114,N_1303);
or U2453 (N_2453,N_1304,N_0);
or U2454 (N_2454,N_232,N_1853);
nand U2455 (N_2455,N_1010,N_1483);
nor U2456 (N_2456,N_777,N_1983);
or U2457 (N_2457,N_38,N_379);
nor U2458 (N_2458,N_1455,N_684);
or U2459 (N_2459,N_1942,N_911);
nand U2460 (N_2460,N_609,N_331);
nor U2461 (N_2461,N_1035,N_824);
nand U2462 (N_2462,N_707,N_1028);
or U2463 (N_2463,N_244,N_1086);
or U2464 (N_2464,N_1524,N_1495);
or U2465 (N_2465,N_599,N_879);
or U2466 (N_2466,N_621,N_752);
nand U2467 (N_2467,N_1187,N_888);
nand U2468 (N_2468,N_1764,N_536);
and U2469 (N_2469,N_156,N_1150);
xor U2470 (N_2470,N_1042,N_1511);
nand U2471 (N_2471,N_1732,N_1577);
nor U2472 (N_2472,N_1949,N_784);
or U2473 (N_2473,N_1386,N_1040);
nand U2474 (N_2474,N_485,N_810);
nor U2475 (N_2475,N_1641,N_1872);
xor U2476 (N_2476,N_1677,N_961);
or U2477 (N_2477,N_200,N_1396);
and U2478 (N_2478,N_515,N_1097);
nand U2479 (N_2479,N_664,N_1640);
nor U2480 (N_2480,N_1340,N_406);
xnor U2481 (N_2481,N_1748,N_1074);
and U2482 (N_2482,N_6,N_1475);
and U2483 (N_2483,N_295,N_589);
or U2484 (N_2484,N_1814,N_691);
or U2485 (N_2485,N_1126,N_1143);
or U2486 (N_2486,N_262,N_1104);
nor U2487 (N_2487,N_1013,N_964);
or U2488 (N_2488,N_56,N_1241);
and U2489 (N_2489,N_385,N_1200);
and U2490 (N_2490,N_894,N_217);
and U2491 (N_2491,N_1792,N_582);
or U2492 (N_2492,N_509,N_1697);
nand U2493 (N_2493,N_886,N_100);
and U2494 (N_2494,N_1039,N_1951);
nand U2495 (N_2495,N_1607,N_351);
nor U2496 (N_2496,N_251,N_1576);
nor U2497 (N_2497,N_145,N_1687);
or U2498 (N_2498,N_362,N_1083);
and U2499 (N_2499,N_1497,N_1085);
and U2500 (N_2500,N_831,N_1654);
nor U2501 (N_2501,N_375,N_17);
or U2502 (N_2502,N_76,N_355);
or U2503 (N_2503,N_1052,N_1908);
or U2504 (N_2504,N_940,N_1116);
xnor U2505 (N_2505,N_922,N_901);
nand U2506 (N_2506,N_1283,N_1408);
nand U2507 (N_2507,N_1375,N_212);
and U2508 (N_2508,N_1891,N_179);
or U2509 (N_2509,N_799,N_387);
nor U2510 (N_2510,N_1138,N_999);
and U2511 (N_2511,N_504,N_1397);
or U2512 (N_2512,N_1966,N_595);
or U2513 (N_2513,N_1474,N_1559);
nor U2514 (N_2514,N_1681,N_292);
nor U2515 (N_2515,N_697,N_921);
or U2516 (N_2516,N_491,N_868);
nor U2517 (N_2517,N_1004,N_1353);
or U2518 (N_2518,N_910,N_400);
or U2519 (N_2519,N_1276,N_1008);
and U2520 (N_2520,N_350,N_1076);
or U2521 (N_2521,N_1789,N_567);
nand U2522 (N_2522,N_1355,N_1573);
or U2523 (N_2523,N_1801,N_919);
and U2524 (N_2524,N_1636,N_439);
or U2525 (N_2525,N_157,N_460);
or U2526 (N_2526,N_26,N_1630);
nor U2527 (N_2527,N_568,N_1881);
nor U2528 (N_2528,N_1978,N_1468);
and U2529 (N_2529,N_75,N_1566);
nor U2530 (N_2530,N_188,N_1805);
and U2531 (N_2531,N_993,N_129);
xor U2532 (N_2532,N_1975,N_1405);
or U2533 (N_2533,N_517,N_762);
nor U2534 (N_2534,N_322,N_1834);
xor U2535 (N_2535,N_882,N_1958);
or U2536 (N_2536,N_1656,N_341);
and U2537 (N_2537,N_1378,N_1673);
or U2538 (N_2538,N_1041,N_319);
or U2539 (N_2539,N_1317,N_1605);
nor U2540 (N_2540,N_628,N_1989);
or U2541 (N_2541,N_1128,N_1345);
nor U2542 (N_2542,N_1322,N_1338);
nor U2543 (N_2543,N_405,N_903);
nand U2544 (N_2544,N_793,N_1618);
nor U2545 (N_2545,N_686,N_560);
and U2546 (N_2546,N_223,N_423);
nand U2547 (N_2547,N_275,N_1601);
nand U2548 (N_2548,N_1952,N_1389);
or U2549 (N_2549,N_1850,N_1790);
or U2550 (N_2550,N_1343,N_524);
nor U2551 (N_2551,N_106,N_692);
nor U2552 (N_2552,N_174,N_291);
and U2553 (N_2553,N_780,N_108);
and U2554 (N_2554,N_1190,N_175);
nand U2555 (N_2555,N_314,N_1450);
nand U2556 (N_2556,N_731,N_1103);
nor U2557 (N_2557,N_1098,N_645);
nor U2558 (N_2558,N_343,N_1970);
nand U2559 (N_2559,N_332,N_1165);
nor U2560 (N_2560,N_1247,N_1252);
nor U2561 (N_2561,N_1739,N_1530);
nand U2562 (N_2562,N_1073,N_1692);
nor U2563 (N_2563,N_1225,N_412);
and U2564 (N_2564,N_838,N_893);
or U2565 (N_2565,N_119,N_872);
nor U2566 (N_2566,N_689,N_823);
nand U2567 (N_2567,N_150,N_214);
nand U2568 (N_2568,N_1914,N_1662);
or U2569 (N_2569,N_240,N_511);
and U2570 (N_2570,N_29,N_287);
nor U2571 (N_2571,N_411,N_983);
or U2572 (N_2572,N_1146,N_74);
xor U2573 (N_2573,N_15,N_1310);
and U2574 (N_2574,N_556,N_1120);
or U2575 (N_2575,N_1706,N_1815);
nor U2576 (N_2576,N_1079,N_812);
and U2577 (N_2577,N_916,N_1679);
or U2578 (N_2578,N_1370,N_1686);
nand U2579 (N_2579,N_51,N_605);
and U2580 (N_2580,N_260,N_714);
nand U2581 (N_2581,N_142,N_1185);
nor U2582 (N_2582,N_171,N_1108);
nor U2583 (N_2583,N_1046,N_1883);
nor U2584 (N_2584,N_1906,N_167);
nand U2585 (N_2585,N_446,N_648);
and U2586 (N_2586,N_278,N_1844);
nor U2587 (N_2587,N_1699,N_386);
and U2588 (N_2588,N_1344,N_786);
xnor U2589 (N_2589,N_1439,N_508);
nor U2590 (N_2590,N_297,N_340);
and U2591 (N_2591,N_1876,N_1562);
or U2592 (N_2592,N_283,N_817);
and U2593 (N_2593,N_70,N_1498);
or U2594 (N_2594,N_139,N_463);
nor U2595 (N_2595,N_1369,N_96);
nand U2596 (N_2596,N_1499,N_1180);
and U2597 (N_2597,N_1582,N_1549);
nor U2598 (N_2598,N_1419,N_481);
and U2599 (N_2599,N_1767,N_717);
nor U2600 (N_2600,N_737,N_1950);
nor U2601 (N_2601,N_603,N_1314);
nand U2602 (N_2602,N_541,N_1761);
nand U2603 (N_2603,N_395,N_569);
nand U2604 (N_2604,N_1142,N_1440);
nand U2605 (N_2605,N_666,N_1227);
or U2606 (N_2606,N_448,N_856);
or U2607 (N_2607,N_293,N_611);
nand U2608 (N_2608,N_1334,N_1738);
or U2609 (N_2609,N_128,N_1324);
nand U2610 (N_2610,N_37,N_615);
nand U2611 (N_2611,N_670,N_1644);
or U2612 (N_2612,N_1148,N_1029);
nor U2613 (N_2613,N_499,N_1590);
nor U2614 (N_2614,N_1192,N_365);
and U2615 (N_2615,N_1459,N_1379);
or U2616 (N_2616,N_1943,N_771);
or U2617 (N_2617,N_1099,N_624);
nand U2618 (N_2618,N_1,N_253);
or U2619 (N_2619,N_1845,N_1868);
nor U2620 (N_2620,N_989,N_1773);
nand U2621 (N_2621,N_521,N_1333);
and U2622 (N_2622,N_1414,N_730);
and U2623 (N_2623,N_1867,N_548);
and U2624 (N_2624,N_1312,N_3);
nand U2625 (N_2625,N_981,N_1298);
and U2626 (N_2626,N_1526,N_533);
nor U2627 (N_2627,N_1327,N_1543);
and U2628 (N_2628,N_738,N_97);
nand U2629 (N_2629,N_988,N_1207);
nor U2630 (N_2630,N_1783,N_1437);
nand U2631 (N_2631,N_660,N_1758);
nand U2632 (N_2632,N_867,N_77);
and U2633 (N_2633,N_766,N_1728);
nor U2634 (N_2634,N_757,N_53);
and U2635 (N_2635,N_1995,N_1184);
or U2636 (N_2636,N_58,N_505);
nand U2637 (N_2637,N_136,N_414);
and U2638 (N_2638,N_1368,N_800);
nor U2639 (N_2639,N_1999,N_1725);
and U2640 (N_2640,N_1198,N_294);
nand U2641 (N_2641,N_1018,N_836);
and U2642 (N_2642,N_806,N_501);
nor U2643 (N_2643,N_1182,N_1998);
nor U2644 (N_2644,N_345,N_123);
or U2645 (N_2645,N_1124,N_11);
or U2646 (N_2646,N_802,N_1583);
nand U2647 (N_2647,N_976,N_538);
nand U2648 (N_2648,N_796,N_724);
nor U2649 (N_2649,N_71,N_1321);
nand U2650 (N_2650,N_349,N_1510);
and U2651 (N_2651,N_1023,N_1479);
or U2652 (N_2652,N_1235,N_1243);
nor U2653 (N_2653,N_732,N_1657);
nand U2654 (N_2654,N_382,N_79);
or U2655 (N_2655,N_1806,N_30);
nand U2656 (N_2656,N_1901,N_14);
or U2657 (N_2657,N_466,N_1813);
or U2658 (N_2658,N_1985,N_396);
nor U2659 (N_2659,N_1750,N_393);
nor U2660 (N_2660,N_1752,N_1940);
nor U2661 (N_2661,N_333,N_881);
or U2662 (N_2662,N_822,N_943);
nor U2663 (N_2663,N_1075,N_979);
nand U2664 (N_2664,N_1804,N_912);
nand U2665 (N_2665,N_1068,N_433);
nor U2666 (N_2666,N_849,N_1072);
or U2667 (N_2667,N_592,N_422);
xor U2668 (N_2668,N_1205,N_863);
nor U2669 (N_2669,N_1827,N_1383);
nand U2670 (N_2670,N_1407,N_1737);
nor U2671 (N_2671,N_955,N_1902);
or U2672 (N_2672,N_1929,N_1326);
nor U2673 (N_2673,N_329,N_539);
and U2674 (N_2674,N_1859,N_1716);
nor U2675 (N_2675,N_1101,N_744);
and U2676 (N_2676,N_1216,N_368);
nand U2677 (N_2677,N_1248,N_1452);
or U2678 (N_2678,N_1208,N_8);
and U2679 (N_2679,N_1223,N_1204);
nor U2680 (N_2680,N_829,N_646);
nand U2681 (N_2681,N_1093,N_671);
and U2682 (N_2682,N_1839,N_378);
and U2683 (N_2683,N_221,N_629);
nand U2684 (N_2684,N_1141,N_769);
nand U2685 (N_2685,N_1220,N_1653);
nor U2686 (N_2686,N_1236,N_1647);
and U2687 (N_2687,N_436,N_1820);
nor U2688 (N_2688,N_65,N_1554);
nand U2689 (N_2689,N_1786,N_1580);
or U2690 (N_2690,N_1361,N_798);
nor U2691 (N_2691,N_1167,N_944);
and U2692 (N_2692,N_183,N_1363);
and U2693 (N_2693,N_1371,N_1525);
and U2694 (N_2694,N_338,N_372);
nand U2695 (N_2695,N_1669,N_1749);
nand U2696 (N_2696,N_1864,N_550);
and U2697 (N_2697,N_407,N_496);
and U2698 (N_2698,N_1447,N_211);
nand U2699 (N_2699,N_1413,N_659);
nand U2700 (N_2700,N_176,N_1169);
or U2701 (N_2701,N_269,N_493);
nor U2702 (N_2702,N_591,N_654);
and U2703 (N_2703,N_977,N_1193);
or U2704 (N_2704,N_1690,N_537);
nand U2705 (N_2705,N_1712,N_547);
or U2706 (N_2706,N_1787,N_853);
and U2707 (N_2707,N_1044,N_949);
and U2708 (N_2708,N_1808,N_1084);
nand U2709 (N_2709,N_722,N_1655);
and U2710 (N_2710,N_409,N_1606);
or U2711 (N_2711,N_472,N_1651);
nor U2712 (N_2712,N_1578,N_962);
or U2713 (N_2713,N_1426,N_1715);
and U2714 (N_2714,N_561,N_1301);
xnor U2715 (N_2715,N_984,N_1916);
or U2716 (N_2716,N_1848,N_736);
nand U2717 (N_2717,N_579,N_299);
nand U2718 (N_2718,N_1376,N_498);
nand U2719 (N_2719,N_486,N_1125);
nand U2720 (N_2720,N_1561,N_1147);
xnor U2721 (N_2721,N_1011,N_1183);
or U2722 (N_2722,N_869,N_1586);
or U2723 (N_2723,N_1800,N_62);
nand U2724 (N_2724,N_87,N_1621);
or U2725 (N_2725,N_998,N_91);
nand U2726 (N_2726,N_1109,N_1938);
or U2727 (N_2727,N_1588,N_1533);
and U2728 (N_2728,N_1481,N_398);
or U2729 (N_2729,N_201,N_1754);
or U2730 (N_2730,N_1753,N_1166);
and U2731 (N_2731,N_540,N_392);
nor U2732 (N_2732,N_245,N_1469);
nor U2733 (N_2733,N_39,N_756);
nor U2734 (N_2734,N_1926,N_870);
nor U2735 (N_2735,N_1347,N_369);
or U2736 (N_2736,N_1504,N_1162);
nor U2737 (N_2737,N_932,N_681);
nor U2738 (N_2738,N_1794,N_1202);
or U2739 (N_2739,N_1961,N_1186);
nor U2740 (N_2740,N_779,N_342);
and U2741 (N_2741,N_1429,N_219);
and U2742 (N_2742,N_1212,N_1619);
nor U2743 (N_2743,N_1945,N_754);
or U2744 (N_2744,N_1358,N_1189);
and U2745 (N_2745,N_1156,N_327);
and U2746 (N_2746,N_172,N_1870);
nor U2747 (N_2747,N_733,N_1470);
nand U2748 (N_2748,N_1122,N_705);
or U2749 (N_2749,N_430,N_1259);
nor U2750 (N_2750,N_848,N_46);
nand U2751 (N_2751,N_159,N_750);
or U2752 (N_2752,N_1009,N_152);
and U2753 (N_2753,N_1484,N_742);
or U2754 (N_2754,N_303,N_401);
nor U2755 (N_2755,N_854,N_842);
or U2756 (N_2756,N_1852,N_158);
or U2757 (N_2757,N_1221,N_1473);
or U2758 (N_2758,N_1646,N_1110);
and U2759 (N_2759,N_370,N_434);
and U2760 (N_2760,N_676,N_1137);
nor U2761 (N_2761,N_1887,N_95);
nand U2762 (N_2762,N_1351,N_1050);
and U2763 (N_2763,N_527,N_826);
and U2764 (N_2764,N_1027,N_1650);
nor U2765 (N_2765,N_1037,N_288);
or U2766 (N_2766,N_265,N_160);
nand U2767 (N_2767,N_1960,N_759);
and U2768 (N_2768,N_1703,N_1416);
xor U2769 (N_2769,N_443,N_770);
nor U2770 (N_2770,N_334,N_252);
nor U2771 (N_2771,N_1933,N_1224);
and U2772 (N_2772,N_575,N_248);
and U2773 (N_2773,N_878,N_1197);
nand U2774 (N_2774,N_373,N_140);
nand U2775 (N_2775,N_1054,N_494);
nand U2776 (N_2776,N_1542,N_1460);
or U2777 (N_2777,N_553,N_1527);
nor U2778 (N_2778,N_1620,N_135);
nand U2779 (N_2779,N_557,N_641);
and U2780 (N_2780,N_124,N_877);
nand U2781 (N_2781,N_281,N_1045);
nor U2782 (N_2782,N_1135,N_1610);
and U2783 (N_2783,N_835,N_1145);
nor U2784 (N_2784,N_1069,N_127);
and U2785 (N_2785,N_49,N_1763);
nand U2786 (N_2786,N_1154,N_1751);
nor U2787 (N_2787,N_1858,N_1476);
nand U2788 (N_2788,N_1293,N_873);
and U2789 (N_2789,N_1502,N_1930);
or U2790 (N_2790,N_694,N_435);
or U2791 (N_2791,N_42,N_1398);
or U2792 (N_2792,N_1319,N_324);
nor U2793 (N_2793,N_360,N_1837);
or U2794 (N_2794,N_1903,N_1895);
or U2795 (N_2795,N_805,N_323);
xnor U2796 (N_2796,N_1356,N_184);
or U2797 (N_2797,N_99,N_506);
or U2798 (N_2798,N_945,N_404);
or U2799 (N_2799,N_489,N_388);
and U2800 (N_2800,N_1078,N_1012);
and U2801 (N_2801,N_312,N_513);
and U2802 (N_2802,N_1403,N_190);
nand U2803 (N_2803,N_1665,N_1705);
or U2804 (N_2804,N_1946,N_518);
and U2805 (N_2805,N_1170,N_476);
nor U2806 (N_2806,N_1548,N_526);
or U2807 (N_2807,N_459,N_347);
and U2808 (N_2808,N_542,N_1330);
nand U2809 (N_2809,N_1972,N_924);
and U2810 (N_2810,N_1736,N_1255);
nor U2811 (N_2811,N_134,N_1449);
nand U2812 (N_2812,N_1986,N_532);
nand U2813 (N_2813,N_410,N_182);
and U2814 (N_2814,N_1500,N_583);
xor U2815 (N_2815,N_1913,N_929);
nor U2816 (N_2816,N_1818,N_113);
nand U2817 (N_2817,N_1152,N_923);
nor U2818 (N_2818,N_88,N_801);
nand U2819 (N_2819,N_45,N_1997);
nor U2820 (N_2820,N_743,N_1564);
and U2821 (N_2821,N_1451,N_683);
nand U2822 (N_2822,N_1140,N_687);
and U2823 (N_2823,N_1708,N_1315);
and U2824 (N_2824,N_209,N_792);
nor U2825 (N_2825,N_1866,N_562);
and U2826 (N_2826,N_874,N_1973);
or U2827 (N_2827,N_1491,N_366);
xor U2828 (N_2828,N_1393,N_1415);
nand U2829 (N_2829,N_1733,N_818);
nor U2830 (N_2830,N_1087,N_1409);
nand U2831 (N_2831,N_1438,N_1721);
nand U2832 (N_2832,N_455,N_1019);
or U2833 (N_2833,N_794,N_840);
nand U2834 (N_2834,N_270,N_1536);
nand U2835 (N_2835,N_1082,N_563);
and U2836 (N_2836,N_1987,N_763);
nand U2837 (N_2837,N_751,N_865);
nor U2838 (N_2838,N_1066,N_996);
or U2839 (N_2839,N_27,N_137);
or U2840 (N_2840,N_1714,N_144);
nor U2841 (N_2841,N_1726,N_126);
nor U2842 (N_2842,N_461,N_778);
and U2843 (N_2843,N_1667,N_1467);
nand U2844 (N_2844,N_652,N_721);
or U2845 (N_2845,N_417,N_168);
and U2846 (N_2846,N_1349,N_1846);
and U2847 (N_2847,N_450,N_1325);
or U2848 (N_2848,N_1740,N_740);
and U2849 (N_2849,N_72,N_44);
or U2850 (N_2850,N_1701,N_1528);
nor U2851 (N_2851,N_305,N_1115);
nor U2852 (N_2852,N_1625,N_862);
or U2853 (N_2853,N_1974,N_1831);
and U2854 (N_2854,N_376,N_994);
nand U2855 (N_2855,N_1294,N_187);
and U2856 (N_2856,N_1267,N_1206);
nand U2857 (N_2857,N_447,N_701);
and U2858 (N_2858,N_321,N_1574);
nor U2859 (N_2859,N_939,N_1828);
and U2860 (N_2860,N_875,N_926);
or U2861 (N_2861,N_1400,N_1522);
nor U2862 (N_2862,N_1433,N_102);
nor U2863 (N_2863,N_1550,N_427);
nand U2864 (N_2864,N_1290,N_699);
nor U2865 (N_2865,N_1348,N_490);
nand U2866 (N_2866,N_1318,N_837);
nand U2867 (N_2867,N_1237,N_720);
nor U2868 (N_2868,N_359,N_1457);
and U2869 (N_2869,N_1367,N_1546);
and U2870 (N_2870,N_90,N_825);
nand U2871 (N_2871,N_1265,N_597);
nor U2872 (N_2872,N_1674,N_690);
nand U2873 (N_2873,N_1159,N_1897);
nor U2874 (N_2874,N_1279,N_845);
or U2875 (N_2875,N_1635,N_1422);
and U2876 (N_2876,N_1273,N_788);
or U2877 (N_2877,N_1797,N_719);
nand U2878 (N_2878,N_103,N_602);
or U2879 (N_2879,N_970,N_546);
or U2880 (N_2880,N_1631,N_254);
and U2881 (N_2881,N_1817,N_358);
or U2882 (N_2882,N_32,N_1063);
nand U2883 (N_2883,N_441,N_726);
nor U2884 (N_2884,N_544,N_247);
nor U2885 (N_2885,N_1181,N_474);
nand U2886 (N_2886,N_1285,N_1809);
nor U2887 (N_2887,N_965,N_1411);
and U2888 (N_2888,N_1292,N_672);
nand U2889 (N_2889,N_653,N_577);
or U2890 (N_2890,N_451,N_440);
nand U2891 (N_2891,N_1770,N_1642);
nor U2892 (N_2892,N_277,N_118);
and U2893 (N_2893,N_1875,N_1274);
nor U2894 (N_2894,N_775,N_1784);
or U2895 (N_2895,N_1352,N_668);
nand U2896 (N_2896,N_1531,N_797);
or U2897 (N_2897,N_1105,N_1339);
and U2898 (N_2898,N_207,N_1628);
and U2899 (N_2899,N_429,N_133);
and U2900 (N_2900,N_149,N_978);
nand U2901 (N_2901,N_1717,N_475);
nand U2902 (N_2902,N_224,N_1939);
or U2903 (N_2903,N_1387,N_956);
nor U2904 (N_2904,N_1515,N_1927);
and U2905 (N_2905,N_280,N_1755);
nor U2906 (N_2906,N_1898,N_1980);
and U2907 (N_2907,N_768,N_1861);
and U2908 (N_2908,N_361,N_1291);
nand U2909 (N_2909,N_109,N_1799);
nand U2910 (N_2910,N_1177,N_678);
or U2911 (N_2911,N_1199,N_1917);
nor U2912 (N_2912,N_154,N_905);
and U2913 (N_2913,N_1569,N_1762);
or U2914 (N_2914,N_1638,N_1091);
nor U2915 (N_2915,N_1095,N_852);
nand U2916 (N_2916,N_48,N_883);
and U2917 (N_2917,N_143,N_685);
and U2918 (N_2918,N_120,N_233);
xor U2919 (N_2919,N_445,N_1645);
nand U2920 (N_2920,N_1088,N_1965);
and U2921 (N_2921,N_588,N_458);
nor U2922 (N_2922,N_444,N_1604);
nor U2923 (N_2923,N_696,N_1092);
or U2924 (N_2924,N_1777,N_1406);
nor U2925 (N_2925,N_418,N_570);
or U2926 (N_2926,N_1979,N_1281);
nand U2927 (N_2927,N_92,N_500);
nor U2928 (N_2928,N_452,N_1486);
or U2929 (N_2929,N_1058,N_1307);
and U2930 (N_2930,N_638,N_665);
nor U2931 (N_2931,N_1354,N_620);
nand U2932 (N_2932,N_170,N_1857);
nand U2933 (N_2933,N_1727,N_1955);
nand U2934 (N_2934,N_1909,N_1959);
and U2935 (N_2935,N_791,N_238);
nand U2936 (N_2936,N_274,N_1821);
and U2937 (N_2937,N_1226,N_16);
and U2938 (N_2938,N_1254,N_1296);
nand U2939 (N_2939,N_1306,N_178);
or U2940 (N_2940,N_1782,N_1963);
nor U2941 (N_2941,N_1131,N_1615);
nand U2942 (N_2942,N_354,N_1482);
nand U2943 (N_2943,N_1432,N_1593);
nor U2944 (N_2944,N_1282,N_1373);
and U2945 (N_2945,N_1114,N_1513);
and U2946 (N_2946,N_787,N_1675);
nor U2947 (N_2947,N_1508,N_606);
or U2948 (N_2948,N_153,N_516);
nor U2949 (N_2949,N_927,N_66);
nand U2950 (N_2950,N_1466,N_861);
and U2951 (N_2951,N_1599,N_246);
nor U2952 (N_2952,N_758,N_122);
nor U2953 (N_2953,N_442,N_1659);
or U2954 (N_2954,N_634,N_104);
and U2955 (N_2955,N_1032,N_1879);
or U2956 (N_2956,N_1772,N_1245);
nand U2957 (N_2957,N_973,N_399);
nand U2958 (N_2958,N_1836,N_1976);
nand U2959 (N_2959,N_1168,N_132);
nor U2960 (N_2960,N_1251,N_1731);
nor U2961 (N_2961,N_381,N_1410);
nor U2962 (N_2962,N_950,N_1678);
and U2963 (N_2963,N_864,N_465);
nor U2964 (N_2964,N_1056,N_394);
nor U2965 (N_2965,N_1856,N_1270);
nor U2966 (N_2966,N_1161,N_895);
or U2967 (N_2967,N_633,N_991);
nor U2968 (N_2968,N_887,N_1402);
nor U2969 (N_2969,N_1179,N_1841);
nor U2970 (N_2970,N_1496,N_636);
and U2971 (N_2971,N_1617,N_1658);
nor U2972 (N_2972,N_1969,N_353);
or U2973 (N_2973,N_522,N_1964);
nor U2974 (N_2974,N_1230,N_1024);
and U2975 (N_2975,N_1825,N_1957);
nand U2976 (N_2976,N_1106,N_1132);
or U2977 (N_2977,N_1587,N_1218);
and U2978 (N_2978,N_1111,N_650);
and U2979 (N_2979,N_1464,N_1130);
nor U2980 (N_2980,N_1047,N_1077);
nor U2981 (N_2981,N_173,N_1649);
or U2982 (N_2982,N_1102,N_1565);
nor U2983 (N_2983,N_1855,N_529);
or U2984 (N_2984,N_1514,N_1518);
or U2985 (N_2985,N_86,N_1268);
and U2986 (N_2986,N_261,N_1021);
nand U2987 (N_2987,N_1862,N_1229);
and U2988 (N_2988,N_1155,N_1427);
nand U2989 (N_2989,N_975,N_712);
xnor U2990 (N_2990,N_1652,N_1685);
nor U2991 (N_2991,N_1925,N_130);
nor U2992 (N_2992,N_920,N_953);
nand U2993 (N_2993,N_1489,N_663);
and U2994 (N_2994,N_1707,N_202);
and U2995 (N_2995,N_1478,N_708);
nor U2996 (N_2996,N_952,N_1246);
nand U2997 (N_2997,N_1520,N_1178);
and U2998 (N_2998,N_785,N_1395);
nor U2999 (N_2999,N_194,N_617);
nand U3000 (N_3000,N_887,N_1567);
or U3001 (N_3001,N_1469,N_541);
or U3002 (N_3002,N_1156,N_1434);
nor U3003 (N_3003,N_878,N_827);
and U3004 (N_3004,N_880,N_1477);
nor U3005 (N_3005,N_1225,N_1415);
nor U3006 (N_3006,N_1502,N_1396);
nand U3007 (N_3007,N_1659,N_1163);
and U3008 (N_3008,N_1470,N_1578);
nor U3009 (N_3009,N_684,N_1805);
nand U3010 (N_3010,N_1131,N_61);
or U3011 (N_3011,N_1446,N_325);
or U3012 (N_3012,N_71,N_1468);
nor U3013 (N_3013,N_359,N_662);
or U3014 (N_3014,N_249,N_1082);
and U3015 (N_3015,N_1707,N_1823);
xnor U3016 (N_3016,N_1566,N_1728);
or U3017 (N_3017,N_1784,N_1805);
nor U3018 (N_3018,N_479,N_1991);
nand U3019 (N_3019,N_1214,N_830);
or U3020 (N_3020,N_972,N_1087);
or U3021 (N_3021,N_1168,N_257);
or U3022 (N_3022,N_1494,N_107);
nor U3023 (N_3023,N_1224,N_1009);
nor U3024 (N_3024,N_295,N_505);
or U3025 (N_3025,N_948,N_1099);
or U3026 (N_3026,N_705,N_1751);
xor U3027 (N_3027,N_1561,N_649);
and U3028 (N_3028,N_1446,N_297);
xnor U3029 (N_3029,N_1479,N_978);
nor U3030 (N_3030,N_1666,N_1250);
and U3031 (N_3031,N_1320,N_924);
and U3032 (N_3032,N_849,N_1198);
nand U3033 (N_3033,N_172,N_792);
xnor U3034 (N_3034,N_680,N_1747);
nor U3035 (N_3035,N_1961,N_545);
nor U3036 (N_3036,N_27,N_1458);
or U3037 (N_3037,N_308,N_686);
or U3038 (N_3038,N_1952,N_78);
nand U3039 (N_3039,N_1991,N_342);
and U3040 (N_3040,N_1771,N_1019);
nor U3041 (N_3041,N_779,N_329);
nand U3042 (N_3042,N_1316,N_1975);
nor U3043 (N_3043,N_267,N_802);
nor U3044 (N_3044,N_414,N_383);
or U3045 (N_3045,N_672,N_424);
or U3046 (N_3046,N_576,N_1014);
or U3047 (N_3047,N_1463,N_1007);
nand U3048 (N_3048,N_82,N_1783);
nor U3049 (N_3049,N_797,N_96);
and U3050 (N_3050,N_987,N_1612);
or U3051 (N_3051,N_56,N_186);
or U3052 (N_3052,N_1579,N_1042);
and U3053 (N_3053,N_1109,N_120);
and U3054 (N_3054,N_1245,N_1384);
nor U3055 (N_3055,N_599,N_1012);
nor U3056 (N_3056,N_1226,N_744);
or U3057 (N_3057,N_1228,N_966);
nand U3058 (N_3058,N_210,N_208);
and U3059 (N_3059,N_1694,N_1613);
nand U3060 (N_3060,N_723,N_952);
and U3061 (N_3061,N_473,N_1713);
and U3062 (N_3062,N_1418,N_143);
or U3063 (N_3063,N_670,N_1866);
and U3064 (N_3064,N_577,N_147);
or U3065 (N_3065,N_1842,N_36);
or U3066 (N_3066,N_1341,N_394);
nand U3067 (N_3067,N_630,N_1631);
nand U3068 (N_3068,N_1832,N_187);
or U3069 (N_3069,N_75,N_1776);
and U3070 (N_3070,N_1854,N_1900);
nand U3071 (N_3071,N_1540,N_954);
and U3072 (N_3072,N_1693,N_1929);
and U3073 (N_3073,N_1031,N_1918);
nand U3074 (N_3074,N_1317,N_1935);
nand U3075 (N_3075,N_10,N_709);
or U3076 (N_3076,N_1410,N_768);
and U3077 (N_3077,N_1686,N_1542);
nor U3078 (N_3078,N_796,N_1360);
nand U3079 (N_3079,N_1808,N_1534);
nor U3080 (N_3080,N_479,N_1257);
nor U3081 (N_3081,N_363,N_541);
or U3082 (N_3082,N_866,N_901);
nand U3083 (N_3083,N_1699,N_1995);
nand U3084 (N_3084,N_1430,N_1193);
or U3085 (N_3085,N_481,N_470);
or U3086 (N_3086,N_275,N_1838);
and U3087 (N_3087,N_182,N_645);
nor U3088 (N_3088,N_1346,N_1151);
nand U3089 (N_3089,N_220,N_1702);
and U3090 (N_3090,N_573,N_1977);
or U3091 (N_3091,N_1683,N_1258);
or U3092 (N_3092,N_1106,N_1701);
nor U3093 (N_3093,N_1910,N_1227);
or U3094 (N_3094,N_778,N_1635);
nand U3095 (N_3095,N_928,N_788);
and U3096 (N_3096,N_783,N_1674);
or U3097 (N_3097,N_883,N_1434);
or U3098 (N_3098,N_1655,N_695);
or U3099 (N_3099,N_662,N_285);
or U3100 (N_3100,N_1129,N_216);
or U3101 (N_3101,N_1189,N_375);
nand U3102 (N_3102,N_800,N_458);
and U3103 (N_3103,N_978,N_1534);
nand U3104 (N_3104,N_1950,N_1156);
and U3105 (N_3105,N_45,N_1564);
or U3106 (N_3106,N_958,N_1489);
or U3107 (N_3107,N_60,N_185);
and U3108 (N_3108,N_91,N_830);
and U3109 (N_3109,N_285,N_23);
or U3110 (N_3110,N_1017,N_819);
or U3111 (N_3111,N_1655,N_1904);
nand U3112 (N_3112,N_1108,N_1315);
or U3113 (N_3113,N_404,N_721);
nor U3114 (N_3114,N_1279,N_1523);
and U3115 (N_3115,N_1191,N_117);
nand U3116 (N_3116,N_404,N_924);
or U3117 (N_3117,N_1784,N_887);
xnor U3118 (N_3118,N_190,N_1350);
and U3119 (N_3119,N_635,N_419);
nor U3120 (N_3120,N_129,N_1828);
or U3121 (N_3121,N_4,N_696);
nor U3122 (N_3122,N_750,N_358);
nor U3123 (N_3123,N_1828,N_373);
and U3124 (N_3124,N_1369,N_1221);
or U3125 (N_3125,N_1054,N_936);
or U3126 (N_3126,N_51,N_527);
nor U3127 (N_3127,N_1081,N_1769);
nor U3128 (N_3128,N_1369,N_1129);
nand U3129 (N_3129,N_1018,N_500);
nand U3130 (N_3130,N_1973,N_1820);
nor U3131 (N_3131,N_670,N_598);
nor U3132 (N_3132,N_1809,N_1901);
and U3133 (N_3133,N_723,N_1356);
and U3134 (N_3134,N_934,N_708);
and U3135 (N_3135,N_1318,N_1193);
nor U3136 (N_3136,N_1654,N_1453);
nor U3137 (N_3137,N_1119,N_463);
and U3138 (N_3138,N_1898,N_406);
and U3139 (N_3139,N_1486,N_176);
nor U3140 (N_3140,N_589,N_170);
nand U3141 (N_3141,N_812,N_446);
nand U3142 (N_3142,N_366,N_647);
nor U3143 (N_3143,N_449,N_964);
or U3144 (N_3144,N_427,N_508);
nand U3145 (N_3145,N_1139,N_1937);
nor U3146 (N_3146,N_1089,N_346);
and U3147 (N_3147,N_1164,N_503);
or U3148 (N_3148,N_1277,N_477);
and U3149 (N_3149,N_786,N_1620);
or U3150 (N_3150,N_1564,N_1698);
or U3151 (N_3151,N_533,N_183);
nand U3152 (N_3152,N_1906,N_1623);
or U3153 (N_3153,N_588,N_1121);
nand U3154 (N_3154,N_1828,N_1460);
and U3155 (N_3155,N_589,N_267);
or U3156 (N_3156,N_1993,N_592);
nand U3157 (N_3157,N_61,N_581);
nor U3158 (N_3158,N_1780,N_271);
and U3159 (N_3159,N_1500,N_1515);
xor U3160 (N_3160,N_1578,N_1979);
or U3161 (N_3161,N_1819,N_724);
or U3162 (N_3162,N_877,N_355);
or U3163 (N_3163,N_429,N_1031);
nand U3164 (N_3164,N_743,N_40);
nor U3165 (N_3165,N_1573,N_1931);
and U3166 (N_3166,N_1514,N_923);
nand U3167 (N_3167,N_1149,N_491);
nor U3168 (N_3168,N_1693,N_904);
or U3169 (N_3169,N_1019,N_58);
or U3170 (N_3170,N_490,N_1351);
or U3171 (N_3171,N_1969,N_1207);
or U3172 (N_3172,N_1209,N_721);
and U3173 (N_3173,N_145,N_1561);
nor U3174 (N_3174,N_287,N_1766);
nand U3175 (N_3175,N_728,N_443);
nor U3176 (N_3176,N_65,N_1208);
and U3177 (N_3177,N_1232,N_1022);
xor U3178 (N_3178,N_1967,N_629);
nand U3179 (N_3179,N_1186,N_970);
or U3180 (N_3180,N_836,N_1742);
nor U3181 (N_3181,N_1789,N_326);
or U3182 (N_3182,N_1949,N_1609);
nand U3183 (N_3183,N_500,N_796);
nor U3184 (N_3184,N_1764,N_907);
or U3185 (N_3185,N_851,N_503);
or U3186 (N_3186,N_1450,N_1392);
or U3187 (N_3187,N_1032,N_1630);
and U3188 (N_3188,N_509,N_1421);
and U3189 (N_3189,N_1260,N_353);
nor U3190 (N_3190,N_1638,N_1622);
nor U3191 (N_3191,N_1820,N_795);
nor U3192 (N_3192,N_847,N_1174);
nand U3193 (N_3193,N_345,N_1854);
nor U3194 (N_3194,N_1857,N_1747);
and U3195 (N_3195,N_871,N_15);
nand U3196 (N_3196,N_1193,N_944);
and U3197 (N_3197,N_1321,N_1069);
and U3198 (N_3198,N_971,N_766);
xor U3199 (N_3199,N_604,N_1784);
nor U3200 (N_3200,N_1359,N_1546);
or U3201 (N_3201,N_883,N_1710);
nor U3202 (N_3202,N_933,N_1101);
nor U3203 (N_3203,N_1745,N_17);
or U3204 (N_3204,N_1394,N_1108);
and U3205 (N_3205,N_1730,N_1956);
and U3206 (N_3206,N_227,N_1618);
and U3207 (N_3207,N_1760,N_908);
and U3208 (N_3208,N_1208,N_729);
nor U3209 (N_3209,N_1030,N_1657);
nand U3210 (N_3210,N_1468,N_495);
and U3211 (N_3211,N_1345,N_582);
or U3212 (N_3212,N_443,N_946);
and U3213 (N_3213,N_1375,N_1636);
nor U3214 (N_3214,N_1228,N_804);
nand U3215 (N_3215,N_484,N_1441);
nor U3216 (N_3216,N_487,N_1732);
and U3217 (N_3217,N_67,N_871);
or U3218 (N_3218,N_1353,N_1097);
nand U3219 (N_3219,N_736,N_717);
and U3220 (N_3220,N_1611,N_1752);
xor U3221 (N_3221,N_483,N_402);
nand U3222 (N_3222,N_1706,N_483);
or U3223 (N_3223,N_1351,N_30);
and U3224 (N_3224,N_334,N_1469);
or U3225 (N_3225,N_1582,N_5);
or U3226 (N_3226,N_412,N_1048);
nand U3227 (N_3227,N_1317,N_1895);
nand U3228 (N_3228,N_204,N_167);
nor U3229 (N_3229,N_1150,N_424);
and U3230 (N_3230,N_901,N_1186);
nor U3231 (N_3231,N_1581,N_1225);
nand U3232 (N_3232,N_635,N_1415);
nor U3233 (N_3233,N_1833,N_1812);
or U3234 (N_3234,N_156,N_1871);
nor U3235 (N_3235,N_1828,N_1876);
and U3236 (N_3236,N_1000,N_1933);
or U3237 (N_3237,N_14,N_561);
nor U3238 (N_3238,N_562,N_298);
or U3239 (N_3239,N_278,N_107);
nor U3240 (N_3240,N_1456,N_1326);
and U3241 (N_3241,N_1660,N_465);
or U3242 (N_3242,N_1033,N_508);
nor U3243 (N_3243,N_694,N_491);
and U3244 (N_3244,N_19,N_1276);
or U3245 (N_3245,N_226,N_1509);
or U3246 (N_3246,N_935,N_1944);
nand U3247 (N_3247,N_1125,N_1921);
nand U3248 (N_3248,N_523,N_209);
nand U3249 (N_3249,N_1001,N_1262);
and U3250 (N_3250,N_647,N_797);
and U3251 (N_3251,N_590,N_244);
nor U3252 (N_3252,N_1843,N_1674);
nand U3253 (N_3253,N_631,N_908);
and U3254 (N_3254,N_780,N_1321);
and U3255 (N_3255,N_468,N_382);
and U3256 (N_3256,N_963,N_374);
nor U3257 (N_3257,N_170,N_385);
nand U3258 (N_3258,N_1036,N_384);
nand U3259 (N_3259,N_1427,N_1804);
nand U3260 (N_3260,N_514,N_834);
or U3261 (N_3261,N_1185,N_1701);
nand U3262 (N_3262,N_1644,N_1378);
nor U3263 (N_3263,N_761,N_1228);
and U3264 (N_3264,N_1644,N_1356);
and U3265 (N_3265,N_1452,N_1175);
and U3266 (N_3266,N_1991,N_267);
and U3267 (N_3267,N_68,N_1410);
nand U3268 (N_3268,N_529,N_437);
nor U3269 (N_3269,N_1428,N_1823);
or U3270 (N_3270,N_1851,N_1448);
and U3271 (N_3271,N_1634,N_1518);
nor U3272 (N_3272,N_62,N_569);
and U3273 (N_3273,N_1429,N_1708);
nand U3274 (N_3274,N_522,N_1475);
nor U3275 (N_3275,N_1555,N_474);
nand U3276 (N_3276,N_1605,N_27);
nand U3277 (N_3277,N_1063,N_545);
or U3278 (N_3278,N_744,N_1150);
nor U3279 (N_3279,N_792,N_1854);
and U3280 (N_3280,N_1884,N_1969);
or U3281 (N_3281,N_1353,N_297);
or U3282 (N_3282,N_1921,N_22);
nand U3283 (N_3283,N_1987,N_1660);
and U3284 (N_3284,N_669,N_1710);
nor U3285 (N_3285,N_584,N_1953);
nor U3286 (N_3286,N_1671,N_1440);
and U3287 (N_3287,N_1667,N_1700);
nor U3288 (N_3288,N_1669,N_879);
and U3289 (N_3289,N_72,N_1936);
nor U3290 (N_3290,N_1416,N_1613);
or U3291 (N_3291,N_1334,N_98);
nand U3292 (N_3292,N_344,N_87);
and U3293 (N_3293,N_772,N_475);
nor U3294 (N_3294,N_21,N_1472);
nand U3295 (N_3295,N_49,N_1446);
nand U3296 (N_3296,N_192,N_476);
nor U3297 (N_3297,N_1188,N_1301);
nor U3298 (N_3298,N_1291,N_1126);
or U3299 (N_3299,N_1208,N_1314);
nand U3300 (N_3300,N_692,N_147);
xnor U3301 (N_3301,N_1248,N_1375);
or U3302 (N_3302,N_1947,N_1655);
or U3303 (N_3303,N_491,N_1450);
nor U3304 (N_3304,N_422,N_1592);
and U3305 (N_3305,N_417,N_1355);
or U3306 (N_3306,N_341,N_607);
and U3307 (N_3307,N_1137,N_1334);
nand U3308 (N_3308,N_278,N_304);
nand U3309 (N_3309,N_654,N_954);
nor U3310 (N_3310,N_1535,N_1525);
or U3311 (N_3311,N_924,N_1410);
nand U3312 (N_3312,N_154,N_1413);
and U3313 (N_3313,N_1978,N_364);
nor U3314 (N_3314,N_1592,N_284);
nand U3315 (N_3315,N_1103,N_1115);
nor U3316 (N_3316,N_545,N_1523);
nand U3317 (N_3317,N_709,N_1972);
nand U3318 (N_3318,N_1175,N_1838);
nand U3319 (N_3319,N_843,N_829);
nor U3320 (N_3320,N_1337,N_1405);
or U3321 (N_3321,N_1748,N_1734);
nand U3322 (N_3322,N_1741,N_1828);
xor U3323 (N_3323,N_273,N_1558);
or U3324 (N_3324,N_1632,N_739);
nand U3325 (N_3325,N_1819,N_1747);
nor U3326 (N_3326,N_1408,N_730);
nor U3327 (N_3327,N_1441,N_116);
or U3328 (N_3328,N_1145,N_1196);
or U3329 (N_3329,N_43,N_408);
or U3330 (N_3330,N_1527,N_1969);
and U3331 (N_3331,N_1377,N_81);
xnor U3332 (N_3332,N_1231,N_671);
or U3333 (N_3333,N_1671,N_1034);
xor U3334 (N_3334,N_767,N_1789);
nand U3335 (N_3335,N_1619,N_1021);
nand U3336 (N_3336,N_747,N_1118);
and U3337 (N_3337,N_822,N_1704);
and U3338 (N_3338,N_1263,N_636);
nor U3339 (N_3339,N_1827,N_512);
nor U3340 (N_3340,N_1314,N_925);
nor U3341 (N_3341,N_867,N_17);
xor U3342 (N_3342,N_1472,N_1775);
nand U3343 (N_3343,N_593,N_345);
nor U3344 (N_3344,N_814,N_1182);
nand U3345 (N_3345,N_1515,N_1082);
or U3346 (N_3346,N_152,N_521);
or U3347 (N_3347,N_1535,N_728);
or U3348 (N_3348,N_105,N_894);
nand U3349 (N_3349,N_605,N_1232);
or U3350 (N_3350,N_1994,N_1997);
nor U3351 (N_3351,N_792,N_875);
nand U3352 (N_3352,N_839,N_1645);
nand U3353 (N_3353,N_449,N_428);
nand U3354 (N_3354,N_1639,N_944);
and U3355 (N_3355,N_587,N_508);
or U3356 (N_3356,N_307,N_1636);
and U3357 (N_3357,N_297,N_1931);
nand U3358 (N_3358,N_1241,N_1276);
nand U3359 (N_3359,N_725,N_1844);
nor U3360 (N_3360,N_518,N_294);
nor U3361 (N_3361,N_1182,N_1771);
and U3362 (N_3362,N_1237,N_1525);
or U3363 (N_3363,N_663,N_1419);
or U3364 (N_3364,N_1791,N_368);
nor U3365 (N_3365,N_1962,N_1105);
nor U3366 (N_3366,N_1348,N_394);
nor U3367 (N_3367,N_763,N_925);
or U3368 (N_3368,N_547,N_1415);
or U3369 (N_3369,N_1276,N_756);
xnor U3370 (N_3370,N_270,N_20);
and U3371 (N_3371,N_103,N_529);
nor U3372 (N_3372,N_1800,N_1181);
nand U3373 (N_3373,N_1200,N_1798);
and U3374 (N_3374,N_421,N_1777);
and U3375 (N_3375,N_476,N_172);
nor U3376 (N_3376,N_1773,N_870);
or U3377 (N_3377,N_793,N_887);
or U3378 (N_3378,N_1628,N_1906);
or U3379 (N_3379,N_896,N_415);
or U3380 (N_3380,N_291,N_841);
nor U3381 (N_3381,N_1585,N_850);
xor U3382 (N_3382,N_469,N_1149);
nor U3383 (N_3383,N_1321,N_471);
nor U3384 (N_3384,N_1080,N_247);
and U3385 (N_3385,N_1312,N_182);
or U3386 (N_3386,N_1644,N_767);
nand U3387 (N_3387,N_386,N_1402);
nor U3388 (N_3388,N_823,N_1567);
nand U3389 (N_3389,N_1171,N_800);
or U3390 (N_3390,N_365,N_1591);
or U3391 (N_3391,N_530,N_1027);
nand U3392 (N_3392,N_1366,N_1589);
or U3393 (N_3393,N_1310,N_1303);
nand U3394 (N_3394,N_569,N_1036);
nand U3395 (N_3395,N_1095,N_796);
and U3396 (N_3396,N_1128,N_221);
nor U3397 (N_3397,N_1210,N_980);
nand U3398 (N_3398,N_331,N_499);
and U3399 (N_3399,N_1605,N_778);
or U3400 (N_3400,N_1096,N_528);
nand U3401 (N_3401,N_1109,N_1116);
nor U3402 (N_3402,N_1294,N_675);
nand U3403 (N_3403,N_1065,N_148);
and U3404 (N_3404,N_1284,N_753);
nand U3405 (N_3405,N_564,N_1019);
and U3406 (N_3406,N_1444,N_407);
nand U3407 (N_3407,N_23,N_1616);
or U3408 (N_3408,N_1153,N_459);
or U3409 (N_3409,N_857,N_518);
nand U3410 (N_3410,N_1260,N_782);
nor U3411 (N_3411,N_662,N_1118);
nor U3412 (N_3412,N_1386,N_1300);
or U3413 (N_3413,N_1498,N_1735);
nand U3414 (N_3414,N_1552,N_864);
nand U3415 (N_3415,N_1583,N_198);
and U3416 (N_3416,N_1273,N_1551);
or U3417 (N_3417,N_617,N_1573);
nand U3418 (N_3418,N_795,N_1927);
nand U3419 (N_3419,N_1770,N_533);
and U3420 (N_3420,N_739,N_1287);
nor U3421 (N_3421,N_459,N_1559);
or U3422 (N_3422,N_1264,N_865);
nor U3423 (N_3423,N_1019,N_722);
and U3424 (N_3424,N_1868,N_1605);
and U3425 (N_3425,N_662,N_1405);
or U3426 (N_3426,N_138,N_1107);
and U3427 (N_3427,N_416,N_1074);
nand U3428 (N_3428,N_935,N_686);
nand U3429 (N_3429,N_1132,N_1877);
nand U3430 (N_3430,N_1059,N_33);
xor U3431 (N_3431,N_247,N_1188);
nor U3432 (N_3432,N_416,N_1189);
and U3433 (N_3433,N_1993,N_744);
nor U3434 (N_3434,N_1417,N_883);
nand U3435 (N_3435,N_20,N_1354);
nand U3436 (N_3436,N_1837,N_44);
nor U3437 (N_3437,N_1377,N_193);
nand U3438 (N_3438,N_777,N_1098);
nand U3439 (N_3439,N_1016,N_202);
and U3440 (N_3440,N_1031,N_339);
nand U3441 (N_3441,N_235,N_232);
or U3442 (N_3442,N_316,N_1673);
nor U3443 (N_3443,N_1797,N_837);
xnor U3444 (N_3444,N_1013,N_1914);
and U3445 (N_3445,N_207,N_1941);
nor U3446 (N_3446,N_1813,N_1744);
nor U3447 (N_3447,N_1266,N_722);
nand U3448 (N_3448,N_1842,N_1187);
nor U3449 (N_3449,N_1599,N_1429);
or U3450 (N_3450,N_1299,N_1301);
or U3451 (N_3451,N_837,N_843);
and U3452 (N_3452,N_1870,N_1413);
and U3453 (N_3453,N_506,N_1404);
nand U3454 (N_3454,N_1733,N_923);
and U3455 (N_3455,N_1054,N_759);
nand U3456 (N_3456,N_1171,N_147);
nand U3457 (N_3457,N_443,N_61);
nand U3458 (N_3458,N_1542,N_1982);
xor U3459 (N_3459,N_1637,N_340);
and U3460 (N_3460,N_634,N_177);
nor U3461 (N_3461,N_704,N_1981);
nand U3462 (N_3462,N_108,N_1955);
nand U3463 (N_3463,N_778,N_725);
nand U3464 (N_3464,N_921,N_1115);
nand U3465 (N_3465,N_279,N_102);
or U3466 (N_3466,N_1837,N_948);
and U3467 (N_3467,N_1872,N_641);
nand U3468 (N_3468,N_1692,N_602);
nand U3469 (N_3469,N_111,N_195);
nand U3470 (N_3470,N_1618,N_1002);
nand U3471 (N_3471,N_1938,N_1048);
nand U3472 (N_3472,N_193,N_1153);
nand U3473 (N_3473,N_1337,N_1137);
or U3474 (N_3474,N_1262,N_1530);
or U3475 (N_3475,N_661,N_27);
or U3476 (N_3476,N_1017,N_857);
nor U3477 (N_3477,N_967,N_585);
nand U3478 (N_3478,N_1644,N_224);
nand U3479 (N_3479,N_329,N_1202);
or U3480 (N_3480,N_1952,N_946);
nor U3481 (N_3481,N_829,N_1287);
nand U3482 (N_3482,N_291,N_1074);
and U3483 (N_3483,N_1843,N_1066);
nand U3484 (N_3484,N_258,N_115);
or U3485 (N_3485,N_1290,N_1480);
or U3486 (N_3486,N_152,N_1786);
nor U3487 (N_3487,N_1301,N_981);
nor U3488 (N_3488,N_1757,N_1958);
and U3489 (N_3489,N_1759,N_519);
nand U3490 (N_3490,N_1040,N_641);
and U3491 (N_3491,N_1131,N_442);
nor U3492 (N_3492,N_442,N_1912);
nor U3493 (N_3493,N_494,N_889);
nand U3494 (N_3494,N_1227,N_807);
nor U3495 (N_3495,N_814,N_677);
nand U3496 (N_3496,N_1495,N_1898);
nand U3497 (N_3497,N_202,N_1858);
nand U3498 (N_3498,N_164,N_597);
and U3499 (N_3499,N_1232,N_1746);
or U3500 (N_3500,N_1121,N_1516);
nand U3501 (N_3501,N_520,N_254);
nand U3502 (N_3502,N_1352,N_1800);
nor U3503 (N_3503,N_154,N_76);
nand U3504 (N_3504,N_815,N_1588);
or U3505 (N_3505,N_427,N_405);
nor U3506 (N_3506,N_1243,N_1650);
and U3507 (N_3507,N_1791,N_658);
nor U3508 (N_3508,N_1489,N_1835);
or U3509 (N_3509,N_1942,N_1595);
or U3510 (N_3510,N_1769,N_898);
xor U3511 (N_3511,N_1590,N_588);
nor U3512 (N_3512,N_71,N_774);
and U3513 (N_3513,N_1536,N_1276);
or U3514 (N_3514,N_1196,N_64);
nand U3515 (N_3515,N_243,N_1645);
nand U3516 (N_3516,N_536,N_853);
or U3517 (N_3517,N_768,N_940);
nand U3518 (N_3518,N_612,N_364);
and U3519 (N_3519,N_1361,N_1056);
or U3520 (N_3520,N_452,N_1867);
or U3521 (N_3521,N_1702,N_1256);
and U3522 (N_3522,N_1389,N_1396);
nor U3523 (N_3523,N_2,N_1070);
xor U3524 (N_3524,N_296,N_1946);
or U3525 (N_3525,N_1239,N_352);
nand U3526 (N_3526,N_268,N_741);
nand U3527 (N_3527,N_1013,N_605);
and U3528 (N_3528,N_1427,N_1500);
nor U3529 (N_3529,N_753,N_698);
and U3530 (N_3530,N_981,N_1928);
nand U3531 (N_3531,N_1966,N_763);
nand U3532 (N_3532,N_88,N_1757);
nand U3533 (N_3533,N_1824,N_522);
and U3534 (N_3534,N_1914,N_1596);
or U3535 (N_3535,N_1884,N_1041);
and U3536 (N_3536,N_68,N_101);
nor U3537 (N_3537,N_1519,N_1900);
and U3538 (N_3538,N_656,N_775);
nor U3539 (N_3539,N_148,N_45);
nor U3540 (N_3540,N_8,N_415);
nand U3541 (N_3541,N_667,N_1888);
or U3542 (N_3542,N_1130,N_803);
nor U3543 (N_3543,N_1722,N_791);
nor U3544 (N_3544,N_1182,N_735);
nor U3545 (N_3545,N_642,N_1533);
nand U3546 (N_3546,N_491,N_1183);
nand U3547 (N_3547,N_341,N_239);
or U3548 (N_3548,N_260,N_692);
and U3549 (N_3549,N_1584,N_99);
nor U3550 (N_3550,N_514,N_609);
nor U3551 (N_3551,N_1771,N_202);
or U3552 (N_3552,N_1724,N_1750);
nor U3553 (N_3553,N_57,N_1665);
nand U3554 (N_3554,N_150,N_266);
or U3555 (N_3555,N_788,N_1642);
nor U3556 (N_3556,N_1560,N_200);
nor U3557 (N_3557,N_1475,N_1506);
or U3558 (N_3558,N_174,N_1776);
or U3559 (N_3559,N_1966,N_361);
or U3560 (N_3560,N_709,N_1704);
or U3561 (N_3561,N_869,N_1032);
nand U3562 (N_3562,N_1512,N_1422);
and U3563 (N_3563,N_218,N_475);
and U3564 (N_3564,N_1535,N_1826);
or U3565 (N_3565,N_208,N_1971);
nor U3566 (N_3566,N_374,N_565);
nor U3567 (N_3567,N_1356,N_246);
or U3568 (N_3568,N_57,N_1079);
nor U3569 (N_3569,N_1468,N_1816);
nand U3570 (N_3570,N_320,N_1281);
nand U3571 (N_3571,N_1678,N_1048);
or U3572 (N_3572,N_829,N_1391);
and U3573 (N_3573,N_1506,N_1863);
nor U3574 (N_3574,N_1821,N_1529);
nor U3575 (N_3575,N_416,N_1587);
nand U3576 (N_3576,N_560,N_1097);
nor U3577 (N_3577,N_96,N_992);
nor U3578 (N_3578,N_190,N_849);
nand U3579 (N_3579,N_1238,N_324);
and U3580 (N_3580,N_756,N_400);
nor U3581 (N_3581,N_956,N_144);
and U3582 (N_3582,N_1433,N_1356);
nor U3583 (N_3583,N_218,N_996);
and U3584 (N_3584,N_1219,N_1291);
and U3585 (N_3585,N_902,N_1028);
or U3586 (N_3586,N_1399,N_1790);
nor U3587 (N_3587,N_1315,N_751);
nor U3588 (N_3588,N_727,N_1350);
and U3589 (N_3589,N_793,N_141);
or U3590 (N_3590,N_107,N_1928);
nand U3591 (N_3591,N_206,N_1978);
and U3592 (N_3592,N_1748,N_464);
nor U3593 (N_3593,N_390,N_128);
nor U3594 (N_3594,N_236,N_4);
and U3595 (N_3595,N_44,N_701);
and U3596 (N_3596,N_1914,N_1156);
and U3597 (N_3597,N_27,N_420);
or U3598 (N_3598,N_5,N_409);
nor U3599 (N_3599,N_978,N_401);
or U3600 (N_3600,N_702,N_49);
or U3601 (N_3601,N_1971,N_376);
and U3602 (N_3602,N_348,N_1482);
and U3603 (N_3603,N_634,N_841);
or U3604 (N_3604,N_58,N_726);
nor U3605 (N_3605,N_1135,N_536);
nor U3606 (N_3606,N_160,N_1841);
and U3607 (N_3607,N_1268,N_1115);
or U3608 (N_3608,N_1096,N_968);
nand U3609 (N_3609,N_1018,N_3);
and U3610 (N_3610,N_1212,N_1793);
and U3611 (N_3611,N_870,N_1304);
nor U3612 (N_3612,N_103,N_1570);
and U3613 (N_3613,N_1864,N_246);
or U3614 (N_3614,N_1052,N_610);
nand U3615 (N_3615,N_375,N_980);
nand U3616 (N_3616,N_467,N_184);
nand U3617 (N_3617,N_1376,N_1962);
nand U3618 (N_3618,N_1322,N_569);
nor U3619 (N_3619,N_524,N_985);
nand U3620 (N_3620,N_1466,N_99);
nor U3621 (N_3621,N_1858,N_1039);
nand U3622 (N_3622,N_223,N_1894);
and U3623 (N_3623,N_522,N_1479);
xnor U3624 (N_3624,N_1251,N_553);
nand U3625 (N_3625,N_218,N_1887);
and U3626 (N_3626,N_26,N_1594);
and U3627 (N_3627,N_190,N_106);
nor U3628 (N_3628,N_1337,N_649);
or U3629 (N_3629,N_847,N_1990);
nor U3630 (N_3630,N_1691,N_1361);
and U3631 (N_3631,N_1565,N_41);
xnor U3632 (N_3632,N_1778,N_218);
nand U3633 (N_3633,N_1780,N_329);
nor U3634 (N_3634,N_1295,N_1136);
nor U3635 (N_3635,N_343,N_330);
or U3636 (N_3636,N_1880,N_1327);
nand U3637 (N_3637,N_621,N_973);
and U3638 (N_3638,N_80,N_1186);
nor U3639 (N_3639,N_860,N_647);
nand U3640 (N_3640,N_1770,N_1409);
or U3641 (N_3641,N_971,N_506);
nor U3642 (N_3642,N_1824,N_1629);
xnor U3643 (N_3643,N_1829,N_1431);
nand U3644 (N_3644,N_1096,N_82);
nor U3645 (N_3645,N_1103,N_453);
nand U3646 (N_3646,N_652,N_519);
nand U3647 (N_3647,N_1002,N_876);
or U3648 (N_3648,N_1125,N_259);
nor U3649 (N_3649,N_1219,N_1130);
nor U3650 (N_3650,N_245,N_228);
and U3651 (N_3651,N_1993,N_1221);
xnor U3652 (N_3652,N_689,N_1780);
nand U3653 (N_3653,N_1173,N_787);
or U3654 (N_3654,N_331,N_1978);
or U3655 (N_3655,N_1803,N_1585);
nand U3656 (N_3656,N_1914,N_734);
nand U3657 (N_3657,N_952,N_154);
and U3658 (N_3658,N_220,N_611);
nand U3659 (N_3659,N_47,N_1688);
or U3660 (N_3660,N_1864,N_691);
and U3661 (N_3661,N_1586,N_15);
nor U3662 (N_3662,N_63,N_1348);
nand U3663 (N_3663,N_1736,N_1289);
nor U3664 (N_3664,N_1561,N_1423);
or U3665 (N_3665,N_1020,N_1670);
and U3666 (N_3666,N_1369,N_146);
and U3667 (N_3667,N_851,N_1722);
and U3668 (N_3668,N_1775,N_1113);
or U3669 (N_3669,N_345,N_257);
or U3670 (N_3670,N_1380,N_1117);
nand U3671 (N_3671,N_613,N_389);
nand U3672 (N_3672,N_1957,N_160);
nor U3673 (N_3673,N_1266,N_1133);
and U3674 (N_3674,N_1822,N_1318);
nand U3675 (N_3675,N_386,N_977);
nor U3676 (N_3676,N_698,N_1576);
nand U3677 (N_3677,N_1456,N_370);
or U3678 (N_3678,N_56,N_1286);
nor U3679 (N_3679,N_42,N_1490);
or U3680 (N_3680,N_1690,N_1345);
or U3681 (N_3681,N_850,N_607);
nor U3682 (N_3682,N_717,N_567);
or U3683 (N_3683,N_426,N_1930);
or U3684 (N_3684,N_754,N_956);
nor U3685 (N_3685,N_1595,N_1586);
nand U3686 (N_3686,N_412,N_157);
or U3687 (N_3687,N_1975,N_473);
or U3688 (N_3688,N_643,N_438);
or U3689 (N_3689,N_1271,N_474);
and U3690 (N_3690,N_343,N_1178);
and U3691 (N_3691,N_782,N_807);
nor U3692 (N_3692,N_806,N_588);
nand U3693 (N_3693,N_493,N_1708);
nor U3694 (N_3694,N_1539,N_1002);
nand U3695 (N_3695,N_1557,N_1116);
nand U3696 (N_3696,N_1810,N_861);
nor U3697 (N_3697,N_1872,N_132);
or U3698 (N_3698,N_1735,N_1891);
or U3699 (N_3699,N_1087,N_1893);
or U3700 (N_3700,N_302,N_1265);
and U3701 (N_3701,N_498,N_795);
or U3702 (N_3702,N_982,N_1625);
or U3703 (N_3703,N_719,N_190);
and U3704 (N_3704,N_212,N_1714);
nor U3705 (N_3705,N_718,N_1309);
nand U3706 (N_3706,N_1288,N_485);
or U3707 (N_3707,N_69,N_871);
and U3708 (N_3708,N_344,N_770);
and U3709 (N_3709,N_1855,N_1190);
nor U3710 (N_3710,N_1307,N_404);
and U3711 (N_3711,N_1121,N_1858);
and U3712 (N_3712,N_1454,N_1332);
nand U3713 (N_3713,N_1575,N_139);
nand U3714 (N_3714,N_67,N_728);
nor U3715 (N_3715,N_833,N_465);
or U3716 (N_3716,N_1128,N_1055);
or U3717 (N_3717,N_1890,N_185);
nor U3718 (N_3718,N_172,N_107);
nor U3719 (N_3719,N_1257,N_170);
and U3720 (N_3720,N_1115,N_1239);
nand U3721 (N_3721,N_546,N_415);
nor U3722 (N_3722,N_1060,N_113);
and U3723 (N_3723,N_473,N_515);
nand U3724 (N_3724,N_1366,N_396);
or U3725 (N_3725,N_368,N_556);
nor U3726 (N_3726,N_1304,N_748);
and U3727 (N_3727,N_1256,N_1475);
nand U3728 (N_3728,N_449,N_1643);
or U3729 (N_3729,N_751,N_110);
or U3730 (N_3730,N_470,N_130);
and U3731 (N_3731,N_1229,N_1446);
or U3732 (N_3732,N_98,N_214);
nand U3733 (N_3733,N_585,N_560);
and U3734 (N_3734,N_1649,N_1961);
nand U3735 (N_3735,N_1777,N_1465);
and U3736 (N_3736,N_1688,N_1683);
and U3737 (N_3737,N_913,N_1049);
and U3738 (N_3738,N_793,N_694);
nor U3739 (N_3739,N_220,N_1209);
or U3740 (N_3740,N_1702,N_51);
nor U3741 (N_3741,N_1856,N_888);
nand U3742 (N_3742,N_1965,N_1596);
and U3743 (N_3743,N_1433,N_1825);
nor U3744 (N_3744,N_1550,N_781);
or U3745 (N_3745,N_780,N_1073);
and U3746 (N_3746,N_1879,N_580);
nor U3747 (N_3747,N_155,N_1451);
and U3748 (N_3748,N_661,N_1226);
nand U3749 (N_3749,N_852,N_77);
or U3750 (N_3750,N_750,N_1476);
and U3751 (N_3751,N_65,N_179);
nor U3752 (N_3752,N_840,N_1765);
nor U3753 (N_3753,N_1346,N_1616);
nor U3754 (N_3754,N_380,N_610);
or U3755 (N_3755,N_878,N_1491);
or U3756 (N_3756,N_906,N_559);
nor U3757 (N_3757,N_1099,N_969);
nand U3758 (N_3758,N_917,N_1569);
or U3759 (N_3759,N_1595,N_535);
and U3760 (N_3760,N_1555,N_818);
nand U3761 (N_3761,N_733,N_1116);
and U3762 (N_3762,N_1197,N_749);
nand U3763 (N_3763,N_908,N_664);
and U3764 (N_3764,N_601,N_1705);
or U3765 (N_3765,N_33,N_4);
or U3766 (N_3766,N_502,N_964);
or U3767 (N_3767,N_1104,N_459);
nand U3768 (N_3768,N_194,N_1293);
or U3769 (N_3769,N_950,N_118);
and U3770 (N_3770,N_710,N_1547);
and U3771 (N_3771,N_1667,N_1274);
nor U3772 (N_3772,N_809,N_1744);
or U3773 (N_3773,N_1524,N_1444);
nor U3774 (N_3774,N_995,N_1478);
nor U3775 (N_3775,N_557,N_1234);
nand U3776 (N_3776,N_1777,N_1153);
and U3777 (N_3777,N_100,N_1955);
and U3778 (N_3778,N_248,N_390);
or U3779 (N_3779,N_18,N_413);
nand U3780 (N_3780,N_1810,N_1347);
nor U3781 (N_3781,N_937,N_331);
nand U3782 (N_3782,N_365,N_785);
nor U3783 (N_3783,N_1707,N_1788);
nor U3784 (N_3784,N_743,N_1130);
nand U3785 (N_3785,N_1662,N_1420);
and U3786 (N_3786,N_1512,N_38);
xnor U3787 (N_3787,N_1924,N_1545);
nand U3788 (N_3788,N_1111,N_310);
nor U3789 (N_3789,N_885,N_1033);
nor U3790 (N_3790,N_510,N_840);
nand U3791 (N_3791,N_1687,N_349);
nand U3792 (N_3792,N_1838,N_1433);
nor U3793 (N_3793,N_963,N_1378);
nor U3794 (N_3794,N_31,N_931);
or U3795 (N_3795,N_976,N_1298);
nand U3796 (N_3796,N_153,N_1601);
or U3797 (N_3797,N_754,N_251);
xor U3798 (N_3798,N_1534,N_292);
or U3799 (N_3799,N_827,N_1845);
nor U3800 (N_3800,N_1390,N_909);
nor U3801 (N_3801,N_1871,N_1588);
nor U3802 (N_3802,N_87,N_305);
nand U3803 (N_3803,N_1995,N_603);
nand U3804 (N_3804,N_1633,N_858);
or U3805 (N_3805,N_1485,N_282);
and U3806 (N_3806,N_1941,N_699);
nand U3807 (N_3807,N_1479,N_313);
nand U3808 (N_3808,N_1326,N_563);
nand U3809 (N_3809,N_938,N_845);
nand U3810 (N_3810,N_953,N_1281);
nand U3811 (N_3811,N_616,N_438);
or U3812 (N_3812,N_1413,N_1385);
nor U3813 (N_3813,N_103,N_1837);
nor U3814 (N_3814,N_1864,N_663);
and U3815 (N_3815,N_123,N_105);
and U3816 (N_3816,N_712,N_242);
nand U3817 (N_3817,N_326,N_1225);
nand U3818 (N_3818,N_1162,N_1121);
nor U3819 (N_3819,N_785,N_985);
nand U3820 (N_3820,N_423,N_797);
or U3821 (N_3821,N_1609,N_1274);
or U3822 (N_3822,N_1647,N_1653);
or U3823 (N_3823,N_1789,N_967);
nor U3824 (N_3824,N_258,N_918);
nand U3825 (N_3825,N_1256,N_72);
or U3826 (N_3826,N_103,N_853);
nor U3827 (N_3827,N_243,N_325);
nand U3828 (N_3828,N_1059,N_1520);
and U3829 (N_3829,N_606,N_1890);
or U3830 (N_3830,N_986,N_1924);
nand U3831 (N_3831,N_1634,N_754);
nor U3832 (N_3832,N_1781,N_1289);
nor U3833 (N_3833,N_1955,N_1556);
nand U3834 (N_3834,N_1510,N_551);
or U3835 (N_3835,N_1619,N_1203);
nor U3836 (N_3836,N_281,N_68);
nand U3837 (N_3837,N_1114,N_1881);
or U3838 (N_3838,N_1862,N_1522);
or U3839 (N_3839,N_314,N_1814);
and U3840 (N_3840,N_1625,N_1935);
nor U3841 (N_3841,N_30,N_158);
nor U3842 (N_3842,N_1245,N_1944);
and U3843 (N_3843,N_18,N_619);
nor U3844 (N_3844,N_1476,N_1744);
and U3845 (N_3845,N_1767,N_1745);
nor U3846 (N_3846,N_1200,N_220);
nor U3847 (N_3847,N_1957,N_605);
nor U3848 (N_3848,N_799,N_581);
or U3849 (N_3849,N_1590,N_763);
nor U3850 (N_3850,N_978,N_1608);
and U3851 (N_3851,N_505,N_1518);
or U3852 (N_3852,N_515,N_1760);
xnor U3853 (N_3853,N_1600,N_1104);
or U3854 (N_3854,N_570,N_1490);
nor U3855 (N_3855,N_843,N_186);
or U3856 (N_3856,N_1748,N_1355);
nor U3857 (N_3857,N_1226,N_1724);
nor U3858 (N_3858,N_362,N_1060);
nand U3859 (N_3859,N_1943,N_1512);
and U3860 (N_3860,N_1504,N_1185);
or U3861 (N_3861,N_106,N_1337);
nor U3862 (N_3862,N_1045,N_1167);
nand U3863 (N_3863,N_812,N_986);
nor U3864 (N_3864,N_1695,N_1345);
nor U3865 (N_3865,N_1725,N_1148);
or U3866 (N_3866,N_1602,N_609);
or U3867 (N_3867,N_257,N_1932);
and U3868 (N_3868,N_17,N_492);
or U3869 (N_3869,N_787,N_646);
nand U3870 (N_3870,N_751,N_1530);
and U3871 (N_3871,N_725,N_1071);
nand U3872 (N_3872,N_955,N_941);
or U3873 (N_3873,N_372,N_967);
and U3874 (N_3874,N_552,N_1549);
nor U3875 (N_3875,N_1623,N_1384);
nand U3876 (N_3876,N_1824,N_1689);
nor U3877 (N_3877,N_1479,N_768);
nand U3878 (N_3878,N_874,N_555);
nand U3879 (N_3879,N_1414,N_771);
or U3880 (N_3880,N_1009,N_853);
nand U3881 (N_3881,N_1095,N_161);
nand U3882 (N_3882,N_1702,N_1660);
or U3883 (N_3883,N_1147,N_1460);
nor U3884 (N_3884,N_1877,N_243);
or U3885 (N_3885,N_1244,N_670);
nand U3886 (N_3886,N_353,N_213);
nand U3887 (N_3887,N_65,N_1679);
nand U3888 (N_3888,N_197,N_1924);
or U3889 (N_3889,N_681,N_1744);
nor U3890 (N_3890,N_668,N_1183);
or U3891 (N_3891,N_1801,N_1488);
nand U3892 (N_3892,N_1460,N_995);
nand U3893 (N_3893,N_689,N_905);
nand U3894 (N_3894,N_1757,N_1813);
nand U3895 (N_3895,N_227,N_1904);
nor U3896 (N_3896,N_77,N_1225);
and U3897 (N_3897,N_1341,N_1900);
or U3898 (N_3898,N_338,N_24);
or U3899 (N_3899,N_1469,N_552);
and U3900 (N_3900,N_1425,N_1614);
nor U3901 (N_3901,N_256,N_1789);
nand U3902 (N_3902,N_1404,N_460);
nand U3903 (N_3903,N_893,N_1956);
nor U3904 (N_3904,N_586,N_1166);
or U3905 (N_3905,N_1009,N_178);
nand U3906 (N_3906,N_85,N_734);
and U3907 (N_3907,N_962,N_989);
nor U3908 (N_3908,N_867,N_321);
or U3909 (N_3909,N_1650,N_1041);
nor U3910 (N_3910,N_96,N_98);
and U3911 (N_3911,N_1216,N_711);
nor U3912 (N_3912,N_1553,N_1777);
nand U3913 (N_3913,N_1632,N_494);
or U3914 (N_3914,N_863,N_777);
nand U3915 (N_3915,N_199,N_293);
and U3916 (N_3916,N_275,N_1346);
or U3917 (N_3917,N_430,N_1276);
nand U3918 (N_3918,N_1637,N_1812);
nor U3919 (N_3919,N_924,N_773);
nand U3920 (N_3920,N_1707,N_26);
and U3921 (N_3921,N_1235,N_1021);
and U3922 (N_3922,N_1984,N_1388);
and U3923 (N_3923,N_65,N_1025);
nor U3924 (N_3924,N_1949,N_1307);
and U3925 (N_3925,N_1650,N_1352);
nand U3926 (N_3926,N_1480,N_1024);
nand U3927 (N_3927,N_1560,N_1278);
and U3928 (N_3928,N_784,N_523);
or U3929 (N_3929,N_1237,N_928);
and U3930 (N_3930,N_907,N_1385);
and U3931 (N_3931,N_1784,N_1024);
or U3932 (N_3932,N_216,N_1680);
nand U3933 (N_3933,N_383,N_1519);
and U3934 (N_3934,N_165,N_4);
and U3935 (N_3935,N_981,N_1153);
nor U3936 (N_3936,N_1548,N_1128);
and U3937 (N_3937,N_715,N_1006);
nor U3938 (N_3938,N_1216,N_1133);
and U3939 (N_3939,N_1377,N_744);
nand U3940 (N_3940,N_1176,N_431);
or U3941 (N_3941,N_1000,N_235);
nand U3942 (N_3942,N_828,N_1574);
and U3943 (N_3943,N_458,N_469);
nand U3944 (N_3944,N_1415,N_1074);
nor U3945 (N_3945,N_1066,N_309);
and U3946 (N_3946,N_1213,N_1384);
nor U3947 (N_3947,N_1699,N_1843);
or U3948 (N_3948,N_1413,N_1809);
or U3949 (N_3949,N_4,N_1616);
nor U3950 (N_3950,N_687,N_1716);
nand U3951 (N_3951,N_1198,N_1973);
nand U3952 (N_3952,N_1829,N_732);
or U3953 (N_3953,N_833,N_285);
and U3954 (N_3954,N_1754,N_1311);
nand U3955 (N_3955,N_1721,N_1804);
nand U3956 (N_3956,N_1355,N_1871);
and U3957 (N_3957,N_1945,N_667);
and U3958 (N_3958,N_611,N_715);
nor U3959 (N_3959,N_1189,N_880);
xor U3960 (N_3960,N_430,N_1944);
and U3961 (N_3961,N_1139,N_1731);
or U3962 (N_3962,N_1821,N_663);
or U3963 (N_3963,N_1298,N_1086);
and U3964 (N_3964,N_1342,N_1889);
nand U3965 (N_3965,N_1156,N_1477);
or U3966 (N_3966,N_118,N_929);
or U3967 (N_3967,N_1367,N_614);
nand U3968 (N_3968,N_930,N_1741);
or U3969 (N_3969,N_1033,N_998);
nor U3970 (N_3970,N_500,N_803);
or U3971 (N_3971,N_1027,N_1034);
and U3972 (N_3972,N_846,N_1879);
nand U3973 (N_3973,N_809,N_1913);
xor U3974 (N_3974,N_1965,N_572);
nand U3975 (N_3975,N_1967,N_1201);
nor U3976 (N_3976,N_759,N_67);
nand U3977 (N_3977,N_1608,N_16);
nor U3978 (N_3978,N_1143,N_1697);
nor U3979 (N_3979,N_1750,N_102);
nand U3980 (N_3980,N_316,N_486);
or U3981 (N_3981,N_166,N_1845);
nand U3982 (N_3982,N_762,N_1053);
xnor U3983 (N_3983,N_1116,N_206);
nand U3984 (N_3984,N_135,N_1132);
or U3985 (N_3985,N_1009,N_1885);
or U3986 (N_3986,N_852,N_804);
nand U3987 (N_3987,N_1317,N_1208);
and U3988 (N_3988,N_1821,N_1722);
and U3989 (N_3989,N_1654,N_960);
nand U3990 (N_3990,N_909,N_1252);
nor U3991 (N_3991,N_553,N_1545);
nand U3992 (N_3992,N_1838,N_745);
nand U3993 (N_3993,N_423,N_1123);
or U3994 (N_3994,N_467,N_797);
nand U3995 (N_3995,N_1692,N_783);
or U3996 (N_3996,N_1955,N_67);
and U3997 (N_3997,N_1084,N_1324);
nand U3998 (N_3998,N_1168,N_1911);
nor U3999 (N_3999,N_160,N_1616);
nor U4000 (N_4000,N_2691,N_3893);
and U4001 (N_4001,N_3935,N_2200);
nand U4002 (N_4002,N_3746,N_3003);
nor U4003 (N_4003,N_3250,N_3178);
or U4004 (N_4004,N_3433,N_3048);
nor U4005 (N_4005,N_3744,N_2354);
and U4006 (N_4006,N_3099,N_3999);
or U4007 (N_4007,N_3374,N_3730);
and U4008 (N_4008,N_3014,N_3550);
or U4009 (N_4009,N_3796,N_3964);
or U4010 (N_4010,N_2449,N_3174);
or U4011 (N_4011,N_2380,N_3287);
nor U4012 (N_4012,N_2226,N_3934);
xor U4013 (N_4013,N_2664,N_3850);
nor U4014 (N_4014,N_2580,N_2598);
or U4015 (N_4015,N_2543,N_3584);
or U4016 (N_4016,N_3232,N_3297);
nor U4017 (N_4017,N_3924,N_3764);
xor U4018 (N_4018,N_3337,N_2299);
or U4019 (N_4019,N_2532,N_2952);
or U4020 (N_4020,N_2926,N_2523);
nand U4021 (N_4021,N_2944,N_3668);
nand U4022 (N_4022,N_2044,N_2727);
nand U4023 (N_4023,N_2704,N_3299);
nor U4024 (N_4024,N_2234,N_3423);
nand U4025 (N_4025,N_2818,N_3139);
xor U4026 (N_4026,N_2512,N_2769);
nor U4027 (N_4027,N_2813,N_2486);
or U4028 (N_4028,N_3356,N_2981);
nand U4029 (N_4029,N_2963,N_3911);
or U4030 (N_4030,N_3036,N_2385);
nand U4031 (N_4031,N_3837,N_2622);
nor U4032 (N_4032,N_3150,N_3377);
and U4033 (N_4033,N_2029,N_2173);
nor U4034 (N_4034,N_2911,N_3741);
nand U4035 (N_4035,N_2966,N_3167);
nor U4036 (N_4036,N_3627,N_2329);
nand U4037 (N_4037,N_2849,N_2587);
nor U4038 (N_4038,N_3801,N_3624);
or U4039 (N_4039,N_2953,N_3005);
nor U4040 (N_4040,N_2368,N_3063);
and U4041 (N_4041,N_3520,N_3417);
nor U4042 (N_4042,N_3392,N_2897);
or U4043 (N_4043,N_3159,N_3756);
and U4044 (N_4044,N_3445,N_3515);
or U4045 (N_4045,N_3635,N_2726);
or U4046 (N_4046,N_2799,N_3107);
nor U4047 (N_4047,N_3110,N_3410);
nor U4048 (N_4048,N_2272,N_3858);
nand U4049 (N_4049,N_2005,N_2305);
or U4050 (N_4050,N_3002,N_3696);
and U4051 (N_4051,N_3636,N_3590);
nand U4052 (N_4052,N_2127,N_3630);
nand U4053 (N_4053,N_3658,N_3505);
or U4054 (N_4054,N_3838,N_2274);
or U4055 (N_4055,N_2714,N_2237);
nor U4056 (N_4056,N_2318,N_3484);
nand U4057 (N_4057,N_3200,N_2888);
or U4058 (N_4058,N_2974,N_2663);
and U4059 (N_4059,N_3702,N_2496);
and U4060 (N_4060,N_2035,N_3407);
nor U4061 (N_4061,N_2358,N_3517);
nand U4062 (N_4062,N_2960,N_2093);
nor U4063 (N_4063,N_3189,N_3751);
or U4064 (N_4064,N_2401,N_3739);
nor U4065 (N_4065,N_2141,N_3334);
or U4066 (N_4066,N_2099,N_3901);
nand U4067 (N_4067,N_3686,N_2770);
or U4068 (N_4068,N_2500,N_3710);
and U4069 (N_4069,N_2373,N_2348);
nand U4070 (N_4070,N_3884,N_3346);
nand U4071 (N_4071,N_2494,N_3214);
nor U4072 (N_4072,N_2201,N_3603);
nand U4073 (N_4073,N_2377,N_2690);
nand U4074 (N_4074,N_3195,N_2651);
and U4075 (N_4075,N_2781,N_2484);
or U4076 (N_4076,N_2505,N_3233);
or U4077 (N_4077,N_3643,N_3351);
and U4078 (N_4078,N_2702,N_3476);
nand U4079 (N_4079,N_3615,N_2865);
or U4080 (N_4080,N_3820,N_3817);
nor U4081 (N_4081,N_2748,N_3980);
or U4082 (N_4082,N_3875,N_3365);
or U4083 (N_4083,N_2140,N_2437);
or U4084 (N_4084,N_2294,N_3400);
nand U4085 (N_4085,N_3493,N_2495);
and U4086 (N_4086,N_3146,N_2232);
and U4087 (N_4087,N_2474,N_2681);
nor U4088 (N_4088,N_3712,N_3412);
and U4089 (N_4089,N_2236,N_3454);
nor U4090 (N_4090,N_2108,N_2519);
or U4091 (N_4091,N_2007,N_2961);
nand U4092 (N_4092,N_3951,N_3102);
and U4093 (N_4093,N_3946,N_2398);
and U4094 (N_4094,N_3667,N_2462);
and U4095 (N_4095,N_2788,N_3937);
or U4096 (N_4096,N_2737,N_3116);
nor U4097 (N_4097,N_3352,N_2261);
or U4098 (N_4098,N_3326,N_2107);
nor U4099 (N_4099,N_3275,N_3545);
nor U4100 (N_4100,N_3302,N_2446);
and U4101 (N_4101,N_3944,N_2003);
nor U4102 (N_4102,N_3810,N_3765);
and U4103 (N_4103,N_2216,N_3188);
or U4104 (N_4104,N_3121,N_2697);
or U4105 (N_4105,N_3008,N_3511);
and U4106 (N_4106,N_2665,N_3211);
or U4107 (N_4107,N_3463,N_3750);
and U4108 (N_4108,N_2732,N_2999);
and U4109 (N_4109,N_3570,N_3833);
nand U4110 (N_4110,N_2645,N_3776);
or U4111 (N_4111,N_3248,N_3539);
or U4112 (N_4112,N_2440,N_2508);
nor U4113 (N_4113,N_2939,N_3991);
or U4114 (N_4114,N_2822,N_3115);
or U4115 (N_4115,N_3502,N_2879);
nor U4116 (N_4116,N_2394,N_2555);
nand U4117 (N_4117,N_3580,N_2563);
or U4118 (N_4118,N_2086,N_2364);
nor U4119 (N_4119,N_3851,N_2076);
nor U4120 (N_4120,N_2477,N_2241);
nor U4121 (N_4121,N_2082,N_3191);
and U4122 (N_4122,N_3303,N_3819);
nand U4123 (N_4123,N_2956,N_3632);
and U4124 (N_4124,N_3784,N_3037);
nand U4125 (N_4125,N_2738,N_3728);
nand U4126 (N_4126,N_2103,N_2658);
nand U4127 (N_4127,N_3927,N_2488);
and U4128 (N_4128,N_2964,N_3821);
nor U4129 (N_4129,N_3525,N_3928);
nor U4130 (N_4130,N_3348,N_2632);
nor U4131 (N_4131,N_3140,N_2680);
or U4132 (N_4132,N_2682,N_2264);
nor U4133 (N_4133,N_3488,N_3706);
or U4134 (N_4134,N_2943,N_2672);
nor U4135 (N_4135,N_2202,N_2148);
nand U4136 (N_4136,N_3164,N_2758);
and U4137 (N_4137,N_2686,N_3568);
and U4138 (N_4138,N_2592,N_3129);
or U4139 (N_4139,N_3070,N_3916);
nor U4140 (N_4140,N_2233,N_3309);
nand U4141 (N_4141,N_3477,N_3874);
nand U4142 (N_4142,N_3359,N_2657);
nand U4143 (N_4143,N_2798,N_2612);
or U4144 (N_4144,N_2936,N_3390);
nor U4145 (N_4145,N_3754,N_3152);
nand U4146 (N_4146,N_2190,N_2835);
and U4147 (N_4147,N_3341,N_3300);
and U4148 (N_4148,N_3291,N_3194);
and U4149 (N_4149,N_2659,N_3905);
or U4150 (N_4150,N_3962,N_3384);
nand U4151 (N_4151,N_2608,N_2263);
nand U4152 (N_4152,N_2668,N_3637);
nor U4153 (N_4153,N_3677,N_2742);
or U4154 (N_4154,N_2594,N_2443);
nor U4155 (N_4155,N_2971,N_3700);
nand U4156 (N_4156,N_3006,N_2689);
nor U4157 (N_4157,N_3997,N_3331);
and U4158 (N_4158,N_2175,N_3717);
and U4159 (N_4159,N_3828,N_3599);
or U4160 (N_4160,N_2656,N_2938);
and U4161 (N_4161,N_3486,N_2650);
and U4162 (N_4162,N_3859,N_3576);
nand U4163 (N_4163,N_3544,N_3338);
and U4164 (N_4164,N_2010,N_2558);
or U4165 (N_4165,N_2641,N_2844);
nor U4166 (N_4166,N_3148,N_3797);
nand U4167 (N_4167,N_3362,N_2882);
or U4168 (N_4168,N_2574,N_2688);
nand U4169 (N_4169,N_2796,N_2239);
nor U4170 (N_4170,N_2203,N_2923);
and U4171 (N_4171,N_3715,N_2554);
nor U4172 (N_4172,N_3379,N_3205);
and U4173 (N_4173,N_2070,N_2642);
or U4174 (N_4174,N_2868,N_3687);
nor U4175 (N_4175,N_2420,N_2432);
nor U4176 (N_4176,N_2254,N_2471);
nor U4177 (N_4177,N_2589,N_2470);
nand U4178 (N_4178,N_3060,N_3518);
and U4179 (N_4179,N_2600,N_3665);
or U4180 (N_4180,N_3108,N_3732);
and U4181 (N_4181,N_2165,N_3202);
or U4182 (N_4182,N_3380,N_2230);
nand U4183 (N_4183,N_2766,N_3949);
nand U4184 (N_4184,N_3458,N_3221);
or U4185 (N_4185,N_3973,N_2791);
or U4186 (N_4186,N_3154,N_3906);
or U4187 (N_4187,N_2370,N_3721);
nand U4188 (N_4188,N_2840,N_3311);
nand U4189 (N_4189,N_2434,N_3333);
nor U4190 (N_4190,N_2772,N_2983);
and U4191 (N_4191,N_3674,N_2208);
and U4192 (N_4192,N_3530,N_2083);
nor U4193 (N_4193,N_2666,N_3323);
nand U4194 (N_4194,N_2694,N_3375);
or U4195 (N_4195,N_3039,N_2104);
nor U4196 (N_4196,N_3224,N_2564);
or U4197 (N_4197,N_2466,N_3990);
or U4198 (N_4198,N_2687,N_2814);
nand U4199 (N_4199,N_2307,N_3708);
nand U4200 (N_4200,N_3438,N_3761);
nor U4201 (N_4201,N_2097,N_3370);
or U4202 (N_4202,N_3807,N_3383);
or U4203 (N_4203,N_2899,N_3079);
and U4204 (N_4204,N_2246,N_2152);
or U4205 (N_4205,N_3013,N_2577);
xnor U4206 (N_4206,N_3832,N_3844);
and U4207 (N_4207,N_2638,N_3854);
nand U4208 (N_4208,N_2988,N_2937);
or U4209 (N_4209,N_3219,N_2605);
nand U4210 (N_4210,N_2809,N_3541);
nor U4211 (N_4211,N_3173,N_2615);
and U4212 (N_4212,N_3087,N_3434);
or U4213 (N_4213,N_2970,N_2625);
or U4214 (N_4214,N_3866,N_3342);
and U4215 (N_4215,N_2250,N_3718);
or U4216 (N_4216,N_3056,N_3082);
nor U4217 (N_4217,N_3912,N_3781);
nand U4218 (N_4218,N_3847,N_3314);
and U4219 (N_4219,N_3141,N_3109);
and U4220 (N_4220,N_2881,N_3157);
nand U4221 (N_4221,N_2187,N_2016);
or U4222 (N_4222,N_2800,N_3808);
nand U4223 (N_4223,N_3651,N_3019);
or U4224 (N_4224,N_3986,N_2343);
or U4225 (N_4225,N_2728,N_3888);
and U4226 (N_4226,N_3536,N_2074);
and U4227 (N_4227,N_2447,N_3669);
nor U4228 (N_4228,N_3881,N_2037);
nor U4229 (N_4229,N_3426,N_2479);
or U4230 (N_4230,N_2805,N_3491);
or U4231 (N_4231,N_3162,N_3397);
nor U4232 (N_4232,N_2597,N_3295);
and U4233 (N_4233,N_3245,N_3805);
nor U4234 (N_4234,N_2804,N_3578);
or U4235 (N_4235,N_3534,N_3085);
nand U4236 (N_4236,N_3408,N_3778);
and U4237 (N_4237,N_2174,N_3282);
nor U4238 (N_4238,N_3049,N_3938);
nor U4239 (N_4239,N_3894,N_3077);
and U4240 (N_4240,N_3596,N_2288);
nand U4241 (N_4241,N_2324,N_3614);
and U4242 (N_4242,N_2721,N_2215);
or U4243 (N_4243,N_2273,N_3605);
or U4244 (N_4244,N_2783,N_3126);
xor U4245 (N_4245,N_3274,N_3045);
and U4246 (N_4246,N_2040,N_3579);
and U4247 (N_4247,N_2206,N_3664);
xor U4248 (N_4248,N_3954,N_2538);
nand U4249 (N_4249,N_2993,N_2426);
or U4250 (N_4250,N_3285,N_2620);
and U4251 (N_4251,N_3465,N_2618);
nand U4252 (N_4252,N_2286,N_2795);
or U4253 (N_4253,N_2821,N_2493);
and U4254 (N_4254,N_3487,N_2359);
or U4255 (N_4255,N_2950,N_2321);
and U4256 (N_4256,N_3865,N_3831);
or U4257 (N_4257,N_2375,N_3914);
or U4258 (N_4258,N_2304,N_3293);
or U4259 (N_4259,N_3165,N_2541);
nor U4260 (N_4260,N_3824,N_3573);
or U4261 (N_4261,N_2012,N_2501);
nand U4262 (N_4262,N_2677,N_2147);
and U4263 (N_4263,N_2731,N_2907);
and U4264 (N_4264,N_2675,N_3207);
and U4265 (N_4265,N_3972,N_3294);
and U4266 (N_4266,N_2621,N_3500);
and U4267 (N_4267,N_3009,N_3093);
nor U4268 (N_4268,N_2276,N_2441);
nand U4269 (N_4269,N_2195,N_2958);
or U4270 (N_4270,N_3900,N_2701);
nand U4271 (N_4271,N_2513,N_2075);
or U4272 (N_4272,N_2736,N_2487);
or U4273 (N_4273,N_3197,N_2308);
or U4274 (N_4274,N_2160,N_2145);
and U4275 (N_4275,N_3829,N_2111);
nor U4276 (N_4276,N_2782,N_3507);
nor U4277 (N_4277,N_2674,N_2395);
nor U4278 (N_4278,N_2545,N_3646);
and U4279 (N_4279,N_3255,N_2703);
nor U4280 (N_4280,N_2906,N_3166);
nor U4281 (N_4281,N_2303,N_2894);
nand U4282 (N_4282,N_2717,N_3886);
and U4283 (N_4283,N_2266,N_3308);
and U4284 (N_4284,N_3478,N_2655);
nand U4285 (N_4285,N_3388,N_2604);
or U4286 (N_4286,N_2457,N_3187);
or U4287 (N_4287,N_3074,N_3519);
and U4288 (N_4288,N_3948,N_3853);
and U4289 (N_4289,N_3903,N_2542);
and U4290 (N_4290,N_2314,N_3033);
nor U4291 (N_4291,N_3089,N_3172);
nand U4292 (N_4292,N_3703,N_2480);
and U4293 (N_4293,N_2257,N_2196);
nand U4294 (N_4294,N_2602,N_2415);
or U4295 (N_4295,N_2311,N_2185);
nor U4296 (N_4296,N_3860,N_3548);
nand U4297 (N_4297,N_2403,N_2031);
nand U4298 (N_4298,N_2869,N_2713);
nor U4299 (N_4299,N_3325,N_3176);
or U4300 (N_4300,N_2948,N_3457);
and U4301 (N_4301,N_2718,N_3780);
and U4302 (N_4302,N_3435,N_3775);
or U4303 (N_4303,N_2749,N_3105);
xor U4304 (N_4304,N_3783,N_3527);
and U4305 (N_4305,N_3183,N_3594);
and U4306 (N_4306,N_2427,N_3405);
nand U4307 (N_4307,N_3406,N_2678);
nand U4308 (N_4308,N_2476,N_2180);
or U4309 (N_4309,N_2149,N_3034);
nor U4310 (N_4310,N_3225,N_3321);
nand U4311 (N_4311,N_3208,N_2861);
and U4312 (N_4312,N_2032,N_2371);
nor U4313 (N_4313,N_3184,N_2138);
nand U4314 (N_4314,N_2812,N_3145);
or U4315 (N_4315,N_2617,N_2131);
nand U4316 (N_4316,N_3025,N_2277);
xor U4317 (N_4317,N_3770,N_2928);
or U4318 (N_4318,N_3443,N_2159);
nand U4319 (N_4319,N_2503,N_2352);
nor U4320 (N_4320,N_2546,N_2864);
and U4321 (N_4321,N_3143,N_3030);
nor U4322 (N_4322,N_3798,N_2765);
and U4323 (N_4323,N_3621,N_2867);
or U4324 (N_4324,N_2699,N_3272);
and U4325 (N_4325,N_2134,N_3068);
nor U4326 (N_4326,N_3685,N_3069);
nand U4327 (N_4327,N_3723,N_3170);
nor U4328 (N_4328,N_3987,N_3942);
and U4329 (N_4329,N_2188,N_2309);
nand U4330 (N_4330,N_2862,N_2715);
or U4331 (N_4331,N_3332,N_2301);
or U4332 (N_4332,N_2064,N_2550);
or U4333 (N_4333,N_3998,N_2151);
or U4334 (N_4334,N_3349,N_2402);
nand U4335 (N_4335,N_2177,N_3830);
nor U4336 (N_4336,N_2839,N_3344);
or U4337 (N_4337,N_2036,N_3719);
and U4338 (N_4338,N_2918,N_2539);
or U4339 (N_4339,N_2285,N_3556);
or U4340 (N_4340,N_3779,N_2984);
nor U4341 (N_4341,N_3956,N_3595);
nand U4342 (N_4342,N_3679,N_3041);
or U4343 (N_4343,N_2472,N_3062);
and U4344 (N_4344,N_3575,N_3790);
nor U4345 (N_4345,N_3076,N_3038);
nor U4346 (N_4346,N_2786,N_3451);
and U4347 (N_4347,N_3235,N_3601);
nand U4348 (N_4348,N_3788,N_2062);
and U4349 (N_4349,N_2310,N_2959);
or U4350 (N_4350,N_3524,N_2312);
nor U4351 (N_4351,N_3051,N_3895);
and U4352 (N_4352,N_2586,N_2584);
nand U4353 (N_4353,N_2456,N_3574);
and U4354 (N_4354,N_3023,N_2755);
nand U4355 (N_4355,N_2848,N_2629);
or U4356 (N_4356,N_2172,N_3683);
or U4357 (N_4357,N_3742,N_3566);
nand U4358 (N_4358,N_3609,N_2431);
and U4359 (N_4359,N_2979,N_3538);
and U4360 (N_4360,N_3021,N_3504);
or U4361 (N_4361,N_2350,N_3876);
or U4362 (N_4362,N_2824,N_2968);
xor U4363 (N_4363,N_2876,N_2313);
nor U4364 (N_4364,N_2850,N_3474);
nor U4365 (N_4365,N_3470,N_3498);
nand U4366 (N_4366,N_3823,N_2391);
or U4367 (N_4367,N_3549,N_2199);
and U4368 (N_4368,N_2410,N_3918);
nand U4369 (N_4369,N_3880,N_3149);
nand U4370 (N_4370,N_2381,N_3835);
or U4371 (N_4371,N_3606,N_2213);
or U4372 (N_4372,N_2113,N_3055);
or U4373 (N_4373,N_3695,N_3215);
nor U4374 (N_4374,N_2019,N_2467);
and U4375 (N_4375,N_3136,N_3743);
and U4376 (N_4376,N_2643,N_2679);
or U4377 (N_4377,N_3909,N_2808);
or U4378 (N_4378,N_2549,N_3506);
or U4379 (N_4379,N_3124,N_2771);
or U4380 (N_4380,N_3825,N_3863);
and U4381 (N_4381,N_3398,N_3608);
xor U4382 (N_4382,N_2349,N_2300);
or U4383 (N_4383,N_2435,N_2756);
or U4384 (N_4384,N_2745,N_3872);
or U4385 (N_4385,N_2453,N_2957);
nor U4386 (N_4386,N_3571,N_3612);
nand U4387 (N_4387,N_2802,N_3993);
and U4388 (N_4388,N_2551,N_3662);
or U4389 (N_4389,N_3482,N_2252);
and U4390 (N_4390,N_2763,N_2183);
nand U4391 (N_4391,N_3747,N_3492);
xnor U4392 (N_4392,N_3616,N_2773);
nand U4393 (N_4393,N_3252,N_3192);
or U4394 (N_4394,N_2890,N_2034);
nor U4395 (N_4395,N_3787,N_3682);
or U4396 (N_4396,N_3771,N_3713);
or U4397 (N_4397,N_3024,N_3193);
or U4398 (N_4398,N_3989,N_2369);
xor U4399 (N_4399,N_3620,N_3289);
nand U4400 (N_4400,N_2916,N_3276);
and U4401 (N_4401,N_2123,N_3581);
nor U4402 (N_4402,N_2855,N_2967);
or U4403 (N_4403,N_2038,N_2338);
or U4404 (N_4404,N_3422,N_2017);
nor U4405 (N_4405,N_3926,N_2933);
and U4406 (N_4406,N_2150,N_3846);
and U4407 (N_4407,N_2667,N_3726);
xnor U4408 (N_4408,N_3597,N_2117);
or U4409 (N_4409,N_2499,N_2709);
nand U4410 (N_4410,N_2379,N_2852);
nand U4411 (N_4411,N_3652,N_3315);
or U4412 (N_4412,N_2874,N_2945);
and U4413 (N_4413,N_2225,N_2009);
or U4414 (N_4414,N_2290,N_2826);
nand U4415 (N_4415,N_2041,N_2877);
and U4416 (N_4416,N_3114,N_2063);
xor U4417 (N_4417,N_2105,N_3922);
and U4418 (N_4418,N_2815,N_2198);
nand U4419 (N_4419,N_2739,N_3675);
nor U4420 (N_4420,N_2774,N_2516);
nor U4421 (N_4421,N_2452,N_2684);
nor U4422 (N_4422,N_2296,N_3748);
and U4423 (N_4423,N_3613,N_2298);
and U4424 (N_4424,N_2919,N_2191);
nor U4425 (N_4425,N_2607,N_2652);
nor U4426 (N_4426,N_2644,N_3284);
or U4427 (N_4427,N_2222,N_2553);
nand U4428 (N_4428,N_2520,N_2413);
and U4429 (N_4429,N_3569,N_2167);
and U4430 (N_4430,N_2790,N_2161);
and U4431 (N_4431,N_3218,N_2363);
and U4432 (N_4432,N_2081,N_3681);
and U4433 (N_4433,N_2414,N_3100);
nor U4434 (N_4434,N_3182,N_2224);
nor U4435 (N_4435,N_2946,N_3080);
or U4436 (N_4436,N_3542,N_3064);
nor U4437 (N_4437,N_3011,N_2166);
nand U4438 (N_4438,N_3420,N_3058);
and U4439 (N_4439,N_2834,N_3968);
nand U4440 (N_4440,N_3103,N_3494);
or U4441 (N_4441,N_3104,N_2760);
or U4442 (N_4442,N_2863,N_3057);
and U4443 (N_4443,N_2378,N_3862);
or U4444 (N_4444,N_3401,N_2634);
nor U4445 (N_4445,N_3396,N_2535);
nand U4446 (N_4446,N_2448,N_3631);
and U4447 (N_4447,N_3199,N_3970);
or U4448 (N_4448,N_2220,N_2339);
or U4449 (N_4449,N_2048,N_3971);
xor U4450 (N_4450,N_3249,N_3084);
nand U4451 (N_4451,N_3985,N_2552);
or U4452 (N_4452,N_3065,N_2859);
nor U4453 (N_4453,N_2015,N_3251);
nand U4454 (N_4454,N_2575,N_2837);
or U4455 (N_4455,N_2750,N_2857);
or U4456 (N_4456,N_2954,N_2836);
or U4457 (N_4457,N_2540,N_3204);
and U4458 (N_4458,N_3588,N_2047);
nand U4459 (N_4459,N_2833,N_2235);
or U4460 (N_4460,N_3757,N_3231);
or U4461 (N_4461,N_3020,N_3607);
nand U4462 (N_4462,N_3995,N_2482);
nor U4463 (N_4463,N_3586,N_3424);
nand U4464 (N_4464,N_3345,N_3591);
or U4465 (N_4465,N_3016,N_2210);
and U4466 (N_4466,N_3256,N_3442);
nor U4467 (N_4467,N_3091,N_2640);
nor U4468 (N_4468,N_2171,N_3512);
nand U4469 (N_4469,N_3304,N_2982);
nand U4470 (N_4470,N_3054,N_3793);
nor U4471 (N_4471,N_3887,N_2109);
nand U4472 (N_4472,N_2588,N_2114);
or U4473 (N_4473,N_2705,N_3305);
and U4474 (N_4474,N_3217,N_2884);
and U4475 (N_4475,N_2399,N_3263);
nor U4476 (N_4476,N_3130,N_2898);
and U4477 (N_4477,N_3768,N_2716);
and U4478 (N_4478,N_3125,N_2436);
or U4479 (N_4479,N_2875,N_3532);
xor U4480 (N_4480,N_2570,N_3856);
nand U4481 (N_4481,N_2854,N_2955);
and U4482 (N_4482,N_2920,N_3663);
and U4483 (N_4483,N_3415,N_3240);
nor U4484 (N_4484,N_2267,N_3514);
nor U4485 (N_4485,N_2524,N_2468);
nand U4486 (N_4486,N_2614,N_2061);
nor U4487 (N_4487,N_3095,N_3932);
nand U4488 (N_4488,N_3804,N_3769);
or U4489 (N_4489,N_3690,N_3269);
nand U4490 (N_4490,N_2055,N_3587);
and U4491 (N_4491,N_2491,N_3280);
and U4492 (N_4492,N_3450,N_2930);
nand U4493 (N_4493,N_3959,N_2977);
nand U4494 (N_4494,N_2011,N_3228);
or U4495 (N_4495,N_2280,N_3158);
nor U4496 (N_4496,N_3794,N_3032);
nand U4497 (N_4497,N_3509,N_2387);
nor U4498 (N_4498,N_2393,N_3961);
or U4499 (N_4499,N_3873,N_3447);
or U4500 (N_4500,N_2683,N_2430);
nand U4501 (N_4501,N_2673,N_2376);
and U4502 (N_4502,N_3444,N_3448);
and U4503 (N_4503,N_2170,N_2613);
and U4504 (N_4504,N_3963,N_2810);
and U4505 (N_4505,N_3151,N_3237);
or U4506 (N_4506,N_2408,N_3890);
nor U4507 (N_4507,N_2935,N_2021);
and U4508 (N_4508,N_2412,N_2473);
nor U4509 (N_4509,N_3393,N_2383);
nor U4510 (N_4510,N_2628,N_3967);
nand U4511 (N_4511,N_3262,N_3720);
nand U4512 (N_4512,N_2469,N_2027);
nor U4513 (N_4513,N_3815,N_2619);
or U4514 (N_4514,N_3899,N_2465);
nor U4515 (N_4515,N_2492,N_2909);
nand U4516 (N_4516,N_2806,N_2685);
nand U4517 (N_4517,N_3010,N_2255);
nand U4518 (N_4518,N_3106,N_2088);
or U4519 (N_4519,N_2843,N_2284);
xor U4520 (N_4520,N_2293,N_3740);
and U4521 (N_4521,N_2351,N_3361);
nand U4522 (N_4522,N_2018,N_2382);
nor U4523 (N_4523,N_3456,N_3322);
or U4524 (N_4524,N_2461,N_3112);
or U4525 (N_4525,N_2347,N_3626);
nand U4526 (N_4526,N_3655,N_3622);
nand U4527 (N_4527,N_3117,N_3421);
and U4528 (N_4528,N_2022,N_2325);
or U4529 (N_4529,N_3697,N_3210);
and U4530 (N_4530,N_2596,N_2828);
and U4531 (N_4531,N_2240,N_3567);
xnor U4532 (N_4532,N_2458,N_2985);
nand U4533 (N_4533,N_2744,N_2606);
and U4534 (N_4534,N_2289,N_2342);
or U4535 (N_4535,N_3220,N_3072);
or U4536 (N_4536,N_3698,N_2767);
nand U4537 (N_4537,N_3028,N_3044);
and U4538 (N_4538,N_2326,N_3848);
nand U4539 (N_4539,N_3602,N_3313);
and U4540 (N_4540,N_3047,N_3460);
and U4541 (N_4541,N_3226,N_2856);
or U4542 (N_4542,N_3371,N_3841);
nor U4543 (N_4543,N_3671,N_3246);
nor U4544 (N_4544,N_2566,N_2921);
xor U4545 (N_4545,N_3733,N_2249);
and U4546 (N_4546,N_3098,N_3119);
or U4547 (N_4547,N_3814,N_2302);
nor U4548 (N_4548,N_2217,N_3931);
nand U4549 (N_4549,N_2507,N_3547);
nand U4550 (N_4550,N_2102,N_2259);
and U4551 (N_4551,N_3811,N_3081);
nor U4552 (N_4552,N_2002,N_3449);
nand U4553 (N_4553,N_2039,N_3857);
and U4554 (N_4554,N_3324,N_3638);
nand U4555 (N_4555,N_3554,N_3660);
and U4556 (N_4556,N_3185,N_2846);
nor U4557 (N_4557,N_2438,N_2322);
and U4558 (N_4558,N_3623,N_2209);
or U4559 (N_4559,N_3941,N_2231);
nand U4560 (N_4560,N_3923,N_3722);
or U4561 (N_4561,N_2404,N_3919);
nand U4562 (N_4562,N_2428,N_3882);
and U4563 (N_4563,N_3977,N_2156);
nand U4564 (N_4564,N_3843,N_2842);
or U4565 (N_4565,N_3701,N_2975);
xor U4566 (N_4566,N_2058,N_3773);
nor U4567 (N_4567,N_2845,N_3917);
or U4568 (N_4568,N_2490,N_2424);
and U4569 (N_4569,N_3168,N_3755);
nand U4570 (N_4570,N_3480,N_3403);
or U4571 (N_4571,N_2725,N_3521);
and U4572 (N_4572,N_3984,N_2292);
or U4573 (N_4573,N_3799,N_3339);
and U4574 (N_4574,N_3716,N_3974);
nor U4575 (N_4575,N_3558,N_2902);
and U4576 (N_4576,N_2889,N_2695);
nor U4577 (N_4577,N_2355,N_3475);
and U4578 (N_4578,N_3593,N_3767);
or U4579 (N_4579,N_2268,N_2593);
or U4580 (N_4580,N_2211,N_3113);
nor U4581 (N_4581,N_2578,N_3050);
nand U4582 (N_4582,N_3446,N_2052);
xor U4583 (N_4583,N_3335,N_3628);
and U4584 (N_4584,N_2319,N_3611);
and U4585 (N_4585,N_3529,N_2297);
and U4586 (N_4586,N_3483,N_2636);
or U4587 (N_4587,N_3431,N_3869);
or U4588 (N_4588,N_2595,N_2576);
nand U4589 (N_4589,N_3203,N_2256);
nand U4590 (N_4590,N_3261,N_2518);
nor U4591 (N_4591,N_3138,N_2841);
and U4592 (N_4592,N_3306,N_3589);
and U4593 (N_4593,N_3656,N_3840);
and U4594 (N_4594,N_3413,N_3540);
nor U4595 (N_4595,N_3510,N_3709);
xnor U4596 (N_4596,N_2819,N_3577);
and U4597 (N_4597,N_2228,N_3642);
or U4598 (N_4598,N_3802,N_3496);
nor U4599 (N_4599,N_3355,N_3684);
or U4600 (N_4600,N_3640,N_2901);
or U4601 (N_4601,N_3598,N_2353);
nor U4602 (N_4602,N_3040,N_2942);
nand U4603 (N_4603,N_3389,N_2511);
and U4604 (N_4604,N_3353,N_2416);
nand U4605 (N_4605,N_2459,N_3290);
and U4606 (N_4606,N_2219,N_3001);
or U4607 (N_4607,N_2085,N_2327);
nor U4608 (N_4608,N_2336,N_2253);
and U4609 (N_4609,N_2825,N_2193);
and U4610 (N_4610,N_2823,N_2556);
or U4611 (N_4611,N_2853,N_3485);
and U4612 (N_4612,N_2418,N_2517);
nor U4613 (N_4613,N_2262,N_2847);
nand U4614 (N_4614,N_3915,N_3727);
and U4615 (N_4615,N_2181,N_3913);
nand U4616 (N_4616,N_3693,N_3891);
or U4617 (N_4617,N_3976,N_3639);
nand U4618 (N_4618,N_2820,N_2013);
nand U4619 (N_4619,N_3849,N_3633);
nor U4620 (N_4620,N_2135,N_3357);
and U4621 (N_4621,N_3436,N_2747);
and U4622 (N_4622,N_2972,N_2066);
nand U4623 (N_4623,N_3822,N_2116);
nor U4624 (N_4624,N_2077,N_2335);
nand U4625 (N_4625,N_2278,N_2084);
nand U4626 (N_4626,N_3186,N_2078);
or U4627 (N_4627,N_2761,N_3546);
and U4628 (N_4628,N_2388,N_3513);
nor U4629 (N_4629,N_2929,N_3259);
nand U4630 (N_4630,N_3229,N_3947);
or U4631 (N_4631,N_2992,N_2094);
nand U4632 (N_4632,N_2720,N_3265);
nor U4633 (N_4633,N_2637,N_2433);
nor U4634 (N_4634,N_2860,N_2711);
and U4635 (N_4635,N_3969,N_3645);
or U4636 (N_4636,N_3239,N_3503);
and U4637 (N_4637,N_2729,N_2671);
nor U4638 (N_4638,N_3759,N_3391);
or U4639 (N_4639,N_2947,N_2573);
or U4640 (N_4640,N_3439,N_2707);
nand U4641 (N_4641,N_2421,N_3827);
or U4642 (N_4642,N_3583,N_3992);
and U4643 (N_4643,N_2973,N_3553);
nor U4644 (N_4644,N_2561,N_2050);
or U4645 (N_4645,N_2419,N_3531);
nand U4646 (N_4646,N_3175,N_2754);
nand U4647 (N_4647,N_3092,N_3267);
nor U4648 (N_4648,N_2128,N_2451);
nand U4649 (N_4649,N_3097,N_2248);
and U4650 (N_4650,N_2793,N_2633);
nand U4651 (N_4651,N_3160,N_3067);
or U4652 (N_4652,N_2153,N_2186);
and U4653 (N_4653,N_2986,N_2091);
or U4654 (N_4654,N_3270,N_2125);
or U4655 (N_4655,N_2777,N_3046);
and U4656 (N_4656,N_2178,N_2531);
nor U4657 (N_4657,N_2000,N_2184);
and U4658 (N_4658,N_2341,N_2242);
and U4659 (N_4659,N_2356,N_3387);
or U4660 (N_4660,N_2635,N_3752);
or U4661 (N_4661,N_3135,N_3707);
nand U4662 (N_4662,N_2144,N_3236);
nor U4663 (N_4663,N_2056,N_3271);
or U4664 (N_4664,N_3473,N_2572);
or U4665 (N_4665,N_3366,N_3132);
nand U4666 (N_4666,N_3111,N_3327);
and U4667 (N_4667,N_3404,N_3704);
nand U4668 (N_4668,N_3729,N_2417);
nor U4669 (N_4669,N_2155,N_3216);
and U4670 (N_4670,N_3242,N_2481);
nor U4671 (N_4671,N_2214,N_2776);
or U4672 (N_4672,N_3292,N_3641);
or U4673 (N_4673,N_2162,N_2789);
or U4674 (N_4674,N_2559,N_2397);
nor U4675 (N_4675,N_3198,N_2475);
nor U4676 (N_4676,N_3792,N_3268);
xor U4677 (N_4677,N_2759,N_2332);
nor U4678 (N_4678,N_2182,N_2143);
or U4679 (N_4679,N_3427,N_3430);
nor U4680 (N_4680,N_3118,N_2411);
or U4681 (N_4681,N_2400,N_3254);
nor U4682 (N_4682,N_3562,N_2751);
or U4683 (N_4683,N_3350,N_2934);
or U4684 (N_4684,N_3889,N_3083);
nor U4685 (N_4685,N_2719,N_3711);
and U4686 (N_4686,N_3499,N_3774);
nand U4687 (N_4687,N_3604,N_3260);
nand U4688 (N_4688,N_2316,N_2030);
nand U4689 (N_4689,N_2654,N_3360);
nor U4690 (N_4690,N_2639,N_2265);
or U4691 (N_4691,N_2908,N_2914);
xnor U4692 (N_4692,N_3625,N_3310);
and U4693 (N_4693,N_3061,N_2792);
nor U4694 (N_4694,N_2941,N_3161);
nor U4695 (N_4695,N_2827,N_2372);
nand U4696 (N_4696,N_3378,N_2154);
and U4697 (N_4697,N_3319,N_2892);
and U4698 (N_4698,N_2797,N_3921);
nor U4699 (N_4699,N_3565,N_3481);
or U4700 (N_4700,N_2251,N_2247);
or U4701 (N_4701,N_2390,N_3737);
or U4702 (N_4702,N_2315,N_2871);
nor U4703 (N_4703,N_2940,N_2653);
nand U4704 (N_4704,N_3957,N_3206);
nor U4705 (N_4705,N_3592,N_2976);
or U4706 (N_4706,N_2647,N_2506);
and U4707 (N_4707,N_3834,N_3127);
and U4708 (N_4708,N_3273,N_3714);
or U4709 (N_4709,N_3806,N_3952);
or U4710 (N_4710,N_3373,N_2623);
and U4711 (N_4711,N_3133,N_2124);
nand U4712 (N_4712,N_2042,N_3409);
nor U4713 (N_4713,N_2537,N_2194);
nor U4714 (N_4714,N_3031,N_3312);
nor U4715 (N_4715,N_3812,N_2344);
nor U4716 (N_4716,N_2396,N_3610);
and U4717 (N_4717,N_2912,N_3930);
nand U4718 (N_4718,N_3247,N_2169);
nor U4719 (N_4719,N_2026,N_2360);
nand U4720 (N_4720,N_3120,N_2460);
or U4721 (N_4721,N_3318,N_3266);
nor U4722 (N_4722,N_2829,N_2891);
nor U4723 (N_4723,N_3369,N_3777);
and U4724 (N_4724,N_3425,N_3555);
or U4725 (N_4725,N_2407,N_2115);
or U4726 (N_4726,N_2080,N_3381);
nor U4727 (N_4727,N_2006,N_3018);
nor U4728 (N_4728,N_2092,N_2095);
and U4729 (N_4729,N_2004,N_2096);
nand U4730 (N_4730,N_2547,N_3101);
and U4731 (N_4731,N_3134,N_3559);
or U4732 (N_4732,N_3459,N_2176);
and U4733 (N_4733,N_2994,N_2260);
nand U4734 (N_4734,N_3004,N_3661);
and U4735 (N_4735,N_3177,N_3960);
or U4736 (N_4736,N_2698,N_2014);
or U4737 (N_4737,N_3885,N_3920);
nand U4738 (N_4738,N_3416,N_2275);
nor U4739 (N_4739,N_2662,N_2069);
and U4740 (N_4740,N_3340,N_2780);
nor U4741 (N_4741,N_3760,N_2965);
nor U4742 (N_4742,N_2295,N_2627);
or U4743 (N_4743,N_2227,N_3852);
nor U4744 (N_4744,N_2483,N_2830);
nor U4745 (N_4745,N_2345,N_2870);
nor U4746 (N_4746,N_2464,N_3196);
nor U4747 (N_4747,N_2059,N_3877);
nand U4748 (N_4748,N_3898,N_2616);
nor U4749 (N_4749,N_2450,N_3015);
or U4750 (N_4750,N_2603,N_3758);
or U4751 (N_4751,N_2885,N_2049);
nor U4752 (N_4752,N_3762,N_3012);
or U4753 (N_4753,N_3745,N_2157);
nor U4754 (N_4754,N_3738,N_3864);
or U4755 (N_4755,N_2271,N_3736);
nor U4756 (N_4756,N_3227,N_3533);
and U4757 (N_4757,N_2803,N_3418);
nor U4758 (N_4758,N_2873,N_2710);
and U4759 (N_4759,N_3836,N_2001);
xor U4760 (N_4760,N_3557,N_2676);
nor U4761 (N_4761,N_2526,N_2136);
or U4762 (N_4762,N_2996,N_3213);
nand U4763 (N_4763,N_3489,N_3878);
and U4764 (N_4764,N_3670,N_3472);
nor U4765 (N_4765,N_3301,N_3386);
nor U4766 (N_4766,N_2611,N_2498);
and U4767 (N_4767,N_3088,N_2454);
xor U4768 (N_4768,N_2357,N_2886);
nand U4769 (N_4769,N_3955,N_3563);
nor U4770 (N_4770,N_2529,N_3734);
nand U4771 (N_4771,N_3634,N_3528);
nor U4772 (N_4772,N_3966,N_2567);
nand U4773 (N_4773,N_2023,N_3399);
and U4774 (N_4774,N_3654,N_3094);
nand U4775 (N_4775,N_3364,N_3908);
or U4776 (N_4776,N_3657,N_2624);
and U4777 (N_4777,N_2238,N_2661);
nand U4778 (N_4778,N_2741,N_2980);
xor U4779 (N_4779,N_2591,N_3336);
or U4780 (N_4780,N_2569,N_3678);
or U4781 (N_4781,N_3979,N_2243);
nand U4782 (N_4782,N_3910,N_2910);
nand U4783 (N_4783,N_3329,N_3394);
or U4784 (N_4784,N_3179,N_3653);
or U4785 (N_4785,N_3142,N_3497);
nor U4786 (N_4786,N_3897,N_2340);
nor U4787 (N_4787,N_3800,N_3749);
nand U4788 (N_4788,N_2425,N_3994);
or U4789 (N_4789,N_3982,N_3816);
or U4790 (N_4790,N_2168,N_3672);
or U4791 (N_4791,N_3035,N_3153);
nand U4792 (N_4792,N_2872,N_3561);
and U4793 (N_4793,N_3791,N_2204);
nand U4794 (N_4794,N_2073,N_2544);
or U4795 (N_4795,N_3288,N_2794);
nand U4796 (N_4796,N_3543,N_3223);
nand U4797 (N_4797,N_2333,N_3156);
and U4798 (N_4798,N_3650,N_3789);
nor U4799 (N_4799,N_3316,N_2337);
and U4800 (N_4800,N_3253,N_3372);
and U4801 (N_4801,N_2205,N_3731);
or U4802 (N_4802,N_2346,N_2100);
or U4803 (N_4803,N_3871,N_2089);
or U4804 (N_4804,N_2648,N_3086);
and U4805 (N_4805,N_2579,N_2832);
or U4806 (N_4806,N_3516,N_3868);
or U4807 (N_4807,N_2087,N_2670);
nor U4808 (N_4808,N_3147,N_2112);
nor U4809 (N_4809,N_3059,N_3879);
or U4810 (N_4810,N_3441,N_2568);
nand U4811 (N_4811,N_2525,N_2122);
and U4812 (N_4812,N_2858,N_2051);
and U4813 (N_4813,N_3735,N_2931);
or U4814 (N_4814,N_3075,N_2392);
and U4815 (N_4815,N_3155,N_3981);
nor U4816 (N_4816,N_2978,N_3786);
xor U4817 (N_4817,N_3042,N_3238);
nor U4818 (N_4818,N_2565,N_3466);
or U4819 (N_4819,N_2444,N_2054);
nor U4820 (N_4820,N_3978,N_2053);
or U4821 (N_4821,N_2212,N_2692);
and U4822 (N_4822,N_2179,N_2028);
xor U4823 (N_4823,N_3892,N_2723);
nor U4824 (N_4824,N_2764,N_2962);
and U4825 (N_4825,N_2548,N_2712);
or U4826 (N_4826,N_2463,N_2478);
or U4827 (N_4827,N_3552,N_2609);
nand U4828 (N_4828,N_2132,N_2158);
nor U4829 (N_4829,N_2838,N_2801);
nor U4830 (N_4830,N_2880,N_3950);
or U4831 (N_4831,N_2269,N_2646);
nor U4832 (N_4832,N_2455,N_3842);
nor U4833 (N_4833,N_3385,N_3222);
or U4834 (N_4834,N_2904,N_3122);
or U4835 (N_4835,N_2334,N_3896);
or U4836 (N_4836,N_3171,N_2536);
nand U4837 (N_4837,N_3181,N_2101);
nand U4838 (N_4838,N_3241,N_3724);
or U4839 (N_4839,N_3163,N_2229);
or U4840 (N_4840,N_3395,N_3123);
and U4841 (N_4841,N_2816,N_2733);
and U4842 (N_4842,N_3096,N_2146);
nor U4843 (N_4843,N_2068,N_3347);
nand U4844 (N_4844,N_3467,N_3522);
nor U4845 (N_4845,N_3564,N_2583);
nand U4846 (N_4846,N_2775,N_3867);
nor U4847 (N_4847,N_2932,N_3953);
or U4848 (N_4848,N_3725,N_2660);
and U4849 (N_4849,N_2905,N_2057);
or U4850 (N_4850,N_2118,N_2601);
nand U4851 (N_4851,N_3560,N_3861);
nor U4852 (N_4852,N_3772,N_3988);
and U4853 (N_4853,N_3234,N_3753);
or U4854 (N_4854,N_3330,N_3462);
or U4855 (N_4855,N_3617,N_3939);
or U4856 (N_4856,N_2406,N_2706);
and U4857 (N_4857,N_3965,N_2245);
and U4858 (N_4858,N_2024,N_2033);
and U4859 (N_4859,N_3902,N_2126);
nand U4860 (N_4860,N_2365,N_3453);
nor U4861 (N_4861,N_2991,N_3688);
nand U4862 (N_4862,N_3090,N_3845);
or U4863 (N_4863,N_2331,N_2560);
or U4864 (N_4864,N_3526,N_2757);
or U4865 (N_4865,N_3537,N_3464);
and U4866 (N_4866,N_2696,N_2903);
nand U4867 (N_4867,N_3975,N_2895);
and U4868 (N_4868,N_2367,N_3414);
nand U4869 (N_4869,N_3461,N_3286);
nor U4870 (N_4870,N_2197,N_3257);
or U4871 (N_4871,N_2090,N_3940);
nand U4872 (N_4872,N_2522,N_2752);
nor U4873 (N_4873,N_3307,N_3666);
or U4874 (N_4874,N_3468,N_3680);
nor U4875 (N_4875,N_3278,N_2323);
and U4876 (N_4876,N_3943,N_2025);
nor U4877 (N_4877,N_3958,N_3209);
or U4878 (N_4878,N_2708,N_3904);
nand U4879 (N_4879,N_2221,N_2787);
nor U4880 (N_4880,N_3479,N_2405);
nand U4881 (N_4881,N_2735,N_3363);
and U4882 (N_4882,N_2384,N_2163);
nor U4883 (N_4883,N_2366,N_3452);
nor U4884 (N_4884,N_2361,N_2582);
and U4885 (N_4885,N_2283,N_2534);
nand U4886 (N_4886,N_3298,N_2060);
or U4887 (N_4887,N_3699,N_2071);
and U4888 (N_4888,N_2883,N_2509);
nor U4889 (N_4889,N_3705,N_3907);
and U4890 (N_4890,N_2409,N_2927);
nand U4891 (N_4891,N_3201,N_3279);
or U4892 (N_4892,N_2223,N_2008);
nor U4893 (N_4893,N_2362,N_3676);
or U4894 (N_4894,N_3659,N_3870);
nor U4895 (N_4895,N_2142,N_2374);
or U4896 (N_4896,N_3382,N_3455);
nand U4897 (N_4897,N_3619,N_2504);
or U4898 (N_4898,N_2386,N_3582);
or U4899 (N_4899,N_2098,N_3689);
and U4900 (N_4900,N_3429,N_2740);
and U4901 (N_4901,N_3402,N_2866);
and U4902 (N_4902,N_3813,N_2599);
and U4903 (N_4903,N_2306,N_2485);
nor U4904 (N_4904,N_2527,N_2164);
xnor U4905 (N_4905,N_2807,N_2987);
or U4906 (N_4906,N_2998,N_3600);
nand U4907 (N_4907,N_2389,N_2502);
nor U4908 (N_4908,N_3945,N_3523);
nand U4909 (N_4909,N_3053,N_3296);
nor U4910 (N_4910,N_2328,N_2878);
or U4911 (N_4911,N_3144,N_2320);
nor U4912 (N_4912,N_3230,N_3432);
nand U4913 (N_4913,N_2120,N_2768);
or U4914 (N_4914,N_2072,N_2442);
or U4915 (N_4915,N_2207,N_2626);
nand U4916 (N_4916,N_3983,N_2045);
or U4917 (N_4917,N_2445,N_3283);
or U4918 (N_4918,N_2046,N_2258);
nand U4919 (N_4919,N_2557,N_2137);
or U4920 (N_4920,N_3066,N_3029);
or U4921 (N_4921,N_2610,N_3649);
or U4922 (N_4922,N_2590,N_3212);
nand U4923 (N_4923,N_2133,N_3763);
and U4924 (N_4924,N_3766,N_2900);
and U4925 (N_4925,N_3803,N_2043);
nor U4926 (N_4926,N_3629,N_2291);
and U4927 (N_4927,N_2631,N_3358);
nand U4928 (N_4928,N_3328,N_2106);
or U4929 (N_4929,N_2244,N_2917);
and U4930 (N_4930,N_3437,N_3320);
nor U4931 (N_4931,N_2110,N_2121);
and U4932 (N_4932,N_2915,N_3495);
nand U4933 (N_4933,N_3190,N_3883);
or U4934 (N_4934,N_2785,N_2510);
and U4935 (N_4935,N_2817,N_2317);
or U4936 (N_4936,N_2533,N_3073);
and U4937 (N_4937,N_3354,N_3017);
and U4938 (N_4938,N_3264,N_2649);
nand U4939 (N_4939,N_2734,N_2020);
nand U4940 (N_4940,N_3243,N_3000);
and U4941 (N_4941,N_3137,N_3839);
nor U4942 (N_4942,N_2630,N_3572);
nor U4943 (N_4943,N_2489,N_2784);
and U4944 (N_4944,N_2887,N_3648);
or U4945 (N_4945,N_3535,N_2079);
nor U4946 (N_4946,N_2521,N_3419);
nor U4947 (N_4947,N_2913,N_3647);
nor U4948 (N_4948,N_2119,N_2189);
or U4949 (N_4949,N_2951,N_3809);
nand U4950 (N_4950,N_2811,N_2995);
nor U4951 (N_4951,N_3007,N_3376);
nand U4952 (N_4952,N_3936,N_2693);
or U4953 (N_4953,N_3258,N_2439);
xnor U4954 (N_4954,N_2778,N_3440);
nand U4955 (N_4955,N_2514,N_3933);
and U4956 (N_4956,N_3022,N_2282);
and U4957 (N_4957,N_2423,N_3128);
xnor U4958 (N_4958,N_3367,N_3673);
nand U4959 (N_4959,N_3644,N_3078);
nand U4960 (N_4960,N_3691,N_3052);
or U4961 (N_4961,N_2722,N_3317);
nor U4962 (N_4962,N_2779,N_2724);
nand U4963 (N_4963,N_2730,N_2218);
nor U4964 (N_4964,N_3692,N_3501);
and U4965 (N_4965,N_3782,N_3244);
nor U4966 (N_4966,N_2192,N_2571);
nor U4967 (N_4967,N_3469,N_3281);
xor U4968 (N_4968,N_3585,N_3551);
nor U4969 (N_4969,N_2743,N_2515);
or U4970 (N_4970,N_2753,N_2129);
nand U4971 (N_4971,N_2287,N_2279);
nand U4972 (N_4972,N_2969,N_3277);
nor U4973 (N_4973,N_3343,N_3180);
or U4974 (N_4974,N_2949,N_3490);
or U4975 (N_4975,N_2989,N_3826);
or U4976 (N_4976,N_3929,N_2669);
or U4977 (N_4977,N_3694,N_3855);
nor U4978 (N_4978,N_2700,N_2997);
and U4979 (N_4979,N_2990,N_3368);
or U4980 (N_4980,N_2581,N_3508);
nand U4981 (N_4981,N_3411,N_2562);
nor U4982 (N_4982,N_2746,N_2429);
and U4983 (N_4983,N_3043,N_3795);
nand U4984 (N_4984,N_2422,N_3618);
nand U4985 (N_4985,N_3996,N_2924);
and U4986 (N_4986,N_2530,N_2893);
and U4987 (N_4987,N_2925,N_3785);
and U4988 (N_4988,N_2139,N_2851);
and U4989 (N_4989,N_2922,N_3925);
nor U4990 (N_4990,N_2067,N_3428);
nand U4991 (N_4991,N_2831,N_2330);
and U4992 (N_4992,N_2585,N_2065);
nor U4993 (N_4993,N_2281,N_2270);
and U4994 (N_4994,N_3169,N_3131);
or U4995 (N_4995,N_3818,N_2497);
or U4996 (N_4996,N_2130,N_3026);
or U4997 (N_4997,N_3471,N_2528);
nand U4998 (N_4998,N_3071,N_3027);
nor U4999 (N_4999,N_2896,N_2762);
and U5000 (N_5000,N_2856,N_2960);
or U5001 (N_5001,N_3792,N_3619);
or U5002 (N_5002,N_3551,N_2348);
nand U5003 (N_5003,N_3277,N_3927);
and U5004 (N_5004,N_2237,N_3846);
nor U5005 (N_5005,N_2775,N_3748);
nand U5006 (N_5006,N_2029,N_3147);
or U5007 (N_5007,N_2801,N_2648);
nor U5008 (N_5008,N_2404,N_3112);
or U5009 (N_5009,N_3489,N_3203);
and U5010 (N_5010,N_2616,N_2484);
or U5011 (N_5011,N_2443,N_2100);
nor U5012 (N_5012,N_2680,N_3313);
and U5013 (N_5013,N_2113,N_3163);
nor U5014 (N_5014,N_3468,N_2952);
or U5015 (N_5015,N_3240,N_2115);
or U5016 (N_5016,N_2257,N_2376);
and U5017 (N_5017,N_3368,N_3109);
and U5018 (N_5018,N_3816,N_3254);
or U5019 (N_5019,N_3942,N_2980);
or U5020 (N_5020,N_2600,N_3309);
nand U5021 (N_5021,N_2841,N_2532);
and U5022 (N_5022,N_3274,N_2452);
nand U5023 (N_5023,N_3172,N_3281);
nor U5024 (N_5024,N_3447,N_2084);
nand U5025 (N_5025,N_3660,N_3003);
or U5026 (N_5026,N_2299,N_3268);
nor U5027 (N_5027,N_3405,N_3496);
nor U5028 (N_5028,N_3766,N_2120);
or U5029 (N_5029,N_3926,N_2946);
and U5030 (N_5030,N_3538,N_2366);
nand U5031 (N_5031,N_2139,N_3902);
nand U5032 (N_5032,N_3553,N_2385);
nand U5033 (N_5033,N_2734,N_2954);
nor U5034 (N_5034,N_2250,N_2201);
nand U5035 (N_5035,N_2802,N_3001);
or U5036 (N_5036,N_2984,N_3231);
nor U5037 (N_5037,N_2480,N_2706);
or U5038 (N_5038,N_3407,N_2447);
nor U5039 (N_5039,N_3602,N_3868);
and U5040 (N_5040,N_2886,N_3193);
or U5041 (N_5041,N_3061,N_3676);
or U5042 (N_5042,N_2397,N_3684);
and U5043 (N_5043,N_2042,N_2996);
xnor U5044 (N_5044,N_3018,N_2445);
nor U5045 (N_5045,N_3425,N_2708);
xnor U5046 (N_5046,N_2239,N_3728);
and U5047 (N_5047,N_3214,N_3657);
nor U5048 (N_5048,N_2665,N_3815);
and U5049 (N_5049,N_2553,N_2022);
nand U5050 (N_5050,N_2956,N_2407);
and U5051 (N_5051,N_3625,N_2131);
nand U5052 (N_5052,N_3971,N_3765);
and U5053 (N_5053,N_3635,N_2448);
nor U5054 (N_5054,N_3749,N_2759);
or U5055 (N_5055,N_2464,N_2293);
and U5056 (N_5056,N_3803,N_3823);
and U5057 (N_5057,N_3385,N_2103);
nor U5058 (N_5058,N_2246,N_2320);
nand U5059 (N_5059,N_3432,N_2633);
and U5060 (N_5060,N_3255,N_2024);
nor U5061 (N_5061,N_2272,N_2660);
nor U5062 (N_5062,N_3613,N_3658);
xnor U5063 (N_5063,N_3386,N_2498);
nand U5064 (N_5064,N_2137,N_3797);
or U5065 (N_5065,N_3181,N_2089);
nand U5066 (N_5066,N_2803,N_3517);
and U5067 (N_5067,N_2197,N_3357);
nand U5068 (N_5068,N_3703,N_2857);
or U5069 (N_5069,N_2335,N_2668);
or U5070 (N_5070,N_2757,N_2758);
nand U5071 (N_5071,N_2993,N_2937);
or U5072 (N_5072,N_3290,N_2916);
and U5073 (N_5073,N_2934,N_3495);
nor U5074 (N_5074,N_3804,N_3604);
or U5075 (N_5075,N_2025,N_3670);
or U5076 (N_5076,N_3198,N_3549);
nand U5077 (N_5077,N_2151,N_3768);
nor U5078 (N_5078,N_2740,N_2146);
nand U5079 (N_5079,N_2573,N_2862);
xor U5080 (N_5080,N_2808,N_2989);
nand U5081 (N_5081,N_2195,N_3315);
nand U5082 (N_5082,N_3967,N_2186);
or U5083 (N_5083,N_2696,N_3615);
or U5084 (N_5084,N_2117,N_2876);
nor U5085 (N_5085,N_3864,N_2324);
nor U5086 (N_5086,N_2451,N_2644);
nor U5087 (N_5087,N_3875,N_2037);
nand U5088 (N_5088,N_3140,N_2570);
and U5089 (N_5089,N_2087,N_2019);
nor U5090 (N_5090,N_2770,N_2082);
xor U5091 (N_5091,N_3518,N_3695);
nor U5092 (N_5092,N_3051,N_2004);
nand U5093 (N_5093,N_3784,N_2776);
nand U5094 (N_5094,N_2152,N_2084);
or U5095 (N_5095,N_3292,N_2073);
and U5096 (N_5096,N_3678,N_2757);
nor U5097 (N_5097,N_2723,N_2854);
nand U5098 (N_5098,N_3739,N_2210);
nor U5099 (N_5099,N_3090,N_2302);
and U5100 (N_5100,N_3144,N_2409);
or U5101 (N_5101,N_2131,N_3550);
and U5102 (N_5102,N_2691,N_3989);
or U5103 (N_5103,N_2728,N_2898);
nand U5104 (N_5104,N_3795,N_3418);
nand U5105 (N_5105,N_3191,N_2964);
nand U5106 (N_5106,N_2136,N_3434);
xnor U5107 (N_5107,N_2299,N_3805);
and U5108 (N_5108,N_2630,N_2700);
or U5109 (N_5109,N_2832,N_2586);
or U5110 (N_5110,N_3649,N_3352);
nand U5111 (N_5111,N_3541,N_2034);
nor U5112 (N_5112,N_2009,N_2561);
or U5113 (N_5113,N_2342,N_2248);
or U5114 (N_5114,N_2341,N_3974);
nor U5115 (N_5115,N_2162,N_2206);
and U5116 (N_5116,N_3762,N_3269);
nor U5117 (N_5117,N_2136,N_2350);
or U5118 (N_5118,N_2349,N_3301);
or U5119 (N_5119,N_3341,N_2682);
nand U5120 (N_5120,N_2315,N_2702);
or U5121 (N_5121,N_3829,N_2399);
nand U5122 (N_5122,N_2915,N_2982);
nor U5123 (N_5123,N_2703,N_3778);
and U5124 (N_5124,N_3803,N_3793);
or U5125 (N_5125,N_3104,N_2442);
or U5126 (N_5126,N_2220,N_2470);
and U5127 (N_5127,N_3758,N_2151);
nor U5128 (N_5128,N_3951,N_2251);
nor U5129 (N_5129,N_3690,N_3904);
nor U5130 (N_5130,N_2955,N_3922);
nand U5131 (N_5131,N_3746,N_3969);
and U5132 (N_5132,N_3836,N_3185);
nand U5133 (N_5133,N_2356,N_3749);
nor U5134 (N_5134,N_3606,N_3754);
or U5135 (N_5135,N_2640,N_3485);
nor U5136 (N_5136,N_3394,N_2830);
or U5137 (N_5137,N_3277,N_2198);
nand U5138 (N_5138,N_3278,N_3829);
and U5139 (N_5139,N_3828,N_3890);
nor U5140 (N_5140,N_2454,N_3072);
or U5141 (N_5141,N_2188,N_2089);
or U5142 (N_5142,N_2554,N_2999);
and U5143 (N_5143,N_3774,N_3796);
and U5144 (N_5144,N_3718,N_2373);
or U5145 (N_5145,N_3540,N_3006);
xnor U5146 (N_5146,N_3298,N_3499);
xnor U5147 (N_5147,N_3535,N_2920);
nor U5148 (N_5148,N_3192,N_2687);
or U5149 (N_5149,N_2675,N_3046);
nor U5150 (N_5150,N_2204,N_2438);
or U5151 (N_5151,N_2240,N_3646);
and U5152 (N_5152,N_2322,N_2856);
nand U5153 (N_5153,N_3398,N_2123);
nand U5154 (N_5154,N_3533,N_3541);
nand U5155 (N_5155,N_2893,N_2896);
and U5156 (N_5156,N_3959,N_3713);
nor U5157 (N_5157,N_3303,N_3395);
nand U5158 (N_5158,N_3263,N_2764);
or U5159 (N_5159,N_3024,N_2920);
and U5160 (N_5160,N_2764,N_2278);
nor U5161 (N_5161,N_2956,N_3754);
nor U5162 (N_5162,N_3915,N_3230);
nand U5163 (N_5163,N_2553,N_3700);
and U5164 (N_5164,N_2003,N_2080);
and U5165 (N_5165,N_3059,N_2192);
and U5166 (N_5166,N_2147,N_3039);
nor U5167 (N_5167,N_3112,N_2381);
nor U5168 (N_5168,N_2666,N_3552);
or U5169 (N_5169,N_3098,N_2535);
and U5170 (N_5170,N_2307,N_3721);
nor U5171 (N_5171,N_2979,N_3455);
nor U5172 (N_5172,N_3347,N_3462);
and U5173 (N_5173,N_3318,N_3389);
or U5174 (N_5174,N_2007,N_2723);
or U5175 (N_5175,N_2485,N_3319);
nor U5176 (N_5176,N_3141,N_2322);
or U5177 (N_5177,N_3896,N_3926);
and U5178 (N_5178,N_2517,N_2087);
nor U5179 (N_5179,N_2744,N_2910);
nand U5180 (N_5180,N_2485,N_3169);
nor U5181 (N_5181,N_3433,N_2873);
and U5182 (N_5182,N_3722,N_3924);
and U5183 (N_5183,N_3838,N_2111);
nand U5184 (N_5184,N_3848,N_3368);
nand U5185 (N_5185,N_3341,N_2892);
nor U5186 (N_5186,N_3815,N_3409);
or U5187 (N_5187,N_3247,N_2267);
nor U5188 (N_5188,N_3608,N_2588);
nand U5189 (N_5189,N_3415,N_3011);
nor U5190 (N_5190,N_3082,N_3201);
nand U5191 (N_5191,N_2030,N_3869);
or U5192 (N_5192,N_2161,N_2188);
nor U5193 (N_5193,N_2759,N_3889);
or U5194 (N_5194,N_3806,N_3583);
nor U5195 (N_5195,N_2275,N_2747);
nor U5196 (N_5196,N_3571,N_2051);
or U5197 (N_5197,N_2265,N_2377);
nand U5198 (N_5198,N_3338,N_2016);
or U5199 (N_5199,N_3816,N_2503);
nand U5200 (N_5200,N_2053,N_3116);
and U5201 (N_5201,N_3624,N_3137);
and U5202 (N_5202,N_3690,N_2668);
or U5203 (N_5203,N_3552,N_3078);
nand U5204 (N_5204,N_3996,N_2370);
nor U5205 (N_5205,N_2464,N_2343);
and U5206 (N_5206,N_3144,N_2482);
nand U5207 (N_5207,N_3793,N_3514);
and U5208 (N_5208,N_3680,N_3113);
or U5209 (N_5209,N_3243,N_3629);
nand U5210 (N_5210,N_2624,N_2312);
nor U5211 (N_5211,N_2411,N_2615);
nand U5212 (N_5212,N_2379,N_2642);
or U5213 (N_5213,N_2534,N_3397);
or U5214 (N_5214,N_3920,N_3648);
nor U5215 (N_5215,N_2484,N_3300);
nor U5216 (N_5216,N_2844,N_2494);
nor U5217 (N_5217,N_2967,N_3070);
nor U5218 (N_5218,N_2942,N_2060);
or U5219 (N_5219,N_3177,N_3194);
nand U5220 (N_5220,N_3192,N_3002);
nand U5221 (N_5221,N_2518,N_3344);
or U5222 (N_5222,N_3692,N_2615);
nand U5223 (N_5223,N_2659,N_3937);
nor U5224 (N_5224,N_2942,N_2632);
and U5225 (N_5225,N_3079,N_3334);
nor U5226 (N_5226,N_2948,N_3439);
nor U5227 (N_5227,N_3234,N_3541);
or U5228 (N_5228,N_3651,N_3656);
and U5229 (N_5229,N_3842,N_3086);
nor U5230 (N_5230,N_3103,N_2709);
nand U5231 (N_5231,N_2515,N_3962);
and U5232 (N_5232,N_2116,N_2542);
nand U5233 (N_5233,N_2784,N_3568);
nor U5234 (N_5234,N_3718,N_3976);
xor U5235 (N_5235,N_2721,N_3700);
and U5236 (N_5236,N_2698,N_3151);
and U5237 (N_5237,N_3625,N_3317);
nand U5238 (N_5238,N_2297,N_3603);
or U5239 (N_5239,N_3561,N_2817);
nand U5240 (N_5240,N_3366,N_2621);
or U5241 (N_5241,N_3333,N_2131);
or U5242 (N_5242,N_2099,N_2802);
nor U5243 (N_5243,N_3778,N_3644);
and U5244 (N_5244,N_2622,N_3109);
and U5245 (N_5245,N_2889,N_3946);
nand U5246 (N_5246,N_3088,N_3444);
and U5247 (N_5247,N_2779,N_2609);
nand U5248 (N_5248,N_3609,N_3458);
or U5249 (N_5249,N_3150,N_2792);
nand U5250 (N_5250,N_2781,N_2832);
nor U5251 (N_5251,N_2571,N_2435);
xor U5252 (N_5252,N_3258,N_2456);
or U5253 (N_5253,N_3382,N_2637);
and U5254 (N_5254,N_2083,N_2039);
or U5255 (N_5255,N_2253,N_2387);
or U5256 (N_5256,N_2794,N_3105);
and U5257 (N_5257,N_3342,N_2701);
or U5258 (N_5258,N_2300,N_2330);
nand U5259 (N_5259,N_2277,N_2525);
or U5260 (N_5260,N_3545,N_2360);
nand U5261 (N_5261,N_2644,N_2231);
nor U5262 (N_5262,N_3718,N_3057);
nor U5263 (N_5263,N_2752,N_2203);
and U5264 (N_5264,N_2753,N_2463);
nor U5265 (N_5265,N_3002,N_3136);
or U5266 (N_5266,N_3683,N_3514);
and U5267 (N_5267,N_2077,N_2971);
nand U5268 (N_5268,N_2089,N_3020);
and U5269 (N_5269,N_3710,N_3326);
nor U5270 (N_5270,N_2646,N_3980);
or U5271 (N_5271,N_3282,N_2123);
and U5272 (N_5272,N_2378,N_2319);
nor U5273 (N_5273,N_2173,N_3918);
nand U5274 (N_5274,N_2364,N_2365);
and U5275 (N_5275,N_3036,N_2549);
nor U5276 (N_5276,N_3297,N_2979);
or U5277 (N_5277,N_2820,N_2766);
and U5278 (N_5278,N_3963,N_3385);
and U5279 (N_5279,N_2181,N_2652);
or U5280 (N_5280,N_2714,N_3503);
nor U5281 (N_5281,N_2562,N_2811);
or U5282 (N_5282,N_3771,N_3904);
and U5283 (N_5283,N_2741,N_2129);
or U5284 (N_5284,N_3861,N_3078);
and U5285 (N_5285,N_3847,N_3796);
nor U5286 (N_5286,N_3208,N_3903);
and U5287 (N_5287,N_2401,N_2046);
nand U5288 (N_5288,N_2954,N_3723);
xor U5289 (N_5289,N_2976,N_3928);
or U5290 (N_5290,N_2747,N_2785);
and U5291 (N_5291,N_2226,N_3999);
nor U5292 (N_5292,N_3404,N_3308);
xnor U5293 (N_5293,N_3021,N_3737);
and U5294 (N_5294,N_3335,N_2631);
and U5295 (N_5295,N_3817,N_2188);
nor U5296 (N_5296,N_2569,N_2276);
or U5297 (N_5297,N_2197,N_2652);
nor U5298 (N_5298,N_2626,N_3832);
or U5299 (N_5299,N_2733,N_3961);
nand U5300 (N_5300,N_2956,N_3341);
or U5301 (N_5301,N_3218,N_3797);
nor U5302 (N_5302,N_3449,N_2037);
nand U5303 (N_5303,N_3092,N_2036);
or U5304 (N_5304,N_2956,N_2583);
and U5305 (N_5305,N_3895,N_2663);
and U5306 (N_5306,N_3409,N_3744);
nand U5307 (N_5307,N_2024,N_3404);
or U5308 (N_5308,N_3949,N_2639);
nor U5309 (N_5309,N_2723,N_3032);
nand U5310 (N_5310,N_2705,N_3645);
or U5311 (N_5311,N_2419,N_2780);
nor U5312 (N_5312,N_2618,N_3286);
nor U5313 (N_5313,N_2972,N_3061);
nand U5314 (N_5314,N_2924,N_3886);
nand U5315 (N_5315,N_2126,N_2836);
or U5316 (N_5316,N_2071,N_3341);
and U5317 (N_5317,N_2320,N_2465);
or U5318 (N_5318,N_2967,N_2959);
and U5319 (N_5319,N_2581,N_3644);
and U5320 (N_5320,N_3808,N_2268);
nor U5321 (N_5321,N_3600,N_3330);
nand U5322 (N_5322,N_2194,N_2667);
nand U5323 (N_5323,N_3233,N_3863);
nor U5324 (N_5324,N_3559,N_2613);
or U5325 (N_5325,N_3968,N_2594);
nand U5326 (N_5326,N_3662,N_3338);
or U5327 (N_5327,N_2702,N_2314);
or U5328 (N_5328,N_3042,N_3633);
nand U5329 (N_5329,N_3755,N_3659);
nor U5330 (N_5330,N_2292,N_2393);
nand U5331 (N_5331,N_3142,N_3445);
nand U5332 (N_5332,N_2320,N_3149);
or U5333 (N_5333,N_2474,N_3170);
or U5334 (N_5334,N_3230,N_3222);
or U5335 (N_5335,N_3510,N_2636);
nor U5336 (N_5336,N_2743,N_3881);
nor U5337 (N_5337,N_3366,N_3390);
and U5338 (N_5338,N_2028,N_2843);
or U5339 (N_5339,N_3737,N_2279);
nor U5340 (N_5340,N_3049,N_3778);
nand U5341 (N_5341,N_3311,N_3539);
nand U5342 (N_5342,N_3894,N_3557);
nand U5343 (N_5343,N_3129,N_2942);
or U5344 (N_5344,N_3173,N_2366);
nor U5345 (N_5345,N_3012,N_3565);
or U5346 (N_5346,N_3698,N_2415);
and U5347 (N_5347,N_2038,N_2428);
nand U5348 (N_5348,N_3638,N_2828);
nor U5349 (N_5349,N_3302,N_3971);
nor U5350 (N_5350,N_2630,N_3243);
or U5351 (N_5351,N_2972,N_3894);
and U5352 (N_5352,N_2293,N_3020);
and U5353 (N_5353,N_2600,N_2651);
nand U5354 (N_5354,N_3157,N_2530);
and U5355 (N_5355,N_2103,N_2552);
nor U5356 (N_5356,N_3379,N_3202);
nand U5357 (N_5357,N_2830,N_3163);
nand U5358 (N_5358,N_3822,N_2595);
or U5359 (N_5359,N_3046,N_3826);
nor U5360 (N_5360,N_2196,N_3359);
nor U5361 (N_5361,N_2472,N_2300);
nand U5362 (N_5362,N_2718,N_3462);
and U5363 (N_5363,N_3763,N_3992);
or U5364 (N_5364,N_3868,N_3874);
and U5365 (N_5365,N_2182,N_2811);
and U5366 (N_5366,N_2859,N_3488);
or U5367 (N_5367,N_2809,N_2835);
nor U5368 (N_5368,N_2764,N_3765);
or U5369 (N_5369,N_2706,N_2324);
nor U5370 (N_5370,N_3300,N_2670);
and U5371 (N_5371,N_3593,N_2043);
and U5372 (N_5372,N_3414,N_2343);
nor U5373 (N_5373,N_2375,N_3638);
nor U5374 (N_5374,N_2742,N_2074);
nand U5375 (N_5375,N_3290,N_2660);
nor U5376 (N_5376,N_3180,N_2127);
nand U5377 (N_5377,N_3795,N_3133);
nand U5378 (N_5378,N_3441,N_2998);
nand U5379 (N_5379,N_3264,N_2495);
or U5380 (N_5380,N_2473,N_2071);
nor U5381 (N_5381,N_2137,N_2509);
or U5382 (N_5382,N_3510,N_3579);
or U5383 (N_5383,N_3204,N_3219);
and U5384 (N_5384,N_2743,N_3491);
and U5385 (N_5385,N_3782,N_2322);
nand U5386 (N_5386,N_2058,N_2885);
or U5387 (N_5387,N_2862,N_2641);
and U5388 (N_5388,N_3493,N_2563);
nor U5389 (N_5389,N_3885,N_2251);
nor U5390 (N_5390,N_3384,N_3619);
nand U5391 (N_5391,N_3937,N_3375);
or U5392 (N_5392,N_2059,N_3644);
or U5393 (N_5393,N_2176,N_3160);
nor U5394 (N_5394,N_3694,N_3331);
and U5395 (N_5395,N_2266,N_3812);
nor U5396 (N_5396,N_2572,N_2768);
nor U5397 (N_5397,N_2449,N_2637);
nand U5398 (N_5398,N_2256,N_2396);
and U5399 (N_5399,N_2269,N_2144);
or U5400 (N_5400,N_3691,N_2881);
nand U5401 (N_5401,N_2298,N_3199);
or U5402 (N_5402,N_3249,N_3346);
or U5403 (N_5403,N_2656,N_3710);
and U5404 (N_5404,N_2350,N_2231);
nor U5405 (N_5405,N_2513,N_2966);
nand U5406 (N_5406,N_2203,N_3256);
nand U5407 (N_5407,N_3725,N_3786);
or U5408 (N_5408,N_2520,N_3733);
or U5409 (N_5409,N_2568,N_2340);
xor U5410 (N_5410,N_2948,N_3706);
or U5411 (N_5411,N_2971,N_2133);
and U5412 (N_5412,N_2424,N_3782);
nand U5413 (N_5413,N_3140,N_2778);
or U5414 (N_5414,N_3783,N_3565);
nor U5415 (N_5415,N_3526,N_2101);
and U5416 (N_5416,N_3076,N_2462);
or U5417 (N_5417,N_2275,N_3207);
or U5418 (N_5418,N_2282,N_3592);
or U5419 (N_5419,N_3132,N_2967);
nand U5420 (N_5420,N_3432,N_3129);
nand U5421 (N_5421,N_2372,N_3024);
or U5422 (N_5422,N_2624,N_2339);
or U5423 (N_5423,N_2159,N_3920);
nor U5424 (N_5424,N_2299,N_3520);
nor U5425 (N_5425,N_2422,N_2715);
and U5426 (N_5426,N_3762,N_3248);
and U5427 (N_5427,N_2837,N_3541);
nor U5428 (N_5428,N_2893,N_2810);
or U5429 (N_5429,N_3293,N_2955);
nor U5430 (N_5430,N_2792,N_2338);
nor U5431 (N_5431,N_2423,N_2903);
and U5432 (N_5432,N_3444,N_3071);
nand U5433 (N_5433,N_3706,N_3033);
nand U5434 (N_5434,N_2690,N_3413);
nand U5435 (N_5435,N_3595,N_2754);
nor U5436 (N_5436,N_3022,N_3589);
and U5437 (N_5437,N_3661,N_2077);
nand U5438 (N_5438,N_2105,N_3332);
and U5439 (N_5439,N_3082,N_3387);
nor U5440 (N_5440,N_2496,N_3167);
or U5441 (N_5441,N_3006,N_3806);
and U5442 (N_5442,N_2935,N_2284);
nand U5443 (N_5443,N_2398,N_2512);
nand U5444 (N_5444,N_3834,N_3524);
nand U5445 (N_5445,N_3295,N_2547);
nand U5446 (N_5446,N_3171,N_3387);
nand U5447 (N_5447,N_3423,N_2844);
nand U5448 (N_5448,N_3137,N_2066);
nor U5449 (N_5449,N_3191,N_2447);
or U5450 (N_5450,N_3995,N_2458);
nand U5451 (N_5451,N_3373,N_3151);
nand U5452 (N_5452,N_2311,N_3019);
and U5453 (N_5453,N_3013,N_3204);
nor U5454 (N_5454,N_3833,N_2744);
nor U5455 (N_5455,N_2779,N_2241);
nor U5456 (N_5456,N_3604,N_3386);
nor U5457 (N_5457,N_3363,N_2799);
or U5458 (N_5458,N_2031,N_3985);
nand U5459 (N_5459,N_2024,N_3198);
or U5460 (N_5460,N_2334,N_2997);
nand U5461 (N_5461,N_2550,N_3291);
or U5462 (N_5462,N_2256,N_2514);
and U5463 (N_5463,N_3335,N_3744);
nor U5464 (N_5464,N_3759,N_3840);
and U5465 (N_5465,N_2369,N_2792);
nand U5466 (N_5466,N_2731,N_2502);
nor U5467 (N_5467,N_3822,N_3135);
nor U5468 (N_5468,N_2538,N_3690);
and U5469 (N_5469,N_3191,N_3871);
and U5470 (N_5470,N_3588,N_2953);
and U5471 (N_5471,N_3709,N_2459);
xor U5472 (N_5472,N_2017,N_2699);
nand U5473 (N_5473,N_2389,N_2411);
nand U5474 (N_5474,N_2525,N_2491);
nor U5475 (N_5475,N_2944,N_3415);
nand U5476 (N_5476,N_2344,N_2219);
and U5477 (N_5477,N_2089,N_3313);
nor U5478 (N_5478,N_2475,N_3879);
nand U5479 (N_5479,N_2122,N_3187);
nand U5480 (N_5480,N_2839,N_3908);
nand U5481 (N_5481,N_2155,N_2566);
or U5482 (N_5482,N_3205,N_2822);
and U5483 (N_5483,N_3557,N_2619);
nor U5484 (N_5484,N_2525,N_3542);
nand U5485 (N_5485,N_2125,N_3907);
or U5486 (N_5486,N_3720,N_2166);
nand U5487 (N_5487,N_3404,N_2782);
or U5488 (N_5488,N_2583,N_2589);
nor U5489 (N_5489,N_3776,N_3296);
nor U5490 (N_5490,N_3858,N_2233);
nand U5491 (N_5491,N_2377,N_2170);
and U5492 (N_5492,N_2054,N_2201);
and U5493 (N_5493,N_3965,N_3386);
nor U5494 (N_5494,N_3823,N_3801);
xor U5495 (N_5495,N_3902,N_3452);
or U5496 (N_5496,N_3944,N_2731);
nand U5497 (N_5497,N_3637,N_2113);
nand U5498 (N_5498,N_3842,N_2942);
nand U5499 (N_5499,N_2541,N_2496);
and U5500 (N_5500,N_3258,N_3864);
nor U5501 (N_5501,N_3875,N_3325);
or U5502 (N_5502,N_3533,N_2113);
or U5503 (N_5503,N_2014,N_3470);
or U5504 (N_5504,N_2893,N_2547);
nor U5505 (N_5505,N_3205,N_3083);
nor U5506 (N_5506,N_3129,N_2876);
and U5507 (N_5507,N_3056,N_2616);
nor U5508 (N_5508,N_2692,N_3934);
nand U5509 (N_5509,N_3297,N_3840);
nand U5510 (N_5510,N_2662,N_3206);
nand U5511 (N_5511,N_3959,N_2391);
and U5512 (N_5512,N_2323,N_2683);
or U5513 (N_5513,N_2418,N_3172);
and U5514 (N_5514,N_2968,N_2216);
or U5515 (N_5515,N_2451,N_3604);
or U5516 (N_5516,N_3405,N_2042);
xor U5517 (N_5517,N_2172,N_3038);
and U5518 (N_5518,N_2970,N_2309);
and U5519 (N_5519,N_2566,N_2380);
nand U5520 (N_5520,N_3688,N_3541);
or U5521 (N_5521,N_2014,N_3998);
nor U5522 (N_5522,N_2097,N_2658);
nor U5523 (N_5523,N_2060,N_3185);
nor U5524 (N_5524,N_3289,N_3192);
and U5525 (N_5525,N_3950,N_3476);
or U5526 (N_5526,N_2238,N_2113);
nand U5527 (N_5527,N_3784,N_3160);
and U5528 (N_5528,N_3385,N_2740);
and U5529 (N_5529,N_3480,N_3515);
or U5530 (N_5530,N_3668,N_3068);
or U5531 (N_5531,N_3686,N_2845);
and U5532 (N_5532,N_2407,N_2275);
and U5533 (N_5533,N_3042,N_3123);
and U5534 (N_5534,N_3018,N_3345);
nor U5535 (N_5535,N_3510,N_2453);
nor U5536 (N_5536,N_2998,N_2445);
nand U5537 (N_5537,N_3662,N_3589);
nand U5538 (N_5538,N_2481,N_2691);
or U5539 (N_5539,N_2389,N_3227);
and U5540 (N_5540,N_2252,N_2854);
or U5541 (N_5541,N_3242,N_3149);
nand U5542 (N_5542,N_2930,N_3067);
and U5543 (N_5543,N_2631,N_3735);
and U5544 (N_5544,N_2559,N_3042);
nand U5545 (N_5545,N_3449,N_2127);
and U5546 (N_5546,N_3870,N_3146);
nand U5547 (N_5547,N_3889,N_2110);
and U5548 (N_5548,N_2106,N_2629);
nand U5549 (N_5549,N_2170,N_3648);
or U5550 (N_5550,N_2967,N_2423);
or U5551 (N_5551,N_3277,N_3499);
nor U5552 (N_5552,N_3021,N_2329);
nor U5553 (N_5553,N_3005,N_2824);
and U5554 (N_5554,N_3660,N_2401);
or U5555 (N_5555,N_2061,N_2400);
or U5556 (N_5556,N_2627,N_2153);
or U5557 (N_5557,N_2053,N_2898);
nand U5558 (N_5558,N_2268,N_3533);
or U5559 (N_5559,N_3749,N_2525);
or U5560 (N_5560,N_2470,N_2802);
xor U5561 (N_5561,N_2546,N_3820);
nor U5562 (N_5562,N_3901,N_2332);
nor U5563 (N_5563,N_3019,N_3838);
and U5564 (N_5564,N_2172,N_2342);
or U5565 (N_5565,N_2222,N_2050);
nor U5566 (N_5566,N_3053,N_3494);
or U5567 (N_5567,N_2149,N_3941);
nor U5568 (N_5568,N_2966,N_2951);
or U5569 (N_5569,N_2857,N_3264);
nor U5570 (N_5570,N_2126,N_2521);
or U5571 (N_5571,N_3527,N_2925);
nand U5572 (N_5572,N_3917,N_3424);
nand U5573 (N_5573,N_2562,N_2160);
nand U5574 (N_5574,N_2682,N_2083);
or U5575 (N_5575,N_2979,N_3326);
xnor U5576 (N_5576,N_2708,N_2625);
or U5577 (N_5577,N_3555,N_2501);
nand U5578 (N_5578,N_3193,N_2016);
xor U5579 (N_5579,N_2409,N_3715);
and U5580 (N_5580,N_3691,N_3037);
or U5581 (N_5581,N_2046,N_3426);
nor U5582 (N_5582,N_3614,N_2614);
nor U5583 (N_5583,N_2335,N_3278);
nand U5584 (N_5584,N_3244,N_2052);
or U5585 (N_5585,N_2509,N_2204);
nand U5586 (N_5586,N_2658,N_2151);
or U5587 (N_5587,N_2284,N_3363);
nor U5588 (N_5588,N_2238,N_2834);
or U5589 (N_5589,N_3888,N_2250);
and U5590 (N_5590,N_3954,N_2178);
nand U5591 (N_5591,N_3127,N_3555);
nand U5592 (N_5592,N_3464,N_3792);
and U5593 (N_5593,N_3472,N_2280);
nand U5594 (N_5594,N_3453,N_3538);
nand U5595 (N_5595,N_3449,N_3659);
and U5596 (N_5596,N_3382,N_3154);
nand U5597 (N_5597,N_2277,N_2390);
or U5598 (N_5598,N_3546,N_3686);
or U5599 (N_5599,N_3105,N_3874);
nor U5600 (N_5600,N_3548,N_2191);
and U5601 (N_5601,N_2012,N_3958);
nand U5602 (N_5602,N_2885,N_2939);
and U5603 (N_5603,N_3648,N_3781);
or U5604 (N_5604,N_3937,N_2285);
and U5605 (N_5605,N_2821,N_2527);
nand U5606 (N_5606,N_2089,N_3451);
or U5607 (N_5607,N_2660,N_3857);
nor U5608 (N_5608,N_3759,N_2866);
nor U5609 (N_5609,N_2644,N_3197);
nand U5610 (N_5610,N_2530,N_2485);
or U5611 (N_5611,N_2013,N_3380);
and U5612 (N_5612,N_3268,N_2679);
and U5613 (N_5613,N_2916,N_3008);
and U5614 (N_5614,N_3872,N_3566);
nand U5615 (N_5615,N_2232,N_3410);
and U5616 (N_5616,N_2620,N_2268);
nand U5617 (N_5617,N_2435,N_3010);
nand U5618 (N_5618,N_3696,N_2472);
or U5619 (N_5619,N_3844,N_2629);
and U5620 (N_5620,N_3566,N_3449);
nand U5621 (N_5621,N_2632,N_3909);
nand U5622 (N_5622,N_2344,N_3773);
nor U5623 (N_5623,N_2878,N_2167);
or U5624 (N_5624,N_3105,N_2461);
nor U5625 (N_5625,N_3210,N_3821);
nor U5626 (N_5626,N_3604,N_2286);
and U5627 (N_5627,N_3612,N_2888);
nor U5628 (N_5628,N_3000,N_2327);
nand U5629 (N_5629,N_2402,N_3703);
nand U5630 (N_5630,N_2307,N_2785);
or U5631 (N_5631,N_3070,N_3523);
nor U5632 (N_5632,N_2986,N_2050);
nor U5633 (N_5633,N_3619,N_3827);
nor U5634 (N_5634,N_3944,N_3955);
nor U5635 (N_5635,N_2288,N_2685);
and U5636 (N_5636,N_3749,N_3516);
nand U5637 (N_5637,N_3366,N_3024);
nor U5638 (N_5638,N_3558,N_2691);
nor U5639 (N_5639,N_3108,N_2753);
and U5640 (N_5640,N_3439,N_3525);
xor U5641 (N_5641,N_2645,N_2880);
and U5642 (N_5642,N_3764,N_2739);
or U5643 (N_5643,N_2740,N_2840);
or U5644 (N_5644,N_2858,N_3219);
nand U5645 (N_5645,N_3667,N_3448);
and U5646 (N_5646,N_2717,N_2946);
nor U5647 (N_5647,N_2133,N_3692);
or U5648 (N_5648,N_3054,N_3423);
nand U5649 (N_5649,N_2423,N_3186);
nand U5650 (N_5650,N_2445,N_2443);
nor U5651 (N_5651,N_3216,N_2123);
nand U5652 (N_5652,N_3301,N_3661);
or U5653 (N_5653,N_2842,N_2496);
and U5654 (N_5654,N_2847,N_2705);
and U5655 (N_5655,N_2509,N_3722);
nand U5656 (N_5656,N_2552,N_3739);
nor U5657 (N_5657,N_3263,N_2991);
nor U5658 (N_5658,N_3828,N_2396);
and U5659 (N_5659,N_2313,N_3998);
nand U5660 (N_5660,N_2118,N_2536);
nor U5661 (N_5661,N_3206,N_2385);
xor U5662 (N_5662,N_2800,N_3513);
and U5663 (N_5663,N_2507,N_3415);
and U5664 (N_5664,N_3306,N_3190);
nand U5665 (N_5665,N_2825,N_2555);
nor U5666 (N_5666,N_3512,N_2239);
and U5667 (N_5667,N_3197,N_2146);
and U5668 (N_5668,N_2908,N_2969);
or U5669 (N_5669,N_3819,N_2782);
xnor U5670 (N_5670,N_2719,N_2479);
nand U5671 (N_5671,N_3072,N_3955);
or U5672 (N_5672,N_3681,N_3193);
or U5673 (N_5673,N_2434,N_2208);
nand U5674 (N_5674,N_2459,N_2989);
and U5675 (N_5675,N_2808,N_2302);
nor U5676 (N_5676,N_3620,N_2400);
and U5677 (N_5677,N_3163,N_3090);
or U5678 (N_5678,N_2098,N_3496);
nor U5679 (N_5679,N_2880,N_2672);
and U5680 (N_5680,N_3802,N_2599);
xnor U5681 (N_5681,N_3466,N_2305);
or U5682 (N_5682,N_3396,N_2536);
and U5683 (N_5683,N_2533,N_3294);
and U5684 (N_5684,N_2546,N_2469);
nand U5685 (N_5685,N_2521,N_2620);
nand U5686 (N_5686,N_3969,N_3819);
nor U5687 (N_5687,N_3734,N_2492);
nand U5688 (N_5688,N_3402,N_3329);
nor U5689 (N_5689,N_2502,N_3888);
or U5690 (N_5690,N_3436,N_2875);
or U5691 (N_5691,N_3043,N_2401);
and U5692 (N_5692,N_3819,N_3242);
or U5693 (N_5693,N_3252,N_3646);
and U5694 (N_5694,N_2553,N_3064);
nor U5695 (N_5695,N_3480,N_2258);
nor U5696 (N_5696,N_3164,N_2076);
nor U5697 (N_5697,N_3247,N_3372);
nand U5698 (N_5698,N_3003,N_3898);
nor U5699 (N_5699,N_3645,N_2754);
and U5700 (N_5700,N_3254,N_2840);
or U5701 (N_5701,N_2014,N_2943);
or U5702 (N_5702,N_2779,N_3298);
nand U5703 (N_5703,N_2493,N_2337);
or U5704 (N_5704,N_2128,N_3909);
nand U5705 (N_5705,N_2430,N_3750);
nand U5706 (N_5706,N_2194,N_2888);
and U5707 (N_5707,N_2836,N_3604);
nor U5708 (N_5708,N_3432,N_3910);
nand U5709 (N_5709,N_2465,N_2746);
nand U5710 (N_5710,N_2350,N_3992);
nand U5711 (N_5711,N_3762,N_2046);
or U5712 (N_5712,N_3509,N_3219);
nor U5713 (N_5713,N_3897,N_2077);
and U5714 (N_5714,N_2371,N_2183);
or U5715 (N_5715,N_2035,N_2446);
nand U5716 (N_5716,N_2172,N_2655);
nor U5717 (N_5717,N_2274,N_2422);
and U5718 (N_5718,N_2814,N_2023);
and U5719 (N_5719,N_3236,N_3774);
or U5720 (N_5720,N_2795,N_2734);
nor U5721 (N_5721,N_3580,N_3952);
nor U5722 (N_5722,N_2609,N_3814);
nor U5723 (N_5723,N_3360,N_3396);
or U5724 (N_5724,N_3763,N_2427);
and U5725 (N_5725,N_2524,N_2399);
xor U5726 (N_5726,N_2586,N_3988);
nand U5727 (N_5727,N_2134,N_2020);
nor U5728 (N_5728,N_3881,N_2772);
and U5729 (N_5729,N_3953,N_2885);
nor U5730 (N_5730,N_2567,N_3717);
nand U5731 (N_5731,N_2823,N_2440);
and U5732 (N_5732,N_3793,N_2509);
or U5733 (N_5733,N_3123,N_2309);
nor U5734 (N_5734,N_2731,N_2855);
nand U5735 (N_5735,N_2305,N_2774);
or U5736 (N_5736,N_3078,N_2212);
and U5737 (N_5737,N_2217,N_3523);
nand U5738 (N_5738,N_2253,N_3302);
xor U5739 (N_5739,N_3695,N_3870);
and U5740 (N_5740,N_3936,N_3693);
xor U5741 (N_5741,N_2335,N_2507);
nand U5742 (N_5742,N_3940,N_2478);
or U5743 (N_5743,N_2132,N_3487);
and U5744 (N_5744,N_2359,N_2840);
or U5745 (N_5745,N_3341,N_2230);
or U5746 (N_5746,N_2028,N_2327);
nor U5747 (N_5747,N_2274,N_3667);
or U5748 (N_5748,N_2862,N_2544);
and U5749 (N_5749,N_2745,N_3191);
or U5750 (N_5750,N_2133,N_3809);
or U5751 (N_5751,N_2453,N_2462);
or U5752 (N_5752,N_2509,N_3956);
and U5753 (N_5753,N_2321,N_3282);
or U5754 (N_5754,N_2098,N_2605);
nand U5755 (N_5755,N_2668,N_2420);
or U5756 (N_5756,N_3391,N_3715);
or U5757 (N_5757,N_3660,N_3482);
nor U5758 (N_5758,N_2929,N_2272);
nor U5759 (N_5759,N_3751,N_2294);
nor U5760 (N_5760,N_2720,N_3507);
nor U5761 (N_5761,N_3889,N_3134);
nand U5762 (N_5762,N_2430,N_3904);
nand U5763 (N_5763,N_2529,N_2464);
and U5764 (N_5764,N_3548,N_2384);
nor U5765 (N_5765,N_2618,N_3940);
nor U5766 (N_5766,N_2222,N_2044);
nand U5767 (N_5767,N_3592,N_2909);
or U5768 (N_5768,N_3572,N_3053);
nand U5769 (N_5769,N_3041,N_3654);
or U5770 (N_5770,N_2758,N_3476);
and U5771 (N_5771,N_2123,N_2390);
nand U5772 (N_5772,N_2899,N_2120);
nand U5773 (N_5773,N_3251,N_2597);
nand U5774 (N_5774,N_3269,N_3209);
or U5775 (N_5775,N_3167,N_3727);
or U5776 (N_5776,N_2891,N_2863);
or U5777 (N_5777,N_3261,N_3954);
or U5778 (N_5778,N_3474,N_3322);
nor U5779 (N_5779,N_3707,N_3980);
nor U5780 (N_5780,N_3941,N_2937);
and U5781 (N_5781,N_2312,N_2354);
or U5782 (N_5782,N_3167,N_3670);
nand U5783 (N_5783,N_3460,N_3587);
nor U5784 (N_5784,N_3898,N_2115);
or U5785 (N_5785,N_3176,N_3961);
and U5786 (N_5786,N_3055,N_3123);
or U5787 (N_5787,N_3397,N_2656);
xnor U5788 (N_5788,N_3839,N_2351);
nor U5789 (N_5789,N_3201,N_2524);
and U5790 (N_5790,N_2321,N_2220);
nand U5791 (N_5791,N_2925,N_3077);
xnor U5792 (N_5792,N_2038,N_2206);
or U5793 (N_5793,N_3119,N_2764);
nand U5794 (N_5794,N_3421,N_2194);
nor U5795 (N_5795,N_3420,N_2232);
xnor U5796 (N_5796,N_2820,N_2761);
or U5797 (N_5797,N_2193,N_2083);
and U5798 (N_5798,N_2715,N_3758);
xor U5799 (N_5799,N_2598,N_3245);
nor U5800 (N_5800,N_2665,N_2622);
or U5801 (N_5801,N_3026,N_3001);
nand U5802 (N_5802,N_3692,N_3065);
or U5803 (N_5803,N_2257,N_3858);
nand U5804 (N_5804,N_3106,N_2139);
nor U5805 (N_5805,N_3085,N_2264);
or U5806 (N_5806,N_3977,N_3336);
and U5807 (N_5807,N_2502,N_3728);
or U5808 (N_5808,N_3491,N_3596);
and U5809 (N_5809,N_2849,N_2372);
nand U5810 (N_5810,N_2278,N_3809);
nand U5811 (N_5811,N_3423,N_2669);
nor U5812 (N_5812,N_2521,N_2010);
nand U5813 (N_5813,N_3436,N_2044);
and U5814 (N_5814,N_3341,N_2305);
xnor U5815 (N_5815,N_3000,N_2236);
nand U5816 (N_5816,N_3732,N_3286);
nand U5817 (N_5817,N_3836,N_2622);
or U5818 (N_5818,N_2927,N_2926);
nand U5819 (N_5819,N_2123,N_2721);
nor U5820 (N_5820,N_3405,N_2103);
and U5821 (N_5821,N_2435,N_3373);
or U5822 (N_5822,N_2448,N_2912);
or U5823 (N_5823,N_3723,N_2846);
nor U5824 (N_5824,N_2212,N_2198);
or U5825 (N_5825,N_3430,N_3375);
or U5826 (N_5826,N_2712,N_3700);
and U5827 (N_5827,N_3105,N_3550);
nand U5828 (N_5828,N_2993,N_3956);
and U5829 (N_5829,N_2721,N_2740);
nor U5830 (N_5830,N_3431,N_2469);
nor U5831 (N_5831,N_3995,N_2375);
nor U5832 (N_5832,N_2822,N_3823);
and U5833 (N_5833,N_2463,N_3736);
nor U5834 (N_5834,N_3588,N_2765);
nor U5835 (N_5835,N_3841,N_2400);
nand U5836 (N_5836,N_3916,N_3455);
xor U5837 (N_5837,N_3819,N_2736);
nor U5838 (N_5838,N_3424,N_2114);
and U5839 (N_5839,N_3787,N_2942);
nand U5840 (N_5840,N_2799,N_2465);
and U5841 (N_5841,N_3414,N_2499);
nor U5842 (N_5842,N_3234,N_2499);
and U5843 (N_5843,N_2728,N_3046);
nand U5844 (N_5844,N_3224,N_3384);
nand U5845 (N_5845,N_3028,N_3300);
nor U5846 (N_5846,N_3480,N_2811);
and U5847 (N_5847,N_3691,N_3546);
and U5848 (N_5848,N_2341,N_2361);
and U5849 (N_5849,N_2048,N_3644);
nand U5850 (N_5850,N_2934,N_2913);
nand U5851 (N_5851,N_2992,N_2867);
and U5852 (N_5852,N_2693,N_2832);
or U5853 (N_5853,N_2761,N_3523);
nor U5854 (N_5854,N_3353,N_2858);
nor U5855 (N_5855,N_2719,N_3665);
nor U5856 (N_5856,N_3576,N_3932);
nand U5857 (N_5857,N_3538,N_2050);
and U5858 (N_5858,N_3771,N_3369);
or U5859 (N_5859,N_2162,N_3472);
nand U5860 (N_5860,N_2072,N_2054);
xor U5861 (N_5861,N_2064,N_3887);
or U5862 (N_5862,N_2536,N_2539);
nand U5863 (N_5863,N_2747,N_2804);
or U5864 (N_5864,N_3449,N_3471);
nor U5865 (N_5865,N_3025,N_3389);
nand U5866 (N_5866,N_3404,N_3967);
and U5867 (N_5867,N_2837,N_2584);
or U5868 (N_5868,N_2390,N_3181);
xor U5869 (N_5869,N_3510,N_3611);
or U5870 (N_5870,N_3183,N_2510);
or U5871 (N_5871,N_3452,N_3859);
or U5872 (N_5872,N_3880,N_3259);
or U5873 (N_5873,N_2701,N_3904);
nand U5874 (N_5874,N_2616,N_2503);
nor U5875 (N_5875,N_2364,N_3272);
and U5876 (N_5876,N_2628,N_2563);
nor U5877 (N_5877,N_2702,N_2648);
nor U5878 (N_5878,N_3406,N_3389);
or U5879 (N_5879,N_3903,N_2220);
nand U5880 (N_5880,N_3116,N_3898);
and U5881 (N_5881,N_3338,N_3224);
or U5882 (N_5882,N_3426,N_3610);
nor U5883 (N_5883,N_3299,N_3285);
xnor U5884 (N_5884,N_2499,N_3621);
nand U5885 (N_5885,N_3003,N_3001);
or U5886 (N_5886,N_3516,N_3931);
nor U5887 (N_5887,N_3180,N_3387);
or U5888 (N_5888,N_2387,N_2928);
and U5889 (N_5889,N_3522,N_3379);
nand U5890 (N_5890,N_3958,N_2380);
or U5891 (N_5891,N_2822,N_3798);
and U5892 (N_5892,N_3463,N_3067);
or U5893 (N_5893,N_2696,N_2353);
and U5894 (N_5894,N_3398,N_2481);
nand U5895 (N_5895,N_3922,N_3617);
nand U5896 (N_5896,N_2773,N_3261);
nor U5897 (N_5897,N_3639,N_3584);
nand U5898 (N_5898,N_2671,N_2857);
nor U5899 (N_5899,N_2889,N_3744);
nor U5900 (N_5900,N_3587,N_2781);
nand U5901 (N_5901,N_2505,N_3161);
and U5902 (N_5902,N_2334,N_2818);
nand U5903 (N_5903,N_3458,N_2997);
or U5904 (N_5904,N_3774,N_2631);
nand U5905 (N_5905,N_3760,N_3518);
nand U5906 (N_5906,N_2976,N_3820);
nand U5907 (N_5907,N_2100,N_3782);
nor U5908 (N_5908,N_2560,N_3261);
nor U5909 (N_5909,N_3656,N_3623);
nor U5910 (N_5910,N_3579,N_3578);
and U5911 (N_5911,N_3391,N_3219);
nand U5912 (N_5912,N_3346,N_3219);
nor U5913 (N_5913,N_3140,N_2682);
and U5914 (N_5914,N_3148,N_2116);
or U5915 (N_5915,N_3389,N_3978);
or U5916 (N_5916,N_2501,N_3903);
and U5917 (N_5917,N_2456,N_2763);
nand U5918 (N_5918,N_2096,N_3861);
nand U5919 (N_5919,N_2260,N_3445);
nor U5920 (N_5920,N_3120,N_3304);
nand U5921 (N_5921,N_3689,N_2669);
or U5922 (N_5922,N_2820,N_2666);
nand U5923 (N_5923,N_3262,N_2222);
and U5924 (N_5924,N_2142,N_2055);
and U5925 (N_5925,N_2088,N_2743);
nor U5926 (N_5926,N_2822,N_2145);
nor U5927 (N_5927,N_2252,N_2047);
or U5928 (N_5928,N_3537,N_2656);
nand U5929 (N_5929,N_2792,N_2245);
or U5930 (N_5930,N_3935,N_2322);
nand U5931 (N_5931,N_3180,N_3323);
nand U5932 (N_5932,N_3011,N_3615);
nor U5933 (N_5933,N_2801,N_3360);
nand U5934 (N_5934,N_2544,N_3141);
nand U5935 (N_5935,N_3559,N_3241);
and U5936 (N_5936,N_3848,N_2923);
or U5937 (N_5937,N_2870,N_2623);
or U5938 (N_5938,N_3210,N_3897);
and U5939 (N_5939,N_3373,N_3967);
nand U5940 (N_5940,N_3619,N_3218);
or U5941 (N_5941,N_2835,N_3740);
or U5942 (N_5942,N_2031,N_3735);
or U5943 (N_5943,N_2235,N_2033);
or U5944 (N_5944,N_2874,N_3090);
xor U5945 (N_5945,N_3470,N_3209);
and U5946 (N_5946,N_2296,N_3194);
nand U5947 (N_5947,N_3846,N_3927);
and U5948 (N_5948,N_3872,N_3507);
nand U5949 (N_5949,N_3666,N_3915);
and U5950 (N_5950,N_2270,N_2005);
nand U5951 (N_5951,N_2283,N_3371);
and U5952 (N_5952,N_2282,N_2503);
nand U5953 (N_5953,N_2934,N_3680);
and U5954 (N_5954,N_2590,N_2056);
or U5955 (N_5955,N_3264,N_3536);
nor U5956 (N_5956,N_3920,N_2897);
xnor U5957 (N_5957,N_3984,N_3934);
nand U5958 (N_5958,N_3883,N_3076);
nand U5959 (N_5959,N_2391,N_3342);
nand U5960 (N_5960,N_2741,N_3319);
or U5961 (N_5961,N_3400,N_2427);
nor U5962 (N_5962,N_2202,N_3656);
nor U5963 (N_5963,N_2525,N_2015);
and U5964 (N_5964,N_2813,N_3671);
or U5965 (N_5965,N_2236,N_2519);
or U5966 (N_5966,N_3425,N_2714);
or U5967 (N_5967,N_3348,N_3452);
or U5968 (N_5968,N_3369,N_3950);
or U5969 (N_5969,N_3657,N_2599);
nor U5970 (N_5970,N_3056,N_2998);
or U5971 (N_5971,N_3014,N_3839);
xor U5972 (N_5972,N_3306,N_2080);
nor U5973 (N_5973,N_2108,N_3650);
or U5974 (N_5974,N_2553,N_2148);
nand U5975 (N_5975,N_2526,N_2994);
or U5976 (N_5976,N_2371,N_2355);
and U5977 (N_5977,N_3652,N_3785);
or U5978 (N_5978,N_3569,N_2739);
nor U5979 (N_5979,N_2360,N_2889);
or U5980 (N_5980,N_3336,N_2090);
and U5981 (N_5981,N_2817,N_2117);
nand U5982 (N_5982,N_3765,N_2068);
and U5983 (N_5983,N_2624,N_2640);
and U5984 (N_5984,N_2223,N_3774);
or U5985 (N_5985,N_2250,N_2640);
or U5986 (N_5986,N_2285,N_3873);
or U5987 (N_5987,N_2595,N_3149);
or U5988 (N_5988,N_3091,N_3521);
xor U5989 (N_5989,N_2695,N_3882);
nand U5990 (N_5990,N_3385,N_2414);
and U5991 (N_5991,N_2407,N_3698);
nand U5992 (N_5992,N_2154,N_3033);
nor U5993 (N_5993,N_3817,N_2916);
and U5994 (N_5994,N_2225,N_2132);
and U5995 (N_5995,N_2620,N_2452);
nor U5996 (N_5996,N_2627,N_2659);
nor U5997 (N_5997,N_3166,N_2788);
or U5998 (N_5998,N_3350,N_3096);
nand U5999 (N_5999,N_2297,N_2993);
nand U6000 (N_6000,N_5276,N_5940);
nand U6001 (N_6001,N_5526,N_4898);
nand U6002 (N_6002,N_5970,N_4641);
nor U6003 (N_6003,N_4396,N_4693);
and U6004 (N_6004,N_5546,N_5538);
and U6005 (N_6005,N_4697,N_5464);
or U6006 (N_6006,N_4804,N_4805);
or U6007 (N_6007,N_5404,N_5254);
nor U6008 (N_6008,N_5146,N_4681);
or U6009 (N_6009,N_5859,N_5542);
or U6010 (N_6010,N_4564,N_4537);
nand U6011 (N_6011,N_5716,N_5525);
nor U6012 (N_6012,N_4787,N_4595);
nor U6013 (N_6013,N_5697,N_4116);
and U6014 (N_6014,N_4470,N_4007);
or U6015 (N_6015,N_4074,N_4063);
nor U6016 (N_6016,N_5650,N_4921);
and U6017 (N_6017,N_5127,N_5971);
nor U6018 (N_6018,N_5961,N_5363);
nor U6019 (N_6019,N_4860,N_4411);
nor U6020 (N_6020,N_5810,N_4381);
or U6021 (N_6021,N_5453,N_5067);
nor U6022 (N_6022,N_4746,N_5843);
or U6023 (N_6023,N_4391,N_5459);
and U6024 (N_6024,N_5574,N_5573);
and U6025 (N_6025,N_4633,N_5735);
and U6026 (N_6026,N_4530,N_5962);
or U6027 (N_6027,N_5243,N_5352);
and U6028 (N_6028,N_5693,N_4900);
and U6029 (N_6029,N_5071,N_4496);
or U6030 (N_6030,N_5303,N_5417);
nand U6031 (N_6031,N_4920,N_4150);
and U6032 (N_6032,N_4613,N_5522);
nand U6033 (N_6033,N_5084,N_4687);
nor U6034 (N_6034,N_4549,N_4209);
and U6035 (N_6035,N_5533,N_4977);
or U6036 (N_6036,N_5783,N_4826);
or U6037 (N_6037,N_5823,N_5437);
nand U6038 (N_6038,N_5186,N_5458);
nor U6039 (N_6039,N_4838,N_4745);
nor U6040 (N_6040,N_4081,N_5981);
or U6041 (N_6041,N_4705,N_5428);
and U6042 (N_6042,N_4297,N_4741);
or U6043 (N_6043,N_4713,N_4991);
or U6044 (N_6044,N_4506,N_5733);
and U6045 (N_6045,N_5196,N_4191);
and U6046 (N_6046,N_5696,N_4199);
nand U6047 (N_6047,N_5892,N_4281);
nor U6048 (N_6048,N_4563,N_5681);
or U6049 (N_6049,N_5394,N_5021);
and U6050 (N_6050,N_5909,N_5711);
and U6051 (N_6051,N_4056,N_4660);
and U6052 (N_6052,N_5708,N_4645);
xnor U6053 (N_6053,N_4022,N_4300);
and U6054 (N_6054,N_5110,N_4169);
nand U6055 (N_6055,N_5361,N_4737);
or U6056 (N_6056,N_4485,N_4398);
or U6057 (N_6057,N_5260,N_4243);
nor U6058 (N_6058,N_4088,N_5555);
nand U6059 (N_6059,N_5806,N_4401);
nor U6060 (N_6060,N_4782,N_5866);
and U6061 (N_6061,N_4943,N_5986);
nor U6062 (N_6062,N_5275,N_4064);
nand U6063 (N_6063,N_5956,N_5504);
nand U6064 (N_6064,N_5601,N_4053);
or U6065 (N_6065,N_4791,N_4904);
nand U6066 (N_6066,N_5562,N_5198);
nand U6067 (N_6067,N_4195,N_5614);
nand U6068 (N_6068,N_5801,N_5158);
nor U6069 (N_6069,N_4431,N_4954);
nand U6070 (N_6070,N_5671,N_4380);
nand U6071 (N_6071,N_5807,N_5759);
nand U6072 (N_6072,N_5982,N_5818);
nor U6073 (N_6073,N_4141,N_4334);
or U6074 (N_6074,N_4201,N_5354);
nor U6075 (N_6075,N_4447,N_5532);
or U6076 (N_6076,N_4212,N_4492);
nor U6077 (N_6077,N_4665,N_4780);
or U6078 (N_6078,N_4942,N_5132);
nand U6079 (N_6079,N_5990,N_4200);
nor U6080 (N_6080,N_5025,N_4952);
nand U6081 (N_6081,N_4117,N_5133);
nor U6082 (N_6082,N_5894,N_5092);
xnor U6083 (N_6083,N_4257,N_5090);
nand U6084 (N_6084,N_5151,N_4123);
or U6085 (N_6085,N_5957,N_4129);
or U6086 (N_6086,N_5229,N_4462);
nand U6087 (N_6087,N_5610,N_4285);
or U6088 (N_6088,N_5030,N_4925);
nor U6089 (N_6089,N_4541,N_4649);
or U6090 (N_6090,N_4744,N_4430);
or U6091 (N_6091,N_4365,N_4813);
and U6092 (N_6092,N_4863,N_5934);
and U6093 (N_6093,N_5495,N_4455);
and U6094 (N_6094,N_5491,N_4103);
nor U6095 (N_6095,N_4426,N_5215);
or U6096 (N_6096,N_4717,N_5479);
and U6097 (N_6097,N_5509,N_4254);
nand U6098 (N_6098,N_4956,N_5435);
nor U6099 (N_6099,N_4998,N_5730);
or U6100 (N_6100,N_5753,N_5480);
nor U6101 (N_6101,N_5689,N_5036);
or U6102 (N_6102,N_5670,N_4912);
or U6103 (N_6103,N_5192,N_5489);
and U6104 (N_6104,N_4870,N_5168);
or U6105 (N_6105,N_5618,N_5413);
and U6106 (N_6106,N_5863,N_4301);
and U6107 (N_6107,N_4131,N_4025);
nand U6108 (N_6108,N_4743,N_4054);
and U6109 (N_6109,N_5919,N_4683);
or U6110 (N_6110,N_5377,N_4815);
xor U6111 (N_6111,N_4397,N_5299);
nand U6112 (N_6112,N_4030,N_5703);
nor U6113 (N_6113,N_4983,N_5790);
nor U6114 (N_6114,N_4695,N_4338);
or U6115 (N_6115,N_5855,N_4070);
and U6116 (N_6116,N_5655,N_4501);
nand U6117 (N_6117,N_5821,N_5584);
or U6118 (N_6118,N_5472,N_4679);
and U6119 (N_6119,N_5993,N_4729);
and U6120 (N_6120,N_4266,N_5668);
nand U6121 (N_6121,N_4072,N_5019);
nor U6122 (N_6122,N_4769,N_5266);
nor U6123 (N_6123,N_4119,N_5579);
and U6124 (N_6124,N_4929,N_5302);
and U6125 (N_6125,N_5322,N_4042);
nand U6126 (N_6126,N_5007,N_4189);
and U6127 (N_6127,N_4092,N_4037);
nor U6128 (N_6128,N_5000,N_5969);
and U6129 (N_6129,N_5131,N_5033);
and U6130 (N_6130,N_5627,N_5604);
nand U6131 (N_6131,N_4934,N_4557);
nor U6132 (N_6132,N_4049,N_4640);
nor U6133 (N_6133,N_5461,N_5086);
and U6134 (N_6134,N_4754,N_5297);
nand U6135 (N_6135,N_5054,N_4188);
or U6136 (N_6136,N_5200,N_4614);
or U6137 (N_6137,N_4638,N_4764);
nand U6138 (N_6138,N_4132,N_4786);
nor U6139 (N_6139,N_5028,N_5365);
and U6140 (N_6140,N_4024,N_5193);
xor U6141 (N_6141,N_5085,N_5176);
or U6142 (N_6142,N_4250,N_5093);
and U6143 (N_6143,N_4948,N_5157);
nand U6144 (N_6144,N_5656,N_5315);
and U6145 (N_6145,N_5220,N_5933);
nand U6146 (N_6146,N_4153,N_5713);
and U6147 (N_6147,N_5384,N_4617);
nor U6148 (N_6148,N_4253,N_4521);
nor U6149 (N_6149,N_4663,N_5166);
nand U6150 (N_6150,N_5439,N_5485);
and U6151 (N_6151,N_4124,N_4482);
or U6152 (N_6152,N_5442,N_5184);
and U6153 (N_6153,N_4794,N_4505);
and U6154 (N_6154,N_5122,N_5293);
and U6155 (N_6155,N_4567,N_4963);
nor U6156 (N_6156,N_4477,N_5372);
nand U6157 (N_6157,N_5420,N_5646);
or U6158 (N_6158,N_5106,N_5989);
nor U6159 (N_6159,N_5660,N_5065);
nor U6160 (N_6160,N_5159,N_4938);
or U6161 (N_6161,N_4583,N_5490);
and U6162 (N_6162,N_4644,N_4849);
or U6163 (N_6163,N_4015,N_4524);
or U6164 (N_6164,N_5182,N_5865);
nor U6165 (N_6165,N_5273,N_5597);
or U6166 (N_6166,N_4601,N_4205);
and U6167 (N_6167,N_5864,N_5486);
or U6168 (N_6168,N_5683,N_5207);
and U6169 (N_6169,N_5027,N_5046);
nor U6170 (N_6170,N_5882,N_4476);
nand U6171 (N_6171,N_5916,N_4923);
or U6172 (N_6172,N_4127,N_4185);
nand U6173 (N_6173,N_4386,N_5550);
nor U6174 (N_6174,N_5852,N_4594);
and U6175 (N_6175,N_4709,N_4115);
and U6176 (N_6176,N_4655,N_5252);
nor U6177 (N_6177,N_5272,N_4176);
nand U6178 (N_6178,N_4003,N_4384);
xnor U6179 (N_6179,N_5945,N_4472);
nor U6180 (N_6180,N_4167,N_5487);
or U6181 (N_6181,N_4371,N_5897);
nand U6182 (N_6182,N_5635,N_5400);
nand U6183 (N_6183,N_5399,N_4507);
nand U6184 (N_6184,N_4690,N_4678);
nor U6185 (N_6185,N_5942,N_5457);
and U6186 (N_6186,N_5494,N_4303);
nand U6187 (N_6187,N_4634,N_4722);
nand U6188 (N_6188,N_5976,N_4936);
nand U6189 (N_6189,N_4619,N_5779);
and U6190 (N_6190,N_4891,N_5633);
xor U6191 (N_6191,N_4783,N_4996);
nand U6192 (N_6192,N_5572,N_4359);
or U6193 (N_6193,N_4436,N_4354);
or U6194 (N_6194,N_4779,N_5463);
nand U6195 (N_6195,N_5838,N_4287);
or U6196 (N_6196,N_5125,N_5230);
nor U6197 (N_6197,N_5382,N_5740);
and U6198 (N_6198,N_4930,N_5714);
nand U6199 (N_6199,N_4036,N_4816);
or U6200 (N_6200,N_4945,N_5747);
or U6201 (N_6201,N_4890,N_4913);
nand U6202 (N_6202,N_5763,N_5544);
and U6203 (N_6203,N_4256,N_5985);
nor U6204 (N_6204,N_5163,N_4238);
nand U6205 (N_6205,N_5422,N_5388);
and U6206 (N_6206,N_5850,N_5418);
nand U6207 (N_6207,N_4880,N_5652);
nor U6208 (N_6208,N_4383,N_5621);
and U6209 (N_6209,N_4146,N_5910);
nand U6210 (N_6210,N_5804,N_4158);
nand U6211 (N_6211,N_5760,N_5819);
nand U6212 (N_6212,N_4551,N_5034);
and U6213 (N_6213,N_4822,N_4967);
or U6214 (N_6214,N_5815,N_5172);
or U6215 (N_6215,N_4527,N_4082);
nand U6216 (N_6216,N_4790,N_5124);
nand U6217 (N_6217,N_5732,N_5396);
and U6218 (N_6218,N_5875,N_4284);
or U6219 (N_6219,N_5424,N_4855);
nor U6220 (N_6220,N_5160,N_5954);
nor U6221 (N_6221,N_5212,N_5039);
nand U6222 (N_6222,N_5261,N_5427);
nand U6223 (N_6223,N_5996,N_4953);
nor U6224 (N_6224,N_5419,N_5355);
or U6225 (N_6225,N_5165,N_5911);
nor U6226 (N_6226,N_5925,N_5140);
nand U6227 (N_6227,N_5283,N_5748);
nor U6228 (N_6228,N_5348,N_4667);
nor U6229 (N_6229,N_5290,N_4376);
nor U6230 (N_6230,N_4211,N_4348);
nor U6231 (N_6231,N_4475,N_5698);
nand U6232 (N_6232,N_4484,N_4445);
nand U6233 (N_6233,N_4770,N_4593);
nor U6234 (N_6234,N_4908,N_5280);
nand U6235 (N_6235,N_4226,N_4576);
nor U6236 (N_6236,N_4612,N_5612);
nand U6237 (N_6237,N_5827,N_4407);
nand U6238 (N_6238,N_4801,N_4706);
and U6239 (N_6239,N_5665,N_4701);
or U6240 (N_6240,N_5690,N_5802);
or U6241 (N_6241,N_5073,N_4197);
nand U6242 (N_6242,N_4155,N_4105);
nand U6243 (N_6243,N_4387,N_4424);
nor U6244 (N_6244,N_5104,N_4421);
and U6245 (N_6245,N_5288,N_4444);
nor U6246 (N_6246,N_5374,N_4452);
and U6247 (N_6247,N_5939,N_4811);
and U6248 (N_6248,N_4824,N_4219);
or U6249 (N_6249,N_5586,N_5143);
nor U6250 (N_6250,N_5587,N_5839);
xnor U6251 (N_6251,N_5590,N_5038);
and U6252 (N_6252,N_5245,N_5792);
or U6253 (N_6253,N_5923,N_5944);
nor U6254 (N_6254,N_4029,N_5846);
or U6255 (N_6255,N_4223,N_5318);
and U6256 (N_6256,N_4728,N_4958);
or U6257 (N_6257,N_5626,N_4393);
nor U6258 (N_6258,N_4218,N_4481);
nor U6259 (N_6259,N_4145,N_5906);
nor U6260 (N_6260,N_4494,N_4214);
or U6261 (N_6261,N_5251,N_4572);
nor U6262 (N_6262,N_4460,N_5031);
or U6263 (N_6263,N_4349,N_4394);
and U6264 (N_6264,N_5503,N_5285);
nand U6265 (N_6265,N_5351,N_4261);
and U6266 (N_6266,N_4216,N_5430);
nor U6267 (N_6267,N_4671,N_5178);
and U6268 (N_6268,N_4162,N_5367);
nand U6269 (N_6269,N_4242,N_5726);
nor U6270 (N_6270,N_4159,N_4710);
or U6271 (N_6271,N_5975,N_4997);
nor U6272 (N_6272,N_5069,N_5529);
nor U6273 (N_6273,N_5095,N_5780);
nor U6274 (N_6274,N_4546,N_4275);
nand U6275 (N_6275,N_5861,N_5840);
or U6276 (N_6276,N_4964,N_5265);
nand U6277 (N_6277,N_4206,N_4775);
or U6278 (N_6278,N_5425,N_5171);
nand U6279 (N_6279,N_4172,N_5967);
and U6280 (N_6280,N_4766,N_5258);
and U6281 (N_6281,N_4038,N_5239);
nand U6282 (N_6282,N_5672,N_4885);
and U6283 (N_6283,N_5682,N_5702);
and U6284 (N_6284,N_5530,N_5543);
nor U6285 (N_6285,N_4500,N_5615);
nor U6286 (N_6286,N_5219,N_5210);
and U6287 (N_6287,N_4662,N_5473);
and U6288 (N_6288,N_5551,N_5568);
or U6289 (N_6289,N_4535,N_5515);
nand U6290 (N_6290,N_5235,N_4305);
nor U6291 (N_6291,N_5891,N_5750);
and U6292 (N_6292,N_4165,N_5808);
nor U6293 (N_6293,N_4708,N_5331);
nor U6294 (N_6294,N_4879,N_4843);
nor U6295 (N_6295,N_4802,N_4949);
nor U6296 (N_6296,N_4198,N_4310);
nand U6297 (N_6297,N_4316,N_5605);
nor U6298 (N_6298,N_4555,N_5088);
and U6299 (N_6299,N_4392,N_5772);
and U6300 (N_6300,N_5216,N_4837);
or U6301 (N_6301,N_5994,N_5075);
or U6302 (N_6302,N_4184,N_4360);
or U6303 (N_6303,N_5262,N_4307);
or U6304 (N_6304,N_5599,N_5598);
and U6305 (N_6305,N_5173,N_5421);
nor U6306 (N_6306,N_5842,N_5032);
nand U6307 (N_6307,N_4881,N_5679);
and U6308 (N_6308,N_4590,N_4433);
nand U6309 (N_6309,N_4122,N_4408);
nor U6310 (N_6310,N_5856,N_4539);
nand U6311 (N_6311,N_4096,N_5052);
nand U6312 (N_6312,N_5329,N_5521);
nand U6313 (N_6313,N_5594,N_5185);
xnor U6314 (N_6314,N_4268,N_4732);
nor U6315 (N_6315,N_5582,N_5770);
or U6316 (N_6316,N_5978,N_5246);
xor U6317 (N_6317,N_5510,N_5798);
and U6318 (N_6318,N_4700,N_5816);
xor U6319 (N_6319,N_5121,N_5217);
and U6320 (N_6320,N_4894,N_5247);
or U6321 (N_6321,N_5447,N_4463);
or U6322 (N_6322,N_5500,N_5545);
nor U6323 (N_6323,N_4324,N_4438);
and U6324 (N_6324,N_5402,N_4752);
nor U6325 (N_6325,N_4762,N_5316);
nand U6326 (N_6326,N_4114,N_4186);
nor U6327 (N_6327,N_4298,N_5519);
and U6328 (N_6328,N_5123,N_4137);
and U6329 (N_6329,N_4323,N_5871);
or U6330 (N_6330,N_4556,N_4570);
or U6331 (N_6331,N_5685,N_5883);
or U6332 (N_6332,N_5931,N_4512);
nand U6333 (N_6333,N_5277,N_4988);
nand U6334 (N_6334,N_4536,N_4224);
nand U6335 (N_6335,N_5547,N_4819);
or U6336 (N_6336,N_4418,N_4043);
nor U6337 (N_6337,N_4062,N_4659);
or U6338 (N_6338,N_4058,N_4917);
nor U6339 (N_6339,N_4727,N_4410);
and U6340 (N_6340,N_4367,N_4357);
nor U6341 (N_6341,N_4085,N_5412);
and U6342 (N_6342,N_5003,N_5609);
or U6343 (N_6343,N_5640,N_5403);
nand U6344 (N_6344,N_4026,N_5407);
or U6345 (N_6345,N_4899,N_4130);
nor U6346 (N_6346,N_5869,N_5870);
or U6347 (N_6347,N_4561,N_4178);
and U6348 (N_6348,N_5832,N_4856);
nand U6349 (N_6349,N_4304,N_4987);
and U6350 (N_6350,N_4255,N_4797);
or U6351 (N_6351,N_5536,N_5409);
or U6352 (N_6352,N_4947,N_5965);
and U6353 (N_6353,N_4836,N_4731);
nand U6354 (N_6354,N_4544,N_4499);
or U6355 (N_6355,N_5449,N_5868);
and U6356 (N_6356,N_4399,N_4451);
and U6357 (N_6357,N_5248,N_4571);
or U6358 (N_6358,N_5777,N_4467);
nor U6359 (N_6359,N_4312,N_5773);
or U6360 (N_6360,N_5799,N_4847);
and U6361 (N_6361,N_4635,N_5333);
nand U6362 (N_6362,N_5170,N_4453);
and U6363 (N_6363,N_5233,N_5145);
nor U6364 (N_6364,N_4013,N_4340);
nand U6365 (N_6365,N_5150,N_5886);
or U6366 (N_6366,N_5053,N_5757);
nor U6367 (N_6367,N_5082,N_4345);
or U6368 (N_6368,N_4441,N_5593);
or U6369 (N_6369,N_4757,N_4259);
nor U6370 (N_6370,N_5356,N_5794);
and U6371 (N_6371,N_5712,N_5234);
nand U6372 (N_6372,N_5287,N_4874);
nand U6373 (N_6373,N_4372,N_5398);
nor U6374 (N_6374,N_4134,N_4810);
nand U6375 (N_6375,N_5507,N_5136);
or U6376 (N_6376,N_4069,N_4866);
nand U6377 (N_6377,N_4578,N_4008);
and U6378 (N_6378,N_5410,N_5721);
nor U6379 (N_6379,N_4857,N_4339);
nand U6380 (N_6380,N_4108,N_4631);
xor U6381 (N_6381,N_4985,N_5332);
nand U6382 (N_6382,N_5887,N_4052);
nand U6383 (N_6383,N_4210,N_5174);
and U6384 (N_6384,N_5921,N_5775);
and U6385 (N_6385,N_5765,N_4968);
or U6386 (N_6386,N_5904,N_5624);
or U6387 (N_6387,N_4245,N_5222);
and U6388 (N_6388,N_4151,N_4677);
or U6389 (N_6389,N_4852,N_4887);
and U6390 (N_6390,N_5224,N_4781);
and U6391 (N_6391,N_5321,N_4853);
and U6392 (N_6392,N_4498,N_5596);
nand U6393 (N_6393,N_5769,N_5844);
nor U6394 (N_6394,N_4009,N_5126);
or U6395 (N_6395,N_5817,N_5194);
and U6396 (N_6396,N_5066,N_5873);
nor U6397 (N_6397,N_5669,N_5205);
and U6398 (N_6398,N_5161,N_5860);
and U6399 (N_6399,N_4402,N_5674);
or U6400 (N_6400,N_4632,N_4630);
nor U6401 (N_6401,N_5269,N_4939);
nor U6402 (N_6402,N_4183,N_5386);
and U6403 (N_6403,N_4932,N_4960);
or U6404 (N_6404,N_5440,N_4689);
or U6405 (N_6405,N_4886,N_5050);
and U6406 (N_6406,N_5045,N_4439);
or U6407 (N_6407,N_4286,N_4425);
and U6408 (N_6408,N_4730,N_5636);
nand U6409 (N_6409,N_4280,N_4374);
nor U6410 (N_6410,N_4233,N_5049);
or U6411 (N_6411,N_5936,N_4629);
nand U6412 (N_6412,N_5024,N_4903);
or U6413 (N_6413,N_5040,N_4423);
nor U6414 (N_6414,N_5446,N_4464);
nand U6415 (N_6415,N_4528,N_4370);
nor U6416 (N_6416,N_4771,N_4154);
or U6417 (N_6417,N_4272,N_5401);
and U6418 (N_6418,N_5884,N_4763);
or U6419 (N_6419,N_4249,N_5411);
and U6420 (N_6420,N_5647,N_4414);
nand U6421 (N_6421,N_5959,N_5317);
nand U6422 (N_6422,N_4691,N_5520);
or U6423 (N_6423,N_5687,N_4547);
nor U6424 (N_6424,N_5102,N_5531);
nor U6425 (N_6425,N_4861,N_5236);
nor U6426 (N_6426,N_4066,N_5788);
nor U6427 (N_6427,N_4133,N_5736);
and U6428 (N_6428,N_5513,N_5922);
nor U6429 (N_6429,N_4094,N_5152);
xor U6430 (N_6430,N_4335,N_4704);
nand U6431 (N_6431,N_4461,N_5116);
xor U6432 (N_6432,N_4919,N_4509);
or U6433 (N_6433,N_4760,N_4288);
or U6434 (N_6434,N_5279,N_5096);
nor U6435 (N_6435,N_5414,N_4497);
and U6436 (N_6436,N_5432,N_4672);
or U6437 (N_6437,N_5137,N_5481);
nor U6438 (N_6438,N_4041,N_4006);
nor U6439 (N_6439,N_5537,N_5048);
nor U6440 (N_6440,N_4656,N_5841);
and U6441 (N_6441,N_5629,N_5468);
and U6442 (N_6442,N_5013,N_5080);
nor U6443 (N_6443,N_5357,N_4795);
or U6444 (N_6444,N_4579,N_5998);
or U6445 (N_6445,N_4814,N_4217);
nor U6446 (N_6446,N_4271,N_4876);
nor U6447 (N_6447,N_4718,N_4566);
nor U6448 (N_6448,N_5089,N_5534);
nand U6449 (N_6449,N_4865,N_4180);
nor U6450 (N_6450,N_4742,N_5341);
xor U6451 (N_6451,N_5701,N_5578);
or U6452 (N_6452,N_4282,N_4552);
nand U6453 (N_6453,N_5709,N_5301);
or U6454 (N_6454,N_5988,N_5901);
nor U6455 (N_6455,N_4610,N_5436);
or U6456 (N_6456,N_4283,N_5072);
nand U6457 (N_6457,N_5183,N_5781);
nor U6458 (N_6458,N_4698,N_5270);
xnor U6459 (N_6459,N_5583,N_5334);
nor U6460 (N_6460,N_5314,N_5666);
and U6461 (N_6461,N_4264,N_4168);
or U6462 (N_6462,N_4785,N_4979);
or U6463 (N_6463,N_4896,N_4712);
nor U6464 (N_6464,N_4000,N_5099);
or U6465 (N_6465,N_4543,N_4673);
and U6466 (N_6466,N_4845,N_5567);
and U6467 (N_6467,N_5876,N_4237);
and U6468 (N_6468,N_5395,N_4336);
nand U6469 (N_6469,N_4927,N_4835);
or U6470 (N_6470,N_5180,N_5857);
nand U6471 (N_6471,N_5528,N_5958);
nand U6472 (N_6472,N_5762,N_5115);
and U6473 (N_6473,N_4193,N_4390);
xnor U6474 (N_6474,N_5899,N_4488);
and U6475 (N_6475,N_5675,N_4406);
and U6476 (N_6476,N_4846,N_5813);
nand U6477 (N_6477,N_4653,N_4067);
or U6478 (N_6478,N_4019,N_4799);
nor U6479 (N_6479,N_4738,N_4194);
and U6480 (N_6480,N_4443,N_5787);
nand U6481 (N_6481,N_5606,N_5103);
nand U6482 (N_6482,N_5426,N_4721);
nand U6483 (N_6483,N_4696,N_5619);
and U6484 (N_6484,N_4263,N_5699);
nor U6485 (N_6485,N_5786,N_5878);
nor U6486 (N_6486,N_4525,N_4035);
or U6487 (N_6487,N_4778,N_5035);
nor U6488 (N_6488,N_4841,N_4608);
and U6489 (N_6489,N_5292,N_4664);
nor U6490 (N_6490,N_5613,N_4888);
or U6491 (N_6491,N_4493,N_5077);
or U6492 (N_6492,N_4582,N_5704);
or U6493 (N_6493,N_5493,N_5890);
nand U6494 (N_6494,N_5305,N_4596);
nor U6495 (N_6495,N_4429,N_4676);
and U6496 (N_6496,N_4120,N_5415);
nand U6497 (N_6497,N_5188,N_4346);
and U6498 (N_6498,N_5385,N_4692);
or U6499 (N_6499,N_4735,N_4457);
and U6500 (N_6500,N_5257,N_5938);
and U6501 (N_6501,N_4585,N_4553);
and U6502 (N_6502,N_4331,N_5100);
nor U6503 (N_6503,N_5455,N_5948);
and U6504 (N_6504,N_4828,N_4419);
nand U6505 (N_6505,N_5889,N_4587);
or U6506 (N_6506,N_5164,N_5784);
nor U6507 (N_6507,N_5563,N_4733);
and U6508 (N_6508,N_5754,N_5776);
nor U6509 (N_6509,N_4969,N_5651);
and U6510 (N_6510,N_4495,N_5362);
or U6511 (N_6511,N_5691,N_4327);
and U6512 (N_6512,N_5060,N_4788);
nor U6513 (N_6513,N_5444,N_5187);
nor U6514 (N_6514,N_5637,N_5062);
nand U6515 (N_6515,N_4373,N_5381);
and U6516 (N_6516,N_4318,N_4809);
nand U6517 (N_6517,N_5710,N_4684);
and U6518 (N_6518,N_5416,N_5197);
or U6519 (N_6519,N_4220,N_4364);
or U6520 (N_6520,N_5016,N_4314);
nand U6521 (N_6521,N_4767,N_4651);
nor U6522 (N_6522,N_4652,N_5497);
or U6523 (N_6523,N_4065,N_4916);
nand U6524 (N_6524,N_5469,N_4588);
and U6525 (N_6525,N_4827,N_5423);
or U6526 (N_6526,N_5941,N_4228);
or U6527 (N_6527,N_4171,N_4221);
nor U6528 (N_6528,N_4982,N_4486);
xnor U6529 (N_6529,N_5478,N_5225);
and U6530 (N_6530,N_4661,N_4479);
and U6531 (N_6531,N_5595,N_4918);
or U6532 (N_6532,N_5960,N_4375);
nor U6533 (N_6533,N_4027,N_5129);
nand U6534 (N_6534,N_4293,N_4342);
or U6535 (N_6535,N_4928,N_5078);
or U6536 (N_6536,N_4575,N_4068);
nor U6537 (N_6537,N_5918,N_4208);
xnor U6538 (N_6538,N_5556,N_5138);
nand U6539 (N_6539,N_5896,N_4950);
or U6540 (N_6540,N_5460,N_5253);
and U6541 (N_6541,N_5620,N_4984);
nand U6542 (N_6542,N_5929,N_4844);
or U6543 (N_6543,N_5589,N_5226);
or U6544 (N_6544,N_4569,N_4520);
or U6545 (N_6545,N_4490,N_4970);
xor U6546 (N_6546,N_5508,N_5731);
nor U6547 (N_6547,N_4028,N_5638);
nor U6548 (N_6548,N_5203,N_5667);
nor U6549 (N_6549,N_4296,N_5977);
nor U6550 (N_6550,N_4851,N_5973);
or U6551 (N_6551,N_4315,N_4060);
nor U6552 (N_6552,N_5195,N_4716);
nand U6553 (N_6553,N_5527,N_4147);
xor U6554 (N_6554,N_5707,N_5849);
nor U6555 (N_6555,N_5888,N_4207);
or U6556 (N_6556,N_5570,N_5324);
and U6557 (N_6557,N_4591,N_5368);
nand U6558 (N_6558,N_4341,N_4642);
nand U6559 (N_6559,N_5872,N_4422);
and U6560 (N_6560,N_4658,N_5338);
nor U6561 (N_6561,N_5995,N_4021);
or U6562 (N_6562,N_4044,N_4404);
xor U6563 (N_6563,N_5678,N_4937);
or U6564 (N_6564,N_4412,N_4075);
or U6565 (N_6565,N_5018,N_4616);
or U6566 (N_6566,N_5724,N_4747);
nor U6567 (N_6567,N_4951,N_5512);
or U6568 (N_6568,N_5484,N_4306);
nor U6569 (N_6569,N_4627,N_5256);
nand U6570 (N_6570,N_5079,N_5734);
xnor U6571 (N_6571,N_4106,N_5228);
nand U6572 (N_6572,N_5242,N_4102);
nor U6573 (N_6573,N_4577,N_4478);
xnor U6574 (N_6574,N_4252,N_5756);
or U6575 (N_6575,N_5749,N_5947);
or U6576 (N_6576,N_5343,N_5915);
nor U6577 (N_6577,N_5471,N_4057);
nand U6578 (N_6578,N_4620,N_4993);
or U6579 (N_6579,N_4308,N_4911);
or U6580 (N_6580,N_4449,N_5588);
nor U6581 (N_6581,N_4740,N_5720);
nand U6582 (N_6582,N_5540,N_5558);
nor U6583 (N_6583,N_4955,N_5908);
or U6584 (N_6584,N_4842,N_4179);
nand U6585 (N_6585,N_4363,N_5070);
nand U6586 (N_6586,N_4513,N_5992);
nand U6587 (N_6587,N_4086,N_5118);
nor U6588 (N_6588,N_5014,N_5950);
or U6589 (N_6589,N_5488,N_4832);
or U6590 (N_6590,N_5264,N_4466);
and U6591 (N_6591,N_5625,N_5134);
nand U6592 (N_6592,N_4388,N_4182);
or U6593 (N_6593,N_4514,N_4321);
nand U6594 (N_6594,N_5298,N_5835);
and U6595 (N_6595,N_4012,N_4637);
or U6596 (N_6596,N_4328,N_4100);
and U6597 (N_6597,N_4459,N_5339);
nor U6598 (N_6598,N_5177,N_4961);
nand U6599 (N_6599,N_4164,N_4258);
nor U6600 (N_6600,N_4765,N_4227);
nand U6601 (N_6601,N_5723,N_5295);
or U6602 (N_6602,N_5811,N_5364);
and U6603 (N_6603,N_4251,N_5953);
and U6604 (N_6604,N_5673,N_5162);
nand U6605 (N_6605,N_4005,N_5645);
nor U6606 (N_6606,N_4618,N_4173);
nor U6607 (N_6607,N_5323,N_4039);
or U6608 (N_6608,N_4972,N_4083);
nand U6609 (N_6609,N_5706,N_5715);
or U6610 (N_6610,N_4234,N_5608);
or U6611 (N_6611,N_4529,N_5648);
nor U6612 (N_6612,N_5795,N_5930);
and U6613 (N_6613,N_5289,N_5387);
and U6614 (N_6614,N_5505,N_4440);
nand U6615 (N_6615,N_4059,N_4873);
and U6616 (N_6616,N_5719,N_5676);
nand U6617 (N_6617,N_4758,N_5496);
or U6618 (N_6618,N_5912,N_4260);
nor U6619 (N_6619,N_4538,N_4241);
and U6620 (N_6620,N_5083,N_5803);
nor U6621 (N_6621,N_5068,N_4437);
nand U6622 (N_6622,N_5700,N_4750);
nor U6623 (N_6623,N_4981,N_5221);
and U6624 (N_6624,N_5949,N_4668);
and U6625 (N_6625,N_4279,N_4550);
or U6626 (N_6626,N_4734,N_5026);
or U6627 (N_6627,N_4489,N_5746);
xnor U6628 (N_6628,N_4793,N_4140);
and U6629 (N_6629,N_4702,N_4666);
nand U6630 (N_6630,N_4931,N_4073);
and U6631 (N_6631,N_4565,N_4883);
nand U6632 (N_6632,N_4990,N_5249);
or U6633 (N_6633,N_4196,N_4469);
and U6634 (N_6634,N_5271,N_4622);
and U6635 (N_6635,N_5617,N_5822);
and U6636 (N_6636,N_5539,N_5946);
nand U6637 (N_6637,N_4098,N_4230);
nand U6638 (N_6638,N_4719,N_4333);
and U6639 (N_6639,N_5661,N_5154);
and U6640 (N_6640,N_4914,N_5937);
and U6641 (N_6641,N_4875,N_4909);
nor U6642 (N_6642,N_4639,N_5694);
or U6643 (N_6643,N_4187,N_5793);
or U6644 (N_6644,N_4580,N_4002);
or U6645 (N_6645,N_5935,N_5056);
nand U6646 (N_6646,N_4192,N_4202);
nor U6647 (N_6647,N_5037,N_4773);
nand U6648 (N_6648,N_5649,N_4277);
nor U6649 (N_6649,N_4090,N_4309);
nand U6650 (N_6650,N_4615,N_4011);
nand U6651 (N_6651,N_5465,N_5963);
nand U6652 (N_6652,N_4046,N_4403);
nor U6653 (N_6653,N_5571,N_4071);
nor U6654 (N_6654,N_4175,N_4125);
or U6655 (N_6655,N_4290,N_5767);
and U6656 (N_6656,N_5191,N_4829);
nand U6657 (N_6657,N_4156,N_5680);
nand U6658 (N_6658,N_4821,N_5814);
and U6659 (N_6659,N_5984,N_4974);
and U6660 (N_6660,N_4598,N_4446);
and U6661 (N_6661,N_4518,N_4871);
nand U6662 (N_6662,N_5851,N_4079);
or U6663 (N_6663,N_5581,N_5837);
xor U6664 (N_6664,N_5218,N_4739);
nor U6665 (N_6665,N_4602,N_5450);
nor U6666 (N_6666,N_5743,N_4109);
or U6667 (N_6667,N_4796,N_4311);
nand U6668 (N_6668,N_5326,N_5232);
and U6669 (N_6669,N_5438,N_5286);
nor U6670 (N_6670,N_5360,N_4244);
or U6671 (N_6671,N_4379,N_4519);
nand U6672 (N_6672,N_5903,N_5677);
nand U6673 (N_6673,N_4097,N_5330);
xnor U6674 (N_6674,N_5380,N_5209);
nand U6675 (N_6675,N_4326,N_5156);
nor U6676 (N_6676,N_5755,N_5535);
xnor U6677 (N_6677,N_4215,N_4456);
and U6678 (N_6678,N_4869,N_4685);
nand U6679 (N_6679,N_5569,N_4267);
nand U6680 (N_6680,N_5274,N_4554);
nand U6681 (N_6681,N_4522,N_5926);
and U6682 (N_6682,N_4624,N_5548);
and U6683 (N_6683,N_4959,N_5055);
or U6684 (N_6684,N_4322,N_5862);
and U6685 (N_6685,N_4144,N_4562);
and U6686 (N_6686,N_4087,N_4014);
or U6687 (N_6687,N_4377,N_5462);
and U6688 (N_6688,N_4803,N_5867);
and U6689 (N_6689,N_5237,N_4724);
nor U6690 (N_6690,N_5047,N_5113);
or U6691 (N_6691,N_5117,N_5611);
nand U6692 (N_6692,N_4047,N_5727);
or U6693 (N_6693,N_4093,N_5029);
or U6694 (N_6694,N_4369,N_4772);
xor U6695 (N_6695,N_4774,N_5111);
nor U6696 (N_6696,N_4091,N_5308);
nor U6697 (N_6697,N_4748,N_4204);
or U6698 (N_6698,N_5022,N_4329);
nor U6699 (N_6699,N_5575,N_5796);
nand U6700 (N_6700,N_5214,N_5347);
xnor U6701 (N_6701,N_4944,N_4126);
nand U6702 (N_6702,N_4533,N_5580);
nand U6703 (N_6703,N_4889,N_4901);
or U6704 (N_6704,N_4686,N_4142);
xor U6705 (N_6705,N_5268,N_5366);
xor U6706 (N_6706,N_5023,N_5376);
or U6707 (N_6707,N_5259,N_4825);
nor U6708 (N_6708,N_4291,N_5227);
nand U6709 (N_6709,N_4907,N_5738);
xnor U6710 (N_6710,N_5109,N_4511);
xor U6711 (N_6711,N_4935,N_4833);
or U6712 (N_6712,N_4020,N_4337);
and U6713 (N_6713,N_4040,N_5390);
nor U6714 (N_6714,N_5063,N_4128);
or U6715 (N_6715,N_5310,N_5206);
nand U6716 (N_6716,N_5433,N_5378);
or U6717 (N_6717,N_5800,N_4922);
nor U6718 (N_6718,N_4366,N_5812);
nor U6719 (N_6719,N_5201,N_4798);
nor U6720 (N_6720,N_5831,N_4473);
nor U6721 (N_6721,N_5017,N_5999);
and U6722 (N_6722,N_4274,N_5008);
or U6723 (N_6723,N_4504,N_5658);
and U6724 (N_6724,N_5576,N_5020);
and U6725 (N_6725,N_4262,N_4222);
nor U6726 (N_6726,N_5141,N_5653);
nor U6727 (N_6727,N_5717,N_4295);
and U6728 (N_6728,N_5654,N_5213);
nor U6729 (N_6729,N_5659,N_4353);
nand U6730 (N_6730,N_4625,N_4143);
nor U6731 (N_6731,N_5255,N_4313);
or U6732 (N_6732,N_4118,N_5250);
nand U6733 (N_6733,N_5561,N_5004);
or U6734 (N_6734,N_4675,N_4170);
nor U6735 (N_6735,N_4483,N_4688);
nand U6736 (N_6736,N_4966,N_5267);
or U6737 (N_6737,N_5105,N_5877);
or U6738 (N_6738,N_5345,N_4703);
nor U6739 (N_6739,N_5006,N_5344);
nor U6740 (N_6740,N_5074,N_5845);
nand U6741 (N_6741,N_5320,N_4061);
or U6742 (N_6742,N_5353,N_4607);
or U6743 (N_6743,N_4902,N_5097);
nand U6744 (N_6744,N_5476,N_4078);
nand U6745 (N_6745,N_4654,N_4302);
nand U6746 (N_6746,N_5094,N_4232);
and U6747 (N_6747,N_4586,N_5244);
nor U6748 (N_6748,N_5434,N_4558);
and U6749 (N_6749,N_5337,N_4468);
or U6750 (N_6750,N_4542,N_5358);
or U6751 (N_6751,N_4152,N_5470);
nor U6752 (N_6752,N_4777,N_4427);
nor U6753 (N_6753,N_4135,N_5902);
nand U6754 (N_6754,N_4877,N_5826);
and U6755 (N_6755,N_4892,N_5379);
nor U6756 (N_6756,N_4139,N_4994);
nor U6757 (N_6757,N_4276,N_4048);
or U6758 (N_6758,N_4491,N_5142);
nor U6759 (N_6759,N_5369,N_4160);
or U6760 (N_6760,N_5120,N_4458);
or U6761 (N_6761,N_5688,N_4628);
or U6762 (N_6762,N_5294,N_4840);
or U6763 (N_6763,N_4269,N_4034);
nor U6764 (N_6764,N_4177,N_5475);
xnor U6765 (N_6765,N_5397,N_5686);
nand U6766 (N_6766,N_5914,N_4573);
nor U6767 (N_6767,N_5833,N_5296);
nor U6768 (N_6768,N_5966,N_4516);
and U6769 (N_6769,N_5858,N_5149);
xor U6770 (N_6770,N_4415,N_4753);
and U6771 (N_6771,N_4420,N_5603);
nor U6772 (N_6772,N_5307,N_4351);
or U6773 (N_6773,N_4358,N_5349);
nor U6774 (N_6774,N_5622,N_4435);
and U6775 (N_6775,N_5241,N_5983);
or U6776 (N_6776,N_4502,N_5393);
nor U6777 (N_6777,N_4808,N_5044);
and U6778 (N_6778,N_5043,N_4017);
nand U6779 (N_6779,N_5829,N_5190);
and U6780 (N_6780,N_4163,N_4669);
or U6781 (N_6781,N_5898,N_5391);
nand U6782 (N_6782,N_4589,N_4971);
nand U6783 (N_6783,N_5148,N_4101);
and U6784 (N_6784,N_4095,N_4670);
nand U6785 (N_6785,N_5153,N_5179);
or U6786 (N_6786,N_4382,N_5112);
nand U6787 (N_6787,N_4957,N_5169);
or U6788 (N_6788,N_5518,N_5204);
nor U6789 (N_6789,N_5951,N_5167);
and U6790 (N_6790,N_5559,N_5591);
nor U6791 (N_6791,N_5058,N_4726);
xnor U6792 (N_6792,N_5429,N_5774);
and U6793 (N_6793,N_4864,N_4789);
nor U6794 (N_6794,N_5600,N_4213);
and U6795 (N_6795,N_5336,N_5758);
or U6796 (N_6796,N_4247,N_5306);
or U6797 (N_6797,N_4992,N_5231);
and U6798 (N_6798,N_4995,N_5718);
nor U6799 (N_6799,N_4111,N_5768);
or U6800 (N_6800,N_4089,N_4356);
nor U6801 (N_6801,N_4409,N_5325);
nor U6802 (N_6802,N_4448,N_5098);
nand U6803 (N_6803,N_5371,N_5848);
nand U6804 (N_6804,N_4107,N_5972);
or U6805 (N_6805,N_5010,N_4831);
nor U6806 (N_6806,N_5284,N_5408);
nor U6807 (N_6807,N_4181,N_5881);
and U6808 (N_6808,N_4148,N_5202);
nand U6809 (N_6809,N_5002,N_4926);
and U6810 (N_6810,N_5081,N_4605);
nand U6811 (N_6811,N_4534,N_4818);
and U6812 (N_6812,N_4723,N_5632);
and U6813 (N_6813,N_4759,N_5076);
nor U6814 (N_6814,N_5263,N_5744);
nand U6815 (N_6815,N_4016,N_4715);
or U6816 (N_6816,N_4413,N_4523);
nand U6817 (N_6817,N_4161,N_4650);
and U6818 (N_6818,N_4273,N_4720);
nand U6819 (N_6819,N_4385,N_4895);
nor U6820 (N_6820,N_4510,N_5797);
or U6821 (N_6821,N_4940,N_5327);
or U6822 (N_6822,N_4389,N_4657);
nor U6823 (N_6823,N_4004,N_4320);
nor U6824 (N_6824,N_4807,N_4850);
nor U6825 (N_6825,N_5477,N_4246);
nand U6826 (N_6826,N_5662,N_5874);
and U6827 (N_6827,N_4465,N_4606);
nor U6828 (N_6828,N_4361,N_4999);
or U6829 (N_6829,N_5692,N_4858);
or U6830 (N_6830,N_5643,N_5524);
nand U6831 (N_6831,N_5175,N_5924);
nand U6832 (N_6832,N_5281,N_5498);
and U6833 (N_6833,N_4190,N_4924);
nand U6834 (N_6834,N_5905,N_4975);
nor U6835 (N_6835,N_4905,N_4055);
nand U6836 (N_6836,N_4270,N_5492);
and U6837 (N_6837,N_4292,N_4980);
xor U6838 (N_6838,N_4915,N_4694);
nor U6839 (N_6839,N_4136,N_4416);
and U6840 (N_6840,N_5623,N_5739);
nor U6841 (N_6841,N_5350,N_4581);
or U6842 (N_6842,N_4545,N_4229);
nor U6843 (N_6843,N_5319,N_5927);
and U6844 (N_6844,N_4368,N_5452);
nand U6845 (N_6845,N_4265,N_5552);
or U6846 (N_6846,N_4395,N_4584);
and U6847 (N_6847,N_5309,N_5725);
xor U6848 (N_6848,N_5830,N_5181);
nand U6849 (N_6849,N_4604,N_4001);
nor U6850 (N_6850,N_5644,N_5311);
and U6851 (N_6851,N_5847,N_5782);
nor U6852 (N_6852,N_5913,N_4626);
and U6853 (N_6853,N_5997,N_5107);
and U6854 (N_6854,N_5791,N_5705);
nor U6855 (N_6855,N_4203,N_5130);
nor U6856 (N_6856,N_4010,N_5752);
nand U6857 (N_6857,N_4574,N_5051);
nor U6858 (N_6858,N_5741,N_5566);
nor U6859 (N_6859,N_5139,N_5628);
nor U6860 (N_6860,N_4643,N_5009);
and U6861 (N_6861,N_4112,N_5778);
or U6862 (N_6862,N_4839,N_4854);
nor U6863 (N_6863,N_4714,N_5557);
and U6864 (N_6864,N_4599,N_5501);
nand U6865 (N_6865,N_4299,N_5991);
or U6866 (N_6866,N_5553,N_4515);
nand U6867 (N_6867,N_4859,N_4325);
nor U6868 (N_6868,N_5854,N_5466);
and U6869 (N_6869,N_4946,N_4933);
nand U6870 (N_6870,N_4289,N_5825);
nand U6871 (N_6871,N_5291,N_5312);
nor U6872 (N_6872,N_5657,N_5448);
or U6873 (N_6873,N_5664,N_4434);
or U6874 (N_6874,N_4099,N_5987);
nor U6875 (N_6875,N_5467,N_5853);
and U6876 (N_6876,N_4225,N_4603);
nand U6877 (N_6877,N_4428,N_5549);
and U6878 (N_6878,N_5907,N_5828);
nand U6879 (N_6879,N_4611,N_5223);
or U6880 (N_6880,N_4317,N_4033);
and U6881 (N_6881,N_5451,N_4559);
nor U6882 (N_6882,N_4884,N_4711);
and U6883 (N_6883,N_4834,N_4812);
or U6884 (N_6884,N_5771,N_5885);
or U6885 (N_6885,N_4674,N_4568);
and U6886 (N_6886,N_5695,N_4973);
nand U6887 (N_6887,N_5340,N_5616);
and U6888 (N_6888,N_4174,N_4648);
nor U6889 (N_6889,N_4480,N_5564);
nand U6890 (N_6890,N_5304,N_4018);
nor U6891 (N_6891,N_4330,N_4517);
nor U6892 (N_6892,N_4417,N_4623);
nor U6893 (N_6893,N_4600,N_5392);
and U6894 (N_6894,N_5300,N_4893);
or U6895 (N_6895,N_5359,N_5482);
nand U6896 (N_6896,N_4962,N_5974);
and U6897 (N_6897,N_5764,N_5278);
or U6898 (N_6898,N_5955,N_4897);
nand U6899 (N_6899,N_5059,N_5506);
nand U6900 (N_6900,N_4725,N_5119);
or U6901 (N_6901,N_5607,N_4560);
nor U6902 (N_6902,N_5805,N_5943);
or U6903 (N_6903,N_5057,N_5514);
or U6904 (N_6904,N_4621,N_4965);
nand U6905 (N_6905,N_5634,N_4862);
or U6906 (N_6906,N_5091,N_5108);
nand U6907 (N_6907,N_5375,N_5630);
and U6908 (N_6908,N_5114,N_4609);
and U6909 (N_6909,N_5061,N_5042);
nand U6910 (N_6910,N_4784,N_4792);
or U6911 (N_6911,N_5238,N_4736);
nand U6912 (N_6912,N_4050,N_5155);
nor U6913 (N_6913,N_4531,N_4872);
nor U6914 (N_6914,N_4080,N_4755);
and U6915 (N_6915,N_5663,N_5483);
or U6916 (N_6916,N_5199,N_4362);
nor U6917 (N_6917,N_5474,N_4823);
or U6918 (N_6918,N_5560,N_4352);
nor U6919 (N_6919,N_5932,N_5592);
xor U6920 (N_6920,N_5282,N_4548);
nor U6921 (N_6921,N_4817,N_4442);
nor U6922 (N_6922,N_4707,N_5745);
and U6923 (N_6923,N_4756,N_5631);
nand U6924 (N_6924,N_4878,N_5809);
and U6925 (N_6925,N_4848,N_5135);
nand U6926 (N_6926,N_4149,N_4800);
and U6927 (N_6927,N_5917,N_4906);
nand U6928 (N_6928,N_4749,N_4646);
nor U6929 (N_6929,N_5523,N_5920);
or U6930 (N_6930,N_4294,N_4113);
and U6931 (N_6931,N_4830,N_5751);
or U6932 (N_6932,N_5101,N_5313);
or U6933 (N_6933,N_4978,N_4867);
nand U6934 (N_6934,N_4031,N_5824);
nor U6935 (N_6935,N_4450,N_5064);
nor U6936 (N_6936,N_5041,N_4768);
or U6937 (N_6937,N_4332,N_4597);
nand U6938 (N_6938,N_5980,N_5342);
or U6939 (N_6939,N_4084,N_4432);
and U6940 (N_6940,N_4045,N_4347);
and U6941 (N_6941,N_5511,N_4976);
and U6942 (N_6942,N_4355,N_4680);
nand U6943 (N_6943,N_5968,N_5565);
or U6944 (N_6944,N_4235,N_5789);
nor U6945 (N_6945,N_4761,N_5766);
nand U6946 (N_6946,N_4636,N_4503);
nor U6947 (N_6947,N_4239,N_5785);
nor U6948 (N_6948,N_4343,N_4240);
nand U6949 (N_6949,N_5516,N_4166);
and U6950 (N_6950,N_5879,N_4319);
and U6951 (N_6951,N_5820,N_5389);
and U6952 (N_6952,N_4051,N_4751);
nor U6953 (N_6953,N_5554,N_4400);
and U6954 (N_6954,N_4076,N_5405);
nor U6955 (N_6955,N_4682,N_5722);
nor U6956 (N_6956,N_5431,N_5011);
and U6957 (N_6957,N_4231,N_5328);
nand U6958 (N_6958,N_4104,N_4776);
or U6959 (N_6959,N_4647,N_5577);
and U6960 (N_6960,N_4986,N_5005);
and U6961 (N_6961,N_5979,N_5373);
nand U6962 (N_6962,N_4487,N_4941);
or U6963 (N_6963,N_5128,N_4405);
xor U6964 (N_6964,N_4508,N_4540);
or U6965 (N_6965,N_5456,N_4806);
nor U6966 (N_6966,N_4989,N_4526);
or U6967 (N_6967,N_4077,N_5684);
nand U6968 (N_6968,N_4910,N_5585);
or U6969 (N_6969,N_5012,N_5445);
or U6970 (N_6970,N_5895,N_5001);
and U6971 (N_6971,N_4882,N_4820);
nor U6972 (N_6972,N_4471,N_4344);
and U6973 (N_6973,N_5964,N_4532);
or U6974 (N_6974,N_5928,N_4699);
nand U6975 (N_6975,N_4121,N_5761);
or U6976 (N_6976,N_5443,N_4236);
nor U6977 (N_6977,N_5893,N_5144);
or U6978 (N_6978,N_4474,N_5641);
or U6979 (N_6979,N_5335,N_4023);
nor U6980 (N_6980,N_5742,N_5517);
nor U6981 (N_6981,N_4592,N_5642);
nor U6982 (N_6982,N_5834,N_5208);
and U6983 (N_6983,N_5441,N_5729);
nor U6984 (N_6984,N_5189,N_4157);
or U6985 (N_6985,N_5737,N_4454);
nand U6986 (N_6986,N_4032,N_4248);
nor U6987 (N_6987,N_5502,N_5499);
or U6988 (N_6988,N_5639,N_5211);
or U6989 (N_6989,N_5880,N_5240);
nor U6990 (N_6990,N_5406,N_5836);
nand U6991 (N_6991,N_4278,N_4138);
and U6992 (N_6992,N_5147,N_5900);
and U6993 (N_6993,N_4868,N_5346);
or U6994 (N_6994,N_5015,N_5383);
or U6995 (N_6995,N_4110,N_4378);
nor U6996 (N_6996,N_5952,N_5087);
nor U6997 (N_6997,N_5454,N_5541);
or U6998 (N_6998,N_5370,N_5728);
or U6999 (N_6999,N_4350,N_5602);
or U7000 (N_7000,N_5666,N_5429);
or U7001 (N_7001,N_5732,N_4489);
nor U7002 (N_7002,N_5228,N_4750);
and U7003 (N_7003,N_4703,N_5457);
nand U7004 (N_7004,N_5833,N_5194);
nor U7005 (N_7005,N_4533,N_4592);
nand U7006 (N_7006,N_5026,N_4158);
nand U7007 (N_7007,N_5028,N_4803);
or U7008 (N_7008,N_4686,N_5440);
nor U7009 (N_7009,N_4006,N_5512);
nor U7010 (N_7010,N_4605,N_4535);
nand U7011 (N_7011,N_5139,N_5980);
or U7012 (N_7012,N_5936,N_5073);
or U7013 (N_7013,N_5914,N_5840);
xor U7014 (N_7014,N_4225,N_5328);
nor U7015 (N_7015,N_4742,N_5774);
nand U7016 (N_7016,N_4259,N_4503);
or U7017 (N_7017,N_4321,N_5067);
or U7018 (N_7018,N_4584,N_4413);
and U7019 (N_7019,N_4339,N_5681);
nand U7020 (N_7020,N_5604,N_4750);
and U7021 (N_7021,N_5819,N_4962);
nor U7022 (N_7022,N_4348,N_5416);
or U7023 (N_7023,N_5369,N_5864);
nor U7024 (N_7024,N_4537,N_5821);
or U7025 (N_7025,N_5210,N_4548);
and U7026 (N_7026,N_5335,N_5771);
or U7027 (N_7027,N_5509,N_4929);
nor U7028 (N_7028,N_5007,N_5944);
or U7029 (N_7029,N_4957,N_5777);
nor U7030 (N_7030,N_4467,N_4128);
or U7031 (N_7031,N_5556,N_5367);
or U7032 (N_7032,N_5115,N_5296);
or U7033 (N_7033,N_5350,N_4804);
nand U7034 (N_7034,N_4504,N_5642);
or U7035 (N_7035,N_5451,N_5949);
or U7036 (N_7036,N_4032,N_4393);
or U7037 (N_7037,N_4806,N_4782);
nand U7038 (N_7038,N_5917,N_4817);
or U7039 (N_7039,N_5217,N_4214);
nor U7040 (N_7040,N_4199,N_5894);
nor U7041 (N_7041,N_4927,N_4811);
nand U7042 (N_7042,N_4009,N_4351);
or U7043 (N_7043,N_4173,N_5185);
nor U7044 (N_7044,N_5149,N_5194);
nor U7045 (N_7045,N_5603,N_5736);
or U7046 (N_7046,N_4533,N_5195);
or U7047 (N_7047,N_5487,N_4608);
or U7048 (N_7048,N_5316,N_5122);
and U7049 (N_7049,N_5547,N_5133);
nand U7050 (N_7050,N_4311,N_5491);
nor U7051 (N_7051,N_5079,N_5370);
and U7052 (N_7052,N_4626,N_4345);
and U7053 (N_7053,N_5519,N_4334);
and U7054 (N_7054,N_5376,N_4195);
or U7055 (N_7055,N_4662,N_4887);
nand U7056 (N_7056,N_5073,N_4314);
nand U7057 (N_7057,N_5137,N_5406);
or U7058 (N_7058,N_4224,N_4280);
nand U7059 (N_7059,N_4531,N_4711);
and U7060 (N_7060,N_5393,N_4283);
and U7061 (N_7061,N_4865,N_5037);
nor U7062 (N_7062,N_5797,N_4372);
nand U7063 (N_7063,N_5881,N_5808);
or U7064 (N_7064,N_4669,N_4330);
and U7065 (N_7065,N_5668,N_5494);
nor U7066 (N_7066,N_5926,N_4279);
nor U7067 (N_7067,N_4414,N_4239);
and U7068 (N_7068,N_4882,N_4346);
nand U7069 (N_7069,N_4474,N_4891);
nand U7070 (N_7070,N_5943,N_5575);
nand U7071 (N_7071,N_5140,N_4435);
nand U7072 (N_7072,N_4808,N_5639);
nor U7073 (N_7073,N_4452,N_4130);
and U7074 (N_7074,N_5243,N_5575);
and U7075 (N_7075,N_5377,N_5011);
and U7076 (N_7076,N_4460,N_4808);
nor U7077 (N_7077,N_4212,N_5334);
nor U7078 (N_7078,N_5793,N_4228);
or U7079 (N_7079,N_4568,N_4681);
and U7080 (N_7080,N_5788,N_5740);
nand U7081 (N_7081,N_5678,N_4356);
nand U7082 (N_7082,N_4521,N_5000);
nor U7083 (N_7083,N_5260,N_5642);
or U7084 (N_7084,N_4442,N_4795);
or U7085 (N_7085,N_4028,N_4683);
nand U7086 (N_7086,N_5111,N_5481);
nor U7087 (N_7087,N_5346,N_5945);
nor U7088 (N_7088,N_5861,N_5583);
and U7089 (N_7089,N_5121,N_4130);
or U7090 (N_7090,N_5534,N_5137);
or U7091 (N_7091,N_4831,N_5506);
and U7092 (N_7092,N_4830,N_4356);
or U7093 (N_7093,N_5430,N_4353);
or U7094 (N_7094,N_4141,N_5791);
nor U7095 (N_7095,N_5086,N_4963);
or U7096 (N_7096,N_4035,N_4212);
and U7097 (N_7097,N_5842,N_5266);
or U7098 (N_7098,N_4856,N_4117);
nand U7099 (N_7099,N_4669,N_4181);
xnor U7100 (N_7100,N_4784,N_5217);
or U7101 (N_7101,N_5158,N_5990);
nand U7102 (N_7102,N_4015,N_5612);
and U7103 (N_7103,N_5763,N_4974);
nand U7104 (N_7104,N_4894,N_4976);
and U7105 (N_7105,N_5308,N_4550);
nand U7106 (N_7106,N_5520,N_5693);
and U7107 (N_7107,N_4075,N_4982);
nor U7108 (N_7108,N_4074,N_5696);
xor U7109 (N_7109,N_4493,N_5215);
nor U7110 (N_7110,N_4482,N_4442);
nor U7111 (N_7111,N_4613,N_5682);
or U7112 (N_7112,N_4991,N_5392);
and U7113 (N_7113,N_4682,N_5331);
nor U7114 (N_7114,N_4896,N_4008);
and U7115 (N_7115,N_4344,N_5202);
and U7116 (N_7116,N_5203,N_4845);
or U7117 (N_7117,N_5080,N_5582);
nor U7118 (N_7118,N_5134,N_5459);
nand U7119 (N_7119,N_5433,N_5692);
nor U7120 (N_7120,N_4142,N_4159);
and U7121 (N_7121,N_4309,N_4467);
and U7122 (N_7122,N_4838,N_4240);
and U7123 (N_7123,N_5992,N_5555);
and U7124 (N_7124,N_4036,N_4300);
nand U7125 (N_7125,N_5593,N_4299);
and U7126 (N_7126,N_4942,N_4890);
nand U7127 (N_7127,N_5043,N_5297);
nand U7128 (N_7128,N_5681,N_5257);
nor U7129 (N_7129,N_4508,N_5773);
and U7130 (N_7130,N_4571,N_4854);
nor U7131 (N_7131,N_5198,N_4039);
and U7132 (N_7132,N_4368,N_4625);
and U7133 (N_7133,N_5890,N_5794);
nor U7134 (N_7134,N_4994,N_5351);
nor U7135 (N_7135,N_4096,N_5966);
or U7136 (N_7136,N_4177,N_5194);
nor U7137 (N_7137,N_4918,N_4607);
and U7138 (N_7138,N_4668,N_4730);
nand U7139 (N_7139,N_4933,N_5899);
nand U7140 (N_7140,N_5748,N_5180);
and U7141 (N_7141,N_5651,N_4076);
and U7142 (N_7142,N_5097,N_5354);
or U7143 (N_7143,N_5721,N_5847);
nand U7144 (N_7144,N_4775,N_5493);
nand U7145 (N_7145,N_4799,N_5115);
and U7146 (N_7146,N_5088,N_4938);
nor U7147 (N_7147,N_5040,N_4342);
or U7148 (N_7148,N_5109,N_4877);
nor U7149 (N_7149,N_4176,N_4325);
nand U7150 (N_7150,N_4841,N_4421);
nand U7151 (N_7151,N_4008,N_4417);
nand U7152 (N_7152,N_5534,N_4992);
and U7153 (N_7153,N_5763,N_4474);
nand U7154 (N_7154,N_4046,N_4885);
and U7155 (N_7155,N_5620,N_5406);
or U7156 (N_7156,N_4922,N_4501);
nor U7157 (N_7157,N_5674,N_4786);
and U7158 (N_7158,N_5929,N_5183);
nand U7159 (N_7159,N_4758,N_5838);
nand U7160 (N_7160,N_4312,N_5379);
nand U7161 (N_7161,N_5298,N_4790);
or U7162 (N_7162,N_5212,N_5949);
nor U7163 (N_7163,N_5281,N_4370);
nor U7164 (N_7164,N_4182,N_4198);
nand U7165 (N_7165,N_4167,N_5338);
nor U7166 (N_7166,N_5691,N_5727);
or U7167 (N_7167,N_4954,N_5083);
and U7168 (N_7168,N_4316,N_5908);
and U7169 (N_7169,N_5282,N_5377);
nand U7170 (N_7170,N_5224,N_4275);
nor U7171 (N_7171,N_5893,N_4020);
nand U7172 (N_7172,N_5577,N_5004);
and U7173 (N_7173,N_4293,N_4638);
and U7174 (N_7174,N_4679,N_4735);
nand U7175 (N_7175,N_4738,N_5688);
nor U7176 (N_7176,N_4348,N_5516);
and U7177 (N_7177,N_4459,N_4639);
or U7178 (N_7178,N_5843,N_4107);
and U7179 (N_7179,N_4240,N_4564);
nand U7180 (N_7180,N_5615,N_4965);
or U7181 (N_7181,N_4413,N_4927);
nand U7182 (N_7182,N_4106,N_5042);
nand U7183 (N_7183,N_4563,N_5880);
and U7184 (N_7184,N_5512,N_5026);
nand U7185 (N_7185,N_5617,N_4942);
and U7186 (N_7186,N_5106,N_4946);
and U7187 (N_7187,N_5976,N_5987);
nor U7188 (N_7188,N_4097,N_5204);
or U7189 (N_7189,N_4954,N_5918);
or U7190 (N_7190,N_4056,N_4934);
or U7191 (N_7191,N_4383,N_5475);
and U7192 (N_7192,N_4082,N_4531);
or U7193 (N_7193,N_5095,N_5452);
and U7194 (N_7194,N_4977,N_4900);
nor U7195 (N_7195,N_5765,N_5718);
nor U7196 (N_7196,N_5364,N_4603);
nor U7197 (N_7197,N_5883,N_5599);
nand U7198 (N_7198,N_5579,N_5286);
and U7199 (N_7199,N_5415,N_5861);
nand U7200 (N_7200,N_4634,N_5180);
and U7201 (N_7201,N_5001,N_5279);
and U7202 (N_7202,N_4147,N_5370);
or U7203 (N_7203,N_5842,N_4235);
nor U7204 (N_7204,N_5601,N_4724);
nor U7205 (N_7205,N_5708,N_4537);
and U7206 (N_7206,N_5564,N_4435);
nor U7207 (N_7207,N_4330,N_5866);
and U7208 (N_7208,N_4668,N_4050);
and U7209 (N_7209,N_5459,N_5085);
and U7210 (N_7210,N_4948,N_5378);
or U7211 (N_7211,N_5490,N_5138);
xnor U7212 (N_7212,N_4498,N_4278);
and U7213 (N_7213,N_4899,N_4460);
and U7214 (N_7214,N_5702,N_5844);
nor U7215 (N_7215,N_4004,N_4695);
and U7216 (N_7216,N_5196,N_4445);
and U7217 (N_7217,N_5975,N_5651);
nor U7218 (N_7218,N_4801,N_5973);
nor U7219 (N_7219,N_5552,N_5950);
nand U7220 (N_7220,N_4349,N_4749);
xor U7221 (N_7221,N_4858,N_4110);
nor U7222 (N_7222,N_4685,N_4662);
and U7223 (N_7223,N_5537,N_5244);
or U7224 (N_7224,N_5927,N_5217);
nor U7225 (N_7225,N_4954,N_5041);
xnor U7226 (N_7226,N_4491,N_5992);
and U7227 (N_7227,N_4884,N_5491);
nand U7228 (N_7228,N_5482,N_5581);
nand U7229 (N_7229,N_4799,N_4838);
nand U7230 (N_7230,N_5216,N_4718);
and U7231 (N_7231,N_4031,N_5230);
nand U7232 (N_7232,N_4957,N_5601);
nor U7233 (N_7233,N_4731,N_5436);
and U7234 (N_7234,N_5272,N_4490);
and U7235 (N_7235,N_5174,N_4346);
nor U7236 (N_7236,N_5834,N_4151);
nand U7237 (N_7237,N_5767,N_5526);
and U7238 (N_7238,N_4131,N_5952);
nand U7239 (N_7239,N_4609,N_5423);
nand U7240 (N_7240,N_5476,N_5951);
nor U7241 (N_7241,N_5901,N_4933);
or U7242 (N_7242,N_4447,N_4319);
nand U7243 (N_7243,N_4991,N_5052);
or U7244 (N_7244,N_5851,N_5326);
or U7245 (N_7245,N_4999,N_4088);
and U7246 (N_7246,N_5995,N_4313);
nor U7247 (N_7247,N_5049,N_4884);
nor U7248 (N_7248,N_5033,N_5369);
and U7249 (N_7249,N_4418,N_5043);
or U7250 (N_7250,N_4618,N_5130);
or U7251 (N_7251,N_5919,N_5414);
nor U7252 (N_7252,N_4158,N_4187);
and U7253 (N_7253,N_5050,N_5727);
or U7254 (N_7254,N_5306,N_4738);
or U7255 (N_7255,N_4048,N_4039);
or U7256 (N_7256,N_4025,N_5415);
nand U7257 (N_7257,N_4402,N_4201);
and U7258 (N_7258,N_4607,N_5903);
and U7259 (N_7259,N_4376,N_5367);
nor U7260 (N_7260,N_5520,N_4809);
nand U7261 (N_7261,N_5057,N_5676);
or U7262 (N_7262,N_4473,N_5783);
nand U7263 (N_7263,N_4361,N_4476);
or U7264 (N_7264,N_4911,N_4064);
or U7265 (N_7265,N_4621,N_4084);
nor U7266 (N_7266,N_5059,N_5089);
and U7267 (N_7267,N_5573,N_5018);
and U7268 (N_7268,N_4162,N_5822);
or U7269 (N_7269,N_4563,N_5472);
nor U7270 (N_7270,N_5270,N_5657);
nor U7271 (N_7271,N_4419,N_4352);
or U7272 (N_7272,N_5391,N_4693);
or U7273 (N_7273,N_4223,N_5720);
nand U7274 (N_7274,N_5593,N_5310);
nor U7275 (N_7275,N_5287,N_4870);
or U7276 (N_7276,N_5667,N_5503);
nand U7277 (N_7277,N_5872,N_5776);
or U7278 (N_7278,N_4803,N_5436);
nand U7279 (N_7279,N_5667,N_5551);
nor U7280 (N_7280,N_5628,N_4954);
or U7281 (N_7281,N_4606,N_5258);
nor U7282 (N_7282,N_4293,N_4333);
and U7283 (N_7283,N_4962,N_5658);
and U7284 (N_7284,N_4205,N_4258);
or U7285 (N_7285,N_5914,N_4825);
or U7286 (N_7286,N_5857,N_4364);
or U7287 (N_7287,N_5627,N_5440);
nand U7288 (N_7288,N_4026,N_4043);
nand U7289 (N_7289,N_5275,N_5854);
or U7290 (N_7290,N_4846,N_4386);
and U7291 (N_7291,N_5694,N_4873);
nor U7292 (N_7292,N_4717,N_4753);
and U7293 (N_7293,N_5471,N_4023);
nand U7294 (N_7294,N_5719,N_4449);
or U7295 (N_7295,N_4708,N_5824);
or U7296 (N_7296,N_5618,N_4508);
nor U7297 (N_7297,N_5723,N_4903);
nor U7298 (N_7298,N_4894,N_4077);
nor U7299 (N_7299,N_4519,N_5316);
or U7300 (N_7300,N_5150,N_4570);
nand U7301 (N_7301,N_5896,N_5405);
or U7302 (N_7302,N_4240,N_4154);
nor U7303 (N_7303,N_4899,N_5772);
and U7304 (N_7304,N_5189,N_5900);
nor U7305 (N_7305,N_5349,N_5643);
or U7306 (N_7306,N_4550,N_4995);
or U7307 (N_7307,N_5600,N_5872);
and U7308 (N_7308,N_4580,N_5760);
nor U7309 (N_7309,N_5559,N_4348);
nor U7310 (N_7310,N_5289,N_5026);
or U7311 (N_7311,N_4086,N_4194);
nor U7312 (N_7312,N_5292,N_5224);
nand U7313 (N_7313,N_5244,N_5989);
and U7314 (N_7314,N_5575,N_5955);
and U7315 (N_7315,N_5415,N_4622);
and U7316 (N_7316,N_5151,N_4533);
and U7317 (N_7317,N_4113,N_4794);
and U7318 (N_7318,N_5918,N_5768);
nand U7319 (N_7319,N_5073,N_4104);
or U7320 (N_7320,N_4986,N_4406);
or U7321 (N_7321,N_5618,N_4743);
and U7322 (N_7322,N_5784,N_4463);
nor U7323 (N_7323,N_5152,N_5251);
and U7324 (N_7324,N_5484,N_4613);
nor U7325 (N_7325,N_4088,N_5844);
nand U7326 (N_7326,N_5408,N_5672);
or U7327 (N_7327,N_5919,N_4150);
or U7328 (N_7328,N_4130,N_5759);
or U7329 (N_7329,N_5277,N_4125);
or U7330 (N_7330,N_5030,N_4157);
nor U7331 (N_7331,N_4319,N_5937);
nor U7332 (N_7332,N_4420,N_5215);
and U7333 (N_7333,N_5504,N_5391);
and U7334 (N_7334,N_4120,N_4103);
nor U7335 (N_7335,N_5738,N_4722);
nor U7336 (N_7336,N_4999,N_5928);
or U7337 (N_7337,N_4446,N_5752);
nand U7338 (N_7338,N_4694,N_4578);
nor U7339 (N_7339,N_5699,N_4129);
nand U7340 (N_7340,N_4106,N_5133);
or U7341 (N_7341,N_5747,N_4965);
and U7342 (N_7342,N_4582,N_5048);
or U7343 (N_7343,N_4887,N_4813);
or U7344 (N_7344,N_5481,N_4129);
xnor U7345 (N_7345,N_5229,N_5002);
or U7346 (N_7346,N_4203,N_5331);
and U7347 (N_7347,N_4089,N_5186);
or U7348 (N_7348,N_4614,N_4852);
xnor U7349 (N_7349,N_5327,N_4734);
and U7350 (N_7350,N_5015,N_5593);
nor U7351 (N_7351,N_4959,N_4356);
nor U7352 (N_7352,N_5776,N_5716);
nand U7353 (N_7353,N_4341,N_4148);
nand U7354 (N_7354,N_5733,N_5785);
and U7355 (N_7355,N_5138,N_4270);
nor U7356 (N_7356,N_4273,N_4968);
nor U7357 (N_7357,N_4593,N_4732);
nand U7358 (N_7358,N_5332,N_5782);
nor U7359 (N_7359,N_5905,N_5665);
and U7360 (N_7360,N_5133,N_4418);
or U7361 (N_7361,N_4923,N_4954);
nand U7362 (N_7362,N_5194,N_5307);
and U7363 (N_7363,N_5829,N_4021);
xnor U7364 (N_7364,N_4226,N_5711);
nand U7365 (N_7365,N_5179,N_4309);
nand U7366 (N_7366,N_5910,N_5471);
nor U7367 (N_7367,N_5141,N_5702);
nor U7368 (N_7368,N_4931,N_5139);
and U7369 (N_7369,N_5948,N_4597);
xnor U7370 (N_7370,N_5146,N_5736);
nand U7371 (N_7371,N_4365,N_5288);
nand U7372 (N_7372,N_5704,N_5087);
and U7373 (N_7373,N_4985,N_4254);
or U7374 (N_7374,N_4762,N_5084);
or U7375 (N_7375,N_5061,N_5215);
nand U7376 (N_7376,N_4005,N_5615);
nand U7377 (N_7377,N_5325,N_4999);
nand U7378 (N_7378,N_5170,N_5383);
or U7379 (N_7379,N_5695,N_5162);
nor U7380 (N_7380,N_5976,N_4709);
nand U7381 (N_7381,N_5743,N_4431);
or U7382 (N_7382,N_5191,N_5274);
nand U7383 (N_7383,N_4750,N_4920);
or U7384 (N_7384,N_5949,N_5181);
or U7385 (N_7385,N_4072,N_5396);
nand U7386 (N_7386,N_4476,N_5602);
or U7387 (N_7387,N_4502,N_4213);
or U7388 (N_7388,N_4459,N_4366);
or U7389 (N_7389,N_5785,N_4494);
or U7390 (N_7390,N_4264,N_4148);
or U7391 (N_7391,N_5251,N_5549);
and U7392 (N_7392,N_5799,N_4903);
nor U7393 (N_7393,N_4541,N_5047);
and U7394 (N_7394,N_4116,N_5910);
and U7395 (N_7395,N_4360,N_5083);
xnor U7396 (N_7396,N_4080,N_5917);
nand U7397 (N_7397,N_5108,N_5165);
nor U7398 (N_7398,N_4096,N_4906);
nor U7399 (N_7399,N_5604,N_4140);
nor U7400 (N_7400,N_4351,N_5126);
nand U7401 (N_7401,N_4556,N_5341);
and U7402 (N_7402,N_5552,N_5785);
and U7403 (N_7403,N_5689,N_5780);
and U7404 (N_7404,N_5286,N_4653);
nor U7405 (N_7405,N_4697,N_5536);
or U7406 (N_7406,N_5952,N_5147);
or U7407 (N_7407,N_5126,N_4826);
or U7408 (N_7408,N_5284,N_4994);
nor U7409 (N_7409,N_5648,N_4476);
and U7410 (N_7410,N_5052,N_5750);
and U7411 (N_7411,N_5759,N_5912);
nand U7412 (N_7412,N_4442,N_4649);
nor U7413 (N_7413,N_4629,N_4954);
or U7414 (N_7414,N_4714,N_4988);
or U7415 (N_7415,N_5150,N_5767);
nor U7416 (N_7416,N_4798,N_4509);
nor U7417 (N_7417,N_4330,N_5486);
nand U7418 (N_7418,N_4732,N_4714);
and U7419 (N_7419,N_4157,N_4541);
and U7420 (N_7420,N_4393,N_4828);
or U7421 (N_7421,N_5068,N_5066);
and U7422 (N_7422,N_4041,N_5688);
and U7423 (N_7423,N_4123,N_4998);
or U7424 (N_7424,N_4652,N_4127);
and U7425 (N_7425,N_4272,N_4977);
nor U7426 (N_7426,N_4984,N_4834);
nand U7427 (N_7427,N_5463,N_5706);
or U7428 (N_7428,N_4959,N_5900);
or U7429 (N_7429,N_4004,N_4878);
nand U7430 (N_7430,N_5236,N_4734);
nor U7431 (N_7431,N_4802,N_4759);
nor U7432 (N_7432,N_5565,N_5280);
and U7433 (N_7433,N_5964,N_4231);
nand U7434 (N_7434,N_5693,N_5048);
xnor U7435 (N_7435,N_4436,N_4790);
or U7436 (N_7436,N_4244,N_4024);
nand U7437 (N_7437,N_4093,N_4009);
nor U7438 (N_7438,N_5781,N_5481);
nor U7439 (N_7439,N_4142,N_4761);
xor U7440 (N_7440,N_5654,N_5965);
nor U7441 (N_7441,N_4613,N_4404);
or U7442 (N_7442,N_4939,N_4375);
or U7443 (N_7443,N_5348,N_5361);
and U7444 (N_7444,N_4437,N_4554);
nor U7445 (N_7445,N_5699,N_5559);
and U7446 (N_7446,N_4250,N_4994);
and U7447 (N_7447,N_5644,N_5782);
and U7448 (N_7448,N_4931,N_4899);
nand U7449 (N_7449,N_5862,N_4081);
nand U7450 (N_7450,N_5507,N_5326);
and U7451 (N_7451,N_4018,N_5561);
nand U7452 (N_7452,N_4429,N_5860);
nand U7453 (N_7453,N_5686,N_5224);
or U7454 (N_7454,N_4064,N_5661);
and U7455 (N_7455,N_4710,N_4702);
nor U7456 (N_7456,N_5791,N_4567);
nand U7457 (N_7457,N_5245,N_5020);
nand U7458 (N_7458,N_5130,N_4128);
nor U7459 (N_7459,N_5749,N_5880);
and U7460 (N_7460,N_4834,N_5249);
or U7461 (N_7461,N_4074,N_5325);
or U7462 (N_7462,N_4456,N_5003);
or U7463 (N_7463,N_5670,N_5266);
nor U7464 (N_7464,N_4221,N_5998);
and U7465 (N_7465,N_4756,N_4062);
and U7466 (N_7466,N_5858,N_5702);
nand U7467 (N_7467,N_4977,N_5154);
nand U7468 (N_7468,N_5856,N_5642);
nor U7469 (N_7469,N_4249,N_5815);
nand U7470 (N_7470,N_5652,N_4355);
nor U7471 (N_7471,N_5103,N_5532);
or U7472 (N_7472,N_5157,N_5506);
or U7473 (N_7473,N_4427,N_5234);
or U7474 (N_7474,N_4805,N_4159);
and U7475 (N_7475,N_5945,N_4869);
or U7476 (N_7476,N_4700,N_5106);
nor U7477 (N_7477,N_4641,N_4874);
nand U7478 (N_7478,N_5982,N_4485);
or U7479 (N_7479,N_4015,N_4930);
and U7480 (N_7480,N_5784,N_5397);
nor U7481 (N_7481,N_4152,N_5036);
nand U7482 (N_7482,N_4473,N_4191);
nand U7483 (N_7483,N_5866,N_5947);
or U7484 (N_7484,N_4253,N_5675);
xor U7485 (N_7485,N_5564,N_5936);
nor U7486 (N_7486,N_5375,N_5170);
nand U7487 (N_7487,N_5432,N_5698);
or U7488 (N_7488,N_4837,N_5653);
or U7489 (N_7489,N_4318,N_5916);
or U7490 (N_7490,N_5555,N_5939);
and U7491 (N_7491,N_5240,N_4838);
and U7492 (N_7492,N_4077,N_5937);
nor U7493 (N_7493,N_4486,N_4365);
nor U7494 (N_7494,N_4860,N_4531);
and U7495 (N_7495,N_5225,N_5483);
nand U7496 (N_7496,N_4108,N_4476);
and U7497 (N_7497,N_5378,N_4389);
or U7498 (N_7498,N_4288,N_4742);
nor U7499 (N_7499,N_4069,N_4609);
or U7500 (N_7500,N_5499,N_4185);
nand U7501 (N_7501,N_4139,N_4443);
nor U7502 (N_7502,N_4710,N_5376);
nand U7503 (N_7503,N_4514,N_4726);
and U7504 (N_7504,N_4376,N_4119);
nor U7505 (N_7505,N_5445,N_5749);
and U7506 (N_7506,N_5249,N_4598);
nor U7507 (N_7507,N_5487,N_5899);
nor U7508 (N_7508,N_4590,N_5520);
nand U7509 (N_7509,N_5218,N_5749);
nand U7510 (N_7510,N_5306,N_4689);
and U7511 (N_7511,N_5081,N_5076);
nor U7512 (N_7512,N_4823,N_4965);
or U7513 (N_7513,N_4872,N_4422);
or U7514 (N_7514,N_5140,N_5144);
and U7515 (N_7515,N_5257,N_4403);
nand U7516 (N_7516,N_5791,N_5018);
nor U7517 (N_7517,N_5029,N_4125);
nor U7518 (N_7518,N_4556,N_4040);
and U7519 (N_7519,N_5498,N_4472);
or U7520 (N_7520,N_5878,N_4463);
nor U7521 (N_7521,N_4243,N_5917);
nor U7522 (N_7522,N_5582,N_5636);
and U7523 (N_7523,N_4675,N_4425);
nor U7524 (N_7524,N_4004,N_4972);
or U7525 (N_7525,N_5557,N_5661);
and U7526 (N_7526,N_4177,N_4405);
nor U7527 (N_7527,N_4214,N_5405);
nand U7528 (N_7528,N_4270,N_5094);
nand U7529 (N_7529,N_4680,N_4837);
or U7530 (N_7530,N_5743,N_5262);
or U7531 (N_7531,N_4108,N_4480);
nor U7532 (N_7532,N_5310,N_4799);
nor U7533 (N_7533,N_5633,N_5158);
nand U7534 (N_7534,N_5658,N_4414);
nor U7535 (N_7535,N_5771,N_4309);
nor U7536 (N_7536,N_4588,N_5059);
nor U7537 (N_7537,N_5856,N_5444);
xnor U7538 (N_7538,N_4519,N_5355);
nand U7539 (N_7539,N_5041,N_4001);
and U7540 (N_7540,N_5892,N_4828);
nand U7541 (N_7541,N_5607,N_4130);
xor U7542 (N_7542,N_5734,N_5877);
or U7543 (N_7543,N_5759,N_5050);
nor U7544 (N_7544,N_5424,N_4645);
or U7545 (N_7545,N_5555,N_5911);
nor U7546 (N_7546,N_5859,N_5727);
nor U7547 (N_7547,N_4160,N_5955);
nand U7548 (N_7548,N_5062,N_5257);
xnor U7549 (N_7549,N_4823,N_4919);
nor U7550 (N_7550,N_5434,N_4825);
or U7551 (N_7551,N_5056,N_4306);
or U7552 (N_7552,N_4113,N_5978);
nand U7553 (N_7553,N_4592,N_4540);
xnor U7554 (N_7554,N_4874,N_5387);
and U7555 (N_7555,N_4900,N_4824);
nand U7556 (N_7556,N_4526,N_5981);
nor U7557 (N_7557,N_4732,N_5519);
nand U7558 (N_7558,N_4184,N_5709);
and U7559 (N_7559,N_4766,N_4497);
nand U7560 (N_7560,N_5495,N_4609);
or U7561 (N_7561,N_5142,N_5700);
nand U7562 (N_7562,N_5640,N_4998);
nand U7563 (N_7563,N_5862,N_4629);
or U7564 (N_7564,N_4536,N_4930);
nand U7565 (N_7565,N_4381,N_4641);
or U7566 (N_7566,N_4144,N_5190);
or U7567 (N_7567,N_4785,N_4960);
nand U7568 (N_7568,N_5701,N_4121);
nand U7569 (N_7569,N_5728,N_4457);
and U7570 (N_7570,N_4227,N_4880);
nand U7571 (N_7571,N_4013,N_5246);
and U7572 (N_7572,N_4095,N_4401);
nand U7573 (N_7573,N_5871,N_5985);
and U7574 (N_7574,N_5568,N_5547);
nor U7575 (N_7575,N_4498,N_4831);
nand U7576 (N_7576,N_5880,N_5219);
and U7577 (N_7577,N_5633,N_4699);
nand U7578 (N_7578,N_5991,N_5636);
or U7579 (N_7579,N_4614,N_5534);
or U7580 (N_7580,N_4714,N_4889);
and U7581 (N_7581,N_5734,N_4930);
and U7582 (N_7582,N_4153,N_5725);
nor U7583 (N_7583,N_5533,N_4477);
and U7584 (N_7584,N_4488,N_5086);
nor U7585 (N_7585,N_4709,N_5997);
nor U7586 (N_7586,N_4339,N_4852);
nor U7587 (N_7587,N_4424,N_5406);
nand U7588 (N_7588,N_5129,N_4919);
and U7589 (N_7589,N_5517,N_5802);
nand U7590 (N_7590,N_4973,N_4039);
nand U7591 (N_7591,N_5143,N_4903);
nor U7592 (N_7592,N_4526,N_4189);
and U7593 (N_7593,N_4558,N_5090);
or U7594 (N_7594,N_4195,N_4760);
nand U7595 (N_7595,N_4831,N_4038);
nand U7596 (N_7596,N_5054,N_4020);
and U7597 (N_7597,N_4384,N_5834);
nand U7598 (N_7598,N_5698,N_5489);
nor U7599 (N_7599,N_4427,N_4347);
nand U7600 (N_7600,N_4225,N_4926);
or U7601 (N_7601,N_5293,N_4458);
nor U7602 (N_7602,N_4627,N_5604);
and U7603 (N_7603,N_5336,N_5141);
nor U7604 (N_7604,N_5386,N_4213);
or U7605 (N_7605,N_5721,N_4770);
nor U7606 (N_7606,N_4248,N_4194);
or U7607 (N_7607,N_4815,N_4775);
nand U7608 (N_7608,N_5806,N_4416);
nand U7609 (N_7609,N_4058,N_5231);
nor U7610 (N_7610,N_4340,N_5162);
and U7611 (N_7611,N_5941,N_4694);
xnor U7612 (N_7612,N_4157,N_4900);
nor U7613 (N_7613,N_5562,N_4032);
nor U7614 (N_7614,N_5210,N_5489);
or U7615 (N_7615,N_5492,N_4752);
nand U7616 (N_7616,N_5456,N_4349);
or U7617 (N_7617,N_5673,N_4080);
nor U7618 (N_7618,N_5615,N_5836);
or U7619 (N_7619,N_5931,N_5211);
nor U7620 (N_7620,N_5035,N_4845);
nor U7621 (N_7621,N_4171,N_5335);
and U7622 (N_7622,N_5337,N_5272);
or U7623 (N_7623,N_4276,N_4346);
and U7624 (N_7624,N_5264,N_5608);
nand U7625 (N_7625,N_4642,N_5019);
nand U7626 (N_7626,N_4387,N_4610);
nor U7627 (N_7627,N_5125,N_5324);
nand U7628 (N_7628,N_5069,N_5759);
and U7629 (N_7629,N_4807,N_5012);
xnor U7630 (N_7630,N_5459,N_4490);
or U7631 (N_7631,N_4657,N_4738);
or U7632 (N_7632,N_4298,N_5671);
nand U7633 (N_7633,N_4041,N_4423);
or U7634 (N_7634,N_5623,N_4997);
and U7635 (N_7635,N_4471,N_4773);
nand U7636 (N_7636,N_4428,N_5181);
and U7637 (N_7637,N_5865,N_5494);
nand U7638 (N_7638,N_4823,N_4409);
nor U7639 (N_7639,N_5725,N_5543);
nand U7640 (N_7640,N_4771,N_5583);
and U7641 (N_7641,N_5062,N_4135);
and U7642 (N_7642,N_4348,N_5752);
and U7643 (N_7643,N_5587,N_4578);
and U7644 (N_7644,N_4134,N_4014);
nand U7645 (N_7645,N_5894,N_5427);
or U7646 (N_7646,N_5366,N_5453);
nor U7647 (N_7647,N_5933,N_5095);
nand U7648 (N_7648,N_5500,N_5318);
and U7649 (N_7649,N_5328,N_5218);
nor U7650 (N_7650,N_4869,N_5797);
or U7651 (N_7651,N_5475,N_4935);
nand U7652 (N_7652,N_4297,N_5191);
and U7653 (N_7653,N_4720,N_4111);
nand U7654 (N_7654,N_5571,N_4275);
and U7655 (N_7655,N_5531,N_4422);
nor U7656 (N_7656,N_4190,N_5487);
and U7657 (N_7657,N_5188,N_5040);
nor U7658 (N_7658,N_4254,N_5851);
nand U7659 (N_7659,N_5657,N_5452);
nor U7660 (N_7660,N_4162,N_5225);
or U7661 (N_7661,N_5571,N_4188);
or U7662 (N_7662,N_5400,N_4761);
or U7663 (N_7663,N_5457,N_5553);
nor U7664 (N_7664,N_5490,N_5796);
xor U7665 (N_7665,N_5169,N_4577);
and U7666 (N_7666,N_5255,N_4776);
and U7667 (N_7667,N_4729,N_5217);
nor U7668 (N_7668,N_5351,N_5318);
nand U7669 (N_7669,N_4456,N_4838);
nor U7670 (N_7670,N_5099,N_4847);
nand U7671 (N_7671,N_4673,N_5901);
xor U7672 (N_7672,N_4478,N_4302);
and U7673 (N_7673,N_4760,N_4607);
nor U7674 (N_7674,N_4353,N_4513);
or U7675 (N_7675,N_4108,N_5312);
nor U7676 (N_7676,N_5513,N_5708);
and U7677 (N_7677,N_5333,N_4750);
nand U7678 (N_7678,N_5798,N_4413);
or U7679 (N_7679,N_4911,N_4205);
or U7680 (N_7680,N_5188,N_5565);
nor U7681 (N_7681,N_4312,N_4527);
or U7682 (N_7682,N_5889,N_5750);
nand U7683 (N_7683,N_5331,N_5694);
nor U7684 (N_7684,N_4681,N_4816);
xor U7685 (N_7685,N_4267,N_5486);
or U7686 (N_7686,N_4088,N_4182);
nand U7687 (N_7687,N_4261,N_5259);
or U7688 (N_7688,N_5650,N_4001);
xnor U7689 (N_7689,N_4364,N_4826);
nand U7690 (N_7690,N_4366,N_5982);
nand U7691 (N_7691,N_4339,N_4434);
or U7692 (N_7692,N_4183,N_4756);
nand U7693 (N_7693,N_4527,N_5879);
and U7694 (N_7694,N_5025,N_5412);
or U7695 (N_7695,N_4237,N_4084);
nor U7696 (N_7696,N_4025,N_4394);
or U7697 (N_7697,N_5762,N_5949);
or U7698 (N_7698,N_5381,N_4675);
nand U7699 (N_7699,N_5426,N_5817);
nor U7700 (N_7700,N_5356,N_4663);
and U7701 (N_7701,N_5432,N_4093);
nor U7702 (N_7702,N_4563,N_5158);
and U7703 (N_7703,N_5883,N_5585);
nor U7704 (N_7704,N_4275,N_4587);
or U7705 (N_7705,N_4002,N_5271);
nand U7706 (N_7706,N_4437,N_5135);
or U7707 (N_7707,N_4465,N_4705);
nand U7708 (N_7708,N_4696,N_4266);
nand U7709 (N_7709,N_5779,N_5972);
nand U7710 (N_7710,N_5694,N_5308);
and U7711 (N_7711,N_4222,N_4511);
nor U7712 (N_7712,N_5101,N_5712);
nand U7713 (N_7713,N_5658,N_4908);
nand U7714 (N_7714,N_4108,N_5429);
nor U7715 (N_7715,N_5787,N_5052);
nor U7716 (N_7716,N_4807,N_5895);
nor U7717 (N_7717,N_4087,N_5634);
nor U7718 (N_7718,N_5827,N_5431);
nand U7719 (N_7719,N_5224,N_5604);
and U7720 (N_7720,N_4288,N_4222);
nor U7721 (N_7721,N_4982,N_5766);
nor U7722 (N_7722,N_4189,N_4476);
and U7723 (N_7723,N_4887,N_4492);
nor U7724 (N_7724,N_5011,N_4239);
or U7725 (N_7725,N_4738,N_4227);
or U7726 (N_7726,N_5382,N_5661);
or U7727 (N_7727,N_5258,N_5453);
or U7728 (N_7728,N_4474,N_5592);
nor U7729 (N_7729,N_4697,N_4172);
or U7730 (N_7730,N_5505,N_4413);
nor U7731 (N_7731,N_4522,N_4970);
xnor U7732 (N_7732,N_5281,N_5391);
nor U7733 (N_7733,N_4766,N_4928);
nor U7734 (N_7734,N_4722,N_5051);
or U7735 (N_7735,N_4912,N_5163);
nand U7736 (N_7736,N_4427,N_4925);
or U7737 (N_7737,N_5816,N_5355);
nand U7738 (N_7738,N_5403,N_4704);
nor U7739 (N_7739,N_4993,N_5555);
nor U7740 (N_7740,N_4236,N_4193);
and U7741 (N_7741,N_5847,N_5569);
nand U7742 (N_7742,N_4733,N_4090);
and U7743 (N_7743,N_4429,N_5119);
or U7744 (N_7744,N_5070,N_5327);
and U7745 (N_7745,N_4384,N_4755);
xor U7746 (N_7746,N_4545,N_4963);
or U7747 (N_7747,N_5891,N_4815);
nor U7748 (N_7748,N_5680,N_4230);
and U7749 (N_7749,N_4298,N_4911);
nor U7750 (N_7750,N_4305,N_5867);
nor U7751 (N_7751,N_5716,N_4511);
nand U7752 (N_7752,N_5788,N_4285);
and U7753 (N_7753,N_4412,N_4071);
xnor U7754 (N_7754,N_4987,N_4897);
nand U7755 (N_7755,N_5855,N_4708);
nand U7756 (N_7756,N_4040,N_4425);
or U7757 (N_7757,N_4884,N_5088);
and U7758 (N_7758,N_4846,N_4726);
nor U7759 (N_7759,N_5466,N_5165);
nor U7760 (N_7760,N_4275,N_4643);
or U7761 (N_7761,N_4277,N_5743);
nor U7762 (N_7762,N_4679,N_5654);
or U7763 (N_7763,N_5956,N_5048);
or U7764 (N_7764,N_4203,N_5339);
or U7765 (N_7765,N_5440,N_5131);
nor U7766 (N_7766,N_4660,N_5026);
nand U7767 (N_7767,N_4140,N_4378);
nor U7768 (N_7768,N_4206,N_4589);
or U7769 (N_7769,N_4173,N_4988);
or U7770 (N_7770,N_5885,N_5897);
and U7771 (N_7771,N_5041,N_4526);
nor U7772 (N_7772,N_5340,N_4717);
nand U7773 (N_7773,N_5156,N_4585);
nand U7774 (N_7774,N_5553,N_5844);
nand U7775 (N_7775,N_4243,N_4583);
or U7776 (N_7776,N_4736,N_4934);
nor U7777 (N_7777,N_5518,N_5344);
nand U7778 (N_7778,N_5479,N_5036);
and U7779 (N_7779,N_5282,N_5808);
nand U7780 (N_7780,N_4161,N_4781);
or U7781 (N_7781,N_5972,N_5224);
or U7782 (N_7782,N_4803,N_5461);
or U7783 (N_7783,N_4645,N_5143);
nor U7784 (N_7784,N_5607,N_5233);
nand U7785 (N_7785,N_5104,N_4234);
nand U7786 (N_7786,N_4608,N_5670);
nor U7787 (N_7787,N_4675,N_4209);
and U7788 (N_7788,N_5964,N_5480);
nand U7789 (N_7789,N_5783,N_5293);
nor U7790 (N_7790,N_5916,N_4929);
and U7791 (N_7791,N_5896,N_4334);
nor U7792 (N_7792,N_4721,N_5181);
nand U7793 (N_7793,N_4531,N_5431);
nor U7794 (N_7794,N_5241,N_5633);
nor U7795 (N_7795,N_5823,N_4011);
and U7796 (N_7796,N_4683,N_4967);
and U7797 (N_7797,N_4865,N_5997);
or U7798 (N_7798,N_5898,N_4537);
nor U7799 (N_7799,N_5328,N_5167);
or U7800 (N_7800,N_5579,N_4962);
xnor U7801 (N_7801,N_5701,N_5412);
nand U7802 (N_7802,N_4534,N_4587);
or U7803 (N_7803,N_5955,N_5582);
nand U7804 (N_7804,N_5625,N_5792);
and U7805 (N_7805,N_5362,N_4206);
and U7806 (N_7806,N_4108,N_4183);
or U7807 (N_7807,N_4977,N_5510);
nand U7808 (N_7808,N_5127,N_5508);
and U7809 (N_7809,N_5636,N_4567);
nand U7810 (N_7810,N_4662,N_5233);
xnor U7811 (N_7811,N_5638,N_4365);
and U7812 (N_7812,N_5137,N_4133);
nor U7813 (N_7813,N_4462,N_4630);
and U7814 (N_7814,N_4041,N_5629);
and U7815 (N_7815,N_4095,N_5503);
nor U7816 (N_7816,N_4529,N_4224);
nand U7817 (N_7817,N_4808,N_5135);
nor U7818 (N_7818,N_5627,N_4967);
or U7819 (N_7819,N_4081,N_4155);
nor U7820 (N_7820,N_4550,N_5340);
nor U7821 (N_7821,N_4672,N_5464);
nand U7822 (N_7822,N_4253,N_4469);
or U7823 (N_7823,N_4015,N_5580);
or U7824 (N_7824,N_4606,N_5093);
nor U7825 (N_7825,N_4031,N_4581);
nand U7826 (N_7826,N_4389,N_5683);
nor U7827 (N_7827,N_4419,N_5698);
nand U7828 (N_7828,N_4509,N_4079);
xnor U7829 (N_7829,N_4392,N_5256);
nand U7830 (N_7830,N_4037,N_5369);
nor U7831 (N_7831,N_5987,N_4331);
or U7832 (N_7832,N_5423,N_5416);
nor U7833 (N_7833,N_4573,N_5536);
and U7834 (N_7834,N_5397,N_4132);
or U7835 (N_7835,N_4983,N_5881);
nor U7836 (N_7836,N_4873,N_4206);
nor U7837 (N_7837,N_5821,N_4148);
nor U7838 (N_7838,N_4263,N_5310);
or U7839 (N_7839,N_5803,N_5556);
nand U7840 (N_7840,N_4740,N_4413);
and U7841 (N_7841,N_4387,N_4032);
or U7842 (N_7842,N_4464,N_5917);
nor U7843 (N_7843,N_4066,N_4297);
or U7844 (N_7844,N_4031,N_4558);
and U7845 (N_7845,N_5573,N_5941);
and U7846 (N_7846,N_4124,N_5792);
nor U7847 (N_7847,N_4001,N_5334);
and U7848 (N_7848,N_4854,N_4153);
nor U7849 (N_7849,N_5025,N_4700);
or U7850 (N_7850,N_5558,N_4462);
nor U7851 (N_7851,N_4328,N_5586);
nor U7852 (N_7852,N_4173,N_5967);
and U7853 (N_7853,N_5200,N_5845);
or U7854 (N_7854,N_5500,N_5763);
nand U7855 (N_7855,N_5809,N_5514);
nand U7856 (N_7856,N_5231,N_4259);
and U7857 (N_7857,N_5315,N_5776);
or U7858 (N_7858,N_5801,N_5077);
nor U7859 (N_7859,N_4212,N_4659);
nor U7860 (N_7860,N_4213,N_4325);
nor U7861 (N_7861,N_4137,N_4622);
and U7862 (N_7862,N_4313,N_5018);
and U7863 (N_7863,N_4349,N_5155);
and U7864 (N_7864,N_5458,N_5979);
nor U7865 (N_7865,N_4325,N_5407);
nor U7866 (N_7866,N_5223,N_4825);
nor U7867 (N_7867,N_4761,N_5623);
nand U7868 (N_7868,N_5987,N_5016);
nand U7869 (N_7869,N_4857,N_4719);
or U7870 (N_7870,N_4312,N_4767);
and U7871 (N_7871,N_4937,N_4729);
and U7872 (N_7872,N_5605,N_5335);
or U7873 (N_7873,N_5279,N_4131);
nand U7874 (N_7874,N_4945,N_5340);
nand U7875 (N_7875,N_5818,N_4902);
nor U7876 (N_7876,N_5933,N_4699);
nand U7877 (N_7877,N_5054,N_5072);
nor U7878 (N_7878,N_5602,N_4019);
nor U7879 (N_7879,N_5579,N_5527);
and U7880 (N_7880,N_4693,N_4176);
or U7881 (N_7881,N_5111,N_4445);
and U7882 (N_7882,N_5265,N_5691);
or U7883 (N_7883,N_5299,N_4534);
nand U7884 (N_7884,N_5495,N_4839);
nor U7885 (N_7885,N_5823,N_4058);
and U7886 (N_7886,N_5500,N_5913);
and U7887 (N_7887,N_5910,N_4359);
nand U7888 (N_7888,N_5577,N_5278);
nand U7889 (N_7889,N_5600,N_5999);
and U7890 (N_7890,N_5728,N_4414);
nand U7891 (N_7891,N_5624,N_4645);
and U7892 (N_7892,N_5937,N_4665);
nor U7893 (N_7893,N_5449,N_4410);
nand U7894 (N_7894,N_5180,N_4900);
nand U7895 (N_7895,N_4948,N_4487);
and U7896 (N_7896,N_4999,N_4610);
and U7897 (N_7897,N_4785,N_5224);
nand U7898 (N_7898,N_5090,N_4363);
and U7899 (N_7899,N_5213,N_4252);
and U7900 (N_7900,N_5881,N_4510);
nand U7901 (N_7901,N_5709,N_4816);
or U7902 (N_7902,N_5130,N_5055);
or U7903 (N_7903,N_4784,N_5570);
and U7904 (N_7904,N_4818,N_4529);
or U7905 (N_7905,N_4865,N_4812);
and U7906 (N_7906,N_4964,N_5478);
and U7907 (N_7907,N_5743,N_5814);
nand U7908 (N_7908,N_5538,N_4931);
or U7909 (N_7909,N_5392,N_5803);
and U7910 (N_7910,N_5328,N_5714);
and U7911 (N_7911,N_4917,N_5275);
xor U7912 (N_7912,N_4494,N_5871);
or U7913 (N_7913,N_5566,N_5633);
and U7914 (N_7914,N_4590,N_5778);
and U7915 (N_7915,N_5724,N_4908);
nand U7916 (N_7916,N_5042,N_5994);
nand U7917 (N_7917,N_4198,N_5334);
and U7918 (N_7918,N_5557,N_4446);
nand U7919 (N_7919,N_5957,N_4371);
nand U7920 (N_7920,N_5845,N_5635);
and U7921 (N_7921,N_4046,N_5724);
nand U7922 (N_7922,N_5064,N_4339);
or U7923 (N_7923,N_4522,N_5669);
or U7924 (N_7924,N_4120,N_5657);
nor U7925 (N_7925,N_4152,N_4803);
nor U7926 (N_7926,N_4348,N_4143);
nor U7927 (N_7927,N_5618,N_5871);
nor U7928 (N_7928,N_4250,N_5626);
xnor U7929 (N_7929,N_5126,N_5041);
and U7930 (N_7930,N_5327,N_5948);
and U7931 (N_7931,N_4566,N_4054);
nand U7932 (N_7932,N_5815,N_4465);
nor U7933 (N_7933,N_4271,N_4507);
and U7934 (N_7934,N_4420,N_4673);
and U7935 (N_7935,N_5657,N_5068);
and U7936 (N_7936,N_4752,N_5610);
and U7937 (N_7937,N_4501,N_5632);
and U7938 (N_7938,N_5399,N_4023);
nor U7939 (N_7939,N_4151,N_5647);
nand U7940 (N_7940,N_4804,N_4853);
nand U7941 (N_7941,N_5147,N_5136);
nor U7942 (N_7942,N_4063,N_4881);
and U7943 (N_7943,N_4293,N_5138);
nor U7944 (N_7944,N_4177,N_4687);
or U7945 (N_7945,N_4771,N_4266);
nand U7946 (N_7946,N_4247,N_5059);
nand U7947 (N_7947,N_5532,N_4116);
and U7948 (N_7948,N_5387,N_5191);
nor U7949 (N_7949,N_5849,N_5490);
nor U7950 (N_7950,N_4928,N_5646);
xor U7951 (N_7951,N_4620,N_4894);
nand U7952 (N_7952,N_4944,N_5494);
and U7953 (N_7953,N_5522,N_5576);
and U7954 (N_7954,N_4138,N_5789);
or U7955 (N_7955,N_4959,N_5821);
nand U7956 (N_7956,N_5480,N_4535);
and U7957 (N_7957,N_4620,N_5090);
nor U7958 (N_7958,N_4345,N_4087);
nor U7959 (N_7959,N_4415,N_5665);
xnor U7960 (N_7960,N_5750,N_5793);
nor U7961 (N_7961,N_5124,N_5378);
or U7962 (N_7962,N_5759,N_4205);
or U7963 (N_7963,N_4641,N_5940);
nand U7964 (N_7964,N_4288,N_4799);
nor U7965 (N_7965,N_5052,N_4337);
nand U7966 (N_7966,N_4404,N_5819);
nand U7967 (N_7967,N_4129,N_4810);
and U7968 (N_7968,N_5252,N_5663);
nor U7969 (N_7969,N_4206,N_5343);
nor U7970 (N_7970,N_5067,N_4642);
nand U7971 (N_7971,N_4608,N_5480);
nand U7972 (N_7972,N_4656,N_4543);
and U7973 (N_7973,N_4296,N_5471);
xor U7974 (N_7974,N_4565,N_5714);
nand U7975 (N_7975,N_5400,N_4486);
and U7976 (N_7976,N_4517,N_5360);
and U7977 (N_7977,N_5715,N_4070);
and U7978 (N_7978,N_4516,N_4534);
nand U7979 (N_7979,N_4460,N_5753);
and U7980 (N_7980,N_5987,N_5930);
nand U7981 (N_7981,N_4623,N_4802);
nand U7982 (N_7982,N_5208,N_5333);
nor U7983 (N_7983,N_5261,N_5703);
and U7984 (N_7984,N_4776,N_5326);
or U7985 (N_7985,N_4171,N_5803);
nand U7986 (N_7986,N_5812,N_4114);
nand U7987 (N_7987,N_4140,N_4646);
and U7988 (N_7988,N_5312,N_4699);
nand U7989 (N_7989,N_5665,N_5301);
nand U7990 (N_7990,N_5328,N_5764);
or U7991 (N_7991,N_5448,N_4797);
nor U7992 (N_7992,N_4580,N_4548);
and U7993 (N_7993,N_4120,N_4328);
and U7994 (N_7994,N_4535,N_4285);
and U7995 (N_7995,N_5857,N_4018);
and U7996 (N_7996,N_5653,N_5265);
and U7997 (N_7997,N_4832,N_5388);
and U7998 (N_7998,N_4576,N_4079);
nor U7999 (N_7999,N_5071,N_5652);
nand U8000 (N_8000,N_6444,N_6013);
nand U8001 (N_8001,N_6316,N_7776);
nand U8002 (N_8002,N_7669,N_6482);
nand U8003 (N_8003,N_6926,N_6334);
nand U8004 (N_8004,N_7011,N_7818);
nor U8005 (N_8005,N_6380,N_6985);
or U8006 (N_8006,N_7304,N_7805);
or U8007 (N_8007,N_6959,N_7578);
and U8008 (N_8008,N_7725,N_7722);
nand U8009 (N_8009,N_7106,N_6578);
nand U8010 (N_8010,N_6913,N_7091);
nor U8011 (N_8011,N_7813,N_6276);
nor U8012 (N_8012,N_7332,N_6387);
and U8013 (N_8013,N_7317,N_7280);
or U8014 (N_8014,N_6896,N_6282);
xnor U8015 (N_8015,N_7850,N_7568);
and U8016 (N_8016,N_6781,N_7871);
nand U8017 (N_8017,N_6352,N_6818);
nor U8018 (N_8018,N_6751,N_6293);
nor U8019 (N_8019,N_6491,N_6159);
nand U8020 (N_8020,N_7452,N_7630);
and U8021 (N_8021,N_6078,N_6581);
or U8022 (N_8022,N_7369,N_6085);
nor U8023 (N_8023,N_7177,N_7559);
or U8024 (N_8024,N_6880,N_6494);
nor U8025 (N_8025,N_6927,N_6255);
or U8026 (N_8026,N_6562,N_7473);
nor U8027 (N_8027,N_7436,N_6060);
or U8028 (N_8028,N_7979,N_7133);
and U8029 (N_8029,N_7203,N_6800);
or U8030 (N_8030,N_6735,N_7632);
and U8031 (N_8031,N_6804,N_7709);
or U8032 (N_8032,N_7992,N_6826);
nor U8033 (N_8033,N_7763,N_6620);
and U8034 (N_8034,N_6897,N_6991);
nand U8035 (N_8035,N_7853,N_6566);
and U8036 (N_8036,N_6840,N_6279);
nor U8037 (N_8037,N_7583,N_6400);
nand U8038 (N_8038,N_6878,N_6930);
or U8039 (N_8039,N_6260,N_6567);
and U8040 (N_8040,N_7801,N_7527);
nor U8041 (N_8041,N_6161,N_6358);
or U8042 (N_8042,N_7388,N_6730);
nand U8043 (N_8043,N_6673,N_6244);
nand U8044 (N_8044,N_7898,N_6905);
or U8045 (N_8045,N_6442,N_6226);
nor U8046 (N_8046,N_7057,N_7733);
or U8047 (N_8047,N_6597,N_7718);
and U8048 (N_8048,N_6219,N_7924);
nand U8049 (N_8049,N_7385,N_6359);
nand U8050 (N_8050,N_6126,N_7124);
and U8051 (N_8051,N_7900,N_6022);
nand U8052 (N_8052,N_6679,N_7395);
nor U8053 (N_8053,N_6104,N_7208);
and U8054 (N_8054,N_6489,N_7986);
nor U8055 (N_8055,N_7470,N_7235);
nand U8056 (N_8056,N_7370,N_7063);
nand U8057 (N_8057,N_6672,N_7954);
nand U8058 (N_8058,N_7159,N_7475);
xor U8059 (N_8059,N_6114,N_7207);
and U8060 (N_8060,N_6678,N_7381);
and U8061 (N_8061,N_6869,N_7822);
and U8062 (N_8062,N_6846,N_6427);
and U8063 (N_8063,N_7827,N_7740);
and U8064 (N_8064,N_7883,N_6314);
nor U8065 (N_8065,N_6548,N_6275);
nand U8066 (N_8066,N_6656,N_6729);
or U8067 (N_8067,N_6452,N_7111);
and U8068 (N_8068,N_7983,N_6351);
and U8069 (N_8069,N_6245,N_7966);
nand U8070 (N_8070,N_7635,N_6325);
and U8071 (N_8071,N_7026,N_6230);
or U8072 (N_8072,N_6857,N_7188);
nand U8073 (N_8073,N_6005,N_6554);
nand U8074 (N_8074,N_7637,N_6523);
nor U8075 (N_8075,N_6353,N_6668);
nand U8076 (N_8076,N_7686,N_7666);
nand U8077 (N_8077,N_7153,N_6172);
or U8078 (N_8078,N_7779,N_6922);
and U8079 (N_8079,N_7768,N_7661);
nor U8080 (N_8080,N_6041,N_7757);
or U8081 (N_8081,N_6875,N_6757);
and U8082 (N_8082,N_6036,N_7500);
nor U8083 (N_8083,N_6046,N_6158);
nand U8084 (N_8084,N_7432,N_6970);
or U8085 (N_8085,N_6369,N_7166);
and U8086 (N_8086,N_7705,N_7673);
xor U8087 (N_8087,N_7297,N_7771);
or U8088 (N_8088,N_6552,N_7045);
and U8089 (N_8089,N_6399,N_6313);
and U8090 (N_8090,N_6422,N_6394);
nand U8091 (N_8091,N_6328,N_6901);
nor U8092 (N_8092,N_7424,N_7321);
and U8093 (N_8093,N_6278,N_7922);
or U8094 (N_8094,N_7109,N_6899);
nand U8095 (N_8095,N_7114,N_7495);
nand U8096 (N_8096,N_6367,N_7327);
or U8097 (N_8097,N_6054,N_6592);
nand U8098 (N_8098,N_7482,N_6663);
nor U8099 (N_8099,N_7511,N_7950);
nor U8100 (N_8100,N_6039,N_7468);
nand U8101 (N_8101,N_6525,N_6654);
or U8102 (N_8102,N_7942,N_6631);
nand U8103 (N_8103,N_6004,N_6681);
and U8104 (N_8104,N_7622,N_7409);
nor U8105 (N_8105,N_7213,N_6902);
or U8106 (N_8106,N_7278,N_6815);
and U8107 (N_8107,N_7972,N_7078);
and U8108 (N_8108,N_6315,N_6366);
or U8109 (N_8109,N_7070,N_7331);
nor U8110 (N_8110,N_6933,N_6929);
nand U8111 (N_8111,N_7258,N_6608);
or U8112 (N_8112,N_7665,N_6438);
nor U8113 (N_8113,N_7503,N_6090);
and U8114 (N_8114,N_7743,N_7714);
nand U8115 (N_8115,N_7967,N_6253);
nor U8116 (N_8116,N_6856,N_6919);
and U8117 (N_8117,N_7835,N_7789);
or U8118 (N_8118,N_6906,N_6565);
and U8119 (N_8119,N_6629,N_6111);
and U8120 (N_8120,N_6957,N_7997);
and U8121 (N_8121,N_6205,N_6540);
and U8122 (N_8122,N_6512,N_7003);
and U8123 (N_8123,N_6762,N_7759);
and U8124 (N_8124,N_7324,N_7056);
or U8125 (N_8125,N_6938,N_7877);
and U8126 (N_8126,N_7175,N_7033);
and U8127 (N_8127,N_6295,N_7141);
and U8128 (N_8128,N_7593,N_6121);
or U8129 (N_8129,N_7335,N_6257);
and U8130 (N_8130,N_6198,N_7354);
or U8131 (N_8131,N_7150,N_6423);
nor U8132 (N_8132,N_7712,N_7919);
nand U8133 (N_8133,N_6647,N_7224);
and U8134 (N_8134,N_7537,N_6412);
or U8135 (N_8135,N_7562,N_6361);
nor U8136 (N_8136,N_7923,N_6921);
or U8137 (N_8137,N_6945,N_7471);
nor U8138 (N_8138,N_6994,N_7929);
nor U8139 (N_8139,N_6236,N_6479);
nor U8140 (N_8140,N_7732,N_7176);
nor U8141 (N_8141,N_6379,N_6954);
nor U8142 (N_8142,N_7271,N_6553);
nand U8143 (N_8143,N_7683,N_7695);
nor U8144 (N_8144,N_7041,N_6980);
and U8145 (N_8145,N_7667,N_6199);
or U8146 (N_8146,N_6460,N_6884);
and U8147 (N_8147,N_7905,N_6468);
nor U8148 (N_8148,N_7693,N_6675);
and U8149 (N_8149,N_6170,N_7507);
nor U8150 (N_8150,N_7326,N_7544);
or U8151 (N_8151,N_7108,N_6488);
and U8152 (N_8152,N_7754,N_6833);
and U8153 (N_8153,N_7202,N_7526);
and U8154 (N_8154,N_6177,N_6411);
nand U8155 (N_8155,N_7115,N_7623);
nor U8156 (N_8156,N_7832,N_7407);
or U8157 (N_8157,N_6433,N_6827);
nand U8158 (N_8158,N_6975,N_7236);
or U8159 (N_8159,N_7570,N_7659);
or U8160 (N_8160,N_6457,N_7869);
or U8161 (N_8161,N_7819,N_7874);
and U8162 (N_8162,N_7588,N_6775);
nand U8163 (N_8163,N_7497,N_6935);
and U8164 (N_8164,N_6732,N_6434);
nor U8165 (N_8165,N_7183,N_6900);
nand U8166 (N_8166,N_6419,N_6089);
and U8167 (N_8167,N_6375,N_6088);
and U8168 (N_8168,N_7004,N_7741);
nor U8169 (N_8169,N_7301,N_6885);
nand U8170 (N_8170,N_6137,N_7684);
nand U8171 (N_8171,N_6124,N_6753);
nor U8172 (N_8172,N_7677,N_7282);
or U8173 (N_8173,N_6821,N_7811);
nor U8174 (N_8174,N_7426,N_7796);
nand U8175 (N_8175,N_6149,N_7340);
nand U8176 (N_8176,N_6229,N_6813);
nor U8177 (N_8177,N_6551,N_7845);
nand U8178 (N_8178,N_6904,N_6690);
and U8179 (N_8179,N_7682,N_6538);
nor U8180 (N_8180,N_7920,N_7882);
and U8181 (N_8181,N_7716,N_6837);
or U8182 (N_8182,N_6831,N_7038);
or U8183 (N_8183,N_6425,N_7621);
or U8184 (N_8184,N_6007,N_7614);
nand U8185 (N_8185,N_6541,N_7171);
and U8186 (N_8186,N_6923,N_6536);
and U8187 (N_8187,N_7981,N_6333);
nand U8188 (N_8188,N_6232,N_7303);
nor U8189 (N_8189,N_6504,N_6166);
nand U8190 (N_8190,N_7915,N_7427);
nor U8191 (N_8191,N_6105,N_6779);
nand U8192 (N_8192,N_6274,N_6524);
and U8193 (N_8193,N_7903,N_6174);
and U8194 (N_8194,N_7116,N_7194);
and U8195 (N_8195,N_6376,N_6416);
and U8196 (N_8196,N_7008,N_7515);
and U8197 (N_8197,N_7288,N_7040);
and U8198 (N_8198,N_6795,N_7880);
or U8199 (N_8199,N_6705,N_7244);
and U8200 (N_8200,N_7787,N_6382);
or U8201 (N_8201,N_6277,N_6962);
or U8202 (N_8202,N_6402,N_7420);
or U8203 (N_8203,N_7774,N_7248);
or U8204 (N_8204,N_7387,N_7734);
or U8205 (N_8205,N_6388,N_7851);
or U8206 (N_8206,N_7201,N_7308);
and U8207 (N_8207,N_6093,N_7165);
nor U8208 (N_8208,N_7261,N_6360);
nand U8209 (N_8209,N_7058,N_6449);
nand U8210 (N_8210,N_6723,N_6684);
or U8211 (N_8211,N_7664,N_6977);
or U8212 (N_8212,N_7283,N_6183);
or U8213 (N_8213,N_7918,N_7601);
nand U8214 (N_8214,N_6171,N_6129);
and U8215 (N_8215,N_6210,N_7000);
or U8216 (N_8216,N_6758,N_6335);
or U8217 (N_8217,N_6292,N_6799);
and U8218 (N_8218,N_6961,N_7976);
or U8219 (N_8219,N_7161,N_6963);
xnor U8220 (N_8220,N_6577,N_6844);
nand U8221 (N_8221,N_7758,N_7653);
nand U8222 (N_8222,N_6662,N_7222);
nor U8223 (N_8223,N_6814,N_7240);
and U8224 (N_8224,N_7446,N_7361);
nand U8225 (N_8225,N_7160,N_6406);
nand U8226 (N_8226,N_6549,N_7138);
nand U8227 (N_8227,N_6211,N_7274);
nand U8228 (N_8228,N_7036,N_7726);
nor U8229 (N_8229,N_6564,N_7937);
nor U8230 (N_8230,N_7348,N_6644);
xor U8231 (N_8231,N_7136,N_6557);
nor U8232 (N_8232,N_7831,N_7587);
nor U8233 (N_8233,N_6971,N_6786);
or U8234 (N_8234,N_6466,N_7378);
or U8235 (N_8235,N_6863,N_7625);
and U8236 (N_8236,N_6290,N_7650);
or U8237 (N_8237,N_7368,N_7338);
or U8238 (N_8238,N_6591,N_6008);
nor U8239 (N_8239,N_6699,N_6350);
nor U8240 (N_8240,N_6530,N_6234);
nand U8241 (N_8241,N_7480,N_7545);
nand U8242 (N_8242,N_6651,N_7122);
and U8243 (N_8243,N_7199,N_6167);
or U8244 (N_8244,N_7534,N_7394);
or U8245 (N_8245,N_6252,N_6495);
or U8246 (N_8246,N_6239,N_6584);
or U8247 (N_8247,N_6766,N_6499);
or U8248 (N_8248,N_6429,N_7824);
nor U8249 (N_8249,N_7702,N_6881);
nor U8250 (N_8250,N_7467,N_7567);
and U8251 (N_8251,N_7334,N_7724);
or U8252 (N_8252,N_6575,N_7571);
nand U8253 (N_8253,N_7243,N_6306);
nor U8254 (N_8254,N_6430,N_7371);
nor U8255 (N_8255,N_6357,N_7310);
nor U8256 (N_8256,N_7459,N_6685);
nand U8257 (N_8257,N_7681,N_6304);
or U8258 (N_8258,N_7728,N_6016);
nor U8259 (N_8259,N_6269,N_7589);
or U8260 (N_8260,N_6600,N_7252);
and U8261 (N_8261,N_7052,N_6780);
nand U8262 (N_8262,N_6773,N_6958);
and U8263 (N_8263,N_6082,N_6446);
or U8264 (N_8264,N_7277,N_6502);
nand U8265 (N_8265,N_7904,N_7964);
and U8266 (N_8266,N_6969,N_6718);
nand U8267 (N_8267,N_6770,N_6640);
or U8268 (N_8268,N_6218,N_7978);
xnor U8269 (N_8269,N_6972,N_7345);
or U8270 (N_8270,N_7099,N_6667);
nand U8271 (N_8271,N_7064,N_6317);
or U8272 (N_8272,N_6664,N_6555);
nand U8273 (N_8273,N_7891,N_6871);
nor U8274 (N_8274,N_7965,N_6222);
nor U8275 (N_8275,N_6618,N_6931);
nor U8276 (N_8276,N_7085,N_6626);
and U8277 (N_8277,N_7707,N_7305);
nand U8278 (N_8278,N_6738,N_7215);
xor U8279 (N_8279,N_7790,N_7646);
and U8280 (N_8280,N_7602,N_6458);
nand U8281 (N_8281,N_7598,N_6700);
or U8282 (N_8282,N_7356,N_7412);
nor U8283 (N_8283,N_6321,N_7542);
or U8284 (N_8284,N_7281,N_6639);
nor U8285 (N_8285,N_6760,N_6096);
and U8286 (N_8286,N_7913,N_6053);
or U8287 (N_8287,N_7443,N_6537);
and U8288 (N_8288,N_7319,N_6187);
and U8289 (N_8289,N_6212,N_7841);
nor U8290 (N_8290,N_7631,N_6755);
or U8291 (N_8291,N_6836,N_6535);
nor U8292 (N_8292,N_6248,N_6687);
and U8293 (N_8293,N_7087,N_7209);
nor U8294 (N_8294,N_7580,N_7455);
nand U8295 (N_8295,N_6889,N_7023);
nor U8296 (N_8296,N_7619,N_7350);
nand U8297 (N_8297,N_6254,N_7640);
or U8298 (N_8298,N_7017,N_6864);
and U8299 (N_8299,N_7447,N_6478);
or U8300 (N_8300,N_7121,N_7826);
nand U8301 (N_8301,N_7239,N_7051);
or U8302 (N_8302,N_6409,N_6475);
and U8303 (N_8303,N_6368,N_6281);
or U8304 (N_8304,N_6747,N_6038);
nor U8305 (N_8305,N_6903,N_6745);
xor U8306 (N_8306,N_7821,N_6364);
nor U8307 (N_8307,N_7250,N_6055);
and U8308 (N_8308,N_6302,N_7386);
or U8309 (N_8309,N_7961,N_7375);
and U8310 (N_8310,N_7553,N_7896);
and U8311 (N_8311,N_6033,N_7465);
and U8312 (N_8312,N_6365,N_6338);
xnor U8313 (N_8313,N_6754,N_6983);
nand U8314 (N_8314,N_7445,N_7518);
or U8315 (N_8315,N_6120,N_6469);
or U8316 (N_8316,N_7090,N_6076);
or U8317 (N_8317,N_6569,N_7316);
nor U8318 (N_8318,N_6133,N_6204);
nand U8319 (N_8319,N_6189,N_7147);
and U8320 (N_8320,N_7413,N_7043);
nor U8321 (N_8321,N_6062,N_7836);
nand U8322 (N_8322,N_7251,N_6034);
or U8323 (N_8323,N_6470,N_6847);
or U8324 (N_8324,N_6498,N_6162);
or U8325 (N_8325,N_7897,N_6595);
and U8326 (N_8326,N_7009,N_7745);
nand U8327 (N_8327,N_7223,N_7930);
and U8328 (N_8328,N_6653,N_7270);
nand U8329 (N_8329,N_7204,N_6774);
or U8330 (N_8330,N_7807,N_7302);
or U8331 (N_8331,N_7131,N_6807);
and U8332 (N_8332,N_7449,N_6417);
and U8333 (N_8333,N_6135,N_6914);
nand U8334 (N_8334,N_7170,N_7329);
and U8335 (N_8335,N_7313,N_7096);
or U8336 (N_8336,N_7463,N_6558);
nand U8337 (N_8337,N_7067,N_7648);
or U8338 (N_8338,N_7543,N_7508);
nand U8339 (N_8339,N_6920,N_7128);
or U8340 (N_8340,N_7856,N_6015);
nand U8341 (N_8341,N_6431,N_6337);
and U8342 (N_8342,N_7925,N_6996);
nor U8343 (N_8343,N_6098,N_7268);
and U8344 (N_8344,N_7573,N_7945);
xor U8345 (N_8345,N_6023,N_6784);
or U8346 (N_8346,N_6420,N_7440);
nand U8347 (N_8347,N_6480,N_6695);
and U8348 (N_8348,N_7028,N_6691);
or U8349 (N_8349,N_6383,N_6843);
and U8350 (N_8350,N_7264,N_6570);
nand U8351 (N_8351,N_7609,N_7685);
and U8352 (N_8352,N_6697,N_7167);
or U8353 (N_8353,N_7644,N_7007);
nand U8354 (N_8354,N_7249,N_7490);
and U8355 (N_8355,N_7522,N_6816);
nand U8356 (N_8356,N_6231,N_7287);
nand U8357 (N_8357,N_7730,N_6649);
nand U8358 (N_8358,N_7088,N_6440);
nand U8359 (N_8359,N_7939,N_6891);
and U8360 (N_8360,N_6696,N_7618);
nor U8361 (N_8361,N_7047,N_6154);
and U8362 (N_8362,N_7410,N_7325);
nor U8363 (N_8363,N_6107,N_6355);
nand U8364 (N_8364,N_6934,N_7982);
nor U8365 (N_8365,N_7149,N_7504);
nand U8366 (N_8366,N_6772,N_6794);
nor U8367 (N_8367,N_7561,N_6987);
or U8368 (N_8368,N_7328,N_7756);
nor U8369 (N_8369,N_6670,N_6633);
nor U8370 (N_8370,N_6455,N_6539);
or U8371 (N_8371,N_6185,N_6250);
nor U8372 (N_8372,N_7100,N_7834);
nor U8373 (N_8373,N_7408,N_6045);
nand U8374 (N_8374,N_6764,N_6580);
nand U8375 (N_8375,N_6845,N_7989);
or U8376 (N_8376,N_7358,N_7346);
or U8377 (N_8377,N_6835,N_6533);
and U8378 (N_8378,N_7312,N_7357);
or U8379 (N_8379,N_7560,N_7808);
nand U8380 (N_8380,N_7528,N_6401);
nor U8381 (N_8381,N_7590,N_7910);
and U8382 (N_8382,N_6951,N_7608);
nor U8383 (N_8383,N_6209,N_6925);
or U8384 (N_8384,N_7362,N_7323);
nor U8385 (N_8385,N_6638,N_7383);
and U8386 (N_8386,N_6576,N_7066);
or U8387 (N_8387,N_7494,N_6630);
and U8388 (N_8388,N_6063,N_6765);
nor U8389 (N_8389,N_7400,N_6207);
nor U8390 (N_8390,N_6711,N_6037);
or U8391 (N_8391,N_6061,N_6609);
and U8392 (N_8392,N_7713,N_6946);
nor U8393 (N_8393,N_6505,N_6214);
and U8394 (N_8394,N_6395,N_6002);
or U8395 (N_8395,N_7016,N_7987);
nor U8396 (N_8396,N_6165,N_6075);
or U8397 (N_8397,N_7263,N_7963);
nand U8398 (N_8398,N_7262,N_7060);
or U8399 (N_8399,N_6830,N_6153);
or U8400 (N_8400,N_7698,N_7802);
nor U8401 (N_8401,N_6415,N_6599);
nor U8402 (N_8402,N_6228,N_6176);
nor U8403 (N_8403,N_6070,N_7696);
nor U8404 (N_8404,N_7764,N_6169);
nand U8405 (N_8405,N_6955,N_7434);
nor U8406 (N_8406,N_7781,N_6883);
nand U8407 (N_8407,N_7353,N_6142);
nor U8408 (N_8408,N_6267,N_7077);
nor U8409 (N_8409,N_7311,N_7988);
nand U8410 (N_8410,N_7633,N_7013);
nor U8411 (N_8411,N_7286,N_7355);
and U8412 (N_8412,N_6682,N_7688);
nor U8413 (N_8413,N_6966,N_7888);
or U8414 (N_8414,N_7242,N_6606);
and U8415 (N_8415,N_6151,N_6854);
and U8416 (N_8416,N_6027,N_7379);
or U8417 (N_8417,N_6324,N_7864);
or U8418 (N_8418,N_6213,N_6974);
or U8419 (N_8419,N_6462,N_6590);
nand U8420 (N_8420,N_6343,N_7001);
or U8421 (N_8421,N_6140,N_7804);
and U8422 (N_8422,N_7823,N_7479);
and U8423 (N_8423,N_7154,N_7934);
and U8424 (N_8424,N_6916,N_6559);
nand U8425 (N_8425,N_6139,N_7844);
or U8426 (N_8426,N_6693,N_7237);
nand U8427 (N_8427,N_7557,N_6243);
nand U8428 (N_8428,N_7951,N_6838);
and U8429 (N_8429,N_7555,N_7102);
nor U8430 (N_8430,N_7948,N_6490);
or U8431 (N_8431,N_6924,N_7275);
nor U8432 (N_8432,N_6132,N_7428);
nand U8433 (N_8433,N_7848,N_7765);
or U8434 (N_8434,N_7241,N_7024);
xnor U8435 (N_8435,N_7018,N_6636);
nor U8436 (N_8436,N_6393,N_6531);
nand U8437 (N_8437,N_6128,N_7185);
nor U8438 (N_8438,N_7061,N_6323);
nor U8439 (N_8439,N_7720,N_6326);
and U8440 (N_8440,N_7197,N_7652);
nor U8441 (N_8441,N_7592,N_7629);
nor U8442 (N_8442,N_6820,N_6032);
nor U8443 (N_8443,N_7753,N_6701);
nor U8444 (N_8444,N_6021,N_6928);
nand U8445 (N_8445,N_7178,N_6262);
or U8446 (N_8446,N_7069,N_7828);
nand U8447 (N_8447,N_6445,N_6509);
and U8448 (N_8448,N_7914,N_7245);
nand U8449 (N_8449,N_7390,N_6180);
or U8450 (N_8450,N_6156,N_7817);
and U8451 (N_8451,N_6110,N_6381);
or U8452 (N_8452,N_7655,N_7169);
xnor U8453 (N_8453,N_6050,N_7220);
or U8454 (N_8454,N_6615,N_6465);
nor U8455 (N_8455,N_7899,N_7546);
or U8456 (N_8456,N_7892,N_7767);
nand U8457 (N_8457,N_7617,N_6097);
or U8458 (N_8458,N_7307,N_7260);
and U8459 (N_8459,N_6118,N_7489);
nand U8460 (N_8460,N_6703,N_7752);
and U8461 (N_8461,N_6865,N_7405);
or U8462 (N_8462,N_7697,N_7212);
xnor U8463 (N_8463,N_6742,N_6362);
xor U8464 (N_8464,N_7944,N_7579);
nand U8465 (N_8465,N_6404,N_6437);
and U8466 (N_8466,N_7437,N_6208);
or U8467 (N_8467,N_6303,N_6069);
and U8468 (N_8468,N_7461,N_6583);
nor U8469 (N_8469,N_7272,N_7292);
nand U8470 (N_8470,N_6613,N_7678);
and U8471 (N_8471,N_6918,N_7531);
or U8472 (N_8472,N_6235,N_7309);
nor U8473 (N_8473,N_7607,N_6297);
nor U8474 (N_8474,N_7246,N_6095);
and U8475 (N_8475,N_7812,N_7117);
nand U8476 (N_8476,N_7135,N_7123);
nand U8477 (N_8477,N_7620,N_6009);
nand U8478 (N_8478,N_7025,N_7450);
and U8479 (N_8479,N_6761,N_7054);
nand U8480 (N_8480,N_6164,N_7735);
and U8481 (N_8481,N_6942,N_7425);
nand U8482 (N_8482,N_6859,N_7276);
or U8483 (N_8483,N_6301,N_6698);
nor U8484 (N_8484,N_6092,N_6319);
or U8485 (N_8485,N_7613,N_6202);
nand U8486 (N_8486,N_6101,N_7137);
nand U8487 (N_8487,N_7600,N_6743);
and U8488 (N_8488,N_7597,N_6798);
nor U8489 (N_8489,N_7739,N_6624);
or U8490 (N_8490,N_6439,N_7585);
and U8491 (N_8491,N_7322,N_7139);
or U8492 (N_8492,N_6787,N_6407);
and U8493 (N_8493,N_7256,N_7140);
or U8494 (N_8494,N_7985,N_6191);
nor U8495 (N_8495,N_7089,N_6612);
nor U8496 (N_8496,N_6261,N_6716);
and U8497 (N_8497,N_7969,N_6385);
nor U8498 (N_8498,N_7866,N_7059);
nand U8499 (N_8499,N_6877,N_7072);
or U8500 (N_8500,N_7806,N_7029);
or U8501 (N_8501,N_6621,N_6492);
nor U8502 (N_8502,N_7927,N_7049);
or U8503 (N_8503,N_7030,N_6224);
nand U8504 (N_8504,N_7267,N_6713);
and U8505 (N_8505,N_6750,N_7876);
nor U8506 (N_8506,N_7442,N_7861);
nand U8507 (N_8507,N_6671,N_6715);
nor U8508 (N_8508,N_6103,N_6574);
and U8509 (N_8509,N_6585,N_6464);
nand U8510 (N_8510,N_6572,N_7970);
and U8511 (N_8511,N_7854,N_6284);
or U8512 (N_8512,N_6006,N_7541);
nor U8513 (N_8513,N_7984,N_7670);
and U8514 (N_8514,N_6190,N_7676);
nand U8515 (N_8515,N_6119,N_7668);
or U8516 (N_8516,N_6655,N_7015);
and U8517 (N_8517,N_7881,N_6405);
or U8518 (N_8518,N_7098,N_7221);
nand U8519 (N_8519,N_7662,N_7125);
nor U8520 (N_8520,N_6749,N_6978);
nor U8521 (N_8521,N_6179,N_6976);
nand U8522 (N_8522,N_7019,N_6010);
nand U8523 (N_8523,N_7576,N_6907);
and U8524 (N_8524,N_7533,N_6841);
nor U8525 (N_8525,N_6341,N_7034);
or U8526 (N_8526,N_7909,N_7558);
nor U8527 (N_8527,N_7377,N_6767);
nand U8528 (N_8528,N_7285,N_6029);
nor U8529 (N_8529,N_7692,N_6674);
nor U8530 (N_8530,N_7336,N_6759);
or U8531 (N_8531,N_7911,N_7506);
nand U8532 (N_8532,N_7521,N_6193);
nor U8533 (N_8533,N_7569,N_7404);
nand U8534 (N_8534,N_6173,N_6125);
or U8535 (N_8535,N_7298,N_6501);
nor U8536 (N_8536,N_6342,N_7457);
or U8537 (N_8537,N_6748,N_6217);
nor U8538 (N_8538,N_6448,N_6858);
nand U8539 (N_8539,N_7675,N_6811);
nor U8540 (N_8540,N_7663,N_6908);
or U8541 (N_8541,N_7456,N_7778);
and U8542 (N_8542,N_6717,N_6168);
and U8543 (N_8543,N_7483,N_7174);
xor U8544 (N_8544,N_7612,N_7606);
and U8545 (N_8545,N_7391,N_6197);
nor U8546 (N_8546,N_6163,N_7849);
nor U8547 (N_8547,N_7296,N_7946);
and U8548 (N_8548,N_6825,N_6079);
nor U8549 (N_8549,N_6771,N_7727);
and U8550 (N_8550,N_7994,N_6842);
or U8551 (N_8551,N_7129,N_7190);
nor U8552 (N_8552,N_7200,N_7991);
nor U8553 (N_8553,N_6329,N_7118);
nor U8554 (N_8554,N_6339,N_6392);
nor U8555 (N_8555,N_6268,N_6853);
or U8556 (N_8556,N_6157,N_7172);
or U8557 (N_8557,N_6769,N_6299);
nor U8558 (N_8558,N_6589,N_7973);
nand U8559 (N_8559,N_7658,N_7269);
nand U8560 (N_8560,N_6436,N_6265);
nand U8561 (N_8561,N_7940,N_6017);
or U8562 (N_8562,N_6242,N_6056);
or U8563 (N_8563,N_6731,N_6997);
nand U8564 (N_8564,N_6739,N_7502);
nor U8565 (N_8565,N_7755,N_6521);
nand U8566 (N_8566,N_6175,N_6992);
nor U8567 (N_8567,N_6866,N_6291);
nor U8568 (N_8568,N_6432,N_7014);
or U8569 (N_8569,N_7960,N_6074);
and U8570 (N_8570,N_6117,N_6850);
nand U8571 (N_8571,N_7517,N_6752);
nand U8572 (N_8572,N_7144,N_7604);
and U8573 (N_8573,N_7372,N_6131);
or U8574 (N_8574,N_6258,N_6216);
or U8575 (N_8575,N_7596,N_7616);
nor U8576 (N_8576,N_7219,N_7742);
nand U8577 (N_8577,N_7975,N_6824);
or U8578 (N_8578,N_7792,N_7524);
and U8579 (N_8579,N_6702,N_7747);
nand U8580 (N_8580,N_7680,N_6915);
or U8581 (N_8581,N_6832,N_7337);
nor U8582 (N_8582,N_7878,N_7318);
nand U8583 (N_8583,N_6944,N_7498);
nor U8584 (N_8584,N_6981,N_6519);
nand U8585 (N_8585,N_7703,N_6953);
nand U8586 (N_8586,N_6112,N_6937);
nor U8587 (N_8587,N_7895,N_6511);
or U8588 (N_8588,N_6474,N_6263);
and U8589 (N_8589,N_6109,N_6048);
nand U8590 (N_8590,N_7173,N_6413);
nor U8591 (N_8591,N_7112,N_6456);
nand U8592 (N_8592,N_7933,N_7130);
nand U8593 (N_8593,N_7595,N_6408);
or U8594 (N_8594,N_7842,N_6855);
xor U8595 (N_8595,N_6892,N_7206);
nor U8596 (N_8596,N_6186,N_7259);
nor U8597 (N_8597,N_6450,N_6616);
nor U8598 (N_8598,N_7226,N_7478);
or U8599 (N_8599,N_7289,N_6534);
nand U8600 (N_8600,N_6828,N_7519);
and U8601 (N_8601,N_7254,N_6712);
nand U8602 (N_8602,N_6106,N_6378);
nand U8603 (N_8603,N_7641,N_6296);
nand U8604 (N_8604,N_7865,N_7143);
nor U8605 (N_8605,N_6071,N_7931);
nand U8606 (N_8606,N_6330,N_7065);
and U8607 (N_8607,N_7398,N_7351);
nor U8608 (N_8608,N_7751,N_7393);
or U8609 (N_8609,N_6886,N_7674);
nand U8610 (N_8610,N_6513,N_6532);
nand U8611 (N_8611,N_6047,N_7198);
and U8612 (N_8612,N_7671,N_7382);
nor U8613 (N_8613,N_7956,N_6529);
nand U8614 (N_8614,N_6227,N_7529);
or U8615 (N_8615,N_7081,N_7993);
nor U8616 (N_8616,N_7472,N_6952);
nand U8617 (N_8617,N_6588,N_7005);
and U8618 (N_8618,N_6973,N_7093);
or U8619 (N_8619,N_6057,N_6067);
or U8620 (N_8620,N_7211,N_6561);
nor U8621 (N_8621,N_7485,N_6130);
and U8622 (N_8622,N_7397,N_6340);
or U8623 (N_8623,N_6586,N_7228);
xor U8624 (N_8624,N_6203,N_7894);
nor U8625 (N_8625,N_7784,N_6066);
and U8626 (N_8626,N_7075,N_6683);
or U8627 (N_8627,N_7392,N_6563);
and U8628 (N_8628,N_7928,N_7769);
or U8629 (N_8629,N_7402,N_7690);
or U8630 (N_8630,N_7083,N_6689);
and U8631 (N_8631,N_7186,N_7840);
or U8632 (N_8632,N_7884,N_6141);
nor U8633 (N_8633,N_6873,N_7002);
nand U8634 (N_8634,N_6145,N_6949);
nor U8635 (N_8635,N_7477,N_7788);
or U8636 (N_8636,N_7523,N_7384);
and U8637 (N_8637,N_6396,N_7145);
nand U8638 (N_8638,N_6148,N_7484);
or U8639 (N_8639,N_7530,N_6635);
or U8640 (N_8640,N_7510,N_6707);
nor U8641 (N_8641,N_6134,N_6108);
nor U8642 (N_8642,N_6793,N_7902);
or U8643 (N_8643,N_6441,N_7127);
nor U8644 (N_8644,N_6882,N_6287);
nand U8645 (N_8645,N_7603,N_6990);
nor U8646 (N_8646,N_7829,N_6547);
and U8647 (N_8647,N_6628,N_6910);
nor U8648 (N_8648,N_6593,N_7225);
xor U8649 (N_8649,N_6508,N_7349);
nand U8650 (N_8650,N_6246,N_6294);
or U8651 (N_8651,N_6587,N_6515);
or U8652 (N_8652,N_7599,N_6077);
nand U8653 (N_8653,N_7076,N_6073);
and U8654 (N_8654,N_6311,N_6796);
nand U8655 (N_8655,N_6528,N_7917);
or U8656 (N_8656,N_7422,N_6058);
nor U8657 (N_8657,N_6817,N_6573);
nor U8658 (N_8658,N_7889,N_6623);
and U8659 (N_8659,N_7949,N_6386);
nand U8660 (N_8660,N_6956,N_7782);
nand U8661 (N_8661,N_6152,N_7830);
nor U8662 (N_8662,N_6298,N_6256);
or U8663 (N_8663,N_6598,N_6645);
and U8664 (N_8664,N_7053,N_6410);
or U8665 (N_8665,N_6627,N_6676);
or U8666 (N_8666,N_7660,N_7858);
nand U8667 (N_8667,N_6184,N_6040);
or U8668 (N_8668,N_7636,N_6550);
nand U8669 (N_8669,N_6861,N_7187);
or U8670 (N_8670,N_7453,N_6223);
nand U8671 (N_8671,N_7119,N_7214);
and U8672 (N_8672,N_6995,N_6848);
nor U8673 (N_8673,N_6398,N_7314);
nor U8674 (N_8674,N_6714,N_7042);
xor U8675 (N_8675,N_6030,N_6912);
or U8676 (N_8676,N_6641,N_6614);
and U8677 (N_8677,N_7838,N_7363);
nor U8678 (N_8678,N_6461,N_7857);
nor U8679 (N_8679,N_7926,N_6136);
nor U8680 (N_8680,N_7189,N_6989);
and U8681 (N_8681,N_6500,N_7572);
or U8682 (N_8682,N_6031,N_6206);
nand U8683 (N_8683,N_6233,N_7959);
nand U8684 (N_8684,N_6271,N_7330);
nand U8685 (N_8685,N_7750,N_7996);
or U8686 (N_8686,N_6619,N_7628);
or U8687 (N_8687,N_7179,N_6194);
and U8688 (N_8688,N_6322,N_6596);
nor U8689 (N_8689,N_7247,N_6560);
nand U8690 (N_8690,N_7196,N_6790);
or U8691 (N_8691,N_7068,N_7574);
nand U8692 (N_8692,N_7134,N_6603);
nand U8693 (N_8693,N_6094,N_7294);
and U8694 (N_8694,N_6849,N_6657);
xor U8695 (N_8695,N_7101,N_7803);
and U8696 (N_8696,N_6241,N_7156);
and U8697 (N_8697,N_7389,N_6763);
and U8698 (N_8698,N_6879,N_6289);
nand U8699 (N_8699,N_6091,N_7875);
nor U8700 (N_8700,N_6686,N_7365);
and U8701 (N_8701,N_7770,N_7162);
and U8702 (N_8702,N_6042,N_7431);
and U8703 (N_8703,N_7210,N_7279);
nor U8704 (N_8704,N_6087,N_7647);
and U8705 (N_8705,N_7403,N_7885);
or U8706 (N_8706,N_6435,N_6984);
nor U8707 (N_8707,N_6454,N_6719);
and U8708 (N_8708,N_6809,N_7094);
or U8709 (N_8709,N_6862,N_6473);
xnor U8710 (N_8710,N_6116,N_6968);
or U8711 (N_8711,N_7651,N_7535);
nand U8712 (N_8712,N_7738,N_6860);
or U8713 (N_8713,N_6377,N_6485);
nor U8714 (N_8714,N_7797,N_7441);
and U8715 (N_8715,N_7935,N_6785);
nor U8716 (N_8716,N_6336,N_6307);
nor U8717 (N_8717,N_6898,N_7704);
nand U8718 (N_8718,N_6424,N_7611);
or U8719 (N_8719,N_6666,N_7512);
and U8720 (N_8720,N_7615,N_7953);
and U8721 (N_8721,N_7234,N_6270);
and U8722 (N_8722,N_7772,N_6373);
or U8723 (N_8723,N_7870,N_7295);
nand U8724 (N_8724,N_7890,N_6138);
nand U8725 (N_8725,N_6993,N_7341);
nand U8726 (N_8726,N_6518,N_7748);
nand U8727 (N_8727,N_7594,N_6579);
and U8728 (N_8728,N_6451,N_7229);
nand U8729 (N_8729,N_7624,N_7893);
nor U8730 (N_8730,N_7039,N_6285);
nor U8731 (N_8731,N_7380,N_6932);
and U8732 (N_8732,N_6659,N_6607);
and U8733 (N_8733,N_6220,N_6272);
and U8734 (N_8734,N_7414,N_6356);
and U8735 (N_8735,N_7591,N_7126);
nor U8736 (N_8736,N_7342,N_6354);
or U8737 (N_8737,N_7481,N_6273);
nor U8738 (N_8738,N_7762,N_7364);
nor U8739 (N_8739,N_7266,N_7105);
nand U8740 (N_8740,N_7487,N_7577);
and U8741 (N_8741,N_7205,N_6374);
and U8742 (N_8742,N_7672,N_6086);
nor U8743 (N_8743,N_7941,N_7451);
or U8744 (N_8744,N_6288,N_7957);
and U8745 (N_8745,N_6543,N_7113);
nand U8746 (N_8746,N_6834,N_6939);
and U8747 (N_8747,N_6812,N_6428);
and U8748 (N_8748,N_6950,N_6318);
nor U8749 (N_8749,N_6721,N_6472);
nor U8750 (N_8750,N_7021,N_6348);
or U8751 (N_8751,N_7839,N_7366);
nor U8752 (N_8752,N_7947,N_6744);
nor U8753 (N_8753,N_6734,N_6346);
nor U8754 (N_8754,N_6390,N_6517);
and U8755 (N_8755,N_7785,N_7417);
or U8756 (N_8756,N_6384,N_7031);
nor U8757 (N_8757,N_6965,N_7855);
and U8758 (N_8758,N_6084,N_6669);
nand U8759 (N_8759,N_6852,N_6720);
nand U8760 (N_8760,N_7180,N_7816);
or U8761 (N_8761,N_7048,N_7103);
or U8762 (N_8762,N_6601,N_6677);
and U8763 (N_8763,N_7843,N_7233);
or U8764 (N_8764,N_7564,N_6874);
nor U8765 (N_8765,N_6249,N_6363);
nand U8766 (N_8766,N_6028,N_7921);
and U8767 (N_8767,N_7359,N_6722);
and U8768 (N_8768,N_7995,N_7719);
nor U8769 (N_8769,N_6986,N_7488);
nand U8770 (N_8770,N_7293,N_7586);
nand U8771 (N_8771,N_7549,N_7773);
or U8772 (N_8772,N_6520,N_6372);
and U8773 (N_8773,N_7513,N_6310);
nand U8774 (N_8774,N_7376,N_7761);
nor U8775 (N_8775,N_6123,N_7373);
nor U8776 (N_8776,N_6345,N_6266);
and U8777 (N_8777,N_7265,N_6851);
nand U8778 (N_8778,N_7439,N_7097);
nand U8779 (N_8779,N_7999,N_6493);
nand U8780 (N_8780,N_6019,N_6822);
and U8781 (N_8781,N_7438,N_7810);
and U8782 (N_8782,N_6240,N_6788);
and U8783 (N_8783,N_6099,N_6476);
and U8784 (N_8784,N_6737,N_7253);
or U8785 (N_8785,N_6688,N_7496);
nand U8786 (N_8786,N_6648,N_7415);
nand U8787 (N_8787,N_7012,N_7736);
nor U8788 (N_8788,N_6496,N_7230);
or U8789 (N_8789,N_7182,N_7406);
and U8790 (N_8790,N_7932,N_7723);
and U8791 (N_8791,N_7158,N_7777);
or U8792 (N_8792,N_6201,N_7548);
or U8793 (N_8793,N_7847,N_7974);
or U8794 (N_8794,N_6895,N_7168);
or U8795 (N_8795,N_7155,N_6443);
or U8796 (N_8796,N_6000,N_6556);
xor U8797 (N_8797,N_6192,N_6792);
nor U8798 (N_8798,N_7080,N_6819);
xnor U8799 (N_8799,N_6467,N_6147);
and U8800 (N_8800,N_7649,N_7232);
or U8801 (N_8801,N_6611,N_6999);
nor U8802 (N_8802,N_6706,N_7418);
and U8803 (N_8803,N_6344,N_6320);
or U8804 (N_8804,N_7079,N_7859);
and U8805 (N_8805,N_7679,N_7912);
nor U8806 (N_8806,N_7998,N_6768);
nor U8807 (N_8807,N_6967,N_7699);
nand U8808 (N_8808,N_7971,N_6025);
and U8809 (N_8809,N_7315,N_7462);
nor U8810 (N_8810,N_7645,N_7694);
nand U8811 (N_8811,N_7216,N_6544);
and U8812 (N_8812,N_7794,N_6238);
nor U8813 (N_8813,N_7815,N_7231);
or U8814 (N_8814,N_6327,N_6453);
nand U8815 (N_8815,N_6100,N_7775);
nand U8816 (N_8816,N_7968,N_7306);
nor U8817 (N_8817,N_7010,N_6637);
nor U8818 (N_8818,N_6940,N_7721);
or U8819 (N_8819,N_6632,N_6594);
nand U8820 (N_8820,N_7492,N_7691);
nor U8821 (N_8821,N_6660,N_7820);
and U8822 (N_8822,N_7766,N_6522);
xnor U8823 (N_8823,N_6113,N_7191);
nand U8824 (N_8824,N_6988,N_7084);
and U8825 (N_8825,N_6740,N_7474);
and U8826 (N_8826,N_6605,N_6797);
xor U8827 (N_8827,N_6710,N_7547);
nor U8828 (N_8828,N_7444,N_6909);
nor U8829 (N_8829,N_6463,N_7022);
nand U8830 (N_8830,N_7958,N_6789);
nand U8831 (N_8831,N_6064,N_6568);
nand U8832 (N_8832,N_7708,N_6805);
or U8833 (N_8833,N_7783,N_7107);
nand U8834 (N_8834,N_7862,N_6503);
or U8835 (N_8835,N_7565,N_7299);
nor U8836 (N_8836,N_6810,N_7411);
nand U8837 (N_8837,N_7977,N_6483);
and U8838 (N_8838,N_7505,N_7701);
and U8839 (N_8839,N_7540,N_6870);
nor U8840 (N_8840,N_6300,N_7551);
nand U8841 (N_8841,N_7255,N_6911);
or U8842 (N_8842,N_7906,N_7799);
nor U8843 (N_8843,N_7509,N_7656);
and U8844 (N_8844,N_7626,N_6646);
nor U8845 (N_8845,N_6894,N_7706);
and U8846 (N_8846,N_6650,N_6237);
nand U8847 (N_8847,N_6264,N_7627);
or U8848 (N_8848,N_6661,N_6012);
or U8849 (N_8849,N_6709,N_6259);
xnor U8850 (N_8850,N_6115,N_7744);
nand U8851 (N_8851,N_7654,N_6155);
or U8852 (N_8852,N_6196,N_7867);
and U8853 (N_8853,N_6527,N_7493);
or U8854 (N_8854,N_6024,N_7786);
or U8855 (N_8855,N_6868,N_7132);
nor U8856 (N_8856,N_6602,N_6776);
nand U8857 (N_8857,N_7962,N_7062);
and U8858 (N_8858,N_6680,N_6658);
nor U8859 (N_8859,N_6867,N_6941);
or U8860 (N_8860,N_7793,N_7374);
or U8861 (N_8861,N_6643,N_6081);
or U8862 (N_8862,N_7642,N_6546);
and U8863 (N_8863,N_7006,N_7657);
nand U8864 (N_8864,N_6652,N_7020);
nand U8865 (N_8865,N_7737,N_7938);
nand U8866 (N_8866,N_6733,N_6160);
nand U8867 (N_8867,N_7164,N_7689);
and U8868 (N_8868,N_6756,N_7055);
nor U8869 (N_8869,N_6280,N_6247);
and U8870 (N_8870,N_6221,N_6477);
and U8871 (N_8871,N_6035,N_6782);
nor U8872 (N_8872,N_7582,N_6068);
and U8873 (N_8873,N_7486,N_7458);
and U8874 (N_8874,N_7990,N_6803);
and U8875 (N_8875,N_7863,N_7192);
nand U8876 (N_8876,N_6146,N_6052);
and U8877 (N_8877,N_6026,N_6414);
or U8878 (N_8878,N_7610,N_7416);
nand U8879 (N_8879,N_7687,N_7448);
nand U8880 (N_8880,N_6571,N_7333);
and U8881 (N_8881,N_6215,N_6486);
nand U8882 (N_8882,N_6542,N_7584);
or U8883 (N_8883,N_7532,N_6403);
nor U8884 (N_8884,N_7814,N_6065);
nor U8885 (N_8885,N_7872,N_6371);
nor U8886 (N_8886,N_7110,N_7086);
nand U8887 (N_8887,N_7809,N_7430);
or U8888 (N_8888,N_7120,N_7501);
xnor U8889 (N_8889,N_7151,N_7852);
or U8890 (N_8890,N_7195,N_6018);
and U8891 (N_8891,N_6308,N_7795);
and U8892 (N_8892,N_7879,N_6806);
or U8893 (N_8893,N_7157,N_6072);
and U8894 (N_8894,N_6704,N_7396);
or U8895 (N_8895,N_6421,N_7291);
nand U8896 (N_8896,N_6708,N_7731);
nor U8897 (N_8897,N_7218,N_6182);
nor U8898 (N_8898,N_7466,N_6051);
and U8899 (N_8899,N_6225,N_7952);
nor U8900 (N_8900,N_7860,N_6001);
nor U8901 (N_8901,N_6694,N_6044);
or U8902 (N_8902,N_7711,N_6604);
nor U8903 (N_8903,N_6516,N_6484);
or U8904 (N_8904,N_7476,N_6506);
and U8905 (N_8905,N_6011,N_7257);
nor U8906 (N_8906,N_7536,N_6823);
nor U8907 (N_8907,N_7421,N_7873);
and U8908 (N_8908,N_6332,N_6839);
nor U8909 (N_8909,N_6736,N_7433);
nor U8910 (N_8910,N_7035,N_7435);
nor U8911 (N_8911,N_7715,N_7300);
nor U8912 (N_8912,N_6200,N_7846);
or U8913 (N_8913,N_7238,N_6872);
or U8914 (N_8914,N_7046,N_7833);
nand U8915 (N_8915,N_6481,N_6692);
nor U8916 (N_8916,N_7566,N_6471);
and U8917 (N_8917,N_6808,N_7491);
and U8918 (N_8918,N_6497,N_7955);
nor U8919 (N_8919,N_6725,N_7525);
nand U8920 (N_8920,N_7074,N_6059);
nor U8921 (N_8921,N_6080,N_6526);
nand U8922 (N_8922,N_7550,N_7980);
nand U8923 (N_8923,N_7825,N_6622);
nand U8924 (N_8924,N_7552,N_7032);
nand U8925 (N_8925,N_7837,N_7227);
nor U8926 (N_8926,N_7916,N_7464);
or U8927 (N_8927,N_6083,N_7399);
xor U8928 (N_8928,N_7554,N_6943);
or U8929 (N_8929,N_6960,N_6122);
nand U8930 (N_8930,N_7791,N_7146);
and U8931 (N_8931,N_7037,N_7360);
and U8932 (N_8932,N_6514,N_6507);
nand U8933 (N_8933,N_6998,N_7643);
nor U8934 (N_8934,N_6617,N_7605);
or U8935 (N_8935,N_7887,N_7886);
nand U8936 (N_8936,N_6286,N_7419);
or U8937 (N_8937,N_7344,N_6331);
nor U8938 (N_8938,N_6020,N_6888);
nor U8939 (N_8939,N_7343,N_6724);
nor U8940 (N_8940,N_7163,N_7429);
and U8941 (N_8941,N_6309,N_7639);
xor U8942 (N_8942,N_7556,N_6418);
nor U8943 (N_8943,N_7634,N_6312);
nor U8944 (N_8944,N_7901,N_6887);
and U8945 (N_8945,N_6982,N_6389);
and U8946 (N_8946,N_6801,N_6948);
nor U8947 (N_8947,N_7516,N_7520);
or U8948 (N_8948,N_6979,N_7760);
nor U8949 (N_8949,N_6003,N_7082);
and U8950 (N_8950,N_7454,N_7367);
or U8951 (N_8951,N_6746,N_7181);
nor U8952 (N_8952,N_7868,N_6890);
or U8953 (N_8953,N_7514,N_6893);
nor U8954 (N_8954,N_6347,N_7710);
nor U8955 (N_8955,N_6777,N_6195);
nor U8956 (N_8956,N_6936,N_7095);
or U8957 (N_8957,N_6102,N_6349);
and U8958 (N_8958,N_6728,N_6778);
nor U8959 (N_8959,N_6283,N_7104);
and U8960 (N_8960,N_7581,N_6726);
or U8961 (N_8961,N_7469,N_6545);
or U8962 (N_8962,N_7148,N_7184);
or U8963 (N_8963,N_6829,N_6665);
nor U8964 (N_8964,N_6634,N_7073);
or U8965 (N_8965,N_6370,N_6625);
or U8966 (N_8966,N_7936,N_7273);
nand U8967 (N_8967,N_6459,N_6802);
nor U8968 (N_8968,N_6143,N_6391);
and U8969 (N_8969,N_7800,N_7284);
or U8970 (N_8970,N_6447,N_6150);
and U8971 (N_8971,N_6305,N_6426);
nand U8972 (N_8972,N_6181,N_6144);
and U8973 (N_8973,N_7717,N_7638);
and U8974 (N_8974,N_7729,N_7352);
and U8975 (N_8975,N_6964,N_6741);
nand U8976 (N_8976,N_6642,N_7746);
nand U8977 (N_8977,N_7217,N_7193);
nand U8978 (N_8978,N_6791,N_6876);
nand U8979 (N_8979,N_6127,N_7539);
and U8980 (N_8980,N_6397,N_7290);
nor U8981 (N_8981,N_7563,N_7401);
nor U8982 (N_8982,N_6510,N_7044);
nor U8983 (N_8983,N_7423,N_6014);
and U8984 (N_8984,N_7943,N_7142);
nor U8985 (N_8985,N_6043,N_6582);
nor U8986 (N_8986,N_7798,N_6251);
nor U8987 (N_8987,N_6487,N_7050);
nand U8988 (N_8988,N_7339,N_6783);
nand U8989 (N_8989,N_7320,N_6049);
nor U8990 (N_8990,N_6947,N_6917);
or U8991 (N_8991,N_7460,N_6727);
nand U8992 (N_8992,N_7538,N_7907);
nand U8993 (N_8993,N_7071,N_6178);
nand U8994 (N_8994,N_6188,N_6610);
nor U8995 (N_8995,N_7027,N_7749);
nor U8996 (N_8996,N_7575,N_7780);
or U8997 (N_8997,N_7499,N_7152);
nand U8998 (N_8998,N_7908,N_7347);
or U8999 (N_8999,N_7092,N_7700);
or U9000 (N_9000,N_7941,N_7440);
nand U9001 (N_9001,N_6209,N_7164);
nand U9002 (N_9002,N_6438,N_6844);
or U9003 (N_9003,N_6526,N_7479);
xnor U9004 (N_9004,N_6171,N_7235);
or U9005 (N_9005,N_7596,N_6854);
nor U9006 (N_9006,N_6427,N_6413);
nor U9007 (N_9007,N_6960,N_6316);
and U9008 (N_9008,N_7884,N_7408);
nand U9009 (N_9009,N_7834,N_7824);
xor U9010 (N_9010,N_7782,N_7458);
nand U9011 (N_9011,N_6155,N_7938);
and U9012 (N_9012,N_7317,N_6389);
and U9013 (N_9013,N_7353,N_6015);
nand U9014 (N_9014,N_6043,N_6301);
nand U9015 (N_9015,N_6806,N_7156);
or U9016 (N_9016,N_6890,N_6138);
or U9017 (N_9017,N_7955,N_7192);
nand U9018 (N_9018,N_7365,N_7220);
or U9019 (N_9019,N_7360,N_7674);
and U9020 (N_9020,N_7563,N_7881);
nor U9021 (N_9021,N_7976,N_7552);
nand U9022 (N_9022,N_6773,N_6402);
nand U9023 (N_9023,N_6772,N_6408);
or U9024 (N_9024,N_6663,N_6018);
nor U9025 (N_9025,N_7937,N_6345);
nor U9026 (N_9026,N_6276,N_7134);
nand U9027 (N_9027,N_7563,N_7814);
and U9028 (N_9028,N_7285,N_6641);
nand U9029 (N_9029,N_7248,N_7106);
xnor U9030 (N_9030,N_7896,N_7924);
nand U9031 (N_9031,N_7177,N_7245);
nor U9032 (N_9032,N_6269,N_6551);
nor U9033 (N_9033,N_6347,N_6286);
and U9034 (N_9034,N_7983,N_7266);
nand U9035 (N_9035,N_7586,N_7910);
nand U9036 (N_9036,N_6665,N_6333);
nand U9037 (N_9037,N_6681,N_7804);
nand U9038 (N_9038,N_7360,N_6481);
or U9039 (N_9039,N_6198,N_6216);
nor U9040 (N_9040,N_7000,N_6392);
and U9041 (N_9041,N_7508,N_6589);
or U9042 (N_9042,N_7022,N_6681);
nor U9043 (N_9043,N_7590,N_6405);
nor U9044 (N_9044,N_7740,N_7286);
nor U9045 (N_9045,N_7504,N_6953);
nand U9046 (N_9046,N_6313,N_7178);
or U9047 (N_9047,N_7665,N_7272);
nor U9048 (N_9048,N_7702,N_6096);
xor U9049 (N_9049,N_7095,N_6805);
or U9050 (N_9050,N_7379,N_7658);
and U9051 (N_9051,N_7172,N_7383);
nand U9052 (N_9052,N_6754,N_7096);
nand U9053 (N_9053,N_7613,N_7158);
xnor U9054 (N_9054,N_6801,N_7579);
nand U9055 (N_9055,N_7691,N_7815);
nor U9056 (N_9056,N_7901,N_6133);
nand U9057 (N_9057,N_6253,N_6676);
nand U9058 (N_9058,N_6540,N_7095);
nand U9059 (N_9059,N_6782,N_7552);
or U9060 (N_9060,N_7049,N_6392);
nor U9061 (N_9061,N_6234,N_6507);
or U9062 (N_9062,N_7513,N_6436);
and U9063 (N_9063,N_6653,N_7453);
nor U9064 (N_9064,N_7669,N_6380);
nor U9065 (N_9065,N_6234,N_7966);
and U9066 (N_9066,N_6515,N_6377);
and U9067 (N_9067,N_7082,N_6674);
xnor U9068 (N_9068,N_6875,N_6683);
nand U9069 (N_9069,N_6657,N_6045);
and U9070 (N_9070,N_7425,N_7438);
or U9071 (N_9071,N_6993,N_6432);
xor U9072 (N_9072,N_6386,N_7139);
and U9073 (N_9073,N_6582,N_7685);
nor U9074 (N_9074,N_7336,N_7010);
nor U9075 (N_9075,N_7541,N_6237);
nand U9076 (N_9076,N_6467,N_7714);
or U9077 (N_9077,N_7629,N_7132);
nand U9078 (N_9078,N_6300,N_7990);
and U9079 (N_9079,N_7429,N_7188);
nor U9080 (N_9080,N_6450,N_6509);
nor U9081 (N_9081,N_7236,N_6213);
nand U9082 (N_9082,N_6322,N_6786);
and U9083 (N_9083,N_6644,N_6285);
nand U9084 (N_9084,N_6586,N_6487);
nor U9085 (N_9085,N_7839,N_6040);
nand U9086 (N_9086,N_7894,N_7511);
nand U9087 (N_9087,N_6504,N_6237);
nand U9088 (N_9088,N_6380,N_6934);
and U9089 (N_9089,N_6926,N_7284);
and U9090 (N_9090,N_6195,N_6546);
nor U9091 (N_9091,N_6355,N_6138);
and U9092 (N_9092,N_7491,N_6376);
nand U9093 (N_9093,N_6330,N_7584);
xnor U9094 (N_9094,N_7495,N_6480);
or U9095 (N_9095,N_7575,N_7533);
or U9096 (N_9096,N_6069,N_6970);
nor U9097 (N_9097,N_7672,N_7348);
and U9098 (N_9098,N_7795,N_7712);
nand U9099 (N_9099,N_7975,N_7007);
and U9100 (N_9100,N_6450,N_6468);
nand U9101 (N_9101,N_7763,N_6594);
nor U9102 (N_9102,N_7974,N_7747);
or U9103 (N_9103,N_7460,N_7966);
nor U9104 (N_9104,N_7511,N_6045);
nor U9105 (N_9105,N_7765,N_6998);
nor U9106 (N_9106,N_7706,N_7092);
nand U9107 (N_9107,N_6325,N_6295);
or U9108 (N_9108,N_6005,N_7166);
nor U9109 (N_9109,N_6916,N_7726);
nor U9110 (N_9110,N_7465,N_6129);
and U9111 (N_9111,N_7390,N_7901);
nand U9112 (N_9112,N_7269,N_7366);
nor U9113 (N_9113,N_6897,N_7807);
and U9114 (N_9114,N_6451,N_7622);
nand U9115 (N_9115,N_6950,N_7820);
nand U9116 (N_9116,N_7590,N_7581);
or U9117 (N_9117,N_6042,N_7586);
or U9118 (N_9118,N_6393,N_7919);
nor U9119 (N_9119,N_6955,N_6643);
xor U9120 (N_9120,N_6098,N_7166);
nor U9121 (N_9121,N_7075,N_6462);
xnor U9122 (N_9122,N_6852,N_7809);
nor U9123 (N_9123,N_7786,N_7805);
or U9124 (N_9124,N_6819,N_6568);
or U9125 (N_9125,N_6021,N_6229);
or U9126 (N_9126,N_7771,N_6846);
or U9127 (N_9127,N_7356,N_7670);
nand U9128 (N_9128,N_6975,N_6727);
nor U9129 (N_9129,N_6391,N_7701);
nand U9130 (N_9130,N_7243,N_7235);
nor U9131 (N_9131,N_7883,N_6252);
nor U9132 (N_9132,N_6407,N_7421);
nor U9133 (N_9133,N_6790,N_7051);
nand U9134 (N_9134,N_6067,N_6860);
nand U9135 (N_9135,N_6232,N_7095);
xor U9136 (N_9136,N_7216,N_6493);
nand U9137 (N_9137,N_7571,N_6265);
and U9138 (N_9138,N_7669,N_6168);
nor U9139 (N_9139,N_7223,N_6712);
or U9140 (N_9140,N_6335,N_6484);
nor U9141 (N_9141,N_7490,N_6296);
nor U9142 (N_9142,N_7073,N_7832);
or U9143 (N_9143,N_6023,N_6808);
and U9144 (N_9144,N_7565,N_6048);
nand U9145 (N_9145,N_6648,N_6172);
nand U9146 (N_9146,N_7316,N_6832);
nor U9147 (N_9147,N_6436,N_6524);
nor U9148 (N_9148,N_6816,N_7944);
nor U9149 (N_9149,N_6879,N_7701);
or U9150 (N_9150,N_6477,N_6387);
nor U9151 (N_9151,N_7942,N_7101);
nor U9152 (N_9152,N_7242,N_6754);
or U9153 (N_9153,N_6911,N_6002);
and U9154 (N_9154,N_6315,N_7779);
or U9155 (N_9155,N_7270,N_7727);
nor U9156 (N_9156,N_6736,N_7812);
or U9157 (N_9157,N_7340,N_6974);
and U9158 (N_9158,N_6985,N_7680);
xor U9159 (N_9159,N_7120,N_7018);
and U9160 (N_9160,N_6788,N_6625);
and U9161 (N_9161,N_7370,N_6445);
and U9162 (N_9162,N_7373,N_6860);
nor U9163 (N_9163,N_6186,N_6809);
nor U9164 (N_9164,N_6598,N_7200);
or U9165 (N_9165,N_6836,N_6528);
or U9166 (N_9166,N_7039,N_6404);
nor U9167 (N_9167,N_7540,N_7736);
nor U9168 (N_9168,N_6520,N_7709);
xor U9169 (N_9169,N_7544,N_7424);
nor U9170 (N_9170,N_7862,N_7340);
and U9171 (N_9171,N_7976,N_6232);
or U9172 (N_9172,N_7833,N_6864);
or U9173 (N_9173,N_6920,N_6034);
nor U9174 (N_9174,N_6111,N_6799);
nand U9175 (N_9175,N_7634,N_7631);
or U9176 (N_9176,N_6088,N_7719);
or U9177 (N_9177,N_7885,N_7568);
and U9178 (N_9178,N_7778,N_6363);
nor U9179 (N_9179,N_6126,N_6434);
or U9180 (N_9180,N_7235,N_7606);
nor U9181 (N_9181,N_6896,N_7122);
nand U9182 (N_9182,N_7460,N_7333);
and U9183 (N_9183,N_7472,N_6110);
or U9184 (N_9184,N_6436,N_6906);
and U9185 (N_9185,N_7229,N_6176);
nand U9186 (N_9186,N_6150,N_7726);
nor U9187 (N_9187,N_6435,N_6446);
and U9188 (N_9188,N_7110,N_6744);
nor U9189 (N_9189,N_6384,N_7371);
or U9190 (N_9190,N_6076,N_6887);
nor U9191 (N_9191,N_6905,N_7871);
and U9192 (N_9192,N_7967,N_7289);
nor U9193 (N_9193,N_7246,N_6251);
nand U9194 (N_9194,N_7706,N_7853);
xnor U9195 (N_9195,N_7141,N_6097);
or U9196 (N_9196,N_6240,N_7783);
nor U9197 (N_9197,N_6539,N_6339);
nor U9198 (N_9198,N_7689,N_6990);
and U9199 (N_9199,N_6616,N_7850);
nor U9200 (N_9200,N_7598,N_6598);
nor U9201 (N_9201,N_7146,N_7405);
nor U9202 (N_9202,N_7396,N_6718);
or U9203 (N_9203,N_7781,N_6180);
or U9204 (N_9204,N_7193,N_7866);
or U9205 (N_9205,N_6181,N_7800);
nor U9206 (N_9206,N_7599,N_6933);
nor U9207 (N_9207,N_6684,N_6902);
and U9208 (N_9208,N_6305,N_6466);
and U9209 (N_9209,N_6798,N_7129);
or U9210 (N_9210,N_7844,N_7133);
nand U9211 (N_9211,N_7988,N_6359);
nor U9212 (N_9212,N_6394,N_7861);
nor U9213 (N_9213,N_7401,N_7863);
and U9214 (N_9214,N_6233,N_6925);
nand U9215 (N_9215,N_6180,N_7117);
nand U9216 (N_9216,N_6116,N_6868);
and U9217 (N_9217,N_7363,N_6686);
or U9218 (N_9218,N_7445,N_7805);
nor U9219 (N_9219,N_6481,N_7129);
nand U9220 (N_9220,N_6499,N_7350);
nor U9221 (N_9221,N_7536,N_6186);
nand U9222 (N_9222,N_6676,N_6539);
nand U9223 (N_9223,N_6135,N_7678);
and U9224 (N_9224,N_7074,N_6595);
or U9225 (N_9225,N_7209,N_6821);
nand U9226 (N_9226,N_6843,N_7057);
or U9227 (N_9227,N_6257,N_7771);
nand U9228 (N_9228,N_7830,N_6588);
and U9229 (N_9229,N_7813,N_6256);
nand U9230 (N_9230,N_7624,N_6630);
or U9231 (N_9231,N_7021,N_6431);
nand U9232 (N_9232,N_6662,N_6217);
and U9233 (N_9233,N_6715,N_7654);
xnor U9234 (N_9234,N_7141,N_7203);
nor U9235 (N_9235,N_6533,N_7996);
nand U9236 (N_9236,N_6406,N_6312);
or U9237 (N_9237,N_6797,N_7011);
or U9238 (N_9238,N_6585,N_6288);
nand U9239 (N_9239,N_7523,N_6625);
nand U9240 (N_9240,N_6705,N_6902);
nor U9241 (N_9241,N_6863,N_7218);
nand U9242 (N_9242,N_6498,N_6568);
and U9243 (N_9243,N_7524,N_6917);
xor U9244 (N_9244,N_7394,N_7425);
and U9245 (N_9245,N_6142,N_7295);
and U9246 (N_9246,N_7724,N_6589);
or U9247 (N_9247,N_7309,N_6620);
nor U9248 (N_9248,N_7657,N_7127);
nor U9249 (N_9249,N_7183,N_7647);
or U9250 (N_9250,N_7627,N_6037);
or U9251 (N_9251,N_7806,N_7605);
nand U9252 (N_9252,N_7373,N_6372);
nor U9253 (N_9253,N_6644,N_7908);
nand U9254 (N_9254,N_7734,N_6920);
nand U9255 (N_9255,N_6343,N_6479);
nor U9256 (N_9256,N_6410,N_7573);
or U9257 (N_9257,N_7138,N_6436);
nor U9258 (N_9258,N_6490,N_7279);
xnor U9259 (N_9259,N_7244,N_7473);
and U9260 (N_9260,N_6214,N_7857);
nor U9261 (N_9261,N_7562,N_6331);
and U9262 (N_9262,N_6532,N_7694);
and U9263 (N_9263,N_6451,N_6167);
xor U9264 (N_9264,N_7272,N_6244);
nand U9265 (N_9265,N_6485,N_7424);
and U9266 (N_9266,N_6271,N_7421);
nand U9267 (N_9267,N_7281,N_7766);
nand U9268 (N_9268,N_7287,N_6550);
nand U9269 (N_9269,N_7662,N_7640);
nand U9270 (N_9270,N_6032,N_7851);
or U9271 (N_9271,N_6808,N_6835);
or U9272 (N_9272,N_6681,N_6112);
and U9273 (N_9273,N_7717,N_7058);
and U9274 (N_9274,N_7143,N_7340);
nand U9275 (N_9275,N_6564,N_6181);
or U9276 (N_9276,N_7312,N_6884);
and U9277 (N_9277,N_6914,N_6060);
nand U9278 (N_9278,N_6211,N_6779);
and U9279 (N_9279,N_7469,N_7414);
and U9280 (N_9280,N_6621,N_6111);
xor U9281 (N_9281,N_7877,N_6521);
or U9282 (N_9282,N_6010,N_6450);
and U9283 (N_9283,N_7599,N_7880);
nand U9284 (N_9284,N_7885,N_6047);
or U9285 (N_9285,N_6345,N_6709);
and U9286 (N_9286,N_6112,N_7496);
or U9287 (N_9287,N_7115,N_6069);
and U9288 (N_9288,N_7249,N_6895);
nor U9289 (N_9289,N_6592,N_6144);
and U9290 (N_9290,N_7777,N_7758);
and U9291 (N_9291,N_7757,N_6200);
and U9292 (N_9292,N_6787,N_6926);
nand U9293 (N_9293,N_6666,N_7279);
or U9294 (N_9294,N_7444,N_7634);
nand U9295 (N_9295,N_7231,N_7034);
and U9296 (N_9296,N_7601,N_7734);
nor U9297 (N_9297,N_7314,N_7404);
or U9298 (N_9298,N_6011,N_6279);
nand U9299 (N_9299,N_6595,N_6686);
and U9300 (N_9300,N_6055,N_7740);
nand U9301 (N_9301,N_6160,N_7955);
or U9302 (N_9302,N_6553,N_7210);
or U9303 (N_9303,N_6185,N_7047);
and U9304 (N_9304,N_7405,N_6793);
nand U9305 (N_9305,N_7667,N_7898);
nor U9306 (N_9306,N_7678,N_6864);
or U9307 (N_9307,N_7155,N_7671);
xnor U9308 (N_9308,N_6381,N_7874);
and U9309 (N_9309,N_7402,N_6689);
nor U9310 (N_9310,N_7570,N_7875);
and U9311 (N_9311,N_7864,N_6679);
and U9312 (N_9312,N_6198,N_7653);
nor U9313 (N_9313,N_7162,N_7389);
and U9314 (N_9314,N_7105,N_7627);
xor U9315 (N_9315,N_7829,N_6904);
or U9316 (N_9316,N_7301,N_7614);
and U9317 (N_9317,N_7616,N_7013);
or U9318 (N_9318,N_6630,N_7890);
and U9319 (N_9319,N_7941,N_6094);
nand U9320 (N_9320,N_7593,N_6085);
nor U9321 (N_9321,N_7386,N_6629);
or U9322 (N_9322,N_6954,N_6531);
and U9323 (N_9323,N_7683,N_6119);
or U9324 (N_9324,N_7776,N_7563);
or U9325 (N_9325,N_6541,N_7990);
nor U9326 (N_9326,N_6792,N_6071);
and U9327 (N_9327,N_7146,N_6877);
nand U9328 (N_9328,N_6951,N_6586);
and U9329 (N_9329,N_7553,N_7727);
nor U9330 (N_9330,N_6442,N_6323);
and U9331 (N_9331,N_6111,N_7107);
and U9332 (N_9332,N_6681,N_7341);
nand U9333 (N_9333,N_6738,N_7443);
nor U9334 (N_9334,N_7469,N_6812);
nand U9335 (N_9335,N_6122,N_7151);
nor U9336 (N_9336,N_7889,N_7749);
nor U9337 (N_9337,N_7785,N_7937);
nand U9338 (N_9338,N_6276,N_7542);
or U9339 (N_9339,N_7261,N_6290);
or U9340 (N_9340,N_7644,N_7481);
nand U9341 (N_9341,N_7660,N_7534);
or U9342 (N_9342,N_6134,N_7990);
nor U9343 (N_9343,N_7414,N_7319);
or U9344 (N_9344,N_7696,N_7509);
nand U9345 (N_9345,N_6613,N_6499);
nor U9346 (N_9346,N_6789,N_7507);
nor U9347 (N_9347,N_6031,N_6786);
xor U9348 (N_9348,N_6354,N_6188);
and U9349 (N_9349,N_7187,N_6050);
and U9350 (N_9350,N_6517,N_7544);
or U9351 (N_9351,N_6528,N_7412);
nor U9352 (N_9352,N_7124,N_7232);
nor U9353 (N_9353,N_7963,N_6265);
or U9354 (N_9354,N_6931,N_7773);
nand U9355 (N_9355,N_6762,N_6069);
nor U9356 (N_9356,N_7251,N_7735);
xnor U9357 (N_9357,N_7467,N_6662);
and U9358 (N_9358,N_7709,N_7039);
and U9359 (N_9359,N_7477,N_7172);
nor U9360 (N_9360,N_7627,N_7374);
and U9361 (N_9361,N_7810,N_7205);
nand U9362 (N_9362,N_6194,N_6804);
nand U9363 (N_9363,N_6440,N_6657);
or U9364 (N_9364,N_7952,N_7039);
or U9365 (N_9365,N_6991,N_7905);
or U9366 (N_9366,N_6162,N_7292);
and U9367 (N_9367,N_7646,N_6285);
xnor U9368 (N_9368,N_6952,N_7113);
and U9369 (N_9369,N_7340,N_6752);
or U9370 (N_9370,N_7738,N_6818);
nor U9371 (N_9371,N_7613,N_6486);
nand U9372 (N_9372,N_6131,N_6707);
nor U9373 (N_9373,N_6578,N_7300);
and U9374 (N_9374,N_6578,N_7774);
nor U9375 (N_9375,N_7982,N_6957);
nand U9376 (N_9376,N_7983,N_6668);
and U9377 (N_9377,N_7761,N_7155);
or U9378 (N_9378,N_7152,N_6826);
and U9379 (N_9379,N_7351,N_6213);
nand U9380 (N_9380,N_7451,N_7495);
and U9381 (N_9381,N_6206,N_7407);
nor U9382 (N_9382,N_6422,N_6761);
nor U9383 (N_9383,N_6629,N_6337);
nor U9384 (N_9384,N_6045,N_6387);
and U9385 (N_9385,N_7249,N_6268);
or U9386 (N_9386,N_6829,N_6347);
or U9387 (N_9387,N_7900,N_7494);
nor U9388 (N_9388,N_6778,N_6283);
nand U9389 (N_9389,N_7143,N_7536);
nor U9390 (N_9390,N_7641,N_7265);
xnor U9391 (N_9391,N_6122,N_7674);
or U9392 (N_9392,N_6624,N_6222);
nor U9393 (N_9393,N_7577,N_6190);
and U9394 (N_9394,N_7307,N_7200);
nand U9395 (N_9395,N_6643,N_7118);
nand U9396 (N_9396,N_7895,N_6831);
nand U9397 (N_9397,N_7757,N_7419);
or U9398 (N_9398,N_7836,N_6833);
or U9399 (N_9399,N_7224,N_7659);
or U9400 (N_9400,N_6802,N_6606);
nor U9401 (N_9401,N_6253,N_7526);
and U9402 (N_9402,N_7285,N_7677);
nand U9403 (N_9403,N_7902,N_7645);
and U9404 (N_9404,N_7172,N_6475);
or U9405 (N_9405,N_6323,N_7630);
nand U9406 (N_9406,N_7681,N_6960);
nor U9407 (N_9407,N_6777,N_6260);
nor U9408 (N_9408,N_6002,N_7400);
and U9409 (N_9409,N_6359,N_6352);
nor U9410 (N_9410,N_6884,N_6332);
nand U9411 (N_9411,N_7240,N_6480);
nor U9412 (N_9412,N_6478,N_7798);
or U9413 (N_9413,N_6686,N_6209);
nand U9414 (N_9414,N_7748,N_6034);
nor U9415 (N_9415,N_6923,N_7266);
or U9416 (N_9416,N_7074,N_7576);
nor U9417 (N_9417,N_7886,N_6250);
nand U9418 (N_9418,N_6683,N_6226);
and U9419 (N_9419,N_6813,N_7958);
nand U9420 (N_9420,N_6477,N_7373);
or U9421 (N_9421,N_6620,N_6469);
nand U9422 (N_9422,N_7333,N_7212);
nand U9423 (N_9423,N_7669,N_7068);
or U9424 (N_9424,N_7413,N_7270);
or U9425 (N_9425,N_6143,N_7350);
or U9426 (N_9426,N_6485,N_7532);
and U9427 (N_9427,N_6056,N_6588);
nor U9428 (N_9428,N_7984,N_7402);
nor U9429 (N_9429,N_7015,N_7088);
nor U9430 (N_9430,N_7592,N_6507);
or U9431 (N_9431,N_6290,N_6137);
nand U9432 (N_9432,N_6115,N_6816);
nand U9433 (N_9433,N_7315,N_7609);
nor U9434 (N_9434,N_6353,N_6418);
and U9435 (N_9435,N_7035,N_7814);
or U9436 (N_9436,N_7802,N_6750);
and U9437 (N_9437,N_7497,N_7650);
nand U9438 (N_9438,N_6493,N_7058);
or U9439 (N_9439,N_7595,N_6697);
nor U9440 (N_9440,N_7476,N_6904);
nand U9441 (N_9441,N_7134,N_7023);
or U9442 (N_9442,N_7397,N_6266);
nor U9443 (N_9443,N_6418,N_7330);
and U9444 (N_9444,N_6416,N_6565);
nand U9445 (N_9445,N_6151,N_6882);
and U9446 (N_9446,N_6014,N_7041);
nand U9447 (N_9447,N_6592,N_6136);
and U9448 (N_9448,N_7783,N_6679);
and U9449 (N_9449,N_7564,N_7418);
or U9450 (N_9450,N_6706,N_6346);
nor U9451 (N_9451,N_6665,N_7015);
and U9452 (N_9452,N_7169,N_7120);
nor U9453 (N_9453,N_7535,N_6331);
nand U9454 (N_9454,N_6107,N_7131);
nand U9455 (N_9455,N_6945,N_7304);
or U9456 (N_9456,N_6391,N_7914);
nor U9457 (N_9457,N_6169,N_6418);
or U9458 (N_9458,N_7027,N_6318);
nand U9459 (N_9459,N_6046,N_6905);
nand U9460 (N_9460,N_6872,N_6618);
nor U9461 (N_9461,N_6808,N_7558);
and U9462 (N_9462,N_7585,N_6850);
nand U9463 (N_9463,N_6428,N_6315);
xnor U9464 (N_9464,N_7414,N_6207);
or U9465 (N_9465,N_6842,N_6361);
or U9466 (N_9466,N_6300,N_7434);
nand U9467 (N_9467,N_7149,N_7120);
nor U9468 (N_9468,N_6973,N_6734);
or U9469 (N_9469,N_7804,N_7898);
nor U9470 (N_9470,N_7304,N_7797);
and U9471 (N_9471,N_6196,N_6448);
and U9472 (N_9472,N_7227,N_6263);
nand U9473 (N_9473,N_6168,N_7511);
nor U9474 (N_9474,N_7150,N_7653);
and U9475 (N_9475,N_7104,N_7382);
nand U9476 (N_9476,N_6882,N_7197);
nand U9477 (N_9477,N_7609,N_7306);
nand U9478 (N_9478,N_6398,N_6125);
nand U9479 (N_9479,N_6272,N_6614);
nand U9480 (N_9480,N_7798,N_6002);
nor U9481 (N_9481,N_6480,N_7292);
and U9482 (N_9482,N_7388,N_6465);
and U9483 (N_9483,N_6588,N_7976);
and U9484 (N_9484,N_7641,N_6434);
and U9485 (N_9485,N_6570,N_7169);
nand U9486 (N_9486,N_7659,N_6754);
nand U9487 (N_9487,N_7789,N_6683);
or U9488 (N_9488,N_6798,N_7081);
nor U9489 (N_9489,N_7296,N_6339);
or U9490 (N_9490,N_7885,N_6873);
nor U9491 (N_9491,N_7827,N_7864);
nand U9492 (N_9492,N_6663,N_6896);
nand U9493 (N_9493,N_6306,N_7530);
nor U9494 (N_9494,N_7836,N_6738);
and U9495 (N_9495,N_7019,N_6065);
or U9496 (N_9496,N_7003,N_7741);
or U9497 (N_9497,N_6894,N_6236);
nand U9498 (N_9498,N_6840,N_6852);
and U9499 (N_9499,N_7996,N_6721);
or U9500 (N_9500,N_6732,N_7745);
nor U9501 (N_9501,N_7603,N_6859);
nor U9502 (N_9502,N_7623,N_6485);
or U9503 (N_9503,N_6686,N_7650);
or U9504 (N_9504,N_6385,N_7032);
nand U9505 (N_9505,N_7618,N_7136);
or U9506 (N_9506,N_6535,N_7494);
or U9507 (N_9507,N_6411,N_7588);
nor U9508 (N_9508,N_7102,N_7159);
and U9509 (N_9509,N_6914,N_7419);
and U9510 (N_9510,N_6389,N_7895);
and U9511 (N_9511,N_6261,N_6028);
or U9512 (N_9512,N_6463,N_6403);
nor U9513 (N_9513,N_6153,N_6820);
nor U9514 (N_9514,N_6931,N_6199);
nand U9515 (N_9515,N_7593,N_7382);
nor U9516 (N_9516,N_6696,N_7832);
nor U9517 (N_9517,N_6965,N_7624);
nor U9518 (N_9518,N_7385,N_6349);
nor U9519 (N_9519,N_7111,N_7074);
or U9520 (N_9520,N_6751,N_7437);
nor U9521 (N_9521,N_7397,N_7473);
and U9522 (N_9522,N_7493,N_7313);
or U9523 (N_9523,N_7642,N_7702);
and U9524 (N_9524,N_6553,N_7255);
nand U9525 (N_9525,N_6264,N_6530);
nor U9526 (N_9526,N_7382,N_7499);
nor U9527 (N_9527,N_7749,N_7369);
nor U9528 (N_9528,N_7357,N_7750);
nor U9529 (N_9529,N_6265,N_6498);
nor U9530 (N_9530,N_7647,N_6655);
and U9531 (N_9531,N_6837,N_6463);
nand U9532 (N_9532,N_7879,N_6372);
nor U9533 (N_9533,N_6943,N_6548);
and U9534 (N_9534,N_6405,N_6694);
nor U9535 (N_9535,N_6814,N_6738);
or U9536 (N_9536,N_6441,N_7569);
nor U9537 (N_9537,N_6000,N_6641);
nand U9538 (N_9538,N_6680,N_7515);
and U9539 (N_9539,N_7169,N_6632);
and U9540 (N_9540,N_6798,N_7845);
or U9541 (N_9541,N_7828,N_6064);
nor U9542 (N_9542,N_7293,N_6826);
or U9543 (N_9543,N_6266,N_7764);
or U9544 (N_9544,N_6073,N_7824);
and U9545 (N_9545,N_7669,N_6996);
or U9546 (N_9546,N_7598,N_7863);
xor U9547 (N_9547,N_7643,N_6183);
nor U9548 (N_9548,N_6464,N_6530);
or U9549 (N_9549,N_6250,N_7651);
nand U9550 (N_9550,N_6254,N_6286);
or U9551 (N_9551,N_7278,N_6725);
and U9552 (N_9552,N_6894,N_6120);
nand U9553 (N_9553,N_6222,N_6330);
nand U9554 (N_9554,N_6627,N_6991);
nor U9555 (N_9555,N_7749,N_7951);
and U9556 (N_9556,N_6166,N_7686);
and U9557 (N_9557,N_7814,N_7235);
nor U9558 (N_9558,N_6057,N_6842);
and U9559 (N_9559,N_7551,N_6894);
and U9560 (N_9560,N_7751,N_7643);
or U9561 (N_9561,N_7191,N_7092);
nand U9562 (N_9562,N_7691,N_6680);
nand U9563 (N_9563,N_7375,N_6217);
nor U9564 (N_9564,N_7838,N_7160);
nor U9565 (N_9565,N_7303,N_6073);
and U9566 (N_9566,N_7874,N_7140);
nand U9567 (N_9567,N_7873,N_6985);
nor U9568 (N_9568,N_6913,N_6003);
nand U9569 (N_9569,N_7392,N_7734);
nand U9570 (N_9570,N_6568,N_7743);
nor U9571 (N_9571,N_7149,N_7390);
or U9572 (N_9572,N_7637,N_7311);
and U9573 (N_9573,N_7128,N_7576);
nand U9574 (N_9574,N_7499,N_7114);
nor U9575 (N_9575,N_6987,N_7763);
nand U9576 (N_9576,N_6152,N_6496);
nand U9577 (N_9577,N_6903,N_6819);
nand U9578 (N_9578,N_7277,N_6053);
nand U9579 (N_9579,N_7856,N_6725);
and U9580 (N_9580,N_7644,N_7536);
and U9581 (N_9581,N_7207,N_7530);
nand U9582 (N_9582,N_7212,N_6841);
and U9583 (N_9583,N_7981,N_6929);
or U9584 (N_9584,N_7762,N_7173);
nand U9585 (N_9585,N_6091,N_7602);
and U9586 (N_9586,N_7367,N_7812);
nand U9587 (N_9587,N_6571,N_6325);
nand U9588 (N_9588,N_6454,N_7232);
nand U9589 (N_9589,N_6976,N_7139);
nand U9590 (N_9590,N_6169,N_6228);
nor U9591 (N_9591,N_6954,N_7746);
and U9592 (N_9592,N_7764,N_6588);
or U9593 (N_9593,N_7624,N_6231);
or U9594 (N_9594,N_7081,N_6505);
nor U9595 (N_9595,N_7993,N_6555);
or U9596 (N_9596,N_7895,N_6103);
and U9597 (N_9597,N_6684,N_7499);
and U9598 (N_9598,N_7590,N_7701);
nor U9599 (N_9599,N_7467,N_6496);
nor U9600 (N_9600,N_7673,N_7359);
and U9601 (N_9601,N_6825,N_6656);
nand U9602 (N_9602,N_7860,N_7648);
nor U9603 (N_9603,N_7102,N_6798);
or U9604 (N_9604,N_7050,N_6470);
nor U9605 (N_9605,N_6589,N_6698);
nand U9606 (N_9606,N_7610,N_7611);
xnor U9607 (N_9607,N_7020,N_7455);
nand U9608 (N_9608,N_6145,N_6068);
nor U9609 (N_9609,N_6918,N_6700);
and U9610 (N_9610,N_6756,N_6409);
nand U9611 (N_9611,N_7995,N_6381);
nand U9612 (N_9612,N_6732,N_6514);
nor U9613 (N_9613,N_7204,N_7875);
nor U9614 (N_9614,N_7550,N_7557);
nand U9615 (N_9615,N_6857,N_7926);
xnor U9616 (N_9616,N_7087,N_6551);
nand U9617 (N_9617,N_6437,N_7028);
nand U9618 (N_9618,N_7994,N_7857);
nor U9619 (N_9619,N_7770,N_7422);
and U9620 (N_9620,N_6118,N_7168);
or U9621 (N_9621,N_6470,N_6321);
nor U9622 (N_9622,N_7935,N_7802);
or U9623 (N_9623,N_6047,N_6805);
nor U9624 (N_9624,N_7518,N_6855);
xnor U9625 (N_9625,N_7297,N_7633);
or U9626 (N_9626,N_6124,N_6074);
or U9627 (N_9627,N_6099,N_7768);
nand U9628 (N_9628,N_7364,N_7579);
or U9629 (N_9629,N_7537,N_6631);
and U9630 (N_9630,N_6070,N_6421);
and U9631 (N_9631,N_6195,N_7976);
or U9632 (N_9632,N_7618,N_6110);
nor U9633 (N_9633,N_6421,N_6427);
nand U9634 (N_9634,N_6535,N_6436);
and U9635 (N_9635,N_7417,N_6945);
or U9636 (N_9636,N_6900,N_7862);
nand U9637 (N_9637,N_6043,N_7322);
nand U9638 (N_9638,N_6626,N_7536);
and U9639 (N_9639,N_6599,N_7635);
xnor U9640 (N_9640,N_7319,N_7022);
nand U9641 (N_9641,N_7881,N_6520);
and U9642 (N_9642,N_6082,N_7258);
nor U9643 (N_9643,N_6156,N_7820);
nand U9644 (N_9644,N_7962,N_7787);
and U9645 (N_9645,N_7556,N_6336);
and U9646 (N_9646,N_6597,N_6961);
nand U9647 (N_9647,N_7197,N_7530);
or U9648 (N_9648,N_6501,N_6369);
nor U9649 (N_9649,N_7625,N_7062);
nand U9650 (N_9650,N_7279,N_6315);
or U9651 (N_9651,N_6198,N_7370);
nor U9652 (N_9652,N_7765,N_6082);
or U9653 (N_9653,N_6489,N_7092);
and U9654 (N_9654,N_6069,N_7564);
or U9655 (N_9655,N_7025,N_6726);
nor U9656 (N_9656,N_7779,N_6847);
and U9657 (N_9657,N_6124,N_6736);
and U9658 (N_9658,N_6722,N_7420);
nor U9659 (N_9659,N_7182,N_6907);
and U9660 (N_9660,N_7345,N_7389);
or U9661 (N_9661,N_7319,N_6515);
or U9662 (N_9662,N_7359,N_6753);
nor U9663 (N_9663,N_7665,N_6648);
and U9664 (N_9664,N_6451,N_6071);
and U9665 (N_9665,N_7898,N_6548);
or U9666 (N_9666,N_6371,N_7602);
and U9667 (N_9667,N_6344,N_7657);
nand U9668 (N_9668,N_7845,N_6078);
nand U9669 (N_9669,N_6144,N_7590);
nand U9670 (N_9670,N_7610,N_6236);
or U9671 (N_9671,N_6084,N_7522);
nand U9672 (N_9672,N_7868,N_6485);
nor U9673 (N_9673,N_7024,N_7089);
and U9674 (N_9674,N_6882,N_7649);
or U9675 (N_9675,N_7199,N_7647);
nand U9676 (N_9676,N_7334,N_7379);
and U9677 (N_9677,N_6749,N_7018);
nor U9678 (N_9678,N_7696,N_6562);
and U9679 (N_9679,N_7041,N_6804);
nor U9680 (N_9680,N_7388,N_7997);
nand U9681 (N_9681,N_7337,N_6317);
or U9682 (N_9682,N_7739,N_6200);
nand U9683 (N_9683,N_6049,N_6107);
and U9684 (N_9684,N_7360,N_7161);
nand U9685 (N_9685,N_7451,N_7771);
nor U9686 (N_9686,N_7282,N_6665);
nor U9687 (N_9687,N_7669,N_6129);
nor U9688 (N_9688,N_6280,N_7614);
nand U9689 (N_9689,N_7242,N_7178);
nor U9690 (N_9690,N_7267,N_6533);
nand U9691 (N_9691,N_7400,N_7734);
or U9692 (N_9692,N_6062,N_7120);
and U9693 (N_9693,N_7316,N_7707);
xor U9694 (N_9694,N_6190,N_7727);
or U9695 (N_9695,N_7048,N_7779);
and U9696 (N_9696,N_7691,N_7203);
xnor U9697 (N_9697,N_7209,N_7869);
nor U9698 (N_9698,N_6423,N_7584);
nor U9699 (N_9699,N_7483,N_7808);
and U9700 (N_9700,N_6343,N_6377);
xnor U9701 (N_9701,N_7338,N_6712);
nor U9702 (N_9702,N_7676,N_6448);
and U9703 (N_9703,N_6136,N_6482);
and U9704 (N_9704,N_6087,N_6441);
nand U9705 (N_9705,N_7849,N_7325);
or U9706 (N_9706,N_7251,N_6715);
nor U9707 (N_9707,N_6777,N_6693);
nor U9708 (N_9708,N_6365,N_7942);
nand U9709 (N_9709,N_7390,N_7636);
and U9710 (N_9710,N_7196,N_7944);
nand U9711 (N_9711,N_6886,N_6301);
nand U9712 (N_9712,N_6829,N_7805);
nand U9713 (N_9713,N_6842,N_7980);
and U9714 (N_9714,N_7751,N_7283);
nor U9715 (N_9715,N_6384,N_6351);
nor U9716 (N_9716,N_7934,N_6135);
nand U9717 (N_9717,N_6884,N_7483);
or U9718 (N_9718,N_6319,N_6563);
nor U9719 (N_9719,N_7543,N_6780);
nand U9720 (N_9720,N_6419,N_6527);
and U9721 (N_9721,N_6689,N_6010);
and U9722 (N_9722,N_6172,N_6728);
nand U9723 (N_9723,N_7080,N_6331);
or U9724 (N_9724,N_6495,N_6128);
or U9725 (N_9725,N_6775,N_7732);
and U9726 (N_9726,N_7529,N_6372);
nor U9727 (N_9727,N_7147,N_6020);
or U9728 (N_9728,N_7103,N_7916);
nor U9729 (N_9729,N_7538,N_7721);
and U9730 (N_9730,N_7415,N_6888);
nor U9731 (N_9731,N_6857,N_7246);
nor U9732 (N_9732,N_7547,N_6678);
nand U9733 (N_9733,N_7823,N_7698);
nand U9734 (N_9734,N_7093,N_7002);
nand U9735 (N_9735,N_7402,N_7148);
nand U9736 (N_9736,N_7228,N_7984);
or U9737 (N_9737,N_6482,N_6248);
nor U9738 (N_9738,N_7615,N_7325);
or U9739 (N_9739,N_7720,N_6582);
or U9740 (N_9740,N_7180,N_7318);
and U9741 (N_9741,N_6353,N_6088);
and U9742 (N_9742,N_7694,N_7794);
or U9743 (N_9743,N_6607,N_6097);
and U9744 (N_9744,N_6320,N_6165);
nor U9745 (N_9745,N_6834,N_6993);
nor U9746 (N_9746,N_6659,N_7446);
or U9747 (N_9747,N_6512,N_6149);
nor U9748 (N_9748,N_6292,N_7058);
and U9749 (N_9749,N_6156,N_6556);
nor U9750 (N_9750,N_6224,N_7104);
or U9751 (N_9751,N_6635,N_7884);
nor U9752 (N_9752,N_7944,N_6779);
or U9753 (N_9753,N_6812,N_7810);
and U9754 (N_9754,N_6258,N_6903);
nand U9755 (N_9755,N_7421,N_7659);
nand U9756 (N_9756,N_6257,N_6418);
nand U9757 (N_9757,N_6856,N_6295);
or U9758 (N_9758,N_6315,N_7646);
nor U9759 (N_9759,N_6134,N_7686);
nor U9760 (N_9760,N_7724,N_6999);
xor U9761 (N_9761,N_7212,N_7045);
nor U9762 (N_9762,N_7559,N_7408);
nand U9763 (N_9763,N_7097,N_6745);
and U9764 (N_9764,N_6577,N_7168);
xor U9765 (N_9765,N_7540,N_7131);
or U9766 (N_9766,N_6188,N_7913);
nand U9767 (N_9767,N_6542,N_7058);
nor U9768 (N_9768,N_6971,N_6924);
or U9769 (N_9769,N_7810,N_7905);
nand U9770 (N_9770,N_6094,N_7677);
or U9771 (N_9771,N_6996,N_7411);
nor U9772 (N_9772,N_7947,N_6545);
nand U9773 (N_9773,N_6974,N_7337);
nor U9774 (N_9774,N_7172,N_6115);
and U9775 (N_9775,N_7120,N_7859);
nor U9776 (N_9776,N_7307,N_6668);
and U9777 (N_9777,N_7884,N_6573);
and U9778 (N_9778,N_7902,N_7612);
nor U9779 (N_9779,N_7462,N_6243);
and U9780 (N_9780,N_7866,N_7228);
nor U9781 (N_9781,N_7304,N_6653);
nor U9782 (N_9782,N_6962,N_6562);
xnor U9783 (N_9783,N_6018,N_7166);
or U9784 (N_9784,N_7856,N_7195);
or U9785 (N_9785,N_6333,N_6671);
nand U9786 (N_9786,N_7802,N_6667);
nand U9787 (N_9787,N_6993,N_7783);
and U9788 (N_9788,N_6328,N_6118);
nor U9789 (N_9789,N_7331,N_6137);
and U9790 (N_9790,N_6209,N_6978);
nor U9791 (N_9791,N_6941,N_6796);
nand U9792 (N_9792,N_6711,N_7953);
nor U9793 (N_9793,N_6190,N_6235);
or U9794 (N_9794,N_7674,N_6509);
or U9795 (N_9795,N_6665,N_7938);
nand U9796 (N_9796,N_7413,N_7294);
or U9797 (N_9797,N_7369,N_6655);
and U9798 (N_9798,N_7867,N_6056);
and U9799 (N_9799,N_6153,N_6884);
or U9800 (N_9800,N_7213,N_7045);
or U9801 (N_9801,N_7217,N_6781);
or U9802 (N_9802,N_6603,N_7113);
nor U9803 (N_9803,N_7856,N_7804);
or U9804 (N_9804,N_6070,N_7510);
nor U9805 (N_9805,N_7215,N_7681);
nand U9806 (N_9806,N_7880,N_7575);
or U9807 (N_9807,N_6212,N_6651);
nand U9808 (N_9808,N_7217,N_6278);
nand U9809 (N_9809,N_6956,N_6459);
nand U9810 (N_9810,N_7670,N_6306);
and U9811 (N_9811,N_6566,N_7309);
and U9812 (N_9812,N_7511,N_6876);
and U9813 (N_9813,N_6673,N_7621);
or U9814 (N_9814,N_7875,N_7235);
and U9815 (N_9815,N_7412,N_6299);
and U9816 (N_9816,N_7570,N_7534);
nand U9817 (N_9817,N_7720,N_7641);
nand U9818 (N_9818,N_7693,N_7155);
and U9819 (N_9819,N_6315,N_6959);
nor U9820 (N_9820,N_7512,N_6421);
nor U9821 (N_9821,N_6225,N_6221);
nand U9822 (N_9822,N_7267,N_7055);
or U9823 (N_9823,N_7395,N_6321);
nand U9824 (N_9824,N_7450,N_7231);
or U9825 (N_9825,N_7346,N_6491);
nand U9826 (N_9826,N_6925,N_6710);
or U9827 (N_9827,N_7463,N_7156);
or U9828 (N_9828,N_6075,N_6932);
and U9829 (N_9829,N_7356,N_6350);
nor U9830 (N_9830,N_6144,N_6907);
xor U9831 (N_9831,N_7023,N_6358);
or U9832 (N_9832,N_7812,N_6237);
and U9833 (N_9833,N_6499,N_6911);
and U9834 (N_9834,N_6595,N_7664);
or U9835 (N_9835,N_6917,N_6359);
and U9836 (N_9836,N_6717,N_7320);
or U9837 (N_9837,N_7331,N_6718);
or U9838 (N_9838,N_7131,N_6093);
or U9839 (N_9839,N_7725,N_7259);
and U9840 (N_9840,N_7984,N_6057);
nor U9841 (N_9841,N_7197,N_6898);
and U9842 (N_9842,N_7267,N_6144);
and U9843 (N_9843,N_7581,N_7343);
nor U9844 (N_9844,N_6225,N_6837);
or U9845 (N_9845,N_7284,N_6184);
nand U9846 (N_9846,N_7864,N_7039);
or U9847 (N_9847,N_7379,N_7793);
nand U9848 (N_9848,N_7634,N_6751);
and U9849 (N_9849,N_6254,N_6558);
nand U9850 (N_9850,N_6922,N_7500);
and U9851 (N_9851,N_6822,N_7440);
or U9852 (N_9852,N_7407,N_6931);
nand U9853 (N_9853,N_7290,N_7144);
and U9854 (N_9854,N_6596,N_6666);
and U9855 (N_9855,N_7410,N_7896);
nand U9856 (N_9856,N_7665,N_6040);
nor U9857 (N_9857,N_7740,N_6024);
or U9858 (N_9858,N_6154,N_7163);
nand U9859 (N_9859,N_7111,N_6241);
and U9860 (N_9860,N_6121,N_7482);
or U9861 (N_9861,N_7661,N_6882);
nor U9862 (N_9862,N_7578,N_7277);
nand U9863 (N_9863,N_6583,N_7708);
nor U9864 (N_9864,N_6540,N_7282);
nor U9865 (N_9865,N_6290,N_7016);
and U9866 (N_9866,N_6479,N_6605);
nor U9867 (N_9867,N_7295,N_7869);
and U9868 (N_9868,N_7793,N_7331);
nor U9869 (N_9869,N_6373,N_7957);
nor U9870 (N_9870,N_7714,N_7397);
nand U9871 (N_9871,N_6207,N_6661);
or U9872 (N_9872,N_7032,N_6802);
nor U9873 (N_9873,N_7602,N_6528);
xor U9874 (N_9874,N_7803,N_6980);
nand U9875 (N_9875,N_7177,N_7765);
and U9876 (N_9876,N_7188,N_7939);
and U9877 (N_9877,N_7024,N_7671);
and U9878 (N_9878,N_7511,N_7868);
or U9879 (N_9879,N_6441,N_6515);
and U9880 (N_9880,N_7666,N_6160);
nand U9881 (N_9881,N_6195,N_7273);
nor U9882 (N_9882,N_7221,N_6046);
nand U9883 (N_9883,N_7881,N_6132);
nand U9884 (N_9884,N_6509,N_6612);
nand U9885 (N_9885,N_7486,N_6410);
nor U9886 (N_9886,N_6672,N_7739);
and U9887 (N_9887,N_6099,N_7253);
or U9888 (N_9888,N_7197,N_6186);
and U9889 (N_9889,N_6419,N_6597);
nor U9890 (N_9890,N_7288,N_7093);
or U9891 (N_9891,N_6732,N_6358);
nand U9892 (N_9892,N_6094,N_6304);
or U9893 (N_9893,N_7173,N_6616);
nor U9894 (N_9894,N_7148,N_7459);
nor U9895 (N_9895,N_6173,N_6149);
nor U9896 (N_9896,N_6255,N_6391);
and U9897 (N_9897,N_6037,N_7855);
nand U9898 (N_9898,N_7685,N_6333);
or U9899 (N_9899,N_6227,N_6317);
or U9900 (N_9900,N_7562,N_6612);
and U9901 (N_9901,N_7648,N_7095);
and U9902 (N_9902,N_7082,N_6418);
nor U9903 (N_9903,N_7514,N_6886);
or U9904 (N_9904,N_6090,N_7122);
and U9905 (N_9905,N_7318,N_6047);
or U9906 (N_9906,N_6214,N_7202);
or U9907 (N_9907,N_6845,N_6464);
or U9908 (N_9908,N_6771,N_7470);
or U9909 (N_9909,N_7664,N_6736);
nor U9910 (N_9910,N_6022,N_7596);
nand U9911 (N_9911,N_7882,N_6368);
nor U9912 (N_9912,N_7197,N_7575);
nor U9913 (N_9913,N_7398,N_7541);
and U9914 (N_9914,N_6583,N_6291);
nand U9915 (N_9915,N_7167,N_6838);
nand U9916 (N_9916,N_7800,N_6890);
nor U9917 (N_9917,N_6961,N_7215);
nand U9918 (N_9918,N_7110,N_6882);
nand U9919 (N_9919,N_7734,N_6455);
or U9920 (N_9920,N_6005,N_6715);
nor U9921 (N_9921,N_7924,N_7489);
nand U9922 (N_9922,N_7848,N_6771);
nand U9923 (N_9923,N_7849,N_7505);
or U9924 (N_9924,N_7263,N_6562);
nor U9925 (N_9925,N_7066,N_6855);
or U9926 (N_9926,N_7267,N_7339);
nand U9927 (N_9927,N_6341,N_7124);
nand U9928 (N_9928,N_6450,N_6773);
nor U9929 (N_9929,N_6343,N_6011);
or U9930 (N_9930,N_6569,N_7308);
and U9931 (N_9931,N_7973,N_7594);
and U9932 (N_9932,N_6483,N_7278);
nor U9933 (N_9933,N_7374,N_7539);
nand U9934 (N_9934,N_6117,N_7077);
nand U9935 (N_9935,N_7641,N_6760);
and U9936 (N_9936,N_6950,N_6269);
nand U9937 (N_9937,N_6836,N_6656);
and U9938 (N_9938,N_6126,N_7366);
nor U9939 (N_9939,N_7006,N_6927);
or U9940 (N_9940,N_7816,N_7279);
or U9941 (N_9941,N_6551,N_7526);
nor U9942 (N_9942,N_7198,N_7818);
or U9943 (N_9943,N_6241,N_7889);
nor U9944 (N_9944,N_6061,N_7061);
nor U9945 (N_9945,N_7692,N_6269);
and U9946 (N_9946,N_7404,N_6758);
nand U9947 (N_9947,N_7489,N_6160);
nand U9948 (N_9948,N_7166,N_7429);
nand U9949 (N_9949,N_7646,N_6612);
nor U9950 (N_9950,N_6060,N_7153);
or U9951 (N_9951,N_6662,N_6010);
and U9952 (N_9952,N_6790,N_6714);
and U9953 (N_9953,N_7403,N_7394);
nand U9954 (N_9954,N_6181,N_6715);
or U9955 (N_9955,N_7057,N_6872);
and U9956 (N_9956,N_6266,N_7636);
or U9957 (N_9957,N_7861,N_6706);
and U9958 (N_9958,N_7594,N_7643);
nor U9959 (N_9959,N_6054,N_7825);
nor U9960 (N_9960,N_6949,N_7352);
and U9961 (N_9961,N_6473,N_7885);
or U9962 (N_9962,N_7205,N_7924);
or U9963 (N_9963,N_6331,N_7255);
nand U9964 (N_9964,N_7594,N_7881);
nor U9965 (N_9965,N_7207,N_7833);
nor U9966 (N_9966,N_6536,N_7887);
and U9967 (N_9967,N_6598,N_6039);
or U9968 (N_9968,N_7353,N_6588);
or U9969 (N_9969,N_6396,N_7922);
nand U9970 (N_9970,N_6331,N_7881);
nand U9971 (N_9971,N_6904,N_7379);
or U9972 (N_9972,N_6042,N_7455);
nand U9973 (N_9973,N_6367,N_6342);
and U9974 (N_9974,N_7230,N_7083);
nor U9975 (N_9975,N_6018,N_6425);
nand U9976 (N_9976,N_6308,N_7905);
and U9977 (N_9977,N_6071,N_6971);
nor U9978 (N_9978,N_6882,N_7274);
or U9979 (N_9979,N_7149,N_7834);
nand U9980 (N_9980,N_7505,N_6198);
or U9981 (N_9981,N_6441,N_6895);
and U9982 (N_9982,N_6176,N_7432);
xnor U9983 (N_9983,N_6594,N_6060);
and U9984 (N_9984,N_6896,N_6950);
nor U9985 (N_9985,N_7017,N_6650);
nor U9986 (N_9986,N_7536,N_6613);
and U9987 (N_9987,N_6758,N_7324);
and U9988 (N_9988,N_6126,N_7928);
nor U9989 (N_9989,N_7256,N_7991);
xor U9990 (N_9990,N_7602,N_6539);
nor U9991 (N_9991,N_7046,N_7923);
nand U9992 (N_9992,N_6363,N_7981);
nand U9993 (N_9993,N_7993,N_6278);
and U9994 (N_9994,N_6870,N_7886);
nand U9995 (N_9995,N_7976,N_7731);
nor U9996 (N_9996,N_6867,N_7297);
or U9997 (N_9997,N_7105,N_6264);
or U9998 (N_9998,N_7636,N_7972);
nand U9999 (N_9999,N_7030,N_6383);
and UO_0 (O_0,N_9480,N_8809);
nand UO_1 (O_1,N_8208,N_8826);
nor UO_2 (O_2,N_8403,N_9322);
nand UO_3 (O_3,N_8358,N_8005);
or UO_4 (O_4,N_9460,N_9061);
or UO_5 (O_5,N_9450,N_9409);
or UO_6 (O_6,N_8489,N_9751);
and UO_7 (O_7,N_9295,N_9729);
and UO_8 (O_8,N_8877,N_9581);
xor UO_9 (O_9,N_8598,N_9529);
or UO_10 (O_10,N_9445,N_9973);
and UO_11 (O_11,N_9692,N_9411);
or UO_12 (O_12,N_8028,N_8189);
and UO_13 (O_13,N_9434,N_9586);
nor UO_14 (O_14,N_8265,N_9668);
or UO_15 (O_15,N_9827,N_8769);
or UO_16 (O_16,N_8740,N_9536);
nor UO_17 (O_17,N_8046,N_8052);
xor UO_18 (O_18,N_8402,N_9300);
or UO_19 (O_19,N_8612,N_8931);
nor UO_20 (O_20,N_9404,N_8716);
nor UO_21 (O_21,N_8406,N_8920);
nor UO_22 (O_22,N_9190,N_8311);
and UO_23 (O_23,N_8910,N_8272);
and UO_24 (O_24,N_8602,N_8805);
nor UO_25 (O_25,N_8381,N_8034);
nor UO_26 (O_26,N_9792,N_9033);
and UO_27 (O_27,N_8230,N_8173);
nand UO_28 (O_28,N_8971,N_8714);
or UO_29 (O_29,N_9548,N_9654);
and UO_30 (O_30,N_8970,N_8419);
nand UO_31 (O_31,N_8421,N_8625);
nand UO_32 (O_32,N_9745,N_9845);
or UO_33 (O_33,N_8220,N_8290);
and UO_34 (O_34,N_9022,N_9169);
nor UO_35 (O_35,N_8478,N_9876);
or UO_36 (O_36,N_9140,N_9379);
nor UO_37 (O_37,N_8552,N_9209);
or UO_38 (O_38,N_9329,N_9262);
or UO_39 (O_39,N_9429,N_8778);
and UO_40 (O_40,N_8460,N_9086);
or UO_41 (O_41,N_8369,N_9834);
or UO_42 (O_42,N_8747,N_9989);
nor UO_43 (O_43,N_8312,N_9687);
or UO_44 (O_44,N_8422,N_8453);
nand UO_45 (O_45,N_8448,N_9184);
and UO_46 (O_46,N_9165,N_9437);
nand UO_47 (O_47,N_8673,N_8177);
nor UO_48 (O_48,N_9981,N_8913);
nand UO_49 (O_49,N_9503,N_8349);
and UO_50 (O_50,N_8770,N_9921);
nand UO_51 (O_51,N_8065,N_9511);
or UO_52 (O_52,N_9475,N_9768);
or UO_53 (O_53,N_9796,N_8309);
nand UO_54 (O_54,N_8631,N_8895);
nand UO_55 (O_55,N_9131,N_9068);
and UO_56 (O_56,N_8346,N_8860);
nor UO_57 (O_57,N_8500,N_8167);
and UO_58 (O_58,N_8694,N_9621);
nor UO_59 (O_59,N_8325,N_9953);
nand UO_60 (O_60,N_8206,N_8827);
nand UO_61 (O_61,N_8976,N_8952);
and UO_62 (O_62,N_9552,N_8670);
nor UO_63 (O_63,N_8808,N_9594);
nor UO_64 (O_64,N_8532,N_9831);
nand UO_65 (O_65,N_9025,N_9324);
or UO_66 (O_66,N_8343,N_8451);
and UO_67 (O_67,N_9613,N_8266);
nand UO_68 (O_68,N_9498,N_9361);
or UO_69 (O_69,N_8323,N_9484);
or UO_70 (O_70,N_9378,N_8975);
or UO_71 (O_71,N_8407,N_9323);
nor UO_72 (O_72,N_8722,N_9854);
nor UO_73 (O_73,N_8076,N_8530);
nor UO_74 (O_74,N_8519,N_8704);
or UO_75 (O_75,N_8313,N_9234);
nor UO_76 (O_76,N_9114,N_9462);
and UO_77 (O_77,N_9570,N_8446);
nand UO_78 (O_78,N_9542,N_8216);
nor UO_79 (O_79,N_9960,N_9943);
and UO_80 (O_80,N_9384,N_9757);
nand UO_81 (O_81,N_8368,N_9312);
or UO_82 (O_82,N_8118,N_9189);
nor UO_83 (O_83,N_8472,N_8004);
or UO_84 (O_84,N_9043,N_9363);
nor UO_85 (O_85,N_9680,N_8745);
nor UO_86 (O_86,N_8661,N_8329);
or UO_87 (O_87,N_8521,N_8505);
and UO_88 (O_88,N_8541,N_8856);
nor UO_89 (O_89,N_8068,N_8980);
nand UO_90 (O_90,N_8558,N_9439);
or UO_91 (O_91,N_8893,N_8674);
nor UO_92 (O_92,N_9377,N_8752);
and UO_93 (O_93,N_8955,N_9399);
nor UO_94 (O_94,N_8319,N_9206);
nand UO_95 (O_95,N_9521,N_9936);
nand UO_96 (O_96,N_9789,N_9365);
and UO_97 (O_97,N_9269,N_9400);
and UO_98 (O_98,N_9065,N_9701);
and UO_99 (O_99,N_9056,N_9698);
or UO_100 (O_100,N_8385,N_9993);
nor UO_101 (O_101,N_8863,N_8619);
nor UO_102 (O_102,N_8081,N_8512);
nand UO_103 (O_103,N_9583,N_9601);
or UO_104 (O_104,N_9814,N_9125);
nand UO_105 (O_105,N_9546,N_9351);
nand UO_106 (O_106,N_8850,N_9898);
or UO_107 (O_107,N_8760,N_8433);
and UO_108 (O_108,N_9470,N_9500);
nor UO_109 (O_109,N_9622,N_8458);
nand UO_110 (O_110,N_8449,N_8550);
nand UO_111 (O_111,N_9020,N_9087);
nand UO_112 (O_112,N_9275,N_8018);
nor UO_113 (O_113,N_8450,N_8679);
or UO_114 (O_114,N_8183,N_9571);
or UO_115 (O_115,N_8969,N_9011);
nor UO_116 (O_116,N_8599,N_9778);
nand UO_117 (O_117,N_9813,N_8843);
nand UO_118 (O_118,N_8972,N_9651);
or UO_119 (O_119,N_9890,N_9906);
xor UO_120 (O_120,N_8390,N_9971);
or UO_121 (O_121,N_9938,N_8200);
nand UO_122 (O_122,N_8494,N_9468);
and UO_123 (O_123,N_9016,N_9103);
or UO_124 (O_124,N_9655,N_8439);
and UO_125 (O_125,N_9994,N_8201);
nor UO_126 (O_126,N_8398,N_9427);
or UO_127 (O_127,N_9862,N_8776);
and UO_128 (O_128,N_8795,N_9839);
nor UO_129 (O_129,N_9251,N_9504);
nand UO_130 (O_130,N_8732,N_8941);
nand UO_131 (O_131,N_9390,N_9804);
or UO_132 (O_132,N_9072,N_9049);
xor UO_133 (O_133,N_9567,N_8538);
nand UO_134 (O_134,N_9910,N_8264);
nor UO_135 (O_135,N_9802,N_9079);
and UO_136 (O_136,N_9382,N_9539);
or UO_137 (O_137,N_8921,N_8681);
nand UO_138 (O_138,N_9634,N_9332);
and UO_139 (O_139,N_8019,N_9222);
or UO_140 (O_140,N_9638,N_8480);
or UO_141 (O_141,N_9937,N_8288);
nor UO_142 (O_142,N_8090,N_8383);
or UO_143 (O_143,N_9284,N_8693);
and UO_144 (O_144,N_8603,N_8730);
nand UO_145 (O_145,N_9666,N_9782);
and UO_146 (O_146,N_9076,N_9481);
nand UO_147 (O_147,N_8964,N_9465);
nor UO_148 (O_148,N_9502,N_8592);
and UO_149 (O_149,N_9391,N_8687);
or UO_150 (O_150,N_9522,N_9343);
or UO_151 (O_151,N_8900,N_8321);
nand UO_152 (O_152,N_8263,N_8262);
nor UO_153 (O_153,N_8361,N_8959);
or UO_154 (O_154,N_9584,N_9194);
nor UO_155 (O_155,N_9878,N_8581);
nor UO_156 (O_156,N_8531,N_9341);
or UO_157 (O_157,N_9841,N_9760);
or UO_158 (O_158,N_9950,N_9408);
nor UO_159 (O_159,N_8966,N_9909);
and UO_160 (O_160,N_8902,N_9501);
nor UO_161 (O_161,N_8788,N_8036);
nand UO_162 (O_162,N_8217,N_8981);
or UO_163 (O_163,N_9210,N_8838);
nand UO_164 (O_164,N_9456,N_9821);
nor UO_165 (O_165,N_9448,N_9014);
xor UO_166 (O_166,N_9725,N_8481);
and UO_167 (O_167,N_9574,N_9505);
or UO_168 (O_168,N_9164,N_8804);
nor UO_169 (O_169,N_9975,N_8585);
and UO_170 (O_170,N_9733,N_8994);
and UO_171 (O_171,N_8654,N_8237);
or UO_172 (O_172,N_9105,N_8360);
nand UO_173 (O_173,N_8040,N_9315);
nand UO_174 (O_174,N_9035,N_8066);
nor UO_175 (O_175,N_9766,N_9191);
nand UO_176 (O_176,N_9660,N_8491);
or UO_177 (O_177,N_9268,N_8096);
or UO_178 (O_178,N_8250,N_8935);
or UO_179 (O_179,N_9737,N_8767);
or UO_180 (O_180,N_8803,N_9967);
or UO_181 (O_181,N_9815,N_9220);
nor UO_182 (O_182,N_8409,N_9566);
nor UO_183 (O_183,N_8437,N_8465);
or UO_184 (O_184,N_9828,N_8961);
and UO_185 (O_185,N_9888,N_8748);
nand UO_186 (O_186,N_9591,N_8866);
and UO_187 (O_187,N_8009,N_9922);
and UO_188 (O_188,N_8033,N_8156);
or UO_189 (O_189,N_8001,N_8587);
and UO_190 (O_190,N_9182,N_9435);
nor UO_191 (O_191,N_8022,N_9700);
or UO_192 (O_192,N_8088,N_9846);
nand UO_193 (O_193,N_9029,N_8092);
and UO_194 (O_194,N_8639,N_9672);
and UO_195 (O_195,N_9098,N_9678);
and UO_196 (O_196,N_8534,N_9368);
nor UO_197 (O_197,N_9469,N_9127);
nand UO_198 (O_198,N_8873,N_9875);
nand UO_199 (O_199,N_9362,N_9818);
or UO_200 (O_200,N_9036,N_8401);
or UO_201 (O_201,N_8241,N_9152);
or UO_202 (O_202,N_8239,N_8306);
or UO_203 (O_203,N_9181,N_8663);
and UO_204 (O_204,N_9259,N_9402);
xnor UO_205 (O_205,N_8726,N_9139);
and UO_206 (O_206,N_8392,N_8777);
or UO_207 (O_207,N_9482,N_9197);
or UO_208 (O_208,N_9096,N_8622);
nand UO_209 (O_209,N_8172,N_8298);
nand UO_210 (O_210,N_8299,N_8199);
and UO_211 (O_211,N_8915,N_9320);
and UO_212 (O_212,N_8245,N_8436);
or UO_213 (O_213,N_8024,N_8378);
or UO_214 (O_214,N_8037,N_9467);
and UO_215 (O_215,N_8141,N_8317);
and UO_216 (O_216,N_8578,N_9732);
nand UO_217 (O_217,N_8048,N_9855);
and UO_218 (O_218,N_8743,N_9483);
or UO_219 (O_219,N_8934,N_9394);
or UO_220 (O_220,N_8261,N_8563);
nor UO_221 (O_221,N_9596,N_8193);
nor UO_222 (O_222,N_8675,N_8107);
nand UO_223 (O_223,N_8720,N_9649);
or UO_224 (O_224,N_9419,N_8819);
or UO_225 (O_225,N_9556,N_8644);
or UO_226 (O_226,N_8852,N_9941);
nand UO_227 (O_227,N_9066,N_9119);
nor UO_228 (O_228,N_9604,N_9866);
nor UO_229 (O_229,N_9565,N_9280);
or UO_230 (O_230,N_9297,N_9199);
nand UO_231 (O_231,N_8365,N_9298);
nand UO_232 (O_232,N_9137,N_9940);
nor UO_233 (O_233,N_8737,N_9389);
nor UO_234 (O_234,N_9147,N_8468);
or UO_235 (O_235,N_9348,N_9748);
nand UO_236 (O_236,N_8949,N_9924);
and UO_237 (O_237,N_9200,N_9364);
nor UO_238 (O_238,N_9812,N_8601);
or UO_239 (O_239,N_8331,N_8353);
or UO_240 (O_240,N_8648,N_9099);
nor UO_241 (O_241,N_8229,N_9620);
nand UO_242 (O_242,N_9790,N_9058);
xnor UO_243 (O_243,N_8565,N_9245);
and UO_244 (O_244,N_9693,N_9090);
nor UO_245 (O_245,N_8984,N_9532);
and UO_246 (O_246,N_9405,N_8228);
nand UO_247 (O_247,N_9126,N_9699);
nand UO_248 (O_248,N_9830,N_9585);
or UO_249 (O_249,N_8702,N_8665);
nor UO_250 (O_250,N_8080,N_9533);
or UO_251 (O_251,N_8680,N_9681);
or UO_252 (O_252,N_9965,N_9142);
nor UO_253 (O_253,N_9204,N_9861);
and UO_254 (O_254,N_9679,N_9537);
nand UO_255 (O_255,N_8462,N_9289);
and UO_256 (O_256,N_8339,N_8698);
nand UO_257 (O_257,N_9101,N_8425);
nand UO_258 (O_258,N_8870,N_8222);
and UO_259 (O_259,N_9488,N_9263);
or UO_260 (O_260,N_8963,N_9321);
or UO_261 (O_261,N_9715,N_9212);
or UO_262 (O_262,N_8127,N_9746);
or UO_263 (O_263,N_8049,N_8432);
and UO_264 (O_264,N_9826,N_9602);
xnor UO_265 (O_265,N_9920,N_8047);
nor UO_266 (O_266,N_9214,N_9637);
or UO_267 (O_267,N_9352,N_8858);
nand UO_268 (O_268,N_9852,N_8571);
nand UO_269 (O_269,N_9835,N_9392);
nand UO_270 (O_270,N_8053,N_8911);
xor UO_271 (O_271,N_9293,N_8463);
or UO_272 (O_272,N_8103,N_9358);
nor UO_273 (O_273,N_9625,N_8705);
nor UO_274 (O_274,N_9155,N_8937);
nand UO_275 (O_275,N_8474,N_8023);
and UO_276 (O_276,N_8627,N_8170);
or UO_277 (O_277,N_8800,N_9454);
or UO_278 (O_278,N_9247,N_8636);
and UO_279 (O_279,N_8916,N_8525);
and UO_280 (O_280,N_8557,N_9230);
nand UO_281 (O_281,N_8798,N_8912);
nand UO_282 (O_282,N_9547,N_8744);
nand UO_283 (O_283,N_9781,N_8651);
and UO_284 (O_284,N_8123,N_8613);
nand UO_285 (O_285,N_8628,N_9153);
nor UO_286 (O_286,N_9978,N_8851);
and UO_287 (O_287,N_8404,N_8171);
nand UO_288 (O_288,N_9487,N_9253);
nand UO_289 (O_289,N_8485,N_9277);
and UO_290 (O_290,N_9398,N_8834);
and UO_291 (O_291,N_8799,N_8344);
nand UO_292 (O_292,N_8828,N_8400);
nor UO_293 (O_293,N_9684,N_9947);
nor UO_294 (O_294,N_8287,N_9990);
nand UO_295 (O_295,N_8362,N_8182);
nor UO_296 (O_296,N_9935,N_9407);
nand UO_297 (O_297,N_9325,N_8204);
or UO_298 (O_298,N_8932,N_9463);
nor UO_299 (O_299,N_9162,N_9641);
and UO_300 (O_300,N_8464,N_9085);
and UO_301 (O_301,N_9051,N_8946);
or UO_302 (O_302,N_8888,N_8987);
nand UO_303 (O_303,N_8078,N_9929);
xnor UO_304 (O_304,N_9755,N_8492);
or UO_305 (O_305,N_9592,N_9357);
nor UO_306 (O_306,N_9446,N_8836);
and UO_307 (O_307,N_8185,N_9636);
nand UO_308 (O_308,N_8825,N_8475);
nor UO_309 (O_309,N_8985,N_8638);
and UO_310 (O_310,N_9461,N_8653);
nor UO_311 (O_311,N_9492,N_9851);
and UO_312 (O_312,N_8377,N_8611);
nand UO_313 (O_313,N_9572,N_8275);
nor UO_314 (O_314,N_9605,N_8350);
and UO_315 (O_315,N_8035,N_8363);
nand UO_316 (O_316,N_8909,N_8671);
nor UO_317 (O_317,N_9396,N_8389);
and UO_318 (O_318,N_9044,N_9884);
xnor UO_319 (O_319,N_8922,N_9514);
nor UO_320 (O_320,N_9261,N_9508);
and UO_321 (O_321,N_8929,N_9472);
or UO_322 (O_322,N_8499,N_8948);
nor UO_323 (O_323,N_9904,N_9939);
nor UO_324 (O_324,N_8807,N_8067);
xor UO_325 (O_325,N_9414,N_9669);
nand UO_326 (O_326,N_9173,N_9863);
and UO_327 (O_327,N_9186,N_8771);
nand UO_328 (O_328,N_9676,N_8724);
nor UO_329 (O_329,N_9490,N_9728);
nor UO_330 (O_330,N_8597,N_8108);
or UO_331 (O_331,N_8396,N_8278);
and UO_332 (O_332,N_9640,N_9741);
or UO_333 (O_333,N_8027,N_8723);
and UO_334 (O_334,N_8128,N_8927);
or UO_335 (O_335,N_9853,N_9896);
nor UO_336 (O_336,N_8149,N_9930);
nand UO_337 (O_337,N_9850,N_9375);
and UO_338 (O_338,N_9696,N_9318);
or UO_339 (O_339,N_8820,N_8695);
or UO_340 (O_340,N_9403,N_8225);
or UO_341 (O_341,N_9913,N_9296);
and UO_342 (O_342,N_8608,N_8021);
nand UO_343 (O_343,N_8551,N_9387);
and UO_344 (O_344,N_9968,N_9969);
nand UO_345 (O_345,N_8178,N_9758);
or UO_346 (O_346,N_9337,N_8546);
nor UO_347 (O_347,N_8996,N_8509);
nand UO_348 (O_348,N_9833,N_8274);
nor UO_349 (O_349,N_8781,N_8372);
nand UO_350 (O_350,N_8044,N_8332);
nor UO_351 (O_351,N_9150,N_9734);
nor UO_352 (O_352,N_9540,N_8031);
or UO_353 (O_353,N_9276,N_8837);
or UO_354 (O_354,N_9769,N_8712);
nand UO_355 (O_355,N_9037,N_8624);
nand UO_356 (O_356,N_9860,N_9559);
nor UO_357 (O_357,N_8082,N_8190);
or UO_358 (O_358,N_9095,N_9717);
or UO_359 (O_359,N_8561,N_9485);
xor UO_360 (O_360,N_8003,N_8466);
and UO_361 (O_361,N_9371,N_8739);
and UO_362 (O_362,N_8874,N_9639);
or UO_363 (O_363,N_9122,N_8337);
nor UO_364 (O_364,N_8131,N_9120);
or UO_365 (O_365,N_9612,N_8430);
nor UO_366 (O_366,N_9144,N_8568);
nand UO_367 (O_367,N_8297,N_9129);
xnor UO_368 (O_368,N_8169,N_9067);
or UO_369 (O_369,N_9388,N_8901);
and UO_370 (O_370,N_8424,N_8232);
or UO_371 (O_371,N_8709,N_9213);
nor UO_372 (O_372,N_9339,N_8459);
nor UO_373 (O_373,N_9635,N_8366);
nor UO_374 (O_374,N_9376,N_9740);
nand UO_375 (O_375,N_9980,N_8226);
nand UO_376 (O_376,N_8057,N_8861);
nor UO_377 (O_377,N_9349,N_9397);
xnor UO_378 (O_378,N_8584,N_9530);
or UO_379 (O_379,N_9082,N_9359);
and UO_380 (O_380,N_9523,N_8655);
nor UO_381 (O_381,N_8577,N_9946);
nand UO_382 (O_382,N_8320,N_8951);
and UO_383 (O_383,N_8833,N_8741);
or UO_384 (O_384,N_9415,N_8054);
and UO_385 (O_385,N_8559,N_8117);
nand UO_386 (O_386,N_9026,N_8701);
and UO_387 (O_387,N_9515,N_8634);
nand UO_388 (O_388,N_9772,N_9034);
nand UO_389 (O_389,N_9545,N_9242);
nor UO_390 (O_390,N_9690,N_8017);
nand UO_391 (O_391,N_9233,N_8356);
nand UO_392 (O_392,N_8632,N_9535);
nor UO_393 (O_393,N_8209,N_9867);
or UO_394 (O_394,N_9458,N_9235);
nand UO_395 (O_395,N_9319,N_9974);
nand UO_396 (O_396,N_9996,N_9008);
nor UO_397 (O_397,N_9653,N_8277);
nand UO_398 (O_398,N_8642,N_8233);
or UO_399 (O_399,N_9202,N_8097);
or UO_400 (O_400,N_9629,N_9966);
xor UO_401 (O_401,N_9616,N_9917);
nand UO_402 (O_402,N_9154,N_9116);
and UO_403 (O_403,N_9691,N_8965);
nand UO_404 (O_404,N_9976,N_8796);
or UO_405 (O_405,N_9624,N_8881);
nor UO_406 (O_406,N_9039,N_8184);
and UO_407 (O_407,N_9603,N_8471);
or UO_408 (O_408,N_9774,N_9987);
and UO_409 (O_409,N_8734,N_8148);
and UO_410 (O_410,N_8426,N_8305);
nand UO_411 (O_411,N_8574,N_9109);
and UO_412 (O_412,N_8609,N_9983);
or UO_413 (O_413,N_9440,N_9767);
nor UO_414 (O_414,N_9031,N_8939);
or UO_415 (O_415,N_8371,N_9626);
and UO_416 (O_416,N_8676,N_8570);
nor UO_417 (O_417,N_8782,N_8573);
nand UO_418 (O_418,N_8605,N_8684);
nand UO_419 (O_419,N_8572,N_9988);
and UO_420 (O_420,N_8301,N_8536);
and UO_421 (O_421,N_8643,N_8295);
nand UO_422 (O_422,N_9112,N_9704);
or UO_423 (O_423,N_8982,N_9628);
and UO_424 (O_424,N_8496,N_8983);
nor UO_425 (O_425,N_8514,N_9714);
nor UO_426 (O_426,N_8063,N_8077);
or UO_427 (O_427,N_9158,N_8696);
and UO_428 (O_428,N_9274,N_9278);
and UO_429 (O_429,N_8308,N_8844);
and UO_430 (O_430,N_8553,N_9723);
nand UO_431 (O_431,N_9283,N_8318);
or UO_432 (O_432,N_9005,N_8213);
and UO_433 (O_433,N_8215,N_9097);
or UO_434 (O_434,N_9385,N_9306);
or UO_435 (O_435,N_9174,N_9393);
or UO_436 (O_436,N_8115,N_9914);
or UO_437 (O_437,N_9576,N_8083);
or UO_438 (O_438,N_8223,N_8691);
or UO_439 (O_439,N_8212,N_9133);
xnor UO_440 (O_440,N_9719,N_9136);
nand UO_441 (O_441,N_9107,N_9657);
and UO_442 (O_442,N_9824,N_8510);
nand UO_443 (O_443,N_8100,N_8682);
nor UO_444 (O_444,N_9731,N_8391);
nor UO_445 (O_445,N_8977,N_9958);
nand UO_446 (O_446,N_9708,N_8810);
nand UO_447 (O_447,N_9355,N_9104);
and UO_448 (O_448,N_8159,N_8801);
xnor UO_449 (O_449,N_9809,N_9201);
or UO_450 (O_450,N_8099,N_9223);
and UO_451 (O_451,N_8854,N_9370);
or UO_452 (O_452,N_8236,N_8150);
nor UO_453 (O_453,N_9840,N_8015);
and UO_454 (O_454,N_8418,N_9178);
nand UO_455 (O_455,N_9911,N_9631);
or UO_456 (O_456,N_8629,N_8785);
and UO_457 (O_457,N_9239,N_9023);
nand UO_458 (O_458,N_9868,N_9281);
nand UO_459 (O_459,N_8956,N_8630);
or UO_460 (O_460,N_9004,N_9009);
nor UO_461 (O_461,N_9892,N_9926);
nand UO_462 (O_462,N_9425,N_9143);
nand UO_463 (O_463,N_9557,N_8990);
nand UO_464 (O_464,N_8566,N_9054);
nand UO_465 (O_465,N_9942,N_9963);
xor UO_466 (O_466,N_8058,N_9015);
nand UO_467 (O_467,N_9648,N_9286);
nand UO_468 (O_468,N_8174,N_8635);
and UO_469 (O_469,N_8919,N_8667);
and UO_470 (O_470,N_8252,N_8069);
and UO_471 (O_471,N_9443,N_8750);
or UO_472 (O_472,N_8615,N_8163);
or UO_473 (O_473,N_8853,N_8125);
and UO_474 (O_474,N_8614,N_8756);
nand UO_475 (O_475,N_8754,N_8379);
nand UO_476 (O_476,N_8555,N_9519);
nor UO_477 (O_477,N_8268,N_8410);
or UO_478 (O_478,N_9771,N_9619);
or UO_479 (O_479,N_9611,N_8656);
or UO_480 (O_480,N_9919,N_8710);
and UO_481 (O_481,N_9527,N_8840);
nor UO_482 (O_482,N_9510,N_9724);
nand UO_483 (O_483,N_9476,N_9897);
or UO_484 (O_484,N_9334,N_9822);
or UO_485 (O_485,N_8428,N_8293);
and UO_486 (O_486,N_8657,N_8529);
nor UO_487 (O_487,N_8133,N_9811);
nand UO_488 (O_488,N_8195,N_9113);
and UO_489 (O_489,N_8084,N_9479);
and UO_490 (O_490,N_9736,N_9420);
and UO_491 (O_491,N_8452,N_9650);
and UO_492 (O_492,N_8070,N_8898);
xor UO_493 (O_493,N_8246,N_9730);
nand UO_494 (O_494,N_8122,N_8119);
and UO_495 (O_495,N_9588,N_8013);
nor UO_496 (O_496,N_8116,N_9360);
nand UO_497 (O_497,N_9806,N_9171);
and UO_498 (O_498,N_8388,N_8486);
nor UO_499 (O_499,N_9441,N_9160);
and UO_500 (O_500,N_9372,N_8936);
nor UO_501 (O_501,N_8445,N_9491);
and UO_502 (O_502,N_9671,N_9328);
or UO_503 (O_503,N_9264,N_9577);
or UO_504 (O_504,N_9549,N_8393);
or UO_505 (O_505,N_8590,N_9313);
nor UO_506 (O_506,N_9682,N_8593);
and UO_507 (O_507,N_8279,N_9123);
and UO_508 (O_508,N_9002,N_8417);
nor UO_509 (O_509,N_9340,N_8136);
nor UO_510 (O_510,N_9243,N_9383);
and UO_511 (O_511,N_8896,N_8940);
or UO_512 (O_512,N_8968,N_8958);
and UO_513 (O_513,N_9452,N_8073);
nand UO_514 (O_514,N_9260,N_8890);
and UO_515 (O_515,N_8658,N_9062);
nand UO_516 (O_516,N_8140,N_8580);
nand UO_517 (O_517,N_9052,N_8121);
nand UO_518 (O_518,N_9013,N_9436);
and UO_519 (O_519,N_9957,N_8506);
nor UO_520 (O_520,N_8690,N_9183);
nand UO_521 (O_521,N_8089,N_9664);
or UO_522 (O_522,N_9573,N_8556);
nand UO_523 (O_523,N_9907,N_8194);
or UO_524 (O_524,N_8025,N_9899);
or UO_525 (O_525,N_8364,N_8899);
or UO_526 (O_526,N_8386,N_8528);
nor UO_527 (O_527,N_8294,N_9513);
and UO_528 (O_528,N_9024,N_9000);
nand UO_529 (O_529,N_9785,N_8539);
or UO_530 (O_530,N_9817,N_9003);
and UO_531 (O_531,N_9721,N_9224);
or UO_532 (O_532,N_8677,N_9010);
nor UO_533 (O_533,N_8707,N_9894);
nand UO_534 (O_534,N_8259,N_9175);
or UO_535 (O_535,N_8729,N_8050);
nor UO_536 (O_536,N_9444,N_8280);
or UO_537 (O_537,N_8749,N_9722);
and UO_538 (O_538,N_9187,N_9045);
and UO_539 (O_539,N_8104,N_9028);
nor UO_540 (O_540,N_8649,N_8924);
nor UO_541 (O_541,N_8006,N_9335);
nor UO_542 (O_542,N_9949,N_8412);
or UO_543 (O_543,N_8868,N_9238);
or UO_544 (O_544,N_9972,N_8218);
nand UO_545 (O_545,N_8328,N_9232);
xnor UO_546 (O_546,N_8224,N_9538);
and UO_547 (O_547,N_8824,N_9857);
xor UO_548 (O_548,N_8882,N_8647);
nand UO_549 (O_549,N_8533,N_9918);
nand UO_550 (O_550,N_8095,N_9568);
and UO_551 (O_551,N_9083,N_8061);
or UO_552 (O_552,N_9266,N_9249);
nand UO_553 (O_553,N_9196,N_9810);
xnor UO_554 (O_554,N_8251,N_9793);
nor UO_555 (O_555,N_9218,N_8904);
nor UO_556 (O_556,N_8746,N_8012);
xor UO_557 (O_557,N_9132,N_9984);
nand UO_558 (O_558,N_9710,N_9327);
or UO_559 (O_559,N_8869,N_9674);
nor UO_560 (O_560,N_9630,N_9455);
nand UO_561 (O_561,N_8132,N_9354);
or UO_562 (O_562,N_8032,N_8269);
and UO_563 (O_563,N_9595,N_9659);
or UO_564 (O_564,N_9241,N_8457);
and UO_565 (O_565,N_9346,N_9686);
nor UO_566 (O_566,N_8508,N_8302);
nor UO_567 (O_567,N_8210,N_8646);
nor UO_568 (O_568,N_8456,N_9226);
nand UO_569 (O_569,N_8848,N_9718);
or UO_570 (O_570,N_8960,N_9254);
nand UO_571 (O_571,N_9551,N_9432);
nor UO_572 (O_572,N_9881,N_8908);
or UO_573 (O_573,N_8780,N_8316);
nor UO_574 (O_574,N_8235,N_9134);
and UO_575 (O_575,N_8993,N_8219);
or UO_576 (O_576,N_8461,N_8548);
nor UO_577 (O_577,N_9986,N_9074);
or UO_578 (O_578,N_8501,N_8124);
nor UO_579 (O_579,N_8887,N_8517);
or UO_580 (O_580,N_8692,N_9712);
nand UO_581 (O_581,N_8303,N_8764);
nand UO_582 (O_582,N_8490,N_9221);
nor UO_583 (O_583,N_9166,N_8079);
nor UO_584 (O_584,N_9331,N_8405);
nand UO_585 (O_585,N_9410,N_9786);
nor UO_586 (O_586,N_8014,N_9423);
and UO_587 (O_587,N_9027,N_9070);
nor UO_588 (O_588,N_9211,N_8055);
and UO_589 (O_589,N_9703,N_8664);
or UO_590 (O_590,N_8711,N_8340);
or UO_591 (O_591,N_9727,N_9229);
nand UO_592 (O_592,N_9598,N_9562);
nor UO_593 (O_593,N_8192,N_8165);
nand UO_594 (O_594,N_8718,N_8281);
or UO_595 (O_595,N_9453,N_9418);
and UO_596 (O_596,N_8637,N_8455);
nand UO_597 (O_597,N_9749,N_9257);
nand UO_598 (O_598,N_8821,N_8444);
nand UO_599 (O_599,N_8285,N_9705);
or UO_600 (O_600,N_9424,N_9739);
nand UO_601 (O_601,N_9520,N_9170);
or UO_602 (O_602,N_9227,N_9747);
or UO_603 (O_603,N_8060,N_8753);
or UO_604 (O_604,N_8144,N_8179);
nor UO_605 (O_605,N_9047,N_9645);
nor UO_606 (O_606,N_9270,N_9580);
nor UO_607 (O_607,N_8814,N_9784);
nand UO_608 (O_608,N_9761,N_8616);
nand UO_609 (O_609,N_8715,N_8020);
or UO_610 (O_610,N_9050,N_9999);
nor UO_611 (O_611,N_9889,N_9167);
nand UO_612 (O_612,N_8370,N_8375);
and UO_613 (O_613,N_8652,N_8242);
nand UO_614 (O_614,N_9954,N_9089);
nor UO_615 (O_615,N_9486,N_9891);
nor UO_616 (O_616,N_8026,N_9554);
or UO_617 (O_617,N_8540,N_9848);
and UO_618 (O_618,N_8113,N_8699);
and UO_619 (O_619,N_8947,N_9380);
and UO_620 (O_620,N_9964,N_9092);
nor UO_621 (O_621,N_8059,N_9555);
and UO_622 (O_622,N_9516,N_8668);
nor UO_623 (O_623,N_8085,N_9299);
nand UO_624 (O_624,N_9073,N_8816);
nor UO_625 (O_625,N_9466,N_8434);
or UO_626 (O_626,N_8045,N_9288);
and UO_627 (O_627,N_8091,N_8591);
nor UO_628 (O_628,N_8071,N_9135);
and UO_629 (O_629,N_8562,N_9271);
or UO_630 (O_630,N_9646,N_8633);
or UO_631 (O_631,N_9106,N_8011);
or UO_632 (O_632,N_8146,N_8479);
or UO_633 (O_633,N_8341,N_8575);
nor UO_634 (O_634,N_9720,N_8168);
nand UO_635 (O_635,N_8056,N_9302);
and UO_636 (O_636,N_8382,N_8271);
and UO_637 (O_637,N_9689,N_9317);
nor UO_638 (O_638,N_9311,N_8974);
and UO_639 (O_639,N_9148,N_9597);
nor UO_640 (O_640,N_8736,N_8074);
nor UO_641 (O_641,N_8891,N_9961);
and UO_642 (O_642,N_8495,N_8697);
nand UO_643 (O_643,N_8126,N_8016);
and UO_644 (O_644,N_8007,N_9869);
and UO_645 (O_645,N_8686,N_8162);
nand UO_646 (O_646,N_8243,N_8894);
xor UO_647 (O_647,N_9992,N_8596);
nand UO_648 (O_648,N_8867,N_8041);
and UO_649 (O_649,N_9912,N_8138);
nor UO_650 (O_650,N_8822,N_9159);
or UO_651 (O_651,N_8883,N_9041);
or UO_652 (O_652,N_9744,N_9735);
and UO_653 (O_653,N_8589,N_8157);
and UO_654 (O_654,N_9742,N_9244);
nor UO_655 (O_655,N_8504,N_9030);
nor UO_656 (O_656,N_8846,N_8830);
nor UO_657 (O_657,N_8440,N_8885);
nor UO_658 (O_658,N_9563,N_8010);
or UO_659 (O_659,N_8483,N_9798);
nor UO_660 (O_660,N_9198,N_9787);
nor UO_661 (O_661,N_8689,N_9477);
nor UO_662 (O_662,N_9895,N_9632);
or UO_663 (O_663,N_9932,N_9779);
nand UO_664 (O_664,N_8196,N_9303);
or UO_665 (O_665,N_9893,N_9803);
and UO_666 (O_666,N_8105,N_8997);
and UO_667 (O_667,N_8524,N_9373);
nand UO_668 (O_668,N_9697,N_9948);
nor UO_669 (O_669,N_9205,N_9195);
and UO_670 (O_670,N_9179,N_9820);
or UO_671 (O_671,N_8260,N_9428);
xnor UO_672 (O_672,N_8062,N_9808);
or UO_673 (O_673,N_8221,N_8258);
or UO_674 (O_674,N_8238,N_9995);
and UO_675 (O_675,N_9716,N_9188);
or UO_676 (O_676,N_8114,N_8477);
nor UO_677 (O_677,N_8988,N_8569);
nor UO_678 (O_678,N_8962,N_9623);
nand UO_679 (O_679,N_9561,N_8203);
and UO_680 (O_680,N_9763,N_9600);
and UO_681 (O_681,N_9108,N_8075);
nand UO_682 (O_682,N_9780,N_8286);
and UO_683 (O_683,N_9886,N_8527);
or UO_684 (O_684,N_9473,N_8583);
nor UO_685 (O_685,N_8153,N_9847);
or UO_686 (O_686,N_9381,N_9267);
and UO_687 (O_687,N_8234,N_9304);
nor UO_688 (O_688,N_9057,N_9240);
nand UO_689 (O_689,N_9908,N_9246);
nand UO_690 (O_690,N_9677,N_9055);
or UO_691 (O_691,N_9447,N_8064);
or UO_692 (O_692,N_9608,N_8797);
and UO_693 (O_693,N_8249,N_8979);
and UO_694 (O_694,N_9738,N_9063);
nand UO_695 (O_695,N_8989,N_8413);
nand UO_696 (O_696,N_9059,N_9711);
or UO_697 (O_697,N_9081,N_9694);
nor UO_698 (O_698,N_8735,N_9702);
nor UO_699 (O_699,N_8791,N_8000);
nand UO_700 (O_700,N_9934,N_8914);
and UO_701 (O_701,N_8845,N_8784);
nor UO_702 (O_702,N_8621,N_8411);
nand UO_703 (O_703,N_8351,N_8352);
nor UO_704 (O_704,N_9882,N_9225);
or UO_705 (O_705,N_8467,N_9558);
nand UO_706 (O_706,N_8879,N_8296);
and UO_707 (O_707,N_8442,N_9675);
or UO_708 (O_708,N_8135,N_8586);
and UO_709 (O_709,N_8384,N_9310);
or UO_710 (O_710,N_8214,N_8547);
or UO_711 (O_711,N_9080,N_9858);
and UO_712 (O_712,N_8129,N_8164);
and UO_713 (O_713,N_9754,N_8137);
nand UO_714 (O_714,N_8607,N_8779);
nor UO_715 (O_715,N_9617,N_8488);
nor UO_716 (O_716,N_9762,N_8180);
nor UO_717 (O_717,N_9493,N_9816);
nor UO_718 (O_718,N_8112,N_9111);
nor UO_719 (O_719,N_8139,N_9865);
nand UO_720 (O_720,N_8256,N_8470);
nor UO_721 (O_721,N_9885,N_9837);
nor UO_722 (O_722,N_9256,N_8560);
or UO_723 (O_723,N_9985,N_9449);
nor UO_724 (O_724,N_9314,N_8943);
nand UO_725 (O_725,N_9709,N_8367);
and UO_726 (O_726,N_8441,N_8427);
and UO_727 (O_727,N_8786,N_8276);
or UO_728 (O_728,N_8380,N_9001);
nand UO_729 (O_729,N_8347,N_9872);
nand UO_730 (O_730,N_8865,N_8755);
nand UO_731 (O_731,N_9962,N_9040);
nor UO_732 (O_732,N_9345,N_8151);
xor UO_733 (O_733,N_8549,N_8884);
and UO_734 (O_734,N_8579,N_9330);
nand UO_735 (O_735,N_9203,N_8700);
nor UO_736 (O_736,N_9945,N_9509);
or UO_737 (O_737,N_9880,N_9442);
or UO_738 (O_738,N_8211,N_8257);
nor UO_739 (O_739,N_8542,N_9290);
or UO_740 (O_740,N_8373,N_9756);
nand UO_741 (O_741,N_8923,N_9255);
xnor UO_742 (O_742,N_8327,N_9607);
or UO_743 (O_743,N_9670,N_9575);
nand UO_744 (O_744,N_8957,N_8207);
or UO_745 (O_745,N_9130,N_8155);
and UO_746 (O_746,N_8240,N_8706);
xor UO_747 (O_747,N_8292,N_9431);
or UO_748 (O_748,N_9859,N_9791);
and UO_749 (O_749,N_9078,N_8928);
and UO_750 (O_750,N_9258,N_9176);
nand UO_751 (O_751,N_9998,N_9753);
or UO_752 (O_752,N_9350,N_9982);
and UO_753 (O_753,N_9707,N_8354);
nand UO_754 (O_754,N_8886,N_9927);
and UO_755 (O_755,N_9593,N_8892);
and UO_756 (O_756,N_9775,N_9783);
or UO_757 (O_757,N_8765,N_8520);
or UO_758 (O_758,N_8315,N_9138);
and UO_759 (O_759,N_8191,N_8284);
nand UO_760 (O_760,N_8145,N_9706);
nor UO_761 (O_761,N_8158,N_9590);
nand UO_762 (O_762,N_9644,N_9713);
nor UO_763 (O_763,N_8416,N_8793);
nor UO_764 (O_764,N_9272,N_9336);
xnor UO_765 (O_765,N_8503,N_9825);
or UO_766 (O_766,N_8110,N_8773);
nand UO_767 (O_767,N_9726,N_8348);
nor UO_768 (O_768,N_9589,N_8789);
and UO_769 (O_769,N_8198,N_9156);
nand UO_770 (O_770,N_8289,N_8267);
or UO_771 (O_771,N_8839,N_8545);
or UO_772 (O_772,N_9543,N_8731);
and UO_773 (O_773,N_9925,N_9531);
or UO_774 (O_774,N_8582,N_8725);
nor UO_775 (O_775,N_9524,N_9507);
nand UO_776 (O_776,N_8620,N_9997);
xor UO_777 (O_777,N_9915,N_8093);
or UO_778 (O_778,N_9064,N_8282);
or UO_779 (O_779,N_8511,N_8859);
nand UO_780 (O_780,N_9366,N_9743);
and UO_781 (O_781,N_9903,N_8154);
and UO_782 (O_782,N_9883,N_9606);
and UO_783 (O_783,N_8376,N_9569);
nor UO_784 (O_784,N_8526,N_8443);
nor UO_785 (O_785,N_8395,N_9525);
and UO_786 (O_786,N_9124,N_8143);
nor UO_787 (O_787,N_8666,N_8942);
nor UO_788 (O_788,N_8254,N_8802);
nor UO_789 (O_789,N_8493,N_8469);
or UO_790 (O_790,N_9301,N_9614);
nor UO_791 (O_791,N_8333,N_9795);
nor UO_792 (O_792,N_8595,N_8880);
nor UO_793 (O_793,N_9849,N_8815);
xor UO_794 (O_794,N_8906,N_9075);
and UO_795 (O_795,N_9344,N_8166);
nand UO_796 (O_796,N_8307,N_8270);
nor UO_797 (O_797,N_9838,N_8669);
and UO_798 (O_798,N_9902,N_8917);
nand UO_799 (O_799,N_8357,N_9141);
and UO_800 (O_800,N_8554,N_8202);
or UO_801 (O_801,N_9395,N_8338);
or UO_802 (O_802,N_8187,N_9578);
or UO_803 (O_803,N_9955,N_9870);
and UO_804 (O_804,N_9873,N_9627);
or UO_805 (O_805,N_8497,N_8420);
and UO_806 (O_806,N_9856,N_8763);
and UO_807 (O_807,N_8447,N_9665);
nand UO_808 (O_808,N_8650,N_8102);
or UO_809 (O_809,N_9192,N_8197);
xnor UO_810 (O_810,N_8832,N_8176);
or UO_811 (O_811,N_9877,N_8604);
nor UO_812 (O_812,N_9309,N_8761);
and UO_813 (O_813,N_8787,N_8564);
and UO_814 (O_814,N_9933,N_9499);
xnor UO_815 (O_815,N_9185,N_9951);
and UO_816 (O_816,N_9438,N_9017);
nand UO_817 (O_817,N_9046,N_8662);
or UO_818 (O_818,N_9291,N_9829);
or UO_819 (O_819,N_9285,N_8106);
and UO_820 (O_820,N_8387,N_9534);
nor UO_821 (O_821,N_9018,N_8925);
nand UO_822 (O_822,N_9773,N_9163);
and UO_823 (O_823,N_9663,N_9843);
nor UO_824 (O_824,N_9091,N_9356);
nor UO_825 (O_825,N_8002,N_9282);
nor UO_826 (O_826,N_8998,N_8247);
xor UO_827 (O_827,N_8841,N_8484);
nand UO_828 (O_828,N_8967,N_9265);
nor UO_829 (O_829,N_8938,N_9471);
nand UO_830 (O_830,N_8355,N_9977);
nand UO_831 (O_831,N_9832,N_8336);
and UO_832 (O_832,N_9842,N_9110);
xnor UO_833 (O_833,N_8728,N_9928);
and UO_834 (O_834,N_8161,N_9207);
and UO_835 (O_835,N_8231,N_9871);
nand UO_836 (O_836,N_9326,N_8719);
nand UO_837 (O_837,N_8507,N_8641);
xor UO_838 (O_838,N_9618,N_9765);
nand UO_839 (O_839,N_9656,N_8283);
nand UO_840 (O_840,N_8147,N_9560);
nand UO_841 (O_841,N_8374,N_9294);
or UO_842 (O_842,N_8335,N_8130);
or UO_843 (O_843,N_9019,N_9550);
nand UO_844 (O_844,N_9879,N_9652);
nor UO_845 (O_845,N_9128,N_8864);
nor UO_846 (O_846,N_8008,N_9219);
nand UO_847 (O_847,N_8543,N_8291);
and UO_848 (O_848,N_9797,N_8473);
nor UO_849 (O_849,N_9250,N_9228);
and UO_850 (O_850,N_8072,N_9673);
xor UO_851 (O_851,N_9658,N_8933);
nor UO_852 (O_852,N_8905,N_8659);
and UO_853 (O_853,N_8812,N_8862);
or UO_854 (O_854,N_9252,N_8408);
nor UO_855 (O_855,N_9308,N_8855);
nand UO_856 (O_856,N_9952,N_9430);
xor UO_857 (O_857,N_9338,N_9038);
nand UO_858 (O_858,N_9094,N_9874);
or UO_859 (O_859,N_9764,N_9900);
nor UO_860 (O_860,N_8101,N_9662);
or UO_861 (O_861,N_8759,N_9084);
or UO_862 (O_862,N_8244,N_9506);
or UO_863 (O_863,N_8876,N_8813);
nand UO_864 (O_864,N_8253,N_8897);
or UO_865 (O_865,N_9517,N_8482);
nand UO_866 (O_866,N_9248,N_8109);
nor UO_867 (O_867,N_8829,N_8610);
nor UO_868 (O_868,N_8953,N_9237);
or UO_869 (O_869,N_9805,N_9695);
nand UO_870 (O_870,N_8790,N_8087);
nand UO_871 (O_871,N_8806,N_8435);
nor UO_872 (O_872,N_8918,N_8227);
nand UO_873 (O_873,N_8576,N_9102);
nand UO_874 (O_874,N_8322,N_8513);
or UO_875 (O_875,N_8098,N_8774);
nor UO_876 (O_876,N_9145,N_9077);
or UO_877 (O_877,N_8522,N_8094);
nor UO_878 (O_878,N_9117,N_8672);
nor UO_879 (O_879,N_9071,N_9667);
or UO_880 (O_880,N_9216,N_8431);
nand UO_881 (O_881,N_9752,N_8086);
and UO_882 (O_882,N_9121,N_8160);
and UO_883 (O_883,N_8043,N_9374);
or UO_884 (O_884,N_9386,N_8476);
nor UO_885 (O_885,N_8849,N_9823);
or UO_886 (O_886,N_9956,N_8618);
nor UO_887 (O_887,N_9457,N_9369);
nor UO_888 (O_888,N_8248,N_8397);
and UO_889 (O_889,N_9788,N_9916);
nor UO_890 (O_890,N_8205,N_8186);
or UO_891 (O_891,N_9100,N_9564);
or UO_892 (O_892,N_9579,N_8871);
nand UO_893 (O_893,N_8300,N_8758);
nor UO_894 (O_894,N_8324,N_9146);
or UO_895 (O_895,N_9643,N_9217);
or UO_896 (O_896,N_8175,N_8487);
or UO_897 (O_897,N_8775,N_8617);
or UO_898 (O_898,N_9759,N_8423);
and UO_899 (O_899,N_8995,N_9287);
or UO_900 (O_900,N_8314,N_9347);
xnor UO_901 (O_901,N_8817,N_8930);
or UO_902 (O_902,N_9451,N_8660);
and UO_903 (O_903,N_9495,N_8708);
nor UO_904 (O_904,N_9421,N_8645);
nand UO_905 (O_905,N_8818,N_9118);
nand UO_906 (O_906,N_9541,N_9528);
nor UO_907 (O_907,N_9115,N_9615);
nor UO_908 (O_908,N_9151,N_9905);
or UO_909 (O_909,N_8342,N_9231);
nand UO_910 (O_910,N_9959,N_9474);
or UO_911 (O_911,N_9794,N_8999);
or UO_912 (O_912,N_8042,N_9042);
nor UO_913 (O_913,N_8842,N_9970);
nand UO_914 (O_914,N_8111,N_9582);
nor UO_915 (O_915,N_9776,N_8640);
or UO_916 (O_916,N_8518,N_8903);
nand UO_917 (O_917,N_9609,N_8857);
nand UO_918 (O_918,N_9799,N_9157);
nor UO_919 (O_919,N_8875,N_9413);
and UO_920 (O_920,N_9307,N_9292);
nor UO_921 (O_921,N_9494,N_9093);
nor UO_922 (O_922,N_8626,N_8181);
nand UO_923 (O_923,N_9406,N_9193);
nand UO_924 (O_924,N_8273,N_9770);
nand UO_925 (O_925,N_9012,N_8414);
and UO_926 (O_926,N_8039,N_8134);
nand UO_927 (O_927,N_8304,N_8688);
or UO_928 (O_928,N_9599,N_9168);
nor UO_929 (O_929,N_8142,N_9401);
nor UO_930 (O_930,N_8685,N_8721);
nand UO_931 (O_931,N_9518,N_9417);
or UO_932 (O_932,N_8594,N_8768);
and UO_933 (O_933,N_9172,N_9464);
nor UO_934 (O_934,N_8359,N_9021);
and UO_935 (O_935,N_9526,N_8978);
or UO_936 (O_936,N_9305,N_8835);
and UO_937 (O_937,N_8567,N_8588);
and UO_938 (O_938,N_9177,N_8330);
nand UO_939 (O_939,N_9688,N_8030);
or UO_940 (O_940,N_9931,N_8394);
and UO_941 (O_941,N_9844,N_8429);
nor UO_942 (O_942,N_8399,N_8703);
nand UO_943 (O_943,N_9422,N_8986);
and UO_944 (O_944,N_8811,N_8188);
nand UO_945 (O_945,N_9048,N_8954);
nand UO_946 (O_946,N_9807,N_8973);
nand UO_947 (O_947,N_9750,N_9426);
nor UO_948 (O_948,N_9088,N_8766);
and UO_949 (O_949,N_8310,N_8038);
nand UO_950 (O_950,N_8623,N_8872);
or UO_951 (O_951,N_8523,N_9633);
nor UO_952 (O_952,N_8334,N_9685);
or UO_953 (O_953,N_9836,N_8606);
nor UO_954 (O_954,N_8907,N_9661);
or UO_955 (O_955,N_8678,N_8683);
nand UO_956 (O_956,N_9459,N_9478);
or UO_957 (O_957,N_9236,N_9007);
nor UO_958 (O_958,N_9512,N_9801);
nand UO_959 (O_959,N_9273,N_9819);
nand UO_960 (O_960,N_9149,N_8992);
and UO_961 (O_961,N_8733,N_9553);
and UO_962 (O_962,N_9777,N_9053);
nand UO_963 (O_963,N_9215,N_9610);
and UO_964 (O_964,N_9416,N_8498);
nand UO_965 (O_965,N_8792,N_9333);
nor UO_966 (O_966,N_9800,N_8772);
and UO_967 (O_967,N_9497,N_8713);
nand UO_968 (O_968,N_8537,N_9279);
or UO_969 (O_969,N_8944,N_8742);
and UO_970 (O_970,N_8415,N_8029);
nand UO_971 (O_971,N_9647,N_9544);
or UO_972 (O_972,N_8152,N_9032);
or UO_973 (O_973,N_8255,N_8438);
nand UO_974 (O_974,N_8945,N_9683);
nand UO_975 (O_975,N_9353,N_9979);
and UO_976 (O_976,N_8717,N_8326);
and UO_977 (O_977,N_9887,N_8751);
or UO_978 (O_978,N_8889,N_9316);
and UO_979 (O_979,N_9433,N_9208);
or UO_980 (O_980,N_9901,N_8738);
nor UO_981 (O_981,N_9069,N_8847);
nand UO_982 (O_982,N_9496,N_8831);
nand UO_983 (O_983,N_9367,N_8535);
and UO_984 (O_984,N_8727,N_8454);
or UO_985 (O_985,N_8345,N_9864);
and UO_986 (O_986,N_9489,N_9006);
or UO_987 (O_987,N_8991,N_9060);
or UO_988 (O_988,N_9944,N_8823);
or UO_989 (O_989,N_8783,N_8515);
nor UO_990 (O_990,N_9587,N_8120);
nand UO_991 (O_991,N_9161,N_8516);
nor UO_992 (O_992,N_9412,N_8544);
and UO_993 (O_993,N_8926,N_8878);
nor UO_994 (O_994,N_8051,N_8757);
or UO_995 (O_995,N_8600,N_9991);
or UO_996 (O_996,N_9342,N_9180);
and UO_997 (O_997,N_8950,N_8794);
and UO_998 (O_998,N_9642,N_9923);
and UO_999 (O_999,N_8502,N_8762);
nand UO_1000 (O_1000,N_8931,N_9155);
and UO_1001 (O_1001,N_8350,N_9760);
nor UO_1002 (O_1002,N_8292,N_8253);
or UO_1003 (O_1003,N_9823,N_9006);
nor UO_1004 (O_1004,N_8361,N_8271);
xor UO_1005 (O_1005,N_8213,N_9235);
and UO_1006 (O_1006,N_9166,N_8929);
nor UO_1007 (O_1007,N_9694,N_8236);
and UO_1008 (O_1008,N_9771,N_9417);
nand UO_1009 (O_1009,N_8347,N_8837);
or UO_1010 (O_1010,N_8328,N_8735);
nor UO_1011 (O_1011,N_8685,N_8507);
and UO_1012 (O_1012,N_8161,N_9993);
or UO_1013 (O_1013,N_9420,N_9627);
nor UO_1014 (O_1014,N_8959,N_8183);
and UO_1015 (O_1015,N_8459,N_8054);
or UO_1016 (O_1016,N_8819,N_8924);
and UO_1017 (O_1017,N_9173,N_8455);
and UO_1018 (O_1018,N_8177,N_8542);
nand UO_1019 (O_1019,N_8654,N_8278);
nor UO_1020 (O_1020,N_8912,N_8643);
or UO_1021 (O_1021,N_9123,N_9043);
nand UO_1022 (O_1022,N_8875,N_8858);
nand UO_1023 (O_1023,N_9773,N_8661);
nand UO_1024 (O_1024,N_9008,N_8325);
nor UO_1025 (O_1025,N_9153,N_9430);
nor UO_1026 (O_1026,N_9507,N_9015);
or UO_1027 (O_1027,N_8518,N_9474);
nor UO_1028 (O_1028,N_8728,N_9952);
nor UO_1029 (O_1029,N_8397,N_8533);
and UO_1030 (O_1030,N_9561,N_8741);
or UO_1031 (O_1031,N_8345,N_8269);
nor UO_1032 (O_1032,N_8967,N_9473);
and UO_1033 (O_1033,N_9382,N_8233);
nand UO_1034 (O_1034,N_8547,N_8591);
nand UO_1035 (O_1035,N_8955,N_8905);
or UO_1036 (O_1036,N_8644,N_9633);
and UO_1037 (O_1037,N_9957,N_9771);
and UO_1038 (O_1038,N_8266,N_8114);
or UO_1039 (O_1039,N_9687,N_9567);
nor UO_1040 (O_1040,N_8996,N_9706);
or UO_1041 (O_1041,N_9309,N_9420);
and UO_1042 (O_1042,N_9363,N_8668);
nor UO_1043 (O_1043,N_8295,N_8278);
nor UO_1044 (O_1044,N_8773,N_8148);
or UO_1045 (O_1045,N_8183,N_8031);
nor UO_1046 (O_1046,N_8663,N_9191);
nor UO_1047 (O_1047,N_9038,N_8456);
and UO_1048 (O_1048,N_8278,N_9528);
or UO_1049 (O_1049,N_9929,N_9156);
nor UO_1050 (O_1050,N_8870,N_8994);
and UO_1051 (O_1051,N_9739,N_9048);
and UO_1052 (O_1052,N_9577,N_8992);
nand UO_1053 (O_1053,N_9775,N_9716);
nor UO_1054 (O_1054,N_8718,N_9932);
xor UO_1055 (O_1055,N_9051,N_9194);
nor UO_1056 (O_1056,N_8647,N_9167);
nand UO_1057 (O_1057,N_8684,N_8890);
nand UO_1058 (O_1058,N_9788,N_9404);
or UO_1059 (O_1059,N_8303,N_8720);
nand UO_1060 (O_1060,N_8814,N_8883);
nand UO_1061 (O_1061,N_8820,N_9463);
or UO_1062 (O_1062,N_8805,N_8589);
nand UO_1063 (O_1063,N_9351,N_9525);
nand UO_1064 (O_1064,N_9164,N_8564);
or UO_1065 (O_1065,N_9763,N_9919);
and UO_1066 (O_1066,N_8421,N_9612);
and UO_1067 (O_1067,N_9759,N_9610);
nand UO_1068 (O_1068,N_8748,N_8590);
nand UO_1069 (O_1069,N_8846,N_9931);
nand UO_1070 (O_1070,N_9035,N_9946);
nor UO_1071 (O_1071,N_8839,N_9380);
nor UO_1072 (O_1072,N_8281,N_9511);
nand UO_1073 (O_1073,N_8088,N_9426);
or UO_1074 (O_1074,N_8438,N_9632);
nor UO_1075 (O_1075,N_9344,N_9555);
nand UO_1076 (O_1076,N_8895,N_8196);
and UO_1077 (O_1077,N_8228,N_8051);
or UO_1078 (O_1078,N_8301,N_9101);
or UO_1079 (O_1079,N_8948,N_9681);
nor UO_1080 (O_1080,N_8829,N_9533);
or UO_1081 (O_1081,N_8519,N_8167);
and UO_1082 (O_1082,N_9362,N_8476);
nor UO_1083 (O_1083,N_9993,N_9376);
or UO_1084 (O_1084,N_9134,N_9184);
nand UO_1085 (O_1085,N_9564,N_9639);
or UO_1086 (O_1086,N_9571,N_9104);
nor UO_1087 (O_1087,N_9071,N_8953);
and UO_1088 (O_1088,N_9759,N_8645);
and UO_1089 (O_1089,N_9808,N_8227);
or UO_1090 (O_1090,N_9070,N_9153);
nand UO_1091 (O_1091,N_8144,N_9454);
and UO_1092 (O_1092,N_9500,N_8035);
or UO_1093 (O_1093,N_9078,N_8020);
nand UO_1094 (O_1094,N_8186,N_8015);
and UO_1095 (O_1095,N_9485,N_8392);
nand UO_1096 (O_1096,N_8918,N_9002);
nand UO_1097 (O_1097,N_8638,N_8554);
nand UO_1098 (O_1098,N_9420,N_9580);
xnor UO_1099 (O_1099,N_9806,N_8046);
nand UO_1100 (O_1100,N_8674,N_8657);
nand UO_1101 (O_1101,N_9659,N_8051);
or UO_1102 (O_1102,N_9918,N_8067);
or UO_1103 (O_1103,N_8529,N_9957);
nand UO_1104 (O_1104,N_8301,N_9581);
or UO_1105 (O_1105,N_9016,N_9655);
or UO_1106 (O_1106,N_9973,N_9941);
nand UO_1107 (O_1107,N_9457,N_9589);
and UO_1108 (O_1108,N_8965,N_9922);
nand UO_1109 (O_1109,N_9243,N_8397);
and UO_1110 (O_1110,N_8655,N_9356);
and UO_1111 (O_1111,N_8151,N_9902);
nand UO_1112 (O_1112,N_8372,N_9755);
nand UO_1113 (O_1113,N_9054,N_9702);
nor UO_1114 (O_1114,N_9942,N_9443);
nor UO_1115 (O_1115,N_9153,N_8528);
nand UO_1116 (O_1116,N_8332,N_9065);
xnor UO_1117 (O_1117,N_9970,N_9153);
and UO_1118 (O_1118,N_8324,N_9867);
or UO_1119 (O_1119,N_8594,N_8736);
xor UO_1120 (O_1120,N_8032,N_9939);
or UO_1121 (O_1121,N_8857,N_8449);
xnor UO_1122 (O_1122,N_9154,N_8431);
and UO_1123 (O_1123,N_9912,N_9399);
nor UO_1124 (O_1124,N_9692,N_9343);
and UO_1125 (O_1125,N_8556,N_9615);
nor UO_1126 (O_1126,N_9643,N_8612);
nor UO_1127 (O_1127,N_8237,N_8038);
and UO_1128 (O_1128,N_9420,N_9079);
nand UO_1129 (O_1129,N_8995,N_8698);
or UO_1130 (O_1130,N_9516,N_9595);
nor UO_1131 (O_1131,N_9636,N_8135);
and UO_1132 (O_1132,N_8221,N_8627);
and UO_1133 (O_1133,N_8540,N_9530);
nand UO_1134 (O_1134,N_8012,N_8831);
nor UO_1135 (O_1135,N_9713,N_9947);
nor UO_1136 (O_1136,N_8756,N_9484);
nand UO_1137 (O_1137,N_9345,N_8956);
and UO_1138 (O_1138,N_9234,N_8365);
and UO_1139 (O_1139,N_9374,N_8786);
nand UO_1140 (O_1140,N_8470,N_8292);
or UO_1141 (O_1141,N_9267,N_8819);
nor UO_1142 (O_1142,N_8904,N_8255);
nand UO_1143 (O_1143,N_8588,N_8428);
nor UO_1144 (O_1144,N_8988,N_8067);
nor UO_1145 (O_1145,N_9600,N_9361);
nand UO_1146 (O_1146,N_9700,N_9075);
and UO_1147 (O_1147,N_8382,N_8915);
or UO_1148 (O_1148,N_8942,N_9299);
nand UO_1149 (O_1149,N_9054,N_8215);
nor UO_1150 (O_1150,N_8439,N_9850);
nor UO_1151 (O_1151,N_9595,N_8518);
nand UO_1152 (O_1152,N_9194,N_9946);
or UO_1153 (O_1153,N_9213,N_9252);
and UO_1154 (O_1154,N_8623,N_8439);
nand UO_1155 (O_1155,N_9966,N_8900);
nor UO_1156 (O_1156,N_9828,N_8196);
nor UO_1157 (O_1157,N_8488,N_9918);
nor UO_1158 (O_1158,N_9408,N_8676);
nor UO_1159 (O_1159,N_9275,N_9213);
and UO_1160 (O_1160,N_9118,N_9665);
nor UO_1161 (O_1161,N_9282,N_9891);
or UO_1162 (O_1162,N_9370,N_9351);
nor UO_1163 (O_1163,N_8634,N_8774);
nor UO_1164 (O_1164,N_8834,N_8763);
nor UO_1165 (O_1165,N_8339,N_9497);
nor UO_1166 (O_1166,N_9549,N_8944);
or UO_1167 (O_1167,N_8989,N_9263);
or UO_1168 (O_1168,N_8994,N_9623);
nor UO_1169 (O_1169,N_9373,N_8917);
and UO_1170 (O_1170,N_8789,N_9280);
nand UO_1171 (O_1171,N_9013,N_9497);
nor UO_1172 (O_1172,N_8773,N_8014);
xor UO_1173 (O_1173,N_9556,N_8324);
or UO_1174 (O_1174,N_8667,N_8434);
or UO_1175 (O_1175,N_9619,N_9909);
and UO_1176 (O_1176,N_9408,N_8779);
and UO_1177 (O_1177,N_9015,N_8980);
nand UO_1178 (O_1178,N_8254,N_8036);
xor UO_1179 (O_1179,N_9107,N_8221);
and UO_1180 (O_1180,N_8568,N_9347);
or UO_1181 (O_1181,N_8850,N_8256);
nor UO_1182 (O_1182,N_9780,N_9865);
nand UO_1183 (O_1183,N_9018,N_9346);
nor UO_1184 (O_1184,N_8165,N_9872);
or UO_1185 (O_1185,N_9556,N_9673);
nor UO_1186 (O_1186,N_8510,N_8839);
or UO_1187 (O_1187,N_9349,N_9529);
or UO_1188 (O_1188,N_9608,N_8736);
nor UO_1189 (O_1189,N_9136,N_9646);
nand UO_1190 (O_1190,N_9967,N_9882);
nor UO_1191 (O_1191,N_8674,N_8018);
and UO_1192 (O_1192,N_8090,N_9392);
nand UO_1193 (O_1193,N_9338,N_9630);
and UO_1194 (O_1194,N_9694,N_8283);
or UO_1195 (O_1195,N_8097,N_9626);
and UO_1196 (O_1196,N_9396,N_8174);
and UO_1197 (O_1197,N_8887,N_8562);
nand UO_1198 (O_1198,N_9000,N_9618);
or UO_1199 (O_1199,N_8104,N_8893);
nand UO_1200 (O_1200,N_8668,N_8580);
nand UO_1201 (O_1201,N_9676,N_8783);
and UO_1202 (O_1202,N_8010,N_8638);
nand UO_1203 (O_1203,N_8661,N_9881);
or UO_1204 (O_1204,N_8451,N_9522);
and UO_1205 (O_1205,N_8650,N_8754);
and UO_1206 (O_1206,N_9411,N_8853);
nor UO_1207 (O_1207,N_8860,N_8856);
or UO_1208 (O_1208,N_9849,N_8537);
nand UO_1209 (O_1209,N_8323,N_9236);
and UO_1210 (O_1210,N_9367,N_9399);
nor UO_1211 (O_1211,N_9250,N_9104);
or UO_1212 (O_1212,N_9289,N_9699);
nand UO_1213 (O_1213,N_9680,N_8738);
xor UO_1214 (O_1214,N_8295,N_8444);
nor UO_1215 (O_1215,N_8495,N_8823);
nand UO_1216 (O_1216,N_8895,N_9582);
nor UO_1217 (O_1217,N_9489,N_9142);
and UO_1218 (O_1218,N_9917,N_9013);
nor UO_1219 (O_1219,N_9248,N_8793);
nor UO_1220 (O_1220,N_9700,N_8608);
and UO_1221 (O_1221,N_9493,N_8275);
nor UO_1222 (O_1222,N_9343,N_9896);
nand UO_1223 (O_1223,N_9365,N_9526);
and UO_1224 (O_1224,N_9277,N_8033);
and UO_1225 (O_1225,N_8114,N_9582);
xor UO_1226 (O_1226,N_9865,N_9307);
or UO_1227 (O_1227,N_8541,N_8680);
nor UO_1228 (O_1228,N_9171,N_9445);
or UO_1229 (O_1229,N_8875,N_9488);
nand UO_1230 (O_1230,N_8444,N_9150);
nor UO_1231 (O_1231,N_8394,N_9083);
nand UO_1232 (O_1232,N_8260,N_9852);
nor UO_1233 (O_1233,N_9034,N_9880);
and UO_1234 (O_1234,N_9367,N_9324);
or UO_1235 (O_1235,N_9840,N_9119);
nand UO_1236 (O_1236,N_9973,N_8039);
nand UO_1237 (O_1237,N_8135,N_8753);
or UO_1238 (O_1238,N_9114,N_9816);
nor UO_1239 (O_1239,N_8982,N_9590);
and UO_1240 (O_1240,N_9699,N_8875);
nor UO_1241 (O_1241,N_9967,N_8352);
and UO_1242 (O_1242,N_8990,N_9434);
nand UO_1243 (O_1243,N_8186,N_8782);
nand UO_1244 (O_1244,N_8855,N_9728);
and UO_1245 (O_1245,N_9542,N_9531);
nand UO_1246 (O_1246,N_9576,N_9925);
nand UO_1247 (O_1247,N_8713,N_8366);
nor UO_1248 (O_1248,N_8544,N_9031);
xnor UO_1249 (O_1249,N_8248,N_8952);
and UO_1250 (O_1250,N_8689,N_9116);
nand UO_1251 (O_1251,N_8644,N_9151);
nor UO_1252 (O_1252,N_9608,N_8907);
nand UO_1253 (O_1253,N_8822,N_8289);
nand UO_1254 (O_1254,N_8453,N_9343);
or UO_1255 (O_1255,N_9663,N_9528);
nand UO_1256 (O_1256,N_8706,N_8095);
xnor UO_1257 (O_1257,N_8584,N_9851);
nor UO_1258 (O_1258,N_9391,N_8928);
nor UO_1259 (O_1259,N_9626,N_9245);
or UO_1260 (O_1260,N_9021,N_9160);
or UO_1261 (O_1261,N_8319,N_8376);
nand UO_1262 (O_1262,N_9390,N_8618);
or UO_1263 (O_1263,N_8617,N_9093);
nor UO_1264 (O_1264,N_9823,N_8853);
nor UO_1265 (O_1265,N_8700,N_8285);
nand UO_1266 (O_1266,N_9582,N_8369);
or UO_1267 (O_1267,N_8386,N_8575);
and UO_1268 (O_1268,N_8335,N_8838);
nor UO_1269 (O_1269,N_8926,N_8438);
nor UO_1270 (O_1270,N_8292,N_8081);
nand UO_1271 (O_1271,N_9220,N_9633);
nand UO_1272 (O_1272,N_8841,N_8136);
or UO_1273 (O_1273,N_8778,N_8236);
nand UO_1274 (O_1274,N_9785,N_9061);
nor UO_1275 (O_1275,N_9932,N_8273);
and UO_1276 (O_1276,N_9584,N_8010);
nor UO_1277 (O_1277,N_8891,N_9584);
nand UO_1278 (O_1278,N_8794,N_8718);
nand UO_1279 (O_1279,N_9364,N_9862);
xnor UO_1280 (O_1280,N_9484,N_9874);
or UO_1281 (O_1281,N_8657,N_8924);
nand UO_1282 (O_1282,N_9230,N_9192);
or UO_1283 (O_1283,N_9471,N_8046);
nor UO_1284 (O_1284,N_8306,N_8205);
or UO_1285 (O_1285,N_8047,N_8067);
nor UO_1286 (O_1286,N_8773,N_8162);
nor UO_1287 (O_1287,N_9374,N_9391);
and UO_1288 (O_1288,N_9230,N_9029);
nor UO_1289 (O_1289,N_9158,N_9215);
nand UO_1290 (O_1290,N_8560,N_8279);
or UO_1291 (O_1291,N_9117,N_9977);
or UO_1292 (O_1292,N_8811,N_9050);
or UO_1293 (O_1293,N_8555,N_9471);
nor UO_1294 (O_1294,N_8534,N_9257);
and UO_1295 (O_1295,N_8223,N_9401);
nor UO_1296 (O_1296,N_9207,N_9124);
xnor UO_1297 (O_1297,N_8487,N_9817);
and UO_1298 (O_1298,N_9990,N_9900);
nand UO_1299 (O_1299,N_8630,N_9276);
or UO_1300 (O_1300,N_9638,N_8764);
or UO_1301 (O_1301,N_8573,N_8490);
nand UO_1302 (O_1302,N_8040,N_9547);
nor UO_1303 (O_1303,N_8540,N_9775);
nand UO_1304 (O_1304,N_8579,N_9624);
and UO_1305 (O_1305,N_9708,N_8560);
nor UO_1306 (O_1306,N_8957,N_9549);
and UO_1307 (O_1307,N_8701,N_8233);
and UO_1308 (O_1308,N_9333,N_9595);
nor UO_1309 (O_1309,N_9488,N_8742);
nor UO_1310 (O_1310,N_9277,N_8748);
or UO_1311 (O_1311,N_8313,N_8719);
or UO_1312 (O_1312,N_9603,N_9561);
nand UO_1313 (O_1313,N_8991,N_9106);
nor UO_1314 (O_1314,N_9551,N_8577);
nand UO_1315 (O_1315,N_8735,N_8618);
or UO_1316 (O_1316,N_8558,N_9167);
nand UO_1317 (O_1317,N_9925,N_8690);
and UO_1318 (O_1318,N_8838,N_9243);
nor UO_1319 (O_1319,N_9944,N_8598);
and UO_1320 (O_1320,N_9060,N_9721);
nor UO_1321 (O_1321,N_8853,N_9163);
nor UO_1322 (O_1322,N_9845,N_8564);
nor UO_1323 (O_1323,N_8424,N_8666);
nor UO_1324 (O_1324,N_9148,N_8012);
nand UO_1325 (O_1325,N_9955,N_8420);
or UO_1326 (O_1326,N_8995,N_8379);
nor UO_1327 (O_1327,N_8114,N_8696);
nand UO_1328 (O_1328,N_8267,N_8186);
nand UO_1329 (O_1329,N_9151,N_8145);
nor UO_1330 (O_1330,N_8079,N_8117);
nand UO_1331 (O_1331,N_9502,N_8771);
or UO_1332 (O_1332,N_9958,N_9520);
or UO_1333 (O_1333,N_8249,N_8206);
or UO_1334 (O_1334,N_8558,N_9545);
nor UO_1335 (O_1335,N_9065,N_8002);
nor UO_1336 (O_1336,N_8721,N_8460);
or UO_1337 (O_1337,N_9259,N_8535);
and UO_1338 (O_1338,N_9667,N_8380);
and UO_1339 (O_1339,N_8126,N_9305);
nor UO_1340 (O_1340,N_9800,N_8578);
nor UO_1341 (O_1341,N_9539,N_9004);
or UO_1342 (O_1342,N_9745,N_9192);
and UO_1343 (O_1343,N_8808,N_8878);
nor UO_1344 (O_1344,N_9685,N_8143);
nor UO_1345 (O_1345,N_9016,N_8418);
or UO_1346 (O_1346,N_8870,N_9608);
or UO_1347 (O_1347,N_8668,N_9433);
and UO_1348 (O_1348,N_8130,N_9289);
and UO_1349 (O_1349,N_8438,N_9146);
and UO_1350 (O_1350,N_9105,N_9467);
nor UO_1351 (O_1351,N_9022,N_8365);
nor UO_1352 (O_1352,N_8005,N_9439);
or UO_1353 (O_1353,N_9390,N_9434);
or UO_1354 (O_1354,N_8804,N_9389);
nand UO_1355 (O_1355,N_9081,N_9221);
nor UO_1356 (O_1356,N_9243,N_9050);
nand UO_1357 (O_1357,N_8865,N_9019);
and UO_1358 (O_1358,N_8852,N_9631);
nor UO_1359 (O_1359,N_9515,N_8503);
and UO_1360 (O_1360,N_8860,N_8302);
nand UO_1361 (O_1361,N_8972,N_8952);
nor UO_1362 (O_1362,N_8507,N_9192);
nand UO_1363 (O_1363,N_9966,N_8490);
nand UO_1364 (O_1364,N_9184,N_8499);
nand UO_1365 (O_1365,N_8335,N_9293);
and UO_1366 (O_1366,N_9985,N_8653);
and UO_1367 (O_1367,N_8661,N_8696);
or UO_1368 (O_1368,N_9811,N_8355);
nor UO_1369 (O_1369,N_8623,N_9242);
or UO_1370 (O_1370,N_9391,N_8404);
nor UO_1371 (O_1371,N_9108,N_9677);
nor UO_1372 (O_1372,N_8773,N_9298);
nand UO_1373 (O_1373,N_8608,N_8917);
or UO_1374 (O_1374,N_9951,N_9901);
or UO_1375 (O_1375,N_8758,N_9614);
and UO_1376 (O_1376,N_8672,N_9691);
or UO_1377 (O_1377,N_8329,N_8270);
nor UO_1378 (O_1378,N_9208,N_8299);
and UO_1379 (O_1379,N_9418,N_8857);
and UO_1380 (O_1380,N_9764,N_9272);
and UO_1381 (O_1381,N_8449,N_9806);
nand UO_1382 (O_1382,N_9494,N_8429);
nand UO_1383 (O_1383,N_9715,N_9419);
or UO_1384 (O_1384,N_8211,N_9052);
and UO_1385 (O_1385,N_9654,N_8979);
and UO_1386 (O_1386,N_9171,N_9316);
or UO_1387 (O_1387,N_8070,N_9504);
nor UO_1388 (O_1388,N_8894,N_8950);
or UO_1389 (O_1389,N_8422,N_9354);
xor UO_1390 (O_1390,N_8556,N_8849);
and UO_1391 (O_1391,N_8686,N_9412);
nand UO_1392 (O_1392,N_9220,N_9519);
nor UO_1393 (O_1393,N_9445,N_8178);
nor UO_1394 (O_1394,N_9329,N_8470);
xor UO_1395 (O_1395,N_9000,N_8316);
and UO_1396 (O_1396,N_8219,N_8628);
nor UO_1397 (O_1397,N_9993,N_9718);
and UO_1398 (O_1398,N_8712,N_8063);
and UO_1399 (O_1399,N_8634,N_8914);
nand UO_1400 (O_1400,N_8571,N_8252);
and UO_1401 (O_1401,N_8996,N_9520);
nand UO_1402 (O_1402,N_9765,N_8436);
nor UO_1403 (O_1403,N_8145,N_8961);
nand UO_1404 (O_1404,N_9946,N_9457);
and UO_1405 (O_1405,N_8383,N_8303);
nor UO_1406 (O_1406,N_8707,N_8151);
or UO_1407 (O_1407,N_8902,N_8052);
or UO_1408 (O_1408,N_8602,N_9087);
and UO_1409 (O_1409,N_8191,N_8081);
nand UO_1410 (O_1410,N_8943,N_8651);
nand UO_1411 (O_1411,N_8287,N_9051);
xor UO_1412 (O_1412,N_8999,N_8740);
nand UO_1413 (O_1413,N_9612,N_9820);
nand UO_1414 (O_1414,N_9110,N_8449);
and UO_1415 (O_1415,N_9774,N_8034);
nor UO_1416 (O_1416,N_8542,N_9957);
or UO_1417 (O_1417,N_9713,N_9476);
and UO_1418 (O_1418,N_8345,N_9618);
nor UO_1419 (O_1419,N_8663,N_9124);
nor UO_1420 (O_1420,N_8241,N_8955);
and UO_1421 (O_1421,N_8399,N_9492);
or UO_1422 (O_1422,N_9777,N_8798);
and UO_1423 (O_1423,N_8076,N_8743);
nor UO_1424 (O_1424,N_9665,N_9872);
or UO_1425 (O_1425,N_8344,N_9951);
nand UO_1426 (O_1426,N_9469,N_8904);
nor UO_1427 (O_1427,N_9567,N_9249);
or UO_1428 (O_1428,N_9557,N_8578);
and UO_1429 (O_1429,N_8459,N_8047);
nor UO_1430 (O_1430,N_8776,N_9152);
or UO_1431 (O_1431,N_9082,N_9728);
nor UO_1432 (O_1432,N_9873,N_8190);
nand UO_1433 (O_1433,N_9914,N_8759);
xnor UO_1434 (O_1434,N_8798,N_9724);
xnor UO_1435 (O_1435,N_9636,N_9852);
or UO_1436 (O_1436,N_9126,N_8841);
and UO_1437 (O_1437,N_8684,N_8047);
and UO_1438 (O_1438,N_8233,N_8122);
or UO_1439 (O_1439,N_9927,N_8347);
and UO_1440 (O_1440,N_8966,N_9814);
and UO_1441 (O_1441,N_8871,N_8777);
or UO_1442 (O_1442,N_9962,N_9275);
nand UO_1443 (O_1443,N_9039,N_8717);
and UO_1444 (O_1444,N_8668,N_9622);
or UO_1445 (O_1445,N_9687,N_8197);
xnor UO_1446 (O_1446,N_9797,N_8802);
nor UO_1447 (O_1447,N_9574,N_9673);
nor UO_1448 (O_1448,N_8270,N_8636);
or UO_1449 (O_1449,N_9479,N_8212);
nor UO_1450 (O_1450,N_8617,N_9678);
nor UO_1451 (O_1451,N_9511,N_8770);
nand UO_1452 (O_1452,N_9075,N_8701);
or UO_1453 (O_1453,N_8160,N_9420);
nand UO_1454 (O_1454,N_9965,N_9333);
nor UO_1455 (O_1455,N_8541,N_9245);
and UO_1456 (O_1456,N_8884,N_9657);
nor UO_1457 (O_1457,N_8016,N_9676);
or UO_1458 (O_1458,N_9920,N_9049);
nand UO_1459 (O_1459,N_8916,N_8448);
or UO_1460 (O_1460,N_9051,N_9670);
nor UO_1461 (O_1461,N_8767,N_8897);
nand UO_1462 (O_1462,N_9370,N_8310);
nand UO_1463 (O_1463,N_8928,N_8139);
nand UO_1464 (O_1464,N_8054,N_8754);
xnor UO_1465 (O_1465,N_8456,N_8948);
or UO_1466 (O_1466,N_9877,N_9234);
nand UO_1467 (O_1467,N_8600,N_9381);
and UO_1468 (O_1468,N_8784,N_8861);
nand UO_1469 (O_1469,N_9029,N_8125);
nand UO_1470 (O_1470,N_8573,N_8084);
or UO_1471 (O_1471,N_9903,N_9430);
nor UO_1472 (O_1472,N_8821,N_9989);
nand UO_1473 (O_1473,N_9766,N_9558);
nor UO_1474 (O_1474,N_9673,N_9006);
nor UO_1475 (O_1475,N_9749,N_9332);
nor UO_1476 (O_1476,N_9347,N_8939);
nand UO_1477 (O_1477,N_8532,N_9288);
and UO_1478 (O_1478,N_9705,N_8033);
xor UO_1479 (O_1479,N_9099,N_9886);
or UO_1480 (O_1480,N_8993,N_9419);
or UO_1481 (O_1481,N_8996,N_8348);
or UO_1482 (O_1482,N_8183,N_9602);
and UO_1483 (O_1483,N_9382,N_9073);
nand UO_1484 (O_1484,N_8103,N_9105);
nand UO_1485 (O_1485,N_9221,N_9461);
or UO_1486 (O_1486,N_9407,N_9842);
nand UO_1487 (O_1487,N_8790,N_9289);
nand UO_1488 (O_1488,N_8500,N_8995);
nand UO_1489 (O_1489,N_9811,N_8856);
or UO_1490 (O_1490,N_8022,N_9240);
nand UO_1491 (O_1491,N_8757,N_8929);
nor UO_1492 (O_1492,N_8635,N_9734);
nor UO_1493 (O_1493,N_9294,N_8528);
nand UO_1494 (O_1494,N_8962,N_9102);
or UO_1495 (O_1495,N_8427,N_9465);
nand UO_1496 (O_1496,N_8106,N_9719);
or UO_1497 (O_1497,N_9089,N_8680);
nor UO_1498 (O_1498,N_9253,N_9625);
nor UO_1499 (O_1499,N_8942,N_9718);
endmodule